magic
tech sky130A
magscale 1 2
timestamp 1746348191
<< pwell >>
rect 1350 1187 2690 1340
rect 1350 153 1503 1187
rect 2537 153 2690 1187
rect 1350 0 2690 153
rect 2710 1187 4050 1340
rect 2710 153 2863 1187
rect 3897 153 4050 1187
rect 2710 0 4050 153
rect 4070 1187 5410 1340
rect 4070 153 4223 1187
rect 5257 153 5410 1187
rect 4070 0 5410 153
rect 5430 1187 6770 1340
rect 5430 153 5583 1187
rect 6617 153 6770 1187
rect 5430 0 6770 153
rect 6790 1187 8130 1340
rect 6790 153 6943 1187
rect 7977 153 8130 1187
rect 6790 0 8130 153
rect 8150 1187 9490 1340
rect 8150 153 8303 1187
rect 9337 153 9490 1187
rect 8150 0 9490 153
<< nbase >>
rect 1503 153 2537 1187
rect 2863 153 3897 1187
rect 4223 153 5257 1187
rect 5583 153 6617 1187
rect 6943 153 7977 1187
rect 8303 153 9337 1187
<< nmos >>
rect 4490 4360 4610 5160
rect 4690 4360 4810 5160
rect 4890 4360 5010 5160
rect 5090 4360 5210 5160
rect 5290 4360 5410 5160
rect 5490 4360 5610 5160
rect 5690 4360 5810 5160
rect 5890 4360 6010 5160
rect 6090 4360 6210 5160
rect 6290 4360 6410 5160
rect 6490 4360 6610 5160
rect 6690 4360 6810 5160
rect 6890 4360 7010 5160
rect 7090 4360 7210 5160
rect 7290 4360 7410 5160
rect 7490 4360 7610 5160
rect 7690 4360 7810 5160
rect 7890 4360 8010 5160
rect 8090 4360 8210 5160
rect 8290 4360 8410 5160
rect 10410 3960 10440 4360
rect 10660 3960 10690 4360
rect 4530 3450 4650 3850
rect 4730 3450 4850 3850
rect 4930 3450 5050 3850
rect 5130 3450 5250 3850
rect 5330 3450 5450 3850
rect 5530 3450 5650 3850
rect 5890 3450 6010 3850
rect 6090 3450 6210 3850
rect 6290 3450 6410 3850
rect 6490 3450 6610 3850
rect 6690 3450 6810 3850
rect 6890 3450 7010 3850
rect 7250 3450 7370 3850
rect 7450 3450 7570 3850
rect 7650 3450 7770 3850
rect 7850 3450 7970 3850
rect 8050 3450 8170 3850
rect 8250 3450 8370 3850
rect 9290 3460 11290 3660
rect 5210 2840 5330 3040
rect 5410 2840 5530 3040
rect 5610 2840 5730 3040
rect 5810 2840 5930 3040
rect 6010 2840 6130 3040
rect 6210 2840 6330 3040
rect 6570 2840 6690 3040
rect 6770 2840 6890 3040
rect 6970 2840 7090 3040
rect 7170 2840 7290 3040
rect 7370 2840 7490 3040
rect 7570 2840 7690 3040
rect 4730 1690 5530 2490
rect 5610 1690 6410 2490
rect 6490 1690 7290 2490
rect 7370 1690 8170 2490
<< ndiff >>
rect 4410 5130 4490 5160
rect 4410 5090 4430 5130
rect 4470 5090 4490 5130
rect 4410 5030 4490 5090
rect 4410 4990 4430 5030
rect 4470 4990 4490 5030
rect 4410 4930 4490 4990
rect 4410 4890 4430 4930
rect 4470 4890 4490 4930
rect 4410 4830 4490 4890
rect 4410 4790 4430 4830
rect 4470 4790 4490 4830
rect 4410 4730 4490 4790
rect 4410 4690 4430 4730
rect 4470 4690 4490 4730
rect 4410 4630 4490 4690
rect 4410 4590 4430 4630
rect 4470 4590 4490 4630
rect 4410 4530 4490 4590
rect 4410 4490 4430 4530
rect 4470 4490 4490 4530
rect 4410 4430 4490 4490
rect 4410 4390 4430 4430
rect 4470 4390 4490 4430
rect 4410 4360 4490 4390
rect 4610 5130 4690 5160
rect 4610 5090 4630 5130
rect 4670 5090 4690 5130
rect 4610 5030 4690 5090
rect 4610 4990 4630 5030
rect 4670 4990 4690 5030
rect 4610 4930 4690 4990
rect 4610 4890 4630 4930
rect 4670 4890 4690 4930
rect 4610 4830 4690 4890
rect 4610 4790 4630 4830
rect 4670 4790 4690 4830
rect 4610 4730 4690 4790
rect 4610 4690 4630 4730
rect 4670 4690 4690 4730
rect 4610 4630 4690 4690
rect 4610 4590 4630 4630
rect 4670 4590 4690 4630
rect 4610 4530 4690 4590
rect 4610 4490 4630 4530
rect 4670 4490 4690 4530
rect 4610 4430 4690 4490
rect 4610 4390 4630 4430
rect 4670 4390 4690 4430
rect 4610 4360 4690 4390
rect 4810 5130 4890 5160
rect 4810 5090 4830 5130
rect 4870 5090 4890 5130
rect 4810 5030 4890 5090
rect 4810 4990 4830 5030
rect 4870 4990 4890 5030
rect 4810 4930 4890 4990
rect 4810 4890 4830 4930
rect 4870 4890 4890 4930
rect 4810 4830 4890 4890
rect 4810 4790 4830 4830
rect 4870 4790 4890 4830
rect 4810 4730 4890 4790
rect 4810 4690 4830 4730
rect 4870 4690 4890 4730
rect 4810 4630 4890 4690
rect 4810 4590 4830 4630
rect 4870 4590 4890 4630
rect 4810 4530 4890 4590
rect 4810 4490 4830 4530
rect 4870 4490 4890 4530
rect 4810 4430 4890 4490
rect 4810 4390 4830 4430
rect 4870 4390 4890 4430
rect 4810 4360 4890 4390
rect 5010 5130 5090 5160
rect 5010 5090 5030 5130
rect 5070 5090 5090 5130
rect 5010 5030 5090 5090
rect 5010 4990 5030 5030
rect 5070 4990 5090 5030
rect 5010 4930 5090 4990
rect 5010 4890 5030 4930
rect 5070 4890 5090 4930
rect 5010 4830 5090 4890
rect 5010 4790 5030 4830
rect 5070 4790 5090 4830
rect 5010 4730 5090 4790
rect 5010 4690 5030 4730
rect 5070 4690 5090 4730
rect 5010 4630 5090 4690
rect 5010 4590 5030 4630
rect 5070 4590 5090 4630
rect 5010 4530 5090 4590
rect 5010 4490 5030 4530
rect 5070 4490 5090 4530
rect 5010 4430 5090 4490
rect 5010 4390 5030 4430
rect 5070 4390 5090 4430
rect 5010 4360 5090 4390
rect 5210 5130 5290 5160
rect 5210 5090 5230 5130
rect 5270 5090 5290 5130
rect 5210 5030 5290 5090
rect 5210 4990 5230 5030
rect 5270 4990 5290 5030
rect 5210 4930 5290 4990
rect 5210 4890 5230 4930
rect 5270 4890 5290 4930
rect 5210 4830 5290 4890
rect 5210 4790 5230 4830
rect 5270 4790 5290 4830
rect 5210 4730 5290 4790
rect 5210 4690 5230 4730
rect 5270 4690 5290 4730
rect 5210 4630 5290 4690
rect 5210 4590 5230 4630
rect 5270 4590 5290 4630
rect 5210 4530 5290 4590
rect 5210 4490 5230 4530
rect 5270 4490 5290 4530
rect 5210 4430 5290 4490
rect 5210 4390 5230 4430
rect 5270 4390 5290 4430
rect 5210 4360 5290 4390
rect 5410 5130 5490 5160
rect 5410 5090 5430 5130
rect 5470 5090 5490 5130
rect 5410 5030 5490 5090
rect 5410 4990 5430 5030
rect 5470 4990 5490 5030
rect 5410 4930 5490 4990
rect 5410 4890 5430 4930
rect 5470 4890 5490 4930
rect 5410 4830 5490 4890
rect 5410 4790 5430 4830
rect 5470 4790 5490 4830
rect 5410 4730 5490 4790
rect 5410 4690 5430 4730
rect 5470 4690 5490 4730
rect 5410 4630 5490 4690
rect 5410 4590 5430 4630
rect 5470 4590 5490 4630
rect 5410 4530 5490 4590
rect 5410 4490 5430 4530
rect 5470 4490 5490 4530
rect 5410 4430 5490 4490
rect 5410 4390 5430 4430
rect 5470 4390 5490 4430
rect 5410 4360 5490 4390
rect 5610 5130 5690 5160
rect 5610 5090 5630 5130
rect 5670 5090 5690 5130
rect 5610 5030 5690 5090
rect 5610 4990 5630 5030
rect 5670 4990 5690 5030
rect 5610 4930 5690 4990
rect 5610 4890 5630 4930
rect 5670 4890 5690 4930
rect 5610 4830 5690 4890
rect 5610 4790 5630 4830
rect 5670 4790 5690 4830
rect 5610 4730 5690 4790
rect 5610 4690 5630 4730
rect 5670 4690 5690 4730
rect 5610 4630 5690 4690
rect 5610 4590 5630 4630
rect 5670 4590 5690 4630
rect 5610 4530 5690 4590
rect 5610 4490 5630 4530
rect 5670 4490 5690 4530
rect 5610 4430 5690 4490
rect 5610 4390 5630 4430
rect 5670 4390 5690 4430
rect 5610 4360 5690 4390
rect 5810 5130 5890 5160
rect 5810 5090 5830 5130
rect 5870 5090 5890 5130
rect 5810 5030 5890 5090
rect 5810 4990 5830 5030
rect 5870 4990 5890 5030
rect 5810 4930 5890 4990
rect 5810 4890 5830 4930
rect 5870 4890 5890 4930
rect 5810 4830 5890 4890
rect 5810 4790 5830 4830
rect 5870 4790 5890 4830
rect 5810 4730 5890 4790
rect 5810 4690 5830 4730
rect 5870 4690 5890 4730
rect 5810 4630 5890 4690
rect 5810 4590 5830 4630
rect 5870 4590 5890 4630
rect 5810 4530 5890 4590
rect 5810 4490 5830 4530
rect 5870 4490 5890 4530
rect 5810 4430 5890 4490
rect 5810 4390 5830 4430
rect 5870 4390 5890 4430
rect 5810 4360 5890 4390
rect 6010 5130 6090 5160
rect 6010 5090 6030 5130
rect 6070 5090 6090 5130
rect 6010 5030 6090 5090
rect 6010 4990 6030 5030
rect 6070 4990 6090 5030
rect 6010 4930 6090 4990
rect 6010 4890 6030 4930
rect 6070 4890 6090 4930
rect 6010 4830 6090 4890
rect 6010 4790 6030 4830
rect 6070 4790 6090 4830
rect 6010 4730 6090 4790
rect 6010 4690 6030 4730
rect 6070 4690 6090 4730
rect 6010 4630 6090 4690
rect 6010 4590 6030 4630
rect 6070 4590 6090 4630
rect 6010 4530 6090 4590
rect 6010 4490 6030 4530
rect 6070 4490 6090 4530
rect 6010 4430 6090 4490
rect 6010 4390 6030 4430
rect 6070 4390 6090 4430
rect 6010 4360 6090 4390
rect 6210 5130 6290 5160
rect 6210 5090 6230 5130
rect 6270 5090 6290 5130
rect 6210 5030 6290 5090
rect 6210 4990 6230 5030
rect 6270 4990 6290 5030
rect 6210 4930 6290 4990
rect 6210 4890 6230 4930
rect 6270 4890 6290 4930
rect 6210 4830 6290 4890
rect 6210 4790 6230 4830
rect 6270 4790 6290 4830
rect 6210 4730 6290 4790
rect 6210 4690 6230 4730
rect 6270 4690 6290 4730
rect 6210 4630 6290 4690
rect 6210 4590 6230 4630
rect 6270 4590 6290 4630
rect 6210 4530 6290 4590
rect 6210 4490 6230 4530
rect 6270 4490 6290 4530
rect 6210 4430 6290 4490
rect 6210 4390 6230 4430
rect 6270 4390 6290 4430
rect 6210 4360 6290 4390
rect 6410 5130 6490 5160
rect 6410 5090 6430 5130
rect 6470 5090 6490 5130
rect 6410 5030 6490 5090
rect 6410 4990 6430 5030
rect 6470 4990 6490 5030
rect 6410 4930 6490 4990
rect 6410 4890 6430 4930
rect 6470 4890 6490 4930
rect 6410 4830 6490 4890
rect 6410 4790 6430 4830
rect 6470 4790 6490 4830
rect 6410 4730 6490 4790
rect 6410 4690 6430 4730
rect 6470 4690 6490 4730
rect 6410 4630 6490 4690
rect 6410 4590 6430 4630
rect 6470 4590 6490 4630
rect 6410 4530 6490 4590
rect 6410 4490 6430 4530
rect 6470 4490 6490 4530
rect 6410 4430 6490 4490
rect 6410 4390 6430 4430
rect 6470 4390 6490 4430
rect 6410 4360 6490 4390
rect 6610 5130 6690 5160
rect 6610 5090 6630 5130
rect 6670 5090 6690 5130
rect 6610 5030 6690 5090
rect 6610 4990 6630 5030
rect 6670 4990 6690 5030
rect 6610 4930 6690 4990
rect 6610 4890 6630 4930
rect 6670 4890 6690 4930
rect 6610 4830 6690 4890
rect 6610 4790 6630 4830
rect 6670 4790 6690 4830
rect 6610 4730 6690 4790
rect 6610 4690 6630 4730
rect 6670 4690 6690 4730
rect 6610 4630 6690 4690
rect 6610 4590 6630 4630
rect 6670 4590 6690 4630
rect 6610 4530 6690 4590
rect 6610 4490 6630 4530
rect 6670 4490 6690 4530
rect 6610 4430 6690 4490
rect 6610 4390 6630 4430
rect 6670 4390 6690 4430
rect 6610 4360 6690 4390
rect 6810 5130 6890 5160
rect 6810 5090 6830 5130
rect 6870 5090 6890 5130
rect 6810 5030 6890 5090
rect 6810 4990 6830 5030
rect 6870 4990 6890 5030
rect 6810 4930 6890 4990
rect 6810 4890 6830 4930
rect 6870 4890 6890 4930
rect 6810 4830 6890 4890
rect 6810 4790 6830 4830
rect 6870 4790 6890 4830
rect 6810 4730 6890 4790
rect 6810 4690 6830 4730
rect 6870 4690 6890 4730
rect 6810 4630 6890 4690
rect 6810 4590 6830 4630
rect 6870 4590 6890 4630
rect 6810 4530 6890 4590
rect 6810 4490 6830 4530
rect 6870 4490 6890 4530
rect 6810 4430 6890 4490
rect 6810 4390 6830 4430
rect 6870 4390 6890 4430
rect 6810 4360 6890 4390
rect 7010 5130 7090 5160
rect 7010 5090 7030 5130
rect 7070 5090 7090 5130
rect 7010 5030 7090 5090
rect 7010 4990 7030 5030
rect 7070 4990 7090 5030
rect 7010 4930 7090 4990
rect 7010 4890 7030 4930
rect 7070 4890 7090 4930
rect 7010 4830 7090 4890
rect 7010 4790 7030 4830
rect 7070 4790 7090 4830
rect 7010 4730 7090 4790
rect 7010 4690 7030 4730
rect 7070 4690 7090 4730
rect 7010 4630 7090 4690
rect 7010 4590 7030 4630
rect 7070 4590 7090 4630
rect 7010 4530 7090 4590
rect 7010 4490 7030 4530
rect 7070 4490 7090 4530
rect 7010 4430 7090 4490
rect 7010 4390 7030 4430
rect 7070 4390 7090 4430
rect 7010 4360 7090 4390
rect 7210 5130 7290 5160
rect 7210 5090 7230 5130
rect 7270 5090 7290 5130
rect 7210 5030 7290 5090
rect 7210 4990 7230 5030
rect 7270 4990 7290 5030
rect 7210 4930 7290 4990
rect 7210 4890 7230 4930
rect 7270 4890 7290 4930
rect 7210 4830 7290 4890
rect 7210 4790 7230 4830
rect 7270 4790 7290 4830
rect 7210 4730 7290 4790
rect 7210 4690 7230 4730
rect 7270 4690 7290 4730
rect 7210 4630 7290 4690
rect 7210 4590 7230 4630
rect 7270 4590 7290 4630
rect 7210 4530 7290 4590
rect 7210 4490 7230 4530
rect 7270 4490 7290 4530
rect 7210 4430 7290 4490
rect 7210 4390 7230 4430
rect 7270 4390 7290 4430
rect 7210 4360 7290 4390
rect 7410 5130 7490 5160
rect 7410 5090 7430 5130
rect 7470 5090 7490 5130
rect 7410 5030 7490 5090
rect 7410 4990 7430 5030
rect 7470 4990 7490 5030
rect 7410 4930 7490 4990
rect 7410 4890 7430 4930
rect 7470 4890 7490 4930
rect 7410 4830 7490 4890
rect 7410 4790 7430 4830
rect 7470 4790 7490 4830
rect 7410 4730 7490 4790
rect 7410 4690 7430 4730
rect 7470 4690 7490 4730
rect 7410 4630 7490 4690
rect 7410 4590 7430 4630
rect 7470 4590 7490 4630
rect 7410 4530 7490 4590
rect 7410 4490 7430 4530
rect 7470 4490 7490 4530
rect 7410 4430 7490 4490
rect 7410 4390 7430 4430
rect 7470 4390 7490 4430
rect 7410 4360 7490 4390
rect 7610 5130 7690 5160
rect 7610 5090 7630 5130
rect 7670 5090 7690 5130
rect 7610 5030 7690 5090
rect 7610 4990 7630 5030
rect 7670 4990 7690 5030
rect 7610 4930 7690 4990
rect 7610 4890 7630 4930
rect 7670 4890 7690 4930
rect 7610 4830 7690 4890
rect 7610 4790 7630 4830
rect 7670 4790 7690 4830
rect 7610 4730 7690 4790
rect 7610 4690 7630 4730
rect 7670 4690 7690 4730
rect 7610 4630 7690 4690
rect 7610 4590 7630 4630
rect 7670 4590 7690 4630
rect 7610 4530 7690 4590
rect 7610 4490 7630 4530
rect 7670 4490 7690 4530
rect 7610 4430 7690 4490
rect 7610 4390 7630 4430
rect 7670 4390 7690 4430
rect 7610 4360 7690 4390
rect 7810 5130 7890 5160
rect 7810 5090 7830 5130
rect 7870 5090 7890 5130
rect 7810 5030 7890 5090
rect 7810 4990 7830 5030
rect 7870 4990 7890 5030
rect 7810 4930 7890 4990
rect 7810 4890 7830 4930
rect 7870 4890 7890 4930
rect 7810 4830 7890 4890
rect 7810 4790 7830 4830
rect 7870 4790 7890 4830
rect 7810 4730 7890 4790
rect 7810 4690 7830 4730
rect 7870 4690 7890 4730
rect 7810 4630 7890 4690
rect 7810 4590 7830 4630
rect 7870 4590 7890 4630
rect 7810 4530 7890 4590
rect 7810 4490 7830 4530
rect 7870 4490 7890 4530
rect 7810 4430 7890 4490
rect 7810 4390 7830 4430
rect 7870 4390 7890 4430
rect 7810 4360 7890 4390
rect 8010 5130 8090 5160
rect 8010 5090 8030 5130
rect 8070 5090 8090 5130
rect 8010 5030 8090 5090
rect 8010 4990 8030 5030
rect 8070 4990 8090 5030
rect 8010 4930 8090 4990
rect 8010 4890 8030 4930
rect 8070 4890 8090 4930
rect 8010 4830 8090 4890
rect 8010 4790 8030 4830
rect 8070 4790 8090 4830
rect 8010 4730 8090 4790
rect 8010 4690 8030 4730
rect 8070 4690 8090 4730
rect 8010 4630 8090 4690
rect 8010 4590 8030 4630
rect 8070 4590 8090 4630
rect 8010 4530 8090 4590
rect 8010 4490 8030 4530
rect 8070 4490 8090 4530
rect 8010 4430 8090 4490
rect 8010 4390 8030 4430
rect 8070 4390 8090 4430
rect 8010 4360 8090 4390
rect 8210 5130 8290 5160
rect 8210 5090 8230 5130
rect 8270 5090 8290 5130
rect 8210 5030 8290 5090
rect 8210 4990 8230 5030
rect 8270 4990 8290 5030
rect 8210 4930 8290 4990
rect 8210 4890 8230 4930
rect 8270 4890 8290 4930
rect 8210 4830 8290 4890
rect 8210 4790 8230 4830
rect 8270 4790 8290 4830
rect 8210 4730 8290 4790
rect 8210 4690 8230 4730
rect 8270 4690 8290 4730
rect 8210 4630 8290 4690
rect 8210 4590 8230 4630
rect 8270 4590 8290 4630
rect 8210 4530 8290 4590
rect 8210 4490 8230 4530
rect 8270 4490 8290 4530
rect 8210 4430 8290 4490
rect 8210 4390 8230 4430
rect 8270 4390 8290 4430
rect 8210 4360 8290 4390
rect 8410 5130 8490 5160
rect 8410 5090 8430 5130
rect 8470 5090 8490 5130
rect 8410 5030 8490 5090
rect 8410 4990 8430 5030
rect 8470 4990 8490 5030
rect 8410 4930 8490 4990
rect 8410 4890 8430 4930
rect 8470 4890 8490 4930
rect 8410 4830 8490 4890
rect 8410 4790 8430 4830
rect 8470 4790 8490 4830
rect 8410 4730 8490 4790
rect 8410 4690 8430 4730
rect 8470 4690 8490 4730
rect 8410 4630 8490 4690
rect 8410 4590 8430 4630
rect 8470 4590 8490 4630
rect 8410 4530 8490 4590
rect 8410 4490 8430 4530
rect 8470 4490 8490 4530
rect 8410 4430 8490 4490
rect 8410 4390 8430 4430
rect 8470 4390 8490 4430
rect 8410 4360 8490 4390
rect 10330 4330 10410 4360
rect 10330 4290 10350 4330
rect 10390 4290 10410 4330
rect 10330 4230 10410 4290
rect 10330 4190 10350 4230
rect 10390 4190 10410 4230
rect 10330 4130 10410 4190
rect 10330 4090 10350 4130
rect 10390 4090 10410 4130
rect 10330 4030 10410 4090
rect 10330 3990 10350 4030
rect 10390 3990 10410 4030
rect 10330 3960 10410 3990
rect 10440 4330 10520 4360
rect 10440 4290 10460 4330
rect 10500 4290 10520 4330
rect 10440 4230 10520 4290
rect 10440 4190 10460 4230
rect 10500 4190 10520 4230
rect 10440 4130 10520 4190
rect 10440 4090 10460 4130
rect 10500 4090 10520 4130
rect 10440 4030 10520 4090
rect 10440 3990 10460 4030
rect 10500 3990 10520 4030
rect 10440 3960 10520 3990
rect 10580 4330 10660 4360
rect 10580 4290 10600 4330
rect 10640 4290 10660 4330
rect 10580 4230 10660 4290
rect 10580 4190 10600 4230
rect 10640 4190 10660 4230
rect 10580 4130 10660 4190
rect 10580 4090 10600 4130
rect 10640 4090 10660 4130
rect 10580 4030 10660 4090
rect 10580 3990 10600 4030
rect 10640 3990 10660 4030
rect 10580 3960 10660 3990
rect 10690 4330 10770 4360
rect 10690 4290 10710 4330
rect 10750 4290 10770 4330
rect 10690 4230 10770 4290
rect 10690 4190 10710 4230
rect 10750 4190 10770 4230
rect 10690 4130 10770 4190
rect 10690 4090 10710 4130
rect 10750 4090 10770 4130
rect 10690 4030 10770 4090
rect 10690 3990 10710 4030
rect 10750 3990 10770 4030
rect 10690 3960 10770 3990
rect 4450 3820 4530 3850
rect 4450 3780 4470 3820
rect 4510 3780 4530 3820
rect 4450 3720 4530 3780
rect 4450 3680 4470 3720
rect 4510 3680 4530 3720
rect 4450 3620 4530 3680
rect 4450 3580 4470 3620
rect 4510 3580 4530 3620
rect 4450 3520 4530 3580
rect 4450 3480 4470 3520
rect 4510 3480 4530 3520
rect 4450 3450 4530 3480
rect 4650 3820 4730 3850
rect 4650 3780 4670 3820
rect 4710 3780 4730 3820
rect 4650 3720 4730 3780
rect 4650 3680 4670 3720
rect 4710 3680 4730 3720
rect 4650 3620 4730 3680
rect 4650 3580 4670 3620
rect 4710 3580 4730 3620
rect 4650 3520 4730 3580
rect 4650 3480 4670 3520
rect 4710 3480 4730 3520
rect 4650 3450 4730 3480
rect 4850 3820 4930 3850
rect 4850 3780 4870 3820
rect 4910 3780 4930 3820
rect 4850 3720 4930 3780
rect 4850 3680 4870 3720
rect 4910 3680 4930 3720
rect 4850 3620 4930 3680
rect 4850 3580 4870 3620
rect 4910 3580 4930 3620
rect 4850 3520 4930 3580
rect 4850 3480 4870 3520
rect 4910 3480 4930 3520
rect 4850 3450 4930 3480
rect 5050 3820 5130 3850
rect 5050 3780 5070 3820
rect 5110 3780 5130 3820
rect 5050 3720 5130 3780
rect 5050 3680 5070 3720
rect 5110 3680 5130 3720
rect 5050 3620 5130 3680
rect 5050 3580 5070 3620
rect 5110 3580 5130 3620
rect 5050 3520 5130 3580
rect 5050 3480 5070 3520
rect 5110 3480 5130 3520
rect 5050 3450 5130 3480
rect 5250 3820 5330 3850
rect 5250 3780 5270 3820
rect 5310 3780 5330 3820
rect 5250 3720 5330 3780
rect 5250 3680 5270 3720
rect 5310 3680 5330 3720
rect 5250 3620 5330 3680
rect 5250 3580 5270 3620
rect 5310 3580 5330 3620
rect 5250 3520 5330 3580
rect 5250 3480 5270 3520
rect 5310 3480 5330 3520
rect 5250 3450 5330 3480
rect 5450 3820 5530 3850
rect 5450 3780 5470 3820
rect 5510 3780 5530 3820
rect 5450 3720 5530 3780
rect 5450 3680 5470 3720
rect 5510 3680 5530 3720
rect 5450 3620 5530 3680
rect 5450 3580 5470 3620
rect 5510 3580 5530 3620
rect 5450 3520 5530 3580
rect 5450 3480 5470 3520
rect 5510 3480 5530 3520
rect 5450 3450 5530 3480
rect 5650 3820 5730 3850
rect 5810 3820 5890 3850
rect 5650 3780 5670 3820
rect 5710 3780 5730 3820
rect 5810 3780 5830 3820
rect 5870 3780 5890 3820
rect 5650 3720 5730 3780
rect 5810 3720 5890 3780
rect 5650 3680 5670 3720
rect 5710 3680 5730 3720
rect 5810 3680 5830 3720
rect 5870 3680 5890 3720
rect 5650 3620 5730 3680
rect 5810 3620 5890 3680
rect 5650 3580 5670 3620
rect 5710 3580 5730 3620
rect 5810 3580 5830 3620
rect 5870 3580 5890 3620
rect 5650 3520 5730 3580
rect 5810 3520 5890 3580
rect 5650 3480 5670 3520
rect 5710 3480 5730 3520
rect 5810 3480 5830 3520
rect 5870 3480 5890 3520
rect 5650 3450 5730 3480
rect 5810 3450 5890 3480
rect 6010 3820 6090 3850
rect 6010 3780 6030 3820
rect 6070 3780 6090 3820
rect 6010 3720 6090 3780
rect 6010 3680 6030 3720
rect 6070 3680 6090 3720
rect 6010 3620 6090 3680
rect 6010 3580 6030 3620
rect 6070 3580 6090 3620
rect 6010 3520 6090 3580
rect 6010 3480 6030 3520
rect 6070 3480 6090 3520
rect 6010 3450 6090 3480
rect 6210 3820 6290 3850
rect 6210 3780 6230 3820
rect 6270 3780 6290 3820
rect 6210 3720 6290 3780
rect 6210 3680 6230 3720
rect 6270 3680 6290 3720
rect 6210 3620 6290 3680
rect 6210 3580 6230 3620
rect 6270 3580 6290 3620
rect 6210 3520 6290 3580
rect 6210 3480 6230 3520
rect 6270 3480 6290 3520
rect 6210 3450 6290 3480
rect 6410 3820 6490 3850
rect 6410 3780 6430 3820
rect 6470 3780 6490 3820
rect 6410 3720 6490 3780
rect 6410 3680 6430 3720
rect 6470 3680 6490 3720
rect 6410 3620 6490 3680
rect 6410 3580 6430 3620
rect 6470 3580 6490 3620
rect 6410 3520 6490 3580
rect 6410 3480 6430 3520
rect 6470 3480 6490 3520
rect 6410 3450 6490 3480
rect 6610 3820 6690 3850
rect 6610 3780 6630 3820
rect 6670 3780 6690 3820
rect 6610 3720 6690 3780
rect 6610 3680 6630 3720
rect 6670 3680 6690 3720
rect 6610 3620 6690 3680
rect 6610 3580 6630 3620
rect 6670 3580 6690 3620
rect 6610 3520 6690 3580
rect 6610 3480 6630 3520
rect 6670 3480 6690 3520
rect 6610 3450 6690 3480
rect 6810 3820 6890 3850
rect 6810 3780 6830 3820
rect 6870 3780 6890 3820
rect 6810 3720 6890 3780
rect 6810 3680 6830 3720
rect 6870 3680 6890 3720
rect 6810 3620 6890 3680
rect 6810 3580 6830 3620
rect 6870 3580 6890 3620
rect 6810 3520 6890 3580
rect 6810 3480 6830 3520
rect 6870 3480 6890 3520
rect 6810 3450 6890 3480
rect 7010 3820 7090 3850
rect 7170 3820 7250 3850
rect 7010 3780 7030 3820
rect 7070 3780 7090 3820
rect 7170 3780 7190 3820
rect 7230 3780 7250 3820
rect 7010 3720 7090 3780
rect 7170 3720 7250 3780
rect 7010 3680 7030 3720
rect 7070 3680 7090 3720
rect 7170 3680 7190 3720
rect 7230 3680 7250 3720
rect 7010 3620 7090 3680
rect 7170 3620 7250 3680
rect 7010 3580 7030 3620
rect 7070 3580 7090 3620
rect 7170 3580 7190 3620
rect 7230 3580 7250 3620
rect 7010 3520 7090 3580
rect 7170 3520 7250 3580
rect 7010 3480 7030 3520
rect 7070 3480 7090 3520
rect 7170 3480 7190 3520
rect 7230 3480 7250 3520
rect 7010 3450 7090 3480
rect 7170 3450 7250 3480
rect 7370 3820 7450 3850
rect 7370 3780 7390 3820
rect 7430 3780 7450 3820
rect 7370 3720 7450 3780
rect 7370 3680 7390 3720
rect 7430 3680 7450 3720
rect 7370 3620 7450 3680
rect 7370 3580 7390 3620
rect 7430 3580 7450 3620
rect 7370 3520 7450 3580
rect 7370 3480 7390 3520
rect 7430 3480 7450 3520
rect 7370 3450 7450 3480
rect 7570 3820 7650 3850
rect 7570 3780 7590 3820
rect 7630 3780 7650 3820
rect 7570 3720 7650 3780
rect 7570 3680 7590 3720
rect 7630 3680 7650 3720
rect 7570 3620 7650 3680
rect 7570 3580 7590 3620
rect 7630 3580 7650 3620
rect 7570 3520 7650 3580
rect 7570 3480 7590 3520
rect 7630 3480 7650 3520
rect 7570 3450 7650 3480
rect 7770 3820 7850 3850
rect 7770 3780 7790 3820
rect 7830 3780 7850 3820
rect 7770 3720 7850 3780
rect 7770 3680 7790 3720
rect 7830 3680 7850 3720
rect 7770 3620 7850 3680
rect 7770 3580 7790 3620
rect 7830 3580 7850 3620
rect 7770 3520 7850 3580
rect 7770 3480 7790 3520
rect 7830 3480 7850 3520
rect 7770 3450 7850 3480
rect 7970 3820 8050 3850
rect 7970 3780 7990 3820
rect 8030 3780 8050 3820
rect 7970 3720 8050 3780
rect 7970 3680 7990 3720
rect 8030 3680 8050 3720
rect 7970 3620 8050 3680
rect 7970 3580 7990 3620
rect 8030 3580 8050 3620
rect 7970 3520 8050 3580
rect 7970 3480 7990 3520
rect 8030 3480 8050 3520
rect 7970 3450 8050 3480
rect 8170 3820 8250 3850
rect 8170 3780 8190 3820
rect 8230 3780 8250 3820
rect 8170 3720 8250 3780
rect 8170 3680 8190 3720
rect 8230 3680 8250 3720
rect 8170 3620 8250 3680
rect 8170 3580 8190 3620
rect 8230 3580 8250 3620
rect 8170 3520 8250 3580
rect 8170 3480 8190 3520
rect 8230 3480 8250 3520
rect 8170 3450 8250 3480
rect 8370 3820 8450 3850
rect 8370 3780 8390 3820
rect 8430 3780 8450 3820
rect 8370 3720 8450 3780
rect 8370 3680 8390 3720
rect 8430 3680 8450 3720
rect 8370 3620 8450 3680
rect 8370 3580 8390 3620
rect 8430 3580 8450 3620
rect 8370 3520 8450 3580
rect 8370 3480 8390 3520
rect 8430 3480 8450 3520
rect 8370 3450 8450 3480
rect 9210 3630 9290 3660
rect 9210 3590 9230 3630
rect 9270 3590 9290 3630
rect 9210 3530 9290 3590
rect 9210 3490 9230 3530
rect 9270 3490 9290 3530
rect 9210 3460 9290 3490
rect 11290 3630 11370 3660
rect 11290 3590 11310 3630
rect 11350 3590 11370 3630
rect 11290 3530 11370 3590
rect 11290 3490 11310 3530
rect 11350 3490 11370 3530
rect 11290 3460 11370 3490
rect 5130 3010 5210 3040
rect 5130 2970 5150 3010
rect 5190 2970 5210 3010
rect 5130 2910 5210 2970
rect 5130 2870 5150 2910
rect 5190 2870 5210 2910
rect 5130 2840 5210 2870
rect 5330 3010 5410 3040
rect 5330 2970 5350 3010
rect 5390 2970 5410 3010
rect 5330 2910 5410 2970
rect 5330 2870 5350 2910
rect 5390 2870 5410 2910
rect 5330 2840 5410 2870
rect 5530 3010 5610 3040
rect 5530 2970 5550 3010
rect 5590 2970 5610 3010
rect 5530 2910 5610 2970
rect 5530 2870 5550 2910
rect 5590 2870 5610 2910
rect 5530 2840 5610 2870
rect 5730 3010 5810 3040
rect 5730 2970 5750 3010
rect 5790 2970 5810 3010
rect 5730 2910 5810 2970
rect 5730 2870 5750 2910
rect 5790 2870 5810 2910
rect 5730 2840 5810 2870
rect 5930 3010 6010 3040
rect 5930 2970 5950 3010
rect 5990 2970 6010 3010
rect 5930 2910 6010 2970
rect 5930 2870 5950 2910
rect 5990 2870 6010 2910
rect 5930 2840 6010 2870
rect 6130 3010 6210 3040
rect 6130 2970 6150 3010
rect 6190 2970 6210 3010
rect 6130 2910 6210 2970
rect 6130 2870 6150 2910
rect 6190 2870 6210 2910
rect 6130 2840 6210 2870
rect 6330 3010 6410 3040
rect 6490 3010 6570 3040
rect 6330 2970 6350 3010
rect 6390 2970 6410 3010
rect 6490 2970 6510 3010
rect 6550 2970 6570 3010
rect 6330 2910 6410 2970
rect 6490 2910 6570 2970
rect 6330 2870 6350 2910
rect 6390 2870 6410 2910
rect 6490 2870 6510 2910
rect 6550 2870 6570 2910
rect 6330 2840 6410 2870
rect 6490 2840 6570 2870
rect 6690 3010 6770 3040
rect 6690 2970 6710 3010
rect 6750 2970 6770 3010
rect 6690 2910 6770 2970
rect 6690 2870 6710 2910
rect 6750 2870 6770 2910
rect 6690 2840 6770 2870
rect 6890 3010 6970 3040
rect 6890 2970 6910 3010
rect 6950 2970 6970 3010
rect 6890 2910 6970 2970
rect 6890 2870 6910 2910
rect 6950 2870 6970 2910
rect 6890 2840 6970 2870
rect 7090 3010 7170 3040
rect 7090 2970 7110 3010
rect 7150 2970 7170 3010
rect 7090 2910 7170 2970
rect 7090 2870 7110 2910
rect 7150 2870 7170 2910
rect 7090 2840 7170 2870
rect 7290 3010 7370 3040
rect 7290 2970 7310 3010
rect 7350 2970 7370 3010
rect 7290 2910 7370 2970
rect 7290 2870 7310 2910
rect 7350 2870 7370 2910
rect 7290 2840 7370 2870
rect 7490 3010 7570 3040
rect 7490 2970 7510 3010
rect 7550 2970 7570 3010
rect 7490 2910 7570 2970
rect 7490 2870 7510 2910
rect 7550 2870 7570 2910
rect 7490 2840 7570 2870
rect 7690 3010 7770 3040
rect 7690 2970 7710 3010
rect 7750 2970 7770 3010
rect 7690 2910 7770 2970
rect 7690 2870 7710 2910
rect 7750 2870 7770 2910
rect 7690 2840 7770 2870
rect 4650 2460 4730 2490
rect 4650 2420 4670 2460
rect 4710 2420 4730 2460
rect 4650 2360 4730 2420
rect 4650 2320 4670 2360
rect 4710 2320 4730 2360
rect 4650 2260 4730 2320
rect 4650 2220 4670 2260
rect 4710 2220 4730 2260
rect 4650 2160 4730 2220
rect 4650 2120 4670 2160
rect 4710 2120 4730 2160
rect 4650 2060 4730 2120
rect 4650 2020 4670 2060
rect 4710 2020 4730 2060
rect 4650 1960 4730 2020
rect 4650 1920 4670 1960
rect 4710 1920 4730 1960
rect 4650 1860 4730 1920
rect 4650 1820 4670 1860
rect 4710 1820 4730 1860
rect 4650 1760 4730 1820
rect 4650 1720 4670 1760
rect 4710 1720 4730 1760
rect 4650 1690 4730 1720
rect 5530 2460 5610 2490
rect 5530 2420 5550 2460
rect 5590 2420 5610 2460
rect 5530 2360 5610 2420
rect 5530 2320 5550 2360
rect 5590 2320 5610 2360
rect 5530 2260 5610 2320
rect 5530 2220 5550 2260
rect 5590 2220 5610 2260
rect 5530 2160 5610 2220
rect 5530 2120 5550 2160
rect 5590 2120 5610 2160
rect 5530 2060 5610 2120
rect 5530 2020 5550 2060
rect 5590 2020 5610 2060
rect 5530 1960 5610 2020
rect 5530 1920 5550 1960
rect 5590 1920 5610 1960
rect 5530 1860 5610 1920
rect 5530 1820 5550 1860
rect 5590 1820 5610 1860
rect 5530 1760 5610 1820
rect 5530 1720 5550 1760
rect 5590 1720 5610 1760
rect 5530 1690 5610 1720
rect 6410 2460 6490 2490
rect 6410 2420 6430 2460
rect 6470 2420 6490 2460
rect 6410 2360 6490 2420
rect 6410 2320 6430 2360
rect 6470 2320 6490 2360
rect 6410 2260 6490 2320
rect 6410 2220 6430 2260
rect 6470 2220 6490 2260
rect 6410 2160 6490 2220
rect 6410 2120 6430 2160
rect 6470 2120 6490 2160
rect 6410 2060 6490 2120
rect 6410 2020 6430 2060
rect 6470 2020 6490 2060
rect 6410 1960 6490 2020
rect 6410 1920 6430 1960
rect 6470 1920 6490 1960
rect 6410 1860 6490 1920
rect 6410 1820 6430 1860
rect 6470 1820 6490 1860
rect 6410 1760 6490 1820
rect 6410 1720 6430 1760
rect 6470 1720 6490 1760
rect 6410 1690 6490 1720
rect 7290 2460 7370 2490
rect 7290 2420 7310 2460
rect 7350 2420 7370 2460
rect 7290 2360 7370 2420
rect 7290 2320 7310 2360
rect 7350 2320 7370 2360
rect 7290 2260 7370 2320
rect 7290 2220 7310 2260
rect 7350 2220 7370 2260
rect 7290 2160 7370 2220
rect 7290 2120 7310 2160
rect 7350 2120 7370 2160
rect 7290 2060 7370 2120
rect 7290 2020 7310 2060
rect 7350 2020 7370 2060
rect 7290 1960 7370 2020
rect 7290 1920 7310 1960
rect 7350 1920 7370 1960
rect 7290 1860 7370 1920
rect 7290 1820 7310 1860
rect 7350 1820 7370 1860
rect 7290 1760 7370 1820
rect 7290 1720 7310 1760
rect 7350 1720 7370 1760
rect 7290 1690 7370 1720
rect 8170 2460 8250 2490
rect 8170 2420 8190 2460
rect 8230 2420 8250 2460
rect 8170 2360 8250 2420
rect 8170 2320 8190 2360
rect 8230 2320 8250 2360
rect 8170 2260 8250 2320
rect 8170 2220 8190 2260
rect 8230 2220 8250 2260
rect 8170 2160 8250 2220
rect 8170 2120 8190 2160
rect 8230 2120 8250 2160
rect 8170 2060 8250 2120
rect 8170 2020 8190 2060
rect 8230 2020 8250 2060
rect 8170 1960 8250 2020
rect 8170 1920 8190 1960
rect 8230 1920 8250 1960
rect 8170 1860 8250 1920
rect 8170 1820 8190 1860
rect 8230 1820 8250 1860
rect 8170 1760 8250 1820
rect 8170 1720 8190 1760
rect 8230 1720 8250 1760
rect 8170 1690 8250 1720
<< pdiff >>
rect 1680 958 2360 1010
rect 1680 924 1734 958
rect 1768 924 1824 958
rect 1858 924 1914 958
rect 1948 924 2004 958
rect 2038 924 2094 958
rect 2128 924 2184 958
rect 2218 924 2274 958
rect 2308 924 2360 958
rect 1680 868 2360 924
rect 1680 834 1734 868
rect 1768 834 1824 868
rect 1858 834 1914 868
rect 1948 834 2004 868
rect 2038 834 2094 868
rect 2128 834 2184 868
rect 2218 834 2274 868
rect 2308 834 2360 868
rect 1680 778 2360 834
rect 1680 744 1734 778
rect 1768 744 1824 778
rect 1858 744 1914 778
rect 1948 744 2004 778
rect 2038 744 2094 778
rect 2128 744 2184 778
rect 2218 744 2274 778
rect 2308 744 2360 778
rect 1680 688 2360 744
rect 1680 654 1734 688
rect 1768 654 1824 688
rect 1858 654 1914 688
rect 1948 654 2004 688
rect 2038 654 2094 688
rect 2128 654 2184 688
rect 2218 654 2274 688
rect 2308 654 2360 688
rect 1680 598 2360 654
rect 1680 564 1734 598
rect 1768 564 1824 598
rect 1858 564 1914 598
rect 1948 564 2004 598
rect 2038 564 2094 598
rect 2128 564 2184 598
rect 2218 564 2274 598
rect 2308 564 2360 598
rect 1680 508 2360 564
rect 1680 474 1734 508
rect 1768 474 1824 508
rect 1858 474 1914 508
rect 1948 474 2004 508
rect 2038 474 2094 508
rect 2128 474 2184 508
rect 2218 474 2274 508
rect 2308 474 2360 508
rect 1680 418 2360 474
rect 1680 384 1734 418
rect 1768 384 1824 418
rect 1858 384 1914 418
rect 1948 384 2004 418
rect 2038 384 2094 418
rect 2128 384 2184 418
rect 2218 384 2274 418
rect 2308 384 2360 418
rect 1680 330 2360 384
rect 3040 958 3720 1010
rect 3040 924 3094 958
rect 3128 924 3184 958
rect 3218 924 3274 958
rect 3308 924 3364 958
rect 3398 924 3454 958
rect 3488 924 3544 958
rect 3578 924 3634 958
rect 3668 924 3720 958
rect 3040 868 3720 924
rect 3040 834 3094 868
rect 3128 834 3184 868
rect 3218 834 3274 868
rect 3308 834 3364 868
rect 3398 834 3454 868
rect 3488 834 3544 868
rect 3578 834 3634 868
rect 3668 834 3720 868
rect 3040 778 3720 834
rect 3040 744 3094 778
rect 3128 744 3184 778
rect 3218 744 3274 778
rect 3308 744 3364 778
rect 3398 744 3454 778
rect 3488 744 3544 778
rect 3578 744 3634 778
rect 3668 744 3720 778
rect 3040 688 3720 744
rect 3040 654 3094 688
rect 3128 654 3184 688
rect 3218 654 3274 688
rect 3308 654 3364 688
rect 3398 654 3454 688
rect 3488 654 3544 688
rect 3578 654 3634 688
rect 3668 654 3720 688
rect 3040 598 3720 654
rect 3040 564 3094 598
rect 3128 564 3184 598
rect 3218 564 3274 598
rect 3308 564 3364 598
rect 3398 564 3454 598
rect 3488 564 3544 598
rect 3578 564 3634 598
rect 3668 564 3720 598
rect 3040 508 3720 564
rect 3040 474 3094 508
rect 3128 474 3184 508
rect 3218 474 3274 508
rect 3308 474 3364 508
rect 3398 474 3454 508
rect 3488 474 3544 508
rect 3578 474 3634 508
rect 3668 474 3720 508
rect 3040 418 3720 474
rect 3040 384 3094 418
rect 3128 384 3184 418
rect 3218 384 3274 418
rect 3308 384 3364 418
rect 3398 384 3454 418
rect 3488 384 3544 418
rect 3578 384 3634 418
rect 3668 384 3720 418
rect 3040 330 3720 384
rect 4400 958 5080 1010
rect 4400 924 4454 958
rect 4488 924 4544 958
rect 4578 924 4634 958
rect 4668 924 4724 958
rect 4758 924 4814 958
rect 4848 924 4904 958
rect 4938 924 4994 958
rect 5028 924 5080 958
rect 4400 868 5080 924
rect 4400 834 4454 868
rect 4488 834 4544 868
rect 4578 834 4634 868
rect 4668 834 4724 868
rect 4758 834 4814 868
rect 4848 834 4904 868
rect 4938 834 4994 868
rect 5028 834 5080 868
rect 4400 778 5080 834
rect 4400 744 4454 778
rect 4488 744 4544 778
rect 4578 744 4634 778
rect 4668 744 4724 778
rect 4758 744 4814 778
rect 4848 744 4904 778
rect 4938 744 4994 778
rect 5028 744 5080 778
rect 4400 688 5080 744
rect 4400 654 4454 688
rect 4488 654 4544 688
rect 4578 654 4634 688
rect 4668 654 4724 688
rect 4758 654 4814 688
rect 4848 654 4904 688
rect 4938 654 4994 688
rect 5028 654 5080 688
rect 4400 598 5080 654
rect 4400 564 4454 598
rect 4488 564 4544 598
rect 4578 564 4634 598
rect 4668 564 4724 598
rect 4758 564 4814 598
rect 4848 564 4904 598
rect 4938 564 4994 598
rect 5028 564 5080 598
rect 4400 508 5080 564
rect 4400 474 4454 508
rect 4488 474 4544 508
rect 4578 474 4634 508
rect 4668 474 4724 508
rect 4758 474 4814 508
rect 4848 474 4904 508
rect 4938 474 4994 508
rect 5028 474 5080 508
rect 4400 418 5080 474
rect 4400 384 4454 418
rect 4488 384 4544 418
rect 4578 384 4634 418
rect 4668 384 4724 418
rect 4758 384 4814 418
rect 4848 384 4904 418
rect 4938 384 4994 418
rect 5028 384 5080 418
rect 4400 330 5080 384
rect 5760 958 6440 1010
rect 5760 924 5814 958
rect 5848 924 5904 958
rect 5938 924 5994 958
rect 6028 924 6084 958
rect 6118 924 6174 958
rect 6208 924 6264 958
rect 6298 924 6354 958
rect 6388 924 6440 958
rect 5760 868 6440 924
rect 5760 834 5814 868
rect 5848 834 5904 868
rect 5938 834 5994 868
rect 6028 834 6084 868
rect 6118 834 6174 868
rect 6208 834 6264 868
rect 6298 834 6354 868
rect 6388 834 6440 868
rect 5760 778 6440 834
rect 5760 744 5814 778
rect 5848 744 5904 778
rect 5938 744 5994 778
rect 6028 744 6084 778
rect 6118 744 6174 778
rect 6208 744 6264 778
rect 6298 744 6354 778
rect 6388 744 6440 778
rect 5760 688 6440 744
rect 5760 654 5814 688
rect 5848 654 5904 688
rect 5938 654 5994 688
rect 6028 654 6084 688
rect 6118 654 6174 688
rect 6208 654 6264 688
rect 6298 654 6354 688
rect 6388 654 6440 688
rect 5760 598 6440 654
rect 5760 564 5814 598
rect 5848 564 5904 598
rect 5938 564 5994 598
rect 6028 564 6084 598
rect 6118 564 6174 598
rect 6208 564 6264 598
rect 6298 564 6354 598
rect 6388 564 6440 598
rect 5760 508 6440 564
rect 5760 474 5814 508
rect 5848 474 5904 508
rect 5938 474 5994 508
rect 6028 474 6084 508
rect 6118 474 6174 508
rect 6208 474 6264 508
rect 6298 474 6354 508
rect 6388 474 6440 508
rect 5760 418 6440 474
rect 5760 384 5814 418
rect 5848 384 5904 418
rect 5938 384 5994 418
rect 6028 384 6084 418
rect 6118 384 6174 418
rect 6208 384 6264 418
rect 6298 384 6354 418
rect 6388 384 6440 418
rect 5760 330 6440 384
rect 7120 958 7800 1010
rect 7120 924 7174 958
rect 7208 924 7264 958
rect 7298 924 7354 958
rect 7388 924 7444 958
rect 7478 924 7534 958
rect 7568 924 7624 958
rect 7658 924 7714 958
rect 7748 924 7800 958
rect 7120 868 7800 924
rect 7120 834 7174 868
rect 7208 834 7264 868
rect 7298 834 7354 868
rect 7388 834 7444 868
rect 7478 834 7534 868
rect 7568 834 7624 868
rect 7658 834 7714 868
rect 7748 834 7800 868
rect 7120 778 7800 834
rect 7120 744 7174 778
rect 7208 744 7264 778
rect 7298 744 7354 778
rect 7388 744 7444 778
rect 7478 744 7534 778
rect 7568 744 7624 778
rect 7658 744 7714 778
rect 7748 744 7800 778
rect 7120 688 7800 744
rect 7120 654 7174 688
rect 7208 654 7264 688
rect 7298 654 7354 688
rect 7388 654 7444 688
rect 7478 654 7534 688
rect 7568 654 7624 688
rect 7658 654 7714 688
rect 7748 654 7800 688
rect 7120 598 7800 654
rect 7120 564 7174 598
rect 7208 564 7264 598
rect 7298 564 7354 598
rect 7388 564 7444 598
rect 7478 564 7534 598
rect 7568 564 7624 598
rect 7658 564 7714 598
rect 7748 564 7800 598
rect 7120 508 7800 564
rect 7120 474 7174 508
rect 7208 474 7264 508
rect 7298 474 7354 508
rect 7388 474 7444 508
rect 7478 474 7534 508
rect 7568 474 7624 508
rect 7658 474 7714 508
rect 7748 474 7800 508
rect 7120 418 7800 474
rect 7120 384 7174 418
rect 7208 384 7264 418
rect 7298 384 7354 418
rect 7388 384 7444 418
rect 7478 384 7534 418
rect 7568 384 7624 418
rect 7658 384 7714 418
rect 7748 384 7800 418
rect 7120 330 7800 384
rect 8480 958 9160 1010
rect 8480 924 8534 958
rect 8568 924 8624 958
rect 8658 924 8714 958
rect 8748 924 8804 958
rect 8838 924 8894 958
rect 8928 924 8984 958
rect 9018 924 9074 958
rect 9108 924 9160 958
rect 8480 868 9160 924
rect 8480 834 8534 868
rect 8568 834 8624 868
rect 8658 834 8714 868
rect 8748 834 8804 868
rect 8838 834 8894 868
rect 8928 834 8984 868
rect 9018 834 9074 868
rect 9108 834 9160 868
rect 8480 778 9160 834
rect 8480 744 8534 778
rect 8568 744 8624 778
rect 8658 744 8714 778
rect 8748 744 8804 778
rect 8838 744 8894 778
rect 8928 744 8984 778
rect 9018 744 9074 778
rect 9108 744 9160 778
rect 8480 688 9160 744
rect 8480 654 8534 688
rect 8568 654 8624 688
rect 8658 654 8714 688
rect 8748 654 8804 688
rect 8838 654 8894 688
rect 8928 654 8984 688
rect 9018 654 9074 688
rect 9108 654 9160 688
rect 8480 598 9160 654
rect 8480 564 8534 598
rect 8568 564 8624 598
rect 8658 564 8714 598
rect 8748 564 8804 598
rect 8838 564 8894 598
rect 8928 564 8984 598
rect 9018 564 9074 598
rect 9108 564 9160 598
rect 8480 508 9160 564
rect 8480 474 8534 508
rect 8568 474 8624 508
rect 8658 474 8714 508
rect 8748 474 8804 508
rect 8838 474 8894 508
rect 8928 474 8984 508
rect 9018 474 9074 508
rect 9108 474 9160 508
rect 8480 418 9160 474
rect 8480 384 8534 418
rect 8568 384 8624 418
rect 8658 384 8714 418
rect 8748 384 8804 418
rect 8838 384 8894 418
rect 8928 384 8984 418
rect 9018 384 9074 418
rect 9108 384 9160 418
rect 8480 330 9160 384
<< ndiffc >>
rect 4430 5090 4470 5130
rect 4430 4990 4470 5030
rect 4430 4890 4470 4930
rect 4430 4790 4470 4830
rect 4430 4690 4470 4730
rect 4430 4590 4470 4630
rect 4430 4490 4470 4530
rect 4430 4390 4470 4430
rect 4630 5090 4670 5130
rect 4630 4990 4670 5030
rect 4630 4890 4670 4930
rect 4630 4790 4670 4830
rect 4630 4690 4670 4730
rect 4630 4590 4670 4630
rect 4630 4490 4670 4530
rect 4630 4390 4670 4430
rect 4830 5090 4870 5130
rect 4830 4990 4870 5030
rect 4830 4890 4870 4930
rect 4830 4790 4870 4830
rect 4830 4690 4870 4730
rect 4830 4590 4870 4630
rect 4830 4490 4870 4530
rect 4830 4390 4870 4430
rect 5030 5090 5070 5130
rect 5030 4990 5070 5030
rect 5030 4890 5070 4930
rect 5030 4790 5070 4830
rect 5030 4690 5070 4730
rect 5030 4590 5070 4630
rect 5030 4490 5070 4530
rect 5030 4390 5070 4430
rect 5230 5090 5270 5130
rect 5230 4990 5270 5030
rect 5230 4890 5270 4930
rect 5230 4790 5270 4830
rect 5230 4690 5270 4730
rect 5230 4590 5270 4630
rect 5230 4490 5270 4530
rect 5230 4390 5270 4430
rect 5430 5090 5470 5130
rect 5430 4990 5470 5030
rect 5430 4890 5470 4930
rect 5430 4790 5470 4830
rect 5430 4690 5470 4730
rect 5430 4590 5470 4630
rect 5430 4490 5470 4530
rect 5430 4390 5470 4430
rect 5630 5090 5670 5130
rect 5630 4990 5670 5030
rect 5630 4890 5670 4930
rect 5630 4790 5670 4830
rect 5630 4690 5670 4730
rect 5630 4590 5670 4630
rect 5630 4490 5670 4530
rect 5630 4390 5670 4430
rect 5830 5090 5870 5130
rect 5830 4990 5870 5030
rect 5830 4890 5870 4930
rect 5830 4790 5870 4830
rect 5830 4690 5870 4730
rect 5830 4590 5870 4630
rect 5830 4490 5870 4530
rect 5830 4390 5870 4430
rect 6030 5090 6070 5130
rect 6030 4990 6070 5030
rect 6030 4890 6070 4930
rect 6030 4790 6070 4830
rect 6030 4690 6070 4730
rect 6030 4590 6070 4630
rect 6030 4490 6070 4530
rect 6030 4390 6070 4430
rect 6230 5090 6270 5130
rect 6230 4990 6270 5030
rect 6230 4890 6270 4930
rect 6230 4790 6270 4830
rect 6230 4690 6270 4730
rect 6230 4590 6270 4630
rect 6230 4490 6270 4530
rect 6230 4390 6270 4430
rect 6430 5090 6470 5130
rect 6430 4990 6470 5030
rect 6430 4890 6470 4930
rect 6430 4790 6470 4830
rect 6430 4690 6470 4730
rect 6430 4590 6470 4630
rect 6430 4490 6470 4530
rect 6430 4390 6470 4430
rect 6630 5090 6670 5130
rect 6630 4990 6670 5030
rect 6630 4890 6670 4930
rect 6630 4790 6670 4830
rect 6630 4690 6670 4730
rect 6630 4590 6670 4630
rect 6630 4490 6670 4530
rect 6630 4390 6670 4430
rect 6830 5090 6870 5130
rect 6830 4990 6870 5030
rect 6830 4890 6870 4930
rect 6830 4790 6870 4830
rect 6830 4690 6870 4730
rect 6830 4590 6870 4630
rect 6830 4490 6870 4530
rect 6830 4390 6870 4430
rect 7030 5090 7070 5130
rect 7030 4990 7070 5030
rect 7030 4890 7070 4930
rect 7030 4790 7070 4830
rect 7030 4690 7070 4730
rect 7030 4590 7070 4630
rect 7030 4490 7070 4530
rect 7030 4390 7070 4430
rect 7230 5090 7270 5130
rect 7230 4990 7270 5030
rect 7230 4890 7270 4930
rect 7230 4790 7270 4830
rect 7230 4690 7270 4730
rect 7230 4590 7270 4630
rect 7230 4490 7270 4530
rect 7230 4390 7270 4430
rect 7430 5090 7470 5130
rect 7430 4990 7470 5030
rect 7430 4890 7470 4930
rect 7430 4790 7470 4830
rect 7430 4690 7470 4730
rect 7430 4590 7470 4630
rect 7430 4490 7470 4530
rect 7430 4390 7470 4430
rect 7630 5090 7670 5130
rect 7630 4990 7670 5030
rect 7630 4890 7670 4930
rect 7630 4790 7670 4830
rect 7630 4690 7670 4730
rect 7630 4590 7670 4630
rect 7630 4490 7670 4530
rect 7630 4390 7670 4430
rect 7830 5090 7870 5130
rect 7830 4990 7870 5030
rect 7830 4890 7870 4930
rect 7830 4790 7870 4830
rect 7830 4690 7870 4730
rect 7830 4590 7870 4630
rect 7830 4490 7870 4530
rect 7830 4390 7870 4430
rect 8030 5090 8070 5130
rect 8030 4990 8070 5030
rect 8030 4890 8070 4930
rect 8030 4790 8070 4830
rect 8030 4690 8070 4730
rect 8030 4590 8070 4630
rect 8030 4490 8070 4530
rect 8030 4390 8070 4430
rect 8230 5090 8270 5130
rect 8230 4990 8270 5030
rect 8230 4890 8270 4930
rect 8230 4790 8270 4830
rect 8230 4690 8270 4730
rect 8230 4590 8270 4630
rect 8230 4490 8270 4530
rect 8230 4390 8270 4430
rect 8430 5090 8470 5130
rect 8430 4990 8470 5030
rect 8430 4890 8470 4930
rect 8430 4790 8470 4830
rect 8430 4690 8470 4730
rect 8430 4590 8470 4630
rect 8430 4490 8470 4530
rect 8430 4390 8470 4430
rect 10350 4290 10390 4330
rect 10350 4190 10390 4230
rect 10350 4090 10390 4130
rect 10350 3990 10390 4030
rect 10460 4290 10500 4330
rect 10460 4190 10500 4230
rect 10460 4090 10500 4130
rect 10460 3990 10500 4030
rect 10600 4290 10640 4330
rect 10600 4190 10640 4230
rect 10600 4090 10640 4130
rect 10600 3990 10640 4030
rect 10710 4290 10750 4330
rect 10710 4190 10750 4230
rect 10710 4090 10750 4130
rect 10710 3990 10750 4030
rect 4470 3780 4510 3820
rect 4470 3680 4510 3720
rect 4470 3580 4510 3620
rect 4470 3480 4510 3520
rect 4670 3780 4710 3820
rect 4670 3680 4710 3720
rect 4670 3580 4710 3620
rect 4670 3480 4710 3520
rect 4870 3780 4910 3820
rect 4870 3680 4910 3720
rect 4870 3580 4910 3620
rect 4870 3480 4910 3520
rect 5070 3780 5110 3820
rect 5070 3680 5110 3720
rect 5070 3580 5110 3620
rect 5070 3480 5110 3520
rect 5270 3780 5310 3820
rect 5270 3680 5310 3720
rect 5270 3580 5310 3620
rect 5270 3480 5310 3520
rect 5470 3780 5510 3820
rect 5470 3680 5510 3720
rect 5470 3580 5510 3620
rect 5470 3480 5510 3520
rect 5670 3780 5710 3820
rect 5830 3780 5870 3820
rect 5670 3680 5710 3720
rect 5830 3680 5870 3720
rect 5670 3580 5710 3620
rect 5830 3580 5870 3620
rect 5670 3480 5710 3520
rect 5830 3480 5870 3520
rect 6030 3780 6070 3820
rect 6030 3680 6070 3720
rect 6030 3580 6070 3620
rect 6030 3480 6070 3520
rect 6230 3780 6270 3820
rect 6230 3680 6270 3720
rect 6230 3580 6270 3620
rect 6230 3480 6270 3520
rect 6430 3780 6470 3820
rect 6430 3680 6470 3720
rect 6430 3580 6470 3620
rect 6430 3480 6470 3520
rect 6630 3780 6670 3820
rect 6630 3680 6670 3720
rect 6630 3580 6670 3620
rect 6630 3480 6670 3520
rect 6830 3780 6870 3820
rect 6830 3680 6870 3720
rect 6830 3580 6870 3620
rect 6830 3480 6870 3520
rect 7030 3780 7070 3820
rect 7190 3780 7230 3820
rect 7030 3680 7070 3720
rect 7190 3680 7230 3720
rect 7030 3580 7070 3620
rect 7190 3580 7230 3620
rect 7030 3480 7070 3520
rect 7190 3480 7230 3520
rect 7390 3780 7430 3820
rect 7390 3680 7430 3720
rect 7390 3580 7430 3620
rect 7390 3480 7430 3520
rect 7590 3780 7630 3820
rect 7590 3680 7630 3720
rect 7590 3580 7630 3620
rect 7590 3480 7630 3520
rect 7790 3780 7830 3820
rect 7790 3680 7830 3720
rect 7790 3580 7830 3620
rect 7790 3480 7830 3520
rect 7990 3780 8030 3820
rect 7990 3680 8030 3720
rect 7990 3580 8030 3620
rect 7990 3480 8030 3520
rect 8190 3780 8230 3820
rect 8190 3680 8230 3720
rect 8190 3580 8230 3620
rect 8190 3480 8230 3520
rect 8390 3780 8430 3820
rect 8390 3680 8430 3720
rect 8390 3580 8430 3620
rect 8390 3480 8430 3520
rect 9230 3590 9270 3630
rect 9230 3490 9270 3530
rect 11310 3590 11350 3630
rect 11310 3490 11350 3530
rect 5150 2970 5190 3010
rect 5150 2870 5190 2910
rect 5350 2970 5390 3010
rect 5350 2870 5390 2910
rect 5550 2970 5590 3010
rect 5550 2870 5590 2910
rect 5750 2970 5790 3010
rect 5750 2870 5790 2910
rect 5950 2970 5990 3010
rect 5950 2870 5990 2910
rect 6150 2970 6190 3010
rect 6150 2870 6190 2910
rect 6350 2970 6390 3010
rect 6510 2970 6550 3010
rect 6350 2870 6390 2910
rect 6510 2870 6550 2910
rect 6710 2970 6750 3010
rect 6710 2870 6750 2910
rect 6910 2970 6950 3010
rect 6910 2870 6950 2910
rect 7110 2970 7150 3010
rect 7110 2870 7150 2910
rect 7310 2970 7350 3010
rect 7310 2870 7350 2910
rect 7510 2970 7550 3010
rect 7510 2870 7550 2910
rect 7710 2970 7750 3010
rect 7710 2870 7750 2910
rect 4670 2420 4710 2460
rect 4670 2320 4710 2360
rect 4670 2220 4710 2260
rect 4670 2120 4710 2160
rect 4670 2020 4710 2060
rect 4670 1920 4710 1960
rect 4670 1820 4710 1860
rect 4670 1720 4710 1760
rect 5550 2420 5590 2460
rect 5550 2320 5590 2360
rect 5550 2220 5590 2260
rect 5550 2120 5590 2160
rect 5550 2020 5590 2060
rect 5550 1920 5590 1960
rect 5550 1820 5590 1860
rect 5550 1720 5590 1760
rect 6430 2420 6470 2460
rect 6430 2320 6470 2360
rect 6430 2220 6470 2260
rect 6430 2120 6470 2160
rect 6430 2020 6470 2060
rect 6430 1920 6470 1960
rect 6430 1820 6470 1860
rect 6430 1720 6470 1760
rect 7310 2420 7350 2460
rect 7310 2320 7350 2360
rect 7310 2220 7350 2260
rect 7310 2120 7350 2160
rect 7310 2020 7350 2060
rect 7310 1920 7350 1960
rect 7310 1820 7350 1860
rect 7310 1720 7350 1760
rect 8190 2420 8230 2460
rect 8190 2320 8230 2360
rect 8190 2220 8230 2260
rect 8190 2120 8230 2160
rect 8190 2020 8230 2060
rect 8190 1920 8230 1960
rect 8190 1820 8230 1860
rect 8190 1720 8230 1760
<< pdiffc >>
rect 1734 924 1768 958
rect 1824 924 1858 958
rect 1914 924 1948 958
rect 2004 924 2038 958
rect 2094 924 2128 958
rect 2184 924 2218 958
rect 2274 924 2308 958
rect 1734 834 1768 868
rect 1824 834 1858 868
rect 1914 834 1948 868
rect 2004 834 2038 868
rect 2094 834 2128 868
rect 2184 834 2218 868
rect 2274 834 2308 868
rect 1734 744 1768 778
rect 1824 744 1858 778
rect 1914 744 1948 778
rect 2004 744 2038 778
rect 2094 744 2128 778
rect 2184 744 2218 778
rect 2274 744 2308 778
rect 1734 654 1768 688
rect 1824 654 1858 688
rect 1914 654 1948 688
rect 2004 654 2038 688
rect 2094 654 2128 688
rect 2184 654 2218 688
rect 2274 654 2308 688
rect 1734 564 1768 598
rect 1824 564 1858 598
rect 1914 564 1948 598
rect 2004 564 2038 598
rect 2094 564 2128 598
rect 2184 564 2218 598
rect 2274 564 2308 598
rect 1734 474 1768 508
rect 1824 474 1858 508
rect 1914 474 1948 508
rect 2004 474 2038 508
rect 2094 474 2128 508
rect 2184 474 2218 508
rect 2274 474 2308 508
rect 1734 384 1768 418
rect 1824 384 1858 418
rect 1914 384 1948 418
rect 2004 384 2038 418
rect 2094 384 2128 418
rect 2184 384 2218 418
rect 2274 384 2308 418
rect 3094 924 3128 958
rect 3184 924 3218 958
rect 3274 924 3308 958
rect 3364 924 3398 958
rect 3454 924 3488 958
rect 3544 924 3578 958
rect 3634 924 3668 958
rect 3094 834 3128 868
rect 3184 834 3218 868
rect 3274 834 3308 868
rect 3364 834 3398 868
rect 3454 834 3488 868
rect 3544 834 3578 868
rect 3634 834 3668 868
rect 3094 744 3128 778
rect 3184 744 3218 778
rect 3274 744 3308 778
rect 3364 744 3398 778
rect 3454 744 3488 778
rect 3544 744 3578 778
rect 3634 744 3668 778
rect 3094 654 3128 688
rect 3184 654 3218 688
rect 3274 654 3308 688
rect 3364 654 3398 688
rect 3454 654 3488 688
rect 3544 654 3578 688
rect 3634 654 3668 688
rect 3094 564 3128 598
rect 3184 564 3218 598
rect 3274 564 3308 598
rect 3364 564 3398 598
rect 3454 564 3488 598
rect 3544 564 3578 598
rect 3634 564 3668 598
rect 3094 474 3128 508
rect 3184 474 3218 508
rect 3274 474 3308 508
rect 3364 474 3398 508
rect 3454 474 3488 508
rect 3544 474 3578 508
rect 3634 474 3668 508
rect 3094 384 3128 418
rect 3184 384 3218 418
rect 3274 384 3308 418
rect 3364 384 3398 418
rect 3454 384 3488 418
rect 3544 384 3578 418
rect 3634 384 3668 418
rect 4454 924 4488 958
rect 4544 924 4578 958
rect 4634 924 4668 958
rect 4724 924 4758 958
rect 4814 924 4848 958
rect 4904 924 4938 958
rect 4994 924 5028 958
rect 4454 834 4488 868
rect 4544 834 4578 868
rect 4634 834 4668 868
rect 4724 834 4758 868
rect 4814 834 4848 868
rect 4904 834 4938 868
rect 4994 834 5028 868
rect 4454 744 4488 778
rect 4544 744 4578 778
rect 4634 744 4668 778
rect 4724 744 4758 778
rect 4814 744 4848 778
rect 4904 744 4938 778
rect 4994 744 5028 778
rect 4454 654 4488 688
rect 4544 654 4578 688
rect 4634 654 4668 688
rect 4724 654 4758 688
rect 4814 654 4848 688
rect 4904 654 4938 688
rect 4994 654 5028 688
rect 4454 564 4488 598
rect 4544 564 4578 598
rect 4634 564 4668 598
rect 4724 564 4758 598
rect 4814 564 4848 598
rect 4904 564 4938 598
rect 4994 564 5028 598
rect 4454 474 4488 508
rect 4544 474 4578 508
rect 4634 474 4668 508
rect 4724 474 4758 508
rect 4814 474 4848 508
rect 4904 474 4938 508
rect 4994 474 5028 508
rect 4454 384 4488 418
rect 4544 384 4578 418
rect 4634 384 4668 418
rect 4724 384 4758 418
rect 4814 384 4848 418
rect 4904 384 4938 418
rect 4994 384 5028 418
rect 5814 924 5848 958
rect 5904 924 5938 958
rect 5994 924 6028 958
rect 6084 924 6118 958
rect 6174 924 6208 958
rect 6264 924 6298 958
rect 6354 924 6388 958
rect 5814 834 5848 868
rect 5904 834 5938 868
rect 5994 834 6028 868
rect 6084 834 6118 868
rect 6174 834 6208 868
rect 6264 834 6298 868
rect 6354 834 6388 868
rect 5814 744 5848 778
rect 5904 744 5938 778
rect 5994 744 6028 778
rect 6084 744 6118 778
rect 6174 744 6208 778
rect 6264 744 6298 778
rect 6354 744 6388 778
rect 5814 654 5848 688
rect 5904 654 5938 688
rect 5994 654 6028 688
rect 6084 654 6118 688
rect 6174 654 6208 688
rect 6264 654 6298 688
rect 6354 654 6388 688
rect 5814 564 5848 598
rect 5904 564 5938 598
rect 5994 564 6028 598
rect 6084 564 6118 598
rect 6174 564 6208 598
rect 6264 564 6298 598
rect 6354 564 6388 598
rect 5814 474 5848 508
rect 5904 474 5938 508
rect 5994 474 6028 508
rect 6084 474 6118 508
rect 6174 474 6208 508
rect 6264 474 6298 508
rect 6354 474 6388 508
rect 5814 384 5848 418
rect 5904 384 5938 418
rect 5994 384 6028 418
rect 6084 384 6118 418
rect 6174 384 6208 418
rect 6264 384 6298 418
rect 6354 384 6388 418
rect 7174 924 7208 958
rect 7264 924 7298 958
rect 7354 924 7388 958
rect 7444 924 7478 958
rect 7534 924 7568 958
rect 7624 924 7658 958
rect 7714 924 7748 958
rect 7174 834 7208 868
rect 7264 834 7298 868
rect 7354 834 7388 868
rect 7444 834 7478 868
rect 7534 834 7568 868
rect 7624 834 7658 868
rect 7714 834 7748 868
rect 7174 744 7208 778
rect 7264 744 7298 778
rect 7354 744 7388 778
rect 7444 744 7478 778
rect 7534 744 7568 778
rect 7624 744 7658 778
rect 7714 744 7748 778
rect 7174 654 7208 688
rect 7264 654 7298 688
rect 7354 654 7388 688
rect 7444 654 7478 688
rect 7534 654 7568 688
rect 7624 654 7658 688
rect 7714 654 7748 688
rect 7174 564 7208 598
rect 7264 564 7298 598
rect 7354 564 7388 598
rect 7444 564 7478 598
rect 7534 564 7568 598
rect 7624 564 7658 598
rect 7714 564 7748 598
rect 7174 474 7208 508
rect 7264 474 7298 508
rect 7354 474 7388 508
rect 7444 474 7478 508
rect 7534 474 7568 508
rect 7624 474 7658 508
rect 7714 474 7748 508
rect 7174 384 7208 418
rect 7264 384 7298 418
rect 7354 384 7388 418
rect 7444 384 7478 418
rect 7534 384 7568 418
rect 7624 384 7658 418
rect 7714 384 7748 418
rect 8534 924 8568 958
rect 8624 924 8658 958
rect 8714 924 8748 958
rect 8804 924 8838 958
rect 8894 924 8928 958
rect 8984 924 9018 958
rect 9074 924 9108 958
rect 8534 834 8568 868
rect 8624 834 8658 868
rect 8714 834 8748 868
rect 8804 834 8838 868
rect 8894 834 8928 868
rect 8984 834 9018 868
rect 9074 834 9108 868
rect 8534 744 8568 778
rect 8624 744 8658 778
rect 8714 744 8748 778
rect 8804 744 8838 778
rect 8894 744 8928 778
rect 8984 744 9018 778
rect 9074 744 9108 778
rect 8534 654 8568 688
rect 8624 654 8658 688
rect 8714 654 8748 688
rect 8804 654 8838 688
rect 8894 654 8928 688
rect 8984 654 9018 688
rect 9074 654 9108 688
rect 8534 564 8568 598
rect 8624 564 8658 598
rect 8714 564 8748 598
rect 8804 564 8838 598
rect 8894 564 8928 598
rect 8984 564 9018 598
rect 9074 564 9108 598
rect 8534 474 8568 508
rect 8624 474 8658 508
rect 8714 474 8748 508
rect 8804 474 8838 508
rect 8894 474 8928 508
rect 8984 474 9018 508
rect 9074 474 9108 508
rect 8534 384 8568 418
rect 8624 384 8658 418
rect 8714 384 8748 418
rect 8804 384 8838 418
rect 8894 384 8928 418
rect 8984 384 9018 418
rect 9074 384 9108 418
<< psubdiff >>
rect 4330 5130 4410 5160
rect 4330 5090 4350 5130
rect 4390 5090 4410 5130
rect 4330 5030 4410 5090
rect 4330 4990 4350 5030
rect 4390 4990 4410 5030
rect 4330 4930 4410 4990
rect 4330 4890 4350 4930
rect 4390 4890 4410 4930
rect 4330 4830 4410 4890
rect 4330 4790 4350 4830
rect 4390 4790 4410 4830
rect 4330 4730 4410 4790
rect 4330 4690 4350 4730
rect 4390 4690 4410 4730
rect 4330 4630 4410 4690
rect 4330 4590 4350 4630
rect 4390 4590 4410 4630
rect 4330 4530 4410 4590
rect 4330 4490 4350 4530
rect 4390 4490 4410 4530
rect 4330 4430 4410 4490
rect 4330 4390 4350 4430
rect 4390 4390 4410 4430
rect 4330 4360 4410 4390
rect 8490 5130 8570 5160
rect 8490 5090 8510 5130
rect 8550 5090 8570 5130
rect 8490 5030 8570 5090
rect 8490 4990 8510 5030
rect 8550 4990 8570 5030
rect 8490 4930 8570 4990
rect 8490 4890 8510 4930
rect 8550 4890 8570 4930
rect 8490 4830 8570 4890
rect 8490 4790 8510 4830
rect 8550 4790 8570 4830
rect 8490 4730 8570 4790
rect 8490 4690 8510 4730
rect 8550 4690 8570 4730
rect 8490 4630 8570 4690
rect 8490 4590 8510 4630
rect 8550 4590 8570 4630
rect 8490 4530 8570 4590
rect 8490 4490 8510 4530
rect 8550 4490 8570 4530
rect 8490 4430 8570 4490
rect 8490 4390 8510 4430
rect 8550 4390 8570 4430
rect 8490 4360 8570 4390
rect 10250 4330 10330 4360
rect 10250 4290 10270 4330
rect 10310 4290 10330 4330
rect 10250 4230 10330 4290
rect 10250 4190 10270 4230
rect 10310 4190 10330 4230
rect 10250 4130 10330 4190
rect 10250 4090 10270 4130
rect 10310 4090 10330 4130
rect 10250 4030 10330 4090
rect 10250 3990 10270 4030
rect 10310 3990 10330 4030
rect 10250 3960 10330 3990
rect 10770 4330 10850 4360
rect 10770 4290 10790 4330
rect 10830 4290 10850 4330
rect 10770 4230 10850 4290
rect 10770 4190 10790 4230
rect 10830 4190 10850 4230
rect 10770 4130 10850 4190
rect 10770 4090 10790 4130
rect 10830 4090 10850 4130
rect 10770 4030 10850 4090
rect 10770 3990 10790 4030
rect 10830 3990 10850 4030
rect 10770 3960 10850 3990
rect 4370 3820 4450 3850
rect 4370 3780 4390 3820
rect 4430 3780 4450 3820
rect 4370 3720 4450 3780
rect 4370 3680 4390 3720
rect 4430 3680 4450 3720
rect 4370 3620 4450 3680
rect 4370 3580 4390 3620
rect 4430 3580 4450 3620
rect 4370 3520 4450 3580
rect 4370 3480 4390 3520
rect 4430 3480 4450 3520
rect 4370 3450 4450 3480
rect 5730 3820 5810 3850
rect 5730 3780 5750 3820
rect 5790 3780 5810 3820
rect 5730 3720 5810 3780
rect 5730 3680 5750 3720
rect 5790 3680 5810 3720
rect 5730 3620 5810 3680
rect 5730 3580 5750 3620
rect 5790 3580 5810 3620
rect 5730 3520 5810 3580
rect 5730 3480 5750 3520
rect 5790 3480 5810 3520
rect 5730 3450 5810 3480
rect 7090 3820 7170 3850
rect 7090 3780 7110 3820
rect 7150 3780 7170 3820
rect 7090 3720 7170 3780
rect 7090 3680 7110 3720
rect 7150 3680 7170 3720
rect 7090 3620 7170 3680
rect 7090 3580 7110 3620
rect 7150 3580 7170 3620
rect 7090 3520 7170 3580
rect 7090 3480 7110 3520
rect 7150 3480 7170 3520
rect 7090 3450 7170 3480
rect 8450 3820 8530 3850
rect 8450 3780 8470 3820
rect 8510 3780 8530 3820
rect 8450 3720 8530 3780
rect 8450 3680 8470 3720
rect 8510 3680 8530 3720
rect 8450 3620 8530 3680
rect 8450 3580 8470 3620
rect 8510 3580 8530 3620
rect 8450 3520 8530 3580
rect 8450 3480 8470 3520
rect 8510 3480 8530 3520
rect 8450 3450 8530 3480
rect 11370 3630 11450 3660
rect 11370 3590 11390 3630
rect 11430 3590 11450 3630
rect 11370 3530 11450 3590
rect 11370 3490 11390 3530
rect 11430 3490 11450 3530
rect 11370 3460 11450 3490
rect 5050 3010 5130 3040
rect 5050 2970 5070 3010
rect 5110 2970 5130 3010
rect 5050 2910 5130 2970
rect 5050 2870 5070 2910
rect 5110 2870 5130 2910
rect 5050 2840 5130 2870
rect 6410 3010 6490 3040
rect 6410 2970 6430 3010
rect 6470 2970 6490 3010
rect 6410 2910 6490 2970
rect 6410 2870 6430 2910
rect 6470 2870 6490 2910
rect 6410 2840 6490 2870
rect 7770 3010 7850 3040
rect 7770 2970 7790 3010
rect 7830 2970 7850 3010
rect 7770 2910 7850 2970
rect 7770 2870 7790 2910
rect 7830 2870 7850 2910
rect 7770 2840 7850 2870
rect 4570 2460 4650 2490
rect 4570 2420 4590 2460
rect 4630 2420 4650 2460
rect 4570 2360 4650 2420
rect 4570 2320 4590 2360
rect 4630 2320 4650 2360
rect 4570 2260 4650 2320
rect 4570 2220 4590 2260
rect 4630 2220 4650 2260
rect 4570 2160 4650 2220
rect 4570 2120 4590 2160
rect 4630 2120 4650 2160
rect 4570 2060 4650 2120
rect 4570 2020 4590 2060
rect 4630 2020 4650 2060
rect 4570 1960 4650 2020
rect 4570 1920 4590 1960
rect 4630 1920 4650 1960
rect 4570 1860 4650 1920
rect 4570 1820 4590 1860
rect 4630 1820 4650 1860
rect 4570 1760 4650 1820
rect 4570 1720 4590 1760
rect 4630 1720 4650 1760
rect 4570 1690 4650 1720
rect 8250 2460 8330 2490
rect 8250 2420 8270 2460
rect 8310 2420 8330 2460
rect 8250 2360 8330 2420
rect 8250 2320 8270 2360
rect 8310 2320 8330 2360
rect 8250 2260 8330 2320
rect 8250 2220 8270 2260
rect 8310 2220 8330 2260
rect 8250 2160 8330 2220
rect 8250 2120 8270 2160
rect 8310 2120 8330 2160
rect 8250 2060 8330 2120
rect 8250 2020 8270 2060
rect 8310 2020 8330 2060
rect 8250 1960 8330 2020
rect 8250 1920 8270 1960
rect 8310 1920 8330 1960
rect 8250 1860 8330 1920
rect 8250 1820 8270 1860
rect 8310 1820 8330 1860
rect 8250 1760 8330 1820
rect 8250 1720 8270 1760
rect 8310 1720 8330 1760
rect 8250 1690 8330 1720
rect 1376 1279 2664 1314
rect 1376 1256 1506 1279
rect 1376 1222 1410 1256
rect 1444 1245 1506 1256
rect 1540 1245 1596 1279
rect 1630 1245 1686 1279
rect 1720 1245 1776 1279
rect 1810 1245 1866 1279
rect 1900 1245 1956 1279
rect 1990 1245 2046 1279
rect 2080 1245 2136 1279
rect 2170 1245 2226 1279
rect 2260 1245 2316 1279
rect 2350 1245 2406 1279
rect 2440 1245 2496 1279
rect 2530 1256 2664 1279
rect 2530 1245 2597 1256
rect 1444 1222 2597 1245
rect 2631 1222 2664 1256
rect 1376 1213 2664 1222
rect 1376 1166 1477 1213
rect 1376 1132 1410 1166
rect 1444 1132 1477 1166
rect 2563 1166 2664 1213
rect 1376 1076 1477 1132
rect 1376 1042 1410 1076
rect 1444 1042 1477 1076
rect 1376 986 1477 1042
rect 1376 952 1410 986
rect 1444 952 1477 986
rect 1376 896 1477 952
rect 1376 862 1410 896
rect 1444 862 1477 896
rect 1376 806 1477 862
rect 1376 772 1410 806
rect 1444 772 1477 806
rect 1376 716 1477 772
rect 1376 682 1410 716
rect 1444 682 1477 716
rect 1376 626 1477 682
rect 1376 592 1410 626
rect 1444 592 1477 626
rect 1376 536 1477 592
rect 1376 502 1410 536
rect 1444 502 1477 536
rect 1376 446 1477 502
rect 1376 412 1410 446
rect 1444 412 1477 446
rect 1376 356 1477 412
rect 1376 322 1410 356
rect 1444 322 1477 356
rect 1376 266 1477 322
rect 1376 232 1410 266
rect 1444 232 1477 266
rect 1376 176 1477 232
rect 2563 1132 2597 1166
rect 2631 1132 2664 1166
rect 2563 1076 2664 1132
rect 2563 1042 2597 1076
rect 2631 1042 2664 1076
rect 2563 986 2664 1042
rect 2563 952 2597 986
rect 2631 952 2664 986
rect 2563 896 2664 952
rect 2563 862 2597 896
rect 2631 862 2664 896
rect 2563 806 2664 862
rect 2563 772 2597 806
rect 2631 772 2664 806
rect 2563 716 2664 772
rect 2563 682 2597 716
rect 2631 682 2664 716
rect 2563 626 2664 682
rect 2563 592 2597 626
rect 2631 592 2664 626
rect 2563 536 2664 592
rect 2563 502 2597 536
rect 2631 502 2664 536
rect 2563 446 2664 502
rect 2563 412 2597 446
rect 2631 412 2664 446
rect 2563 356 2664 412
rect 2563 322 2597 356
rect 2631 322 2664 356
rect 2563 266 2664 322
rect 2563 232 2597 266
rect 2631 232 2664 266
rect 1376 142 1410 176
rect 1444 142 1477 176
rect 1376 127 1477 142
rect 2563 176 2664 232
rect 2563 142 2597 176
rect 2631 142 2664 176
rect 2563 127 2664 142
rect 1376 92 2664 127
rect 1376 58 1506 92
rect 1540 58 1596 92
rect 1630 58 1686 92
rect 1720 58 1776 92
rect 1810 58 1866 92
rect 1900 58 1956 92
rect 1990 58 2046 92
rect 2080 58 2136 92
rect 2170 58 2226 92
rect 2260 58 2316 92
rect 2350 58 2406 92
rect 2440 58 2496 92
rect 2530 58 2664 92
rect 1376 26 2664 58
rect 2736 1279 4024 1314
rect 2736 1256 2866 1279
rect 2736 1222 2770 1256
rect 2804 1245 2866 1256
rect 2900 1245 2956 1279
rect 2990 1245 3046 1279
rect 3080 1245 3136 1279
rect 3170 1245 3226 1279
rect 3260 1245 3316 1279
rect 3350 1245 3406 1279
rect 3440 1245 3496 1279
rect 3530 1245 3586 1279
rect 3620 1245 3676 1279
rect 3710 1245 3766 1279
rect 3800 1245 3856 1279
rect 3890 1256 4024 1279
rect 3890 1245 3957 1256
rect 2804 1222 3957 1245
rect 3991 1222 4024 1256
rect 2736 1213 4024 1222
rect 2736 1166 2837 1213
rect 2736 1132 2770 1166
rect 2804 1132 2837 1166
rect 3923 1166 4024 1213
rect 2736 1076 2837 1132
rect 2736 1042 2770 1076
rect 2804 1042 2837 1076
rect 2736 986 2837 1042
rect 2736 952 2770 986
rect 2804 952 2837 986
rect 2736 896 2837 952
rect 2736 862 2770 896
rect 2804 862 2837 896
rect 2736 806 2837 862
rect 2736 772 2770 806
rect 2804 772 2837 806
rect 2736 716 2837 772
rect 2736 682 2770 716
rect 2804 682 2837 716
rect 2736 626 2837 682
rect 2736 592 2770 626
rect 2804 592 2837 626
rect 2736 536 2837 592
rect 2736 502 2770 536
rect 2804 502 2837 536
rect 2736 446 2837 502
rect 2736 412 2770 446
rect 2804 412 2837 446
rect 2736 356 2837 412
rect 2736 322 2770 356
rect 2804 322 2837 356
rect 2736 266 2837 322
rect 2736 232 2770 266
rect 2804 232 2837 266
rect 2736 176 2837 232
rect 3923 1132 3957 1166
rect 3991 1132 4024 1166
rect 3923 1076 4024 1132
rect 3923 1042 3957 1076
rect 3991 1042 4024 1076
rect 3923 986 4024 1042
rect 3923 952 3957 986
rect 3991 952 4024 986
rect 3923 896 4024 952
rect 3923 862 3957 896
rect 3991 862 4024 896
rect 3923 806 4024 862
rect 3923 772 3957 806
rect 3991 772 4024 806
rect 3923 716 4024 772
rect 3923 682 3957 716
rect 3991 682 4024 716
rect 3923 626 4024 682
rect 3923 592 3957 626
rect 3991 592 4024 626
rect 3923 536 4024 592
rect 3923 502 3957 536
rect 3991 502 4024 536
rect 3923 446 4024 502
rect 3923 412 3957 446
rect 3991 412 4024 446
rect 3923 356 4024 412
rect 3923 322 3957 356
rect 3991 322 4024 356
rect 3923 266 4024 322
rect 3923 232 3957 266
rect 3991 232 4024 266
rect 2736 142 2770 176
rect 2804 142 2837 176
rect 2736 127 2837 142
rect 3923 176 4024 232
rect 3923 142 3957 176
rect 3991 142 4024 176
rect 3923 127 4024 142
rect 2736 92 4024 127
rect 2736 58 2866 92
rect 2900 58 2956 92
rect 2990 58 3046 92
rect 3080 58 3136 92
rect 3170 58 3226 92
rect 3260 58 3316 92
rect 3350 58 3406 92
rect 3440 58 3496 92
rect 3530 58 3586 92
rect 3620 58 3676 92
rect 3710 58 3766 92
rect 3800 58 3856 92
rect 3890 58 4024 92
rect 2736 26 4024 58
rect 4096 1279 5384 1314
rect 4096 1256 4226 1279
rect 4096 1222 4130 1256
rect 4164 1245 4226 1256
rect 4260 1245 4316 1279
rect 4350 1245 4406 1279
rect 4440 1245 4496 1279
rect 4530 1245 4586 1279
rect 4620 1245 4676 1279
rect 4710 1245 4766 1279
rect 4800 1245 4856 1279
rect 4890 1245 4946 1279
rect 4980 1245 5036 1279
rect 5070 1245 5126 1279
rect 5160 1245 5216 1279
rect 5250 1256 5384 1279
rect 5250 1245 5317 1256
rect 4164 1222 5317 1245
rect 5351 1222 5384 1256
rect 4096 1213 5384 1222
rect 4096 1166 4197 1213
rect 4096 1132 4130 1166
rect 4164 1132 4197 1166
rect 5283 1166 5384 1213
rect 4096 1076 4197 1132
rect 4096 1042 4130 1076
rect 4164 1042 4197 1076
rect 4096 986 4197 1042
rect 4096 952 4130 986
rect 4164 952 4197 986
rect 4096 896 4197 952
rect 4096 862 4130 896
rect 4164 862 4197 896
rect 4096 806 4197 862
rect 4096 772 4130 806
rect 4164 772 4197 806
rect 4096 716 4197 772
rect 4096 682 4130 716
rect 4164 682 4197 716
rect 4096 626 4197 682
rect 4096 592 4130 626
rect 4164 592 4197 626
rect 4096 536 4197 592
rect 4096 502 4130 536
rect 4164 502 4197 536
rect 4096 446 4197 502
rect 4096 412 4130 446
rect 4164 412 4197 446
rect 4096 356 4197 412
rect 4096 322 4130 356
rect 4164 322 4197 356
rect 4096 266 4197 322
rect 4096 232 4130 266
rect 4164 232 4197 266
rect 4096 176 4197 232
rect 5283 1132 5317 1166
rect 5351 1132 5384 1166
rect 5283 1076 5384 1132
rect 5283 1042 5317 1076
rect 5351 1042 5384 1076
rect 5283 986 5384 1042
rect 5283 952 5317 986
rect 5351 952 5384 986
rect 5283 896 5384 952
rect 5283 862 5317 896
rect 5351 862 5384 896
rect 5283 806 5384 862
rect 5283 772 5317 806
rect 5351 772 5384 806
rect 5283 716 5384 772
rect 5283 682 5317 716
rect 5351 682 5384 716
rect 5283 626 5384 682
rect 5283 592 5317 626
rect 5351 592 5384 626
rect 5283 536 5384 592
rect 5283 502 5317 536
rect 5351 502 5384 536
rect 5283 446 5384 502
rect 5283 412 5317 446
rect 5351 412 5384 446
rect 5283 356 5384 412
rect 5283 322 5317 356
rect 5351 322 5384 356
rect 5283 266 5384 322
rect 5283 232 5317 266
rect 5351 232 5384 266
rect 4096 142 4130 176
rect 4164 142 4197 176
rect 4096 127 4197 142
rect 5283 176 5384 232
rect 5283 142 5317 176
rect 5351 142 5384 176
rect 5283 127 5384 142
rect 4096 92 5384 127
rect 4096 58 4226 92
rect 4260 58 4316 92
rect 4350 58 4406 92
rect 4440 58 4496 92
rect 4530 58 4586 92
rect 4620 58 4676 92
rect 4710 58 4766 92
rect 4800 58 4856 92
rect 4890 58 4946 92
rect 4980 58 5036 92
rect 5070 58 5126 92
rect 5160 58 5216 92
rect 5250 58 5384 92
rect 4096 26 5384 58
rect 5456 1279 6744 1314
rect 5456 1256 5586 1279
rect 5456 1222 5490 1256
rect 5524 1245 5586 1256
rect 5620 1245 5676 1279
rect 5710 1245 5766 1279
rect 5800 1245 5856 1279
rect 5890 1245 5946 1279
rect 5980 1245 6036 1279
rect 6070 1245 6126 1279
rect 6160 1245 6216 1279
rect 6250 1245 6306 1279
rect 6340 1245 6396 1279
rect 6430 1245 6486 1279
rect 6520 1245 6576 1279
rect 6610 1256 6744 1279
rect 6610 1245 6677 1256
rect 5524 1222 6677 1245
rect 6711 1222 6744 1256
rect 5456 1213 6744 1222
rect 5456 1166 5557 1213
rect 5456 1132 5490 1166
rect 5524 1132 5557 1166
rect 6643 1166 6744 1213
rect 5456 1076 5557 1132
rect 5456 1042 5490 1076
rect 5524 1042 5557 1076
rect 5456 986 5557 1042
rect 5456 952 5490 986
rect 5524 952 5557 986
rect 5456 896 5557 952
rect 5456 862 5490 896
rect 5524 862 5557 896
rect 5456 806 5557 862
rect 5456 772 5490 806
rect 5524 772 5557 806
rect 5456 716 5557 772
rect 5456 682 5490 716
rect 5524 682 5557 716
rect 5456 626 5557 682
rect 5456 592 5490 626
rect 5524 592 5557 626
rect 5456 536 5557 592
rect 5456 502 5490 536
rect 5524 502 5557 536
rect 5456 446 5557 502
rect 5456 412 5490 446
rect 5524 412 5557 446
rect 5456 356 5557 412
rect 5456 322 5490 356
rect 5524 322 5557 356
rect 5456 266 5557 322
rect 5456 232 5490 266
rect 5524 232 5557 266
rect 5456 176 5557 232
rect 6643 1132 6677 1166
rect 6711 1132 6744 1166
rect 6643 1076 6744 1132
rect 6643 1042 6677 1076
rect 6711 1042 6744 1076
rect 6643 986 6744 1042
rect 6643 952 6677 986
rect 6711 952 6744 986
rect 6643 896 6744 952
rect 6643 862 6677 896
rect 6711 862 6744 896
rect 6643 806 6744 862
rect 6643 772 6677 806
rect 6711 772 6744 806
rect 6643 716 6744 772
rect 6643 682 6677 716
rect 6711 682 6744 716
rect 6643 626 6744 682
rect 6643 592 6677 626
rect 6711 592 6744 626
rect 6643 536 6744 592
rect 6643 502 6677 536
rect 6711 502 6744 536
rect 6643 446 6744 502
rect 6643 412 6677 446
rect 6711 412 6744 446
rect 6643 356 6744 412
rect 6643 322 6677 356
rect 6711 322 6744 356
rect 6643 266 6744 322
rect 6643 232 6677 266
rect 6711 232 6744 266
rect 5456 142 5490 176
rect 5524 142 5557 176
rect 5456 127 5557 142
rect 6643 176 6744 232
rect 6643 142 6677 176
rect 6711 142 6744 176
rect 6643 127 6744 142
rect 5456 92 6744 127
rect 5456 58 5586 92
rect 5620 58 5676 92
rect 5710 58 5766 92
rect 5800 58 5856 92
rect 5890 58 5946 92
rect 5980 58 6036 92
rect 6070 58 6126 92
rect 6160 58 6216 92
rect 6250 58 6306 92
rect 6340 58 6396 92
rect 6430 58 6486 92
rect 6520 58 6576 92
rect 6610 58 6744 92
rect 5456 26 6744 58
rect 6816 1279 8104 1314
rect 6816 1256 6946 1279
rect 6816 1222 6850 1256
rect 6884 1245 6946 1256
rect 6980 1245 7036 1279
rect 7070 1245 7126 1279
rect 7160 1245 7216 1279
rect 7250 1245 7306 1279
rect 7340 1245 7396 1279
rect 7430 1245 7486 1279
rect 7520 1245 7576 1279
rect 7610 1245 7666 1279
rect 7700 1245 7756 1279
rect 7790 1245 7846 1279
rect 7880 1245 7936 1279
rect 7970 1256 8104 1279
rect 7970 1245 8037 1256
rect 6884 1222 8037 1245
rect 8071 1222 8104 1256
rect 6816 1213 8104 1222
rect 6816 1166 6917 1213
rect 6816 1132 6850 1166
rect 6884 1132 6917 1166
rect 8003 1166 8104 1213
rect 6816 1076 6917 1132
rect 6816 1042 6850 1076
rect 6884 1042 6917 1076
rect 6816 986 6917 1042
rect 6816 952 6850 986
rect 6884 952 6917 986
rect 6816 896 6917 952
rect 6816 862 6850 896
rect 6884 862 6917 896
rect 6816 806 6917 862
rect 6816 772 6850 806
rect 6884 772 6917 806
rect 6816 716 6917 772
rect 6816 682 6850 716
rect 6884 682 6917 716
rect 6816 626 6917 682
rect 6816 592 6850 626
rect 6884 592 6917 626
rect 6816 536 6917 592
rect 6816 502 6850 536
rect 6884 502 6917 536
rect 6816 446 6917 502
rect 6816 412 6850 446
rect 6884 412 6917 446
rect 6816 356 6917 412
rect 6816 322 6850 356
rect 6884 322 6917 356
rect 6816 266 6917 322
rect 6816 232 6850 266
rect 6884 232 6917 266
rect 6816 176 6917 232
rect 8003 1132 8037 1166
rect 8071 1132 8104 1166
rect 8003 1076 8104 1132
rect 8003 1042 8037 1076
rect 8071 1042 8104 1076
rect 8003 986 8104 1042
rect 8003 952 8037 986
rect 8071 952 8104 986
rect 8003 896 8104 952
rect 8003 862 8037 896
rect 8071 862 8104 896
rect 8003 806 8104 862
rect 8003 772 8037 806
rect 8071 772 8104 806
rect 8003 716 8104 772
rect 8003 682 8037 716
rect 8071 682 8104 716
rect 8003 626 8104 682
rect 8003 592 8037 626
rect 8071 592 8104 626
rect 8003 536 8104 592
rect 8003 502 8037 536
rect 8071 502 8104 536
rect 8003 446 8104 502
rect 8003 412 8037 446
rect 8071 412 8104 446
rect 8003 356 8104 412
rect 8003 322 8037 356
rect 8071 322 8104 356
rect 8003 266 8104 322
rect 8003 232 8037 266
rect 8071 232 8104 266
rect 6816 142 6850 176
rect 6884 142 6917 176
rect 6816 127 6917 142
rect 8003 176 8104 232
rect 8003 142 8037 176
rect 8071 142 8104 176
rect 8003 127 8104 142
rect 6816 92 8104 127
rect 6816 58 6946 92
rect 6980 58 7036 92
rect 7070 58 7126 92
rect 7160 58 7216 92
rect 7250 58 7306 92
rect 7340 58 7396 92
rect 7430 58 7486 92
rect 7520 58 7576 92
rect 7610 58 7666 92
rect 7700 58 7756 92
rect 7790 58 7846 92
rect 7880 58 7936 92
rect 7970 58 8104 92
rect 6816 26 8104 58
rect 8176 1279 9464 1314
rect 8176 1256 8306 1279
rect 8176 1222 8210 1256
rect 8244 1245 8306 1256
rect 8340 1245 8396 1279
rect 8430 1245 8486 1279
rect 8520 1245 8576 1279
rect 8610 1245 8666 1279
rect 8700 1245 8756 1279
rect 8790 1245 8846 1279
rect 8880 1245 8936 1279
rect 8970 1245 9026 1279
rect 9060 1245 9116 1279
rect 9150 1245 9206 1279
rect 9240 1245 9296 1279
rect 9330 1256 9464 1279
rect 9330 1245 9397 1256
rect 8244 1222 9397 1245
rect 9431 1222 9464 1256
rect 8176 1213 9464 1222
rect 8176 1166 8277 1213
rect 8176 1132 8210 1166
rect 8244 1132 8277 1166
rect 9363 1166 9464 1213
rect 8176 1076 8277 1132
rect 8176 1042 8210 1076
rect 8244 1042 8277 1076
rect 8176 986 8277 1042
rect 8176 952 8210 986
rect 8244 952 8277 986
rect 8176 896 8277 952
rect 8176 862 8210 896
rect 8244 862 8277 896
rect 8176 806 8277 862
rect 8176 772 8210 806
rect 8244 772 8277 806
rect 8176 716 8277 772
rect 8176 682 8210 716
rect 8244 682 8277 716
rect 8176 626 8277 682
rect 8176 592 8210 626
rect 8244 592 8277 626
rect 8176 536 8277 592
rect 8176 502 8210 536
rect 8244 502 8277 536
rect 8176 446 8277 502
rect 8176 412 8210 446
rect 8244 412 8277 446
rect 8176 356 8277 412
rect 8176 322 8210 356
rect 8244 322 8277 356
rect 8176 266 8277 322
rect 8176 232 8210 266
rect 8244 232 8277 266
rect 8176 176 8277 232
rect 9363 1132 9397 1166
rect 9431 1132 9464 1166
rect 9363 1076 9464 1132
rect 9363 1042 9397 1076
rect 9431 1042 9464 1076
rect 9363 986 9464 1042
rect 9363 952 9397 986
rect 9431 952 9464 986
rect 9363 896 9464 952
rect 9363 862 9397 896
rect 9431 862 9464 896
rect 9363 806 9464 862
rect 9363 772 9397 806
rect 9431 772 9464 806
rect 9363 716 9464 772
rect 9363 682 9397 716
rect 9431 682 9464 716
rect 9363 626 9464 682
rect 9363 592 9397 626
rect 9431 592 9464 626
rect 9363 536 9464 592
rect 9363 502 9397 536
rect 9431 502 9464 536
rect 9363 446 9464 502
rect 9363 412 9397 446
rect 9431 412 9464 446
rect 9363 356 9464 412
rect 9363 322 9397 356
rect 9431 322 9464 356
rect 9363 266 9464 322
rect 9363 232 9397 266
rect 9431 232 9464 266
rect 8176 142 8210 176
rect 8244 142 8277 176
rect 8176 127 8277 142
rect 9363 176 9464 232
rect 9363 142 9397 176
rect 9431 142 9464 176
rect 9363 127 9464 142
rect 8176 92 9464 127
rect 8176 58 8306 92
rect 8340 58 8396 92
rect 8430 58 8486 92
rect 8520 58 8576 92
rect 8610 58 8666 92
rect 8700 58 8756 92
rect 8790 58 8846 92
rect 8880 58 8936 92
rect 8970 58 9026 92
rect 9060 58 9116 92
rect 9150 58 9206 92
rect 9240 58 9296 92
rect 9330 58 9464 92
rect 8176 26 9464 58
<< nsubdiff >>
rect 1539 1132 2501 1151
rect 1539 1098 1670 1132
rect 1704 1098 1760 1132
rect 1794 1098 1850 1132
rect 1884 1098 1940 1132
rect 1974 1098 2030 1132
rect 2064 1098 2120 1132
rect 2154 1098 2210 1132
rect 2244 1098 2300 1132
rect 2334 1098 2390 1132
rect 2424 1098 2501 1132
rect 1539 1079 2501 1098
rect 1539 1075 1611 1079
rect 1539 1041 1558 1075
rect 1592 1041 1611 1075
rect 1539 985 1611 1041
rect 2429 1056 2501 1079
rect 2429 1022 2448 1056
rect 2482 1022 2501 1056
rect 1539 951 1558 985
rect 1592 951 1611 985
rect 1539 895 1611 951
rect 1539 861 1558 895
rect 1592 861 1611 895
rect 1539 805 1611 861
rect 1539 771 1558 805
rect 1592 771 1611 805
rect 1539 715 1611 771
rect 1539 681 1558 715
rect 1592 681 1611 715
rect 1539 625 1611 681
rect 1539 591 1558 625
rect 1592 591 1611 625
rect 1539 535 1611 591
rect 1539 501 1558 535
rect 1592 501 1611 535
rect 1539 445 1611 501
rect 1539 411 1558 445
rect 1592 411 1611 445
rect 1539 355 1611 411
rect 1539 321 1558 355
rect 1592 321 1611 355
rect 2429 966 2501 1022
rect 2429 932 2448 966
rect 2482 932 2501 966
rect 2429 876 2501 932
rect 2429 842 2448 876
rect 2482 842 2501 876
rect 2429 786 2501 842
rect 2429 752 2448 786
rect 2482 752 2501 786
rect 2429 696 2501 752
rect 2429 662 2448 696
rect 2482 662 2501 696
rect 2429 606 2501 662
rect 2429 572 2448 606
rect 2482 572 2501 606
rect 2429 516 2501 572
rect 2429 482 2448 516
rect 2482 482 2501 516
rect 2429 426 2501 482
rect 2429 392 2448 426
rect 2482 392 2501 426
rect 2429 336 2501 392
rect 1539 261 1611 321
rect 2429 302 2448 336
rect 2482 302 2501 336
rect 2429 261 2501 302
rect 1539 242 2501 261
rect 1539 208 1636 242
rect 1670 208 1726 242
rect 1760 208 1816 242
rect 1850 208 1906 242
rect 1940 208 1996 242
rect 2030 208 2086 242
rect 2120 208 2176 242
rect 2210 208 2266 242
rect 2300 208 2356 242
rect 2390 208 2501 242
rect 1539 189 2501 208
rect 2899 1132 3861 1151
rect 2899 1098 3030 1132
rect 3064 1098 3120 1132
rect 3154 1098 3210 1132
rect 3244 1098 3300 1132
rect 3334 1098 3390 1132
rect 3424 1098 3480 1132
rect 3514 1098 3570 1132
rect 3604 1098 3660 1132
rect 3694 1098 3750 1132
rect 3784 1098 3861 1132
rect 2899 1079 3861 1098
rect 2899 1075 2971 1079
rect 2899 1041 2918 1075
rect 2952 1041 2971 1075
rect 2899 985 2971 1041
rect 3789 1056 3861 1079
rect 3789 1022 3808 1056
rect 3842 1022 3861 1056
rect 2899 951 2918 985
rect 2952 951 2971 985
rect 2899 895 2971 951
rect 2899 861 2918 895
rect 2952 861 2971 895
rect 2899 805 2971 861
rect 2899 771 2918 805
rect 2952 771 2971 805
rect 2899 715 2971 771
rect 2899 681 2918 715
rect 2952 681 2971 715
rect 2899 625 2971 681
rect 2899 591 2918 625
rect 2952 591 2971 625
rect 2899 535 2971 591
rect 2899 501 2918 535
rect 2952 501 2971 535
rect 2899 445 2971 501
rect 2899 411 2918 445
rect 2952 411 2971 445
rect 2899 355 2971 411
rect 2899 321 2918 355
rect 2952 321 2971 355
rect 3789 966 3861 1022
rect 3789 932 3808 966
rect 3842 932 3861 966
rect 3789 876 3861 932
rect 3789 842 3808 876
rect 3842 842 3861 876
rect 3789 786 3861 842
rect 3789 752 3808 786
rect 3842 752 3861 786
rect 3789 696 3861 752
rect 3789 662 3808 696
rect 3842 662 3861 696
rect 3789 606 3861 662
rect 3789 572 3808 606
rect 3842 572 3861 606
rect 3789 516 3861 572
rect 3789 482 3808 516
rect 3842 482 3861 516
rect 3789 426 3861 482
rect 3789 392 3808 426
rect 3842 392 3861 426
rect 3789 336 3861 392
rect 2899 261 2971 321
rect 3789 302 3808 336
rect 3842 302 3861 336
rect 3789 261 3861 302
rect 2899 242 3861 261
rect 2899 208 2996 242
rect 3030 208 3086 242
rect 3120 208 3176 242
rect 3210 208 3266 242
rect 3300 208 3356 242
rect 3390 208 3446 242
rect 3480 208 3536 242
rect 3570 208 3626 242
rect 3660 208 3716 242
rect 3750 208 3861 242
rect 2899 189 3861 208
rect 4259 1132 5221 1151
rect 4259 1098 4390 1132
rect 4424 1098 4480 1132
rect 4514 1098 4570 1132
rect 4604 1098 4660 1132
rect 4694 1098 4750 1132
rect 4784 1098 4840 1132
rect 4874 1098 4930 1132
rect 4964 1098 5020 1132
rect 5054 1098 5110 1132
rect 5144 1098 5221 1132
rect 4259 1079 5221 1098
rect 4259 1075 4331 1079
rect 4259 1041 4278 1075
rect 4312 1041 4331 1075
rect 4259 985 4331 1041
rect 5149 1056 5221 1079
rect 5149 1022 5168 1056
rect 5202 1022 5221 1056
rect 4259 951 4278 985
rect 4312 951 4331 985
rect 4259 895 4331 951
rect 4259 861 4278 895
rect 4312 861 4331 895
rect 4259 805 4331 861
rect 4259 771 4278 805
rect 4312 771 4331 805
rect 4259 715 4331 771
rect 4259 681 4278 715
rect 4312 681 4331 715
rect 4259 625 4331 681
rect 4259 591 4278 625
rect 4312 591 4331 625
rect 4259 535 4331 591
rect 4259 501 4278 535
rect 4312 501 4331 535
rect 4259 445 4331 501
rect 4259 411 4278 445
rect 4312 411 4331 445
rect 4259 355 4331 411
rect 4259 321 4278 355
rect 4312 321 4331 355
rect 5149 966 5221 1022
rect 5149 932 5168 966
rect 5202 932 5221 966
rect 5149 876 5221 932
rect 5149 842 5168 876
rect 5202 842 5221 876
rect 5149 786 5221 842
rect 5149 752 5168 786
rect 5202 752 5221 786
rect 5149 696 5221 752
rect 5149 662 5168 696
rect 5202 662 5221 696
rect 5149 606 5221 662
rect 5149 572 5168 606
rect 5202 572 5221 606
rect 5149 516 5221 572
rect 5149 482 5168 516
rect 5202 482 5221 516
rect 5149 426 5221 482
rect 5149 392 5168 426
rect 5202 392 5221 426
rect 5149 336 5221 392
rect 4259 261 4331 321
rect 5149 302 5168 336
rect 5202 302 5221 336
rect 5149 261 5221 302
rect 4259 242 5221 261
rect 4259 208 4356 242
rect 4390 208 4446 242
rect 4480 208 4536 242
rect 4570 208 4626 242
rect 4660 208 4716 242
rect 4750 208 4806 242
rect 4840 208 4896 242
rect 4930 208 4986 242
rect 5020 208 5076 242
rect 5110 208 5221 242
rect 4259 189 5221 208
rect 5619 1132 6581 1151
rect 5619 1098 5750 1132
rect 5784 1098 5840 1132
rect 5874 1098 5930 1132
rect 5964 1098 6020 1132
rect 6054 1098 6110 1132
rect 6144 1098 6200 1132
rect 6234 1098 6290 1132
rect 6324 1098 6380 1132
rect 6414 1098 6470 1132
rect 6504 1098 6581 1132
rect 5619 1079 6581 1098
rect 5619 1075 5691 1079
rect 5619 1041 5638 1075
rect 5672 1041 5691 1075
rect 5619 985 5691 1041
rect 6509 1056 6581 1079
rect 6509 1022 6528 1056
rect 6562 1022 6581 1056
rect 5619 951 5638 985
rect 5672 951 5691 985
rect 5619 895 5691 951
rect 5619 861 5638 895
rect 5672 861 5691 895
rect 5619 805 5691 861
rect 5619 771 5638 805
rect 5672 771 5691 805
rect 5619 715 5691 771
rect 5619 681 5638 715
rect 5672 681 5691 715
rect 5619 625 5691 681
rect 5619 591 5638 625
rect 5672 591 5691 625
rect 5619 535 5691 591
rect 5619 501 5638 535
rect 5672 501 5691 535
rect 5619 445 5691 501
rect 5619 411 5638 445
rect 5672 411 5691 445
rect 5619 355 5691 411
rect 5619 321 5638 355
rect 5672 321 5691 355
rect 6509 966 6581 1022
rect 6509 932 6528 966
rect 6562 932 6581 966
rect 6509 876 6581 932
rect 6509 842 6528 876
rect 6562 842 6581 876
rect 6509 786 6581 842
rect 6509 752 6528 786
rect 6562 752 6581 786
rect 6509 696 6581 752
rect 6509 662 6528 696
rect 6562 662 6581 696
rect 6509 606 6581 662
rect 6509 572 6528 606
rect 6562 572 6581 606
rect 6509 516 6581 572
rect 6509 482 6528 516
rect 6562 482 6581 516
rect 6509 426 6581 482
rect 6509 392 6528 426
rect 6562 392 6581 426
rect 6509 336 6581 392
rect 5619 261 5691 321
rect 6509 302 6528 336
rect 6562 302 6581 336
rect 6509 261 6581 302
rect 5619 242 6581 261
rect 5619 208 5716 242
rect 5750 208 5806 242
rect 5840 208 5896 242
rect 5930 208 5986 242
rect 6020 208 6076 242
rect 6110 208 6166 242
rect 6200 208 6256 242
rect 6290 208 6346 242
rect 6380 208 6436 242
rect 6470 208 6581 242
rect 5619 189 6581 208
rect 6979 1132 7941 1151
rect 6979 1098 7110 1132
rect 7144 1098 7200 1132
rect 7234 1098 7290 1132
rect 7324 1098 7380 1132
rect 7414 1098 7470 1132
rect 7504 1098 7560 1132
rect 7594 1098 7650 1132
rect 7684 1098 7740 1132
rect 7774 1098 7830 1132
rect 7864 1098 7941 1132
rect 6979 1079 7941 1098
rect 6979 1075 7051 1079
rect 6979 1041 6998 1075
rect 7032 1041 7051 1075
rect 6979 985 7051 1041
rect 7869 1056 7941 1079
rect 7869 1022 7888 1056
rect 7922 1022 7941 1056
rect 6979 951 6998 985
rect 7032 951 7051 985
rect 6979 895 7051 951
rect 6979 861 6998 895
rect 7032 861 7051 895
rect 6979 805 7051 861
rect 6979 771 6998 805
rect 7032 771 7051 805
rect 6979 715 7051 771
rect 6979 681 6998 715
rect 7032 681 7051 715
rect 6979 625 7051 681
rect 6979 591 6998 625
rect 7032 591 7051 625
rect 6979 535 7051 591
rect 6979 501 6998 535
rect 7032 501 7051 535
rect 6979 445 7051 501
rect 6979 411 6998 445
rect 7032 411 7051 445
rect 6979 355 7051 411
rect 6979 321 6998 355
rect 7032 321 7051 355
rect 7869 966 7941 1022
rect 7869 932 7888 966
rect 7922 932 7941 966
rect 7869 876 7941 932
rect 7869 842 7888 876
rect 7922 842 7941 876
rect 7869 786 7941 842
rect 7869 752 7888 786
rect 7922 752 7941 786
rect 7869 696 7941 752
rect 7869 662 7888 696
rect 7922 662 7941 696
rect 7869 606 7941 662
rect 7869 572 7888 606
rect 7922 572 7941 606
rect 7869 516 7941 572
rect 7869 482 7888 516
rect 7922 482 7941 516
rect 7869 426 7941 482
rect 7869 392 7888 426
rect 7922 392 7941 426
rect 7869 336 7941 392
rect 6979 261 7051 321
rect 7869 302 7888 336
rect 7922 302 7941 336
rect 7869 261 7941 302
rect 6979 242 7941 261
rect 6979 208 7076 242
rect 7110 208 7166 242
rect 7200 208 7256 242
rect 7290 208 7346 242
rect 7380 208 7436 242
rect 7470 208 7526 242
rect 7560 208 7616 242
rect 7650 208 7706 242
rect 7740 208 7796 242
rect 7830 208 7941 242
rect 6979 189 7941 208
rect 8339 1132 9301 1151
rect 8339 1098 8470 1132
rect 8504 1098 8560 1132
rect 8594 1098 8650 1132
rect 8684 1098 8740 1132
rect 8774 1098 8830 1132
rect 8864 1098 8920 1132
rect 8954 1098 9010 1132
rect 9044 1098 9100 1132
rect 9134 1098 9190 1132
rect 9224 1098 9301 1132
rect 8339 1079 9301 1098
rect 8339 1075 8411 1079
rect 8339 1041 8358 1075
rect 8392 1041 8411 1075
rect 8339 985 8411 1041
rect 9229 1056 9301 1079
rect 9229 1022 9248 1056
rect 9282 1022 9301 1056
rect 8339 951 8358 985
rect 8392 951 8411 985
rect 8339 895 8411 951
rect 8339 861 8358 895
rect 8392 861 8411 895
rect 8339 805 8411 861
rect 8339 771 8358 805
rect 8392 771 8411 805
rect 8339 715 8411 771
rect 8339 681 8358 715
rect 8392 681 8411 715
rect 8339 625 8411 681
rect 8339 591 8358 625
rect 8392 591 8411 625
rect 8339 535 8411 591
rect 8339 501 8358 535
rect 8392 501 8411 535
rect 8339 445 8411 501
rect 8339 411 8358 445
rect 8392 411 8411 445
rect 8339 355 8411 411
rect 8339 321 8358 355
rect 8392 321 8411 355
rect 9229 966 9301 1022
rect 9229 932 9248 966
rect 9282 932 9301 966
rect 9229 876 9301 932
rect 9229 842 9248 876
rect 9282 842 9301 876
rect 9229 786 9301 842
rect 9229 752 9248 786
rect 9282 752 9301 786
rect 9229 696 9301 752
rect 9229 662 9248 696
rect 9282 662 9301 696
rect 9229 606 9301 662
rect 9229 572 9248 606
rect 9282 572 9301 606
rect 9229 516 9301 572
rect 9229 482 9248 516
rect 9282 482 9301 516
rect 9229 426 9301 482
rect 9229 392 9248 426
rect 9282 392 9301 426
rect 9229 336 9301 392
rect 8339 261 8411 321
rect 9229 302 9248 336
rect 9282 302 9301 336
rect 9229 261 9301 302
rect 8339 242 9301 261
rect 8339 208 8436 242
rect 8470 208 8526 242
rect 8560 208 8616 242
rect 8650 208 8706 242
rect 8740 208 8796 242
rect 8830 208 8886 242
rect 8920 208 8976 242
rect 9010 208 9066 242
rect 9100 208 9156 242
rect 9190 208 9301 242
rect 8339 189 9301 208
<< psubdiffcont >>
rect 4350 5090 4390 5130
rect 4350 4990 4390 5030
rect 4350 4890 4390 4930
rect 4350 4790 4390 4830
rect 4350 4690 4390 4730
rect 4350 4590 4390 4630
rect 4350 4490 4390 4530
rect 4350 4390 4390 4430
rect 8510 5090 8550 5130
rect 8510 4990 8550 5030
rect 8510 4890 8550 4930
rect 8510 4790 8550 4830
rect 8510 4690 8550 4730
rect 8510 4590 8550 4630
rect 8510 4490 8550 4530
rect 8510 4390 8550 4430
rect 10270 4290 10310 4330
rect 10270 4190 10310 4230
rect 10270 4090 10310 4130
rect 10270 3990 10310 4030
rect 10790 4290 10830 4330
rect 10790 4190 10830 4230
rect 10790 4090 10830 4130
rect 10790 3990 10830 4030
rect 4390 3780 4430 3820
rect 4390 3680 4430 3720
rect 4390 3580 4430 3620
rect 4390 3480 4430 3520
rect 5750 3780 5790 3820
rect 5750 3680 5790 3720
rect 5750 3580 5790 3620
rect 5750 3480 5790 3520
rect 7110 3780 7150 3820
rect 7110 3680 7150 3720
rect 7110 3580 7150 3620
rect 7110 3480 7150 3520
rect 8470 3780 8510 3820
rect 8470 3680 8510 3720
rect 8470 3580 8510 3620
rect 8470 3480 8510 3520
rect 11390 3590 11430 3630
rect 11390 3490 11430 3530
rect 5070 2970 5110 3010
rect 5070 2870 5110 2910
rect 6430 2970 6470 3010
rect 6430 2870 6470 2910
rect 7790 2970 7830 3010
rect 7790 2870 7830 2910
rect 4590 2420 4630 2460
rect 4590 2320 4630 2360
rect 4590 2220 4630 2260
rect 4590 2120 4630 2160
rect 4590 2020 4630 2060
rect 4590 1920 4630 1960
rect 4590 1820 4630 1860
rect 4590 1720 4630 1760
rect 8270 2420 8310 2460
rect 8270 2320 8310 2360
rect 8270 2220 8310 2260
rect 8270 2120 8310 2160
rect 8270 2020 8310 2060
rect 8270 1920 8310 1960
rect 8270 1820 8310 1860
rect 8270 1720 8310 1760
rect 1410 1222 1444 1256
rect 1506 1245 1540 1279
rect 1596 1245 1630 1279
rect 1686 1245 1720 1279
rect 1776 1245 1810 1279
rect 1866 1245 1900 1279
rect 1956 1245 1990 1279
rect 2046 1245 2080 1279
rect 2136 1245 2170 1279
rect 2226 1245 2260 1279
rect 2316 1245 2350 1279
rect 2406 1245 2440 1279
rect 2496 1245 2530 1279
rect 2597 1222 2631 1256
rect 1410 1132 1444 1166
rect 1410 1042 1444 1076
rect 1410 952 1444 986
rect 1410 862 1444 896
rect 1410 772 1444 806
rect 1410 682 1444 716
rect 1410 592 1444 626
rect 1410 502 1444 536
rect 1410 412 1444 446
rect 1410 322 1444 356
rect 1410 232 1444 266
rect 2597 1132 2631 1166
rect 2597 1042 2631 1076
rect 2597 952 2631 986
rect 2597 862 2631 896
rect 2597 772 2631 806
rect 2597 682 2631 716
rect 2597 592 2631 626
rect 2597 502 2631 536
rect 2597 412 2631 446
rect 2597 322 2631 356
rect 2597 232 2631 266
rect 1410 142 1444 176
rect 2597 142 2631 176
rect 1506 58 1540 92
rect 1596 58 1630 92
rect 1686 58 1720 92
rect 1776 58 1810 92
rect 1866 58 1900 92
rect 1956 58 1990 92
rect 2046 58 2080 92
rect 2136 58 2170 92
rect 2226 58 2260 92
rect 2316 58 2350 92
rect 2406 58 2440 92
rect 2496 58 2530 92
rect 2770 1222 2804 1256
rect 2866 1245 2900 1279
rect 2956 1245 2990 1279
rect 3046 1245 3080 1279
rect 3136 1245 3170 1279
rect 3226 1245 3260 1279
rect 3316 1245 3350 1279
rect 3406 1245 3440 1279
rect 3496 1245 3530 1279
rect 3586 1245 3620 1279
rect 3676 1245 3710 1279
rect 3766 1245 3800 1279
rect 3856 1245 3890 1279
rect 3957 1222 3991 1256
rect 2770 1132 2804 1166
rect 2770 1042 2804 1076
rect 2770 952 2804 986
rect 2770 862 2804 896
rect 2770 772 2804 806
rect 2770 682 2804 716
rect 2770 592 2804 626
rect 2770 502 2804 536
rect 2770 412 2804 446
rect 2770 322 2804 356
rect 2770 232 2804 266
rect 3957 1132 3991 1166
rect 3957 1042 3991 1076
rect 3957 952 3991 986
rect 3957 862 3991 896
rect 3957 772 3991 806
rect 3957 682 3991 716
rect 3957 592 3991 626
rect 3957 502 3991 536
rect 3957 412 3991 446
rect 3957 322 3991 356
rect 3957 232 3991 266
rect 2770 142 2804 176
rect 3957 142 3991 176
rect 2866 58 2900 92
rect 2956 58 2990 92
rect 3046 58 3080 92
rect 3136 58 3170 92
rect 3226 58 3260 92
rect 3316 58 3350 92
rect 3406 58 3440 92
rect 3496 58 3530 92
rect 3586 58 3620 92
rect 3676 58 3710 92
rect 3766 58 3800 92
rect 3856 58 3890 92
rect 4130 1222 4164 1256
rect 4226 1245 4260 1279
rect 4316 1245 4350 1279
rect 4406 1245 4440 1279
rect 4496 1245 4530 1279
rect 4586 1245 4620 1279
rect 4676 1245 4710 1279
rect 4766 1245 4800 1279
rect 4856 1245 4890 1279
rect 4946 1245 4980 1279
rect 5036 1245 5070 1279
rect 5126 1245 5160 1279
rect 5216 1245 5250 1279
rect 5317 1222 5351 1256
rect 4130 1132 4164 1166
rect 4130 1042 4164 1076
rect 4130 952 4164 986
rect 4130 862 4164 896
rect 4130 772 4164 806
rect 4130 682 4164 716
rect 4130 592 4164 626
rect 4130 502 4164 536
rect 4130 412 4164 446
rect 4130 322 4164 356
rect 4130 232 4164 266
rect 5317 1132 5351 1166
rect 5317 1042 5351 1076
rect 5317 952 5351 986
rect 5317 862 5351 896
rect 5317 772 5351 806
rect 5317 682 5351 716
rect 5317 592 5351 626
rect 5317 502 5351 536
rect 5317 412 5351 446
rect 5317 322 5351 356
rect 5317 232 5351 266
rect 4130 142 4164 176
rect 5317 142 5351 176
rect 4226 58 4260 92
rect 4316 58 4350 92
rect 4406 58 4440 92
rect 4496 58 4530 92
rect 4586 58 4620 92
rect 4676 58 4710 92
rect 4766 58 4800 92
rect 4856 58 4890 92
rect 4946 58 4980 92
rect 5036 58 5070 92
rect 5126 58 5160 92
rect 5216 58 5250 92
rect 5490 1222 5524 1256
rect 5586 1245 5620 1279
rect 5676 1245 5710 1279
rect 5766 1245 5800 1279
rect 5856 1245 5890 1279
rect 5946 1245 5980 1279
rect 6036 1245 6070 1279
rect 6126 1245 6160 1279
rect 6216 1245 6250 1279
rect 6306 1245 6340 1279
rect 6396 1245 6430 1279
rect 6486 1245 6520 1279
rect 6576 1245 6610 1279
rect 6677 1222 6711 1256
rect 5490 1132 5524 1166
rect 5490 1042 5524 1076
rect 5490 952 5524 986
rect 5490 862 5524 896
rect 5490 772 5524 806
rect 5490 682 5524 716
rect 5490 592 5524 626
rect 5490 502 5524 536
rect 5490 412 5524 446
rect 5490 322 5524 356
rect 5490 232 5524 266
rect 6677 1132 6711 1166
rect 6677 1042 6711 1076
rect 6677 952 6711 986
rect 6677 862 6711 896
rect 6677 772 6711 806
rect 6677 682 6711 716
rect 6677 592 6711 626
rect 6677 502 6711 536
rect 6677 412 6711 446
rect 6677 322 6711 356
rect 6677 232 6711 266
rect 5490 142 5524 176
rect 6677 142 6711 176
rect 5586 58 5620 92
rect 5676 58 5710 92
rect 5766 58 5800 92
rect 5856 58 5890 92
rect 5946 58 5980 92
rect 6036 58 6070 92
rect 6126 58 6160 92
rect 6216 58 6250 92
rect 6306 58 6340 92
rect 6396 58 6430 92
rect 6486 58 6520 92
rect 6576 58 6610 92
rect 6850 1222 6884 1256
rect 6946 1245 6980 1279
rect 7036 1245 7070 1279
rect 7126 1245 7160 1279
rect 7216 1245 7250 1279
rect 7306 1245 7340 1279
rect 7396 1245 7430 1279
rect 7486 1245 7520 1279
rect 7576 1245 7610 1279
rect 7666 1245 7700 1279
rect 7756 1245 7790 1279
rect 7846 1245 7880 1279
rect 7936 1245 7970 1279
rect 8037 1222 8071 1256
rect 6850 1132 6884 1166
rect 6850 1042 6884 1076
rect 6850 952 6884 986
rect 6850 862 6884 896
rect 6850 772 6884 806
rect 6850 682 6884 716
rect 6850 592 6884 626
rect 6850 502 6884 536
rect 6850 412 6884 446
rect 6850 322 6884 356
rect 6850 232 6884 266
rect 8037 1132 8071 1166
rect 8037 1042 8071 1076
rect 8037 952 8071 986
rect 8037 862 8071 896
rect 8037 772 8071 806
rect 8037 682 8071 716
rect 8037 592 8071 626
rect 8037 502 8071 536
rect 8037 412 8071 446
rect 8037 322 8071 356
rect 8037 232 8071 266
rect 6850 142 6884 176
rect 8037 142 8071 176
rect 6946 58 6980 92
rect 7036 58 7070 92
rect 7126 58 7160 92
rect 7216 58 7250 92
rect 7306 58 7340 92
rect 7396 58 7430 92
rect 7486 58 7520 92
rect 7576 58 7610 92
rect 7666 58 7700 92
rect 7756 58 7790 92
rect 7846 58 7880 92
rect 7936 58 7970 92
rect 8210 1222 8244 1256
rect 8306 1245 8340 1279
rect 8396 1245 8430 1279
rect 8486 1245 8520 1279
rect 8576 1245 8610 1279
rect 8666 1245 8700 1279
rect 8756 1245 8790 1279
rect 8846 1245 8880 1279
rect 8936 1245 8970 1279
rect 9026 1245 9060 1279
rect 9116 1245 9150 1279
rect 9206 1245 9240 1279
rect 9296 1245 9330 1279
rect 9397 1222 9431 1256
rect 8210 1132 8244 1166
rect 8210 1042 8244 1076
rect 8210 952 8244 986
rect 8210 862 8244 896
rect 8210 772 8244 806
rect 8210 682 8244 716
rect 8210 592 8244 626
rect 8210 502 8244 536
rect 8210 412 8244 446
rect 8210 322 8244 356
rect 8210 232 8244 266
rect 9397 1132 9431 1166
rect 9397 1042 9431 1076
rect 9397 952 9431 986
rect 9397 862 9431 896
rect 9397 772 9431 806
rect 9397 682 9431 716
rect 9397 592 9431 626
rect 9397 502 9431 536
rect 9397 412 9431 446
rect 9397 322 9431 356
rect 9397 232 9431 266
rect 8210 142 8244 176
rect 9397 142 9431 176
rect 8306 58 8340 92
rect 8396 58 8430 92
rect 8486 58 8520 92
rect 8576 58 8610 92
rect 8666 58 8700 92
rect 8756 58 8790 92
rect 8846 58 8880 92
rect 8936 58 8970 92
rect 9026 58 9060 92
rect 9116 58 9150 92
rect 9206 58 9240 92
rect 9296 58 9330 92
<< nsubdiffcont >>
rect 1670 1098 1704 1132
rect 1760 1098 1794 1132
rect 1850 1098 1884 1132
rect 1940 1098 1974 1132
rect 2030 1098 2064 1132
rect 2120 1098 2154 1132
rect 2210 1098 2244 1132
rect 2300 1098 2334 1132
rect 2390 1098 2424 1132
rect 1558 1041 1592 1075
rect 2448 1022 2482 1056
rect 1558 951 1592 985
rect 1558 861 1592 895
rect 1558 771 1592 805
rect 1558 681 1592 715
rect 1558 591 1592 625
rect 1558 501 1592 535
rect 1558 411 1592 445
rect 1558 321 1592 355
rect 2448 932 2482 966
rect 2448 842 2482 876
rect 2448 752 2482 786
rect 2448 662 2482 696
rect 2448 572 2482 606
rect 2448 482 2482 516
rect 2448 392 2482 426
rect 2448 302 2482 336
rect 1636 208 1670 242
rect 1726 208 1760 242
rect 1816 208 1850 242
rect 1906 208 1940 242
rect 1996 208 2030 242
rect 2086 208 2120 242
rect 2176 208 2210 242
rect 2266 208 2300 242
rect 2356 208 2390 242
rect 3030 1098 3064 1132
rect 3120 1098 3154 1132
rect 3210 1098 3244 1132
rect 3300 1098 3334 1132
rect 3390 1098 3424 1132
rect 3480 1098 3514 1132
rect 3570 1098 3604 1132
rect 3660 1098 3694 1132
rect 3750 1098 3784 1132
rect 2918 1041 2952 1075
rect 3808 1022 3842 1056
rect 2918 951 2952 985
rect 2918 861 2952 895
rect 2918 771 2952 805
rect 2918 681 2952 715
rect 2918 591 2952 625
rect 2918 501 2952 535
rect 2918 411 2952 445
rect 2918 321 2952 355
rect 3808 932 3842 966
rect 3808 842 3842 876
rect 3808 752 3842 786
rect 3808 662 3842 696
rect 3808 572 3842 606
rect 3808 482 3842 516
rect 3808 392 3842 426
rect 3808 302 3842 336
rect 2996 208 3030 242
rect 3086 208 3120 242
rect 3176 208 3210 242
rect 3266 208 3300 242
rect 3356 208 3390 242
rect 3446 208 3480 242
rect 3536 208 3570 242
rect 3626 208 3660 242
rect 3716 208 3750 242
rect 4390 1098 4424 1132
rect 4480 1098 4514 1132
rect 4570 1098 4604 1132
rect 4660 1098 4694 1132
rect 4750 1098 4784 1132
rect 4840 1098 4874 1132
rect 4930 1098 4964 1132
rect 5020 1098 5054 1132
rect 5110 1098 5144 1132
rect 4278 1041 4312 1075
rect 5168 1022 5202 1056
rect 4278 951 4312 985
rect 4278 861 4312 895
rect 4278 771 4312 805
rect 4278 681 4312 715
rect 4278 591 4312 625
rect 4278 501 4312 535
rect 4278 411 4312 445
rect 4278 321 4312 355
rect 5168 932 5202 966
rect 5168 842 5202 876
rect 5168 752 5202 786
rect 5168 662 5202 696
rect 5168 572 5202 606
rect 5168 482 5202 516
rect 5168 392 5202 426
rect 5168 302 5202 336
rect 4356 208 4390 242
rect 4446 208 4480 242
rect 4536 208 4570 242
rect 4626 208 4660 242
rect 4716 208 4750 242
rect 4806 208 4840 242
rect 4896 208 4930 242
rect 4986 208 5020 242
rect 5076 208 5110 242
rect 5750 1098 5784 1132
rect 5840 1098 5874 1132
rect 5930 1098 5964 1132
rect 6020 1098 6054 1132
rect 6110 1098 6144 1132
rect 6200 1098 6234 1132
rect 6290 1098 6324 1132
rect 6380 1098 6414 1132
rect 6470 1098 6504 1132
rect 5638 1041 5672 1075
rect 6528 1022 6562 1056
rect 5638 951 5672 985
rect 5638 861 5672 895
rect 5638 771 5672 805
rect 5638 681 5672 715
rect 5638 591 5672 625
rect 5638 501 5672 535
rect 5638 411 5672 445
rect 5638 321 5672 355
rect 6528 932 6562 966
rect 6528 842 6562 876
rect 6528 752 6562 786
rect 6528 662 6562 696
rect 6528 572 6562 606
rect 6528 482 6562 516
rect 6528 392 6562 426
rect 6528 302 6562 336
rect 5716 208 5750 242
rect 5806 208 5840 242
rect 5896 208 5930 242
rect 5986 208 6020 242
rect 6076 208 6110 242
rect 6166 208 6200 242
rect 6256 208 6290 242
rect 6346 208 6380 242
rect 6436 208 6470 242
rect 7110 1098 7144 1132
rect 7200 1098 7234 1132
rect 7290 1098 7324 1132
rect 7380 1098 7414 1132
rect 7470 1098 7504 1132
rect 7560 1098 7594 1132
rect 7650 1098 7684 1132
rect 7740 1098 7774 1132
rect 7830 1098 7864 1132
rect 6998 1041 7032 1075
rect 7888 1022 7922 1056
rect 6998 951 7032 985
rect 6998 861 7032 895
rect 6998 771 7032 805
rect 6998 681 7032 715
rect 6998 591 7032 625
rect 6998 501 7032 535
rect 6998 411 7032 445
rect 6998 321 7032 355
rect 7888 932 7922 966
rect 7888 842 7922 876
rect 7888 752 7922 786
rect 7888 662 7922 696
rect 7888 572 7922 606
rect 7888 482 7922 516
rect 7888 392 7922 426
rect 7888 302 7922 336
rect 7076 208 7110 242
rect 7166 208 7200 242
rect 7256 208 7290 242
rect 7346 208 7380 242
rect 7436 208 7470 242
rect 7526 208 7560 242
rect 7616 208 7650 242
rect 7706 208 7740 242
rect 7796 208 7830 242
rect 8470 1098 8504 1132
rect 8560 1098 8594 1132
rect 8650 1098 8684 1132
rect 8740 1098 8774 1132
rect 8830 1098 8864 1132
rect 8920 1098 8954 1132
rect 9010 1098 9044 1132
rect 9100 1098 9134 1132
rect 9190 1098 9224 1132
rect 8358 1041 8392 1075
rect 9248 1022 9282 1056
rect 8358 951 8392 985
rect 8358 861 8392 895
rect 8358 771 8392 805
rect 8358 681 8392 715
rect 8358 591 8392 625
rect 8358 501 8392 535
rect 8358 411 8392 445
rect 8358 321 8392 355
rect 9248 932 9282 966
rect 9248 842 9282 876
rect 9248 752 9282 786
rect 9248 662 9282 696
rect 9248 572 9282 606
rect 9248 482 9282 516
rect 9248 392 9282 426
rect 9248 302 9282 336
rect 8436 208 8470 242
rect 8526 208 8560 242
rect 8616 208 8650 242
rect 8706 208 8740 242
rect 8796 208 8830 242
rect 8886 208 8920 242
rect 8976 208 9010 242
rect 9066 208 9100 242
rect 9156 208 9190 242
<< poly >>
rect 4490 5160 4610 5190
rect 4690 5160 4810 5190
rect 4890 5160 5010 5190
rect 5090 5160 5210 5190
rect 5290 5160 5410 5190
rect 5490 5160 5610 5190
rect 5690 5160 5810 5190
rect 5890 5160 6010 5190
rect 6090 5160 6210 5190
rect 6290 5160 6410 5190
rect 6490 5160 6610 5190
rect 6690 5160 6810 5190
rect 6890 5160 7010 5190
rect 7090 5160 7210 5190
rect 7290 5160 7410 5190
rect 7490 5160 7610 5190
rect 7690 5160 7810 5190
rect 7890 5160 8010 5190
rect 8090 5160 8210 5190
rect 8290 5160 8410 5190
rect 10410 4530 10490 4550
rect 10410 4490 10430 4530
rect 10470 4490 10490 4530
rect 10410 4470 10490 4490
rect 10410 4360 10440 4470
rect 10610 4450 10690 4470
rect 10610 4410 10630 4450
rect 10670 4410 10690 4450
rect 10610 4390 10690 4410
rect 10660 4360 10690 4390
rect 4490 4330 4610 4360
rect 4690 4340 4810 4360
rect 4890 4340 5010 4360
rect 5090 4340 5210 4360
rect 5290 4340 5410 4360
rect 5490 4340 5610 4360
rect 5690 4340 5810 4360
rect 5890 4340 6010 4360
rect 6090 4340 6210 4360
rect 6290 4340 6410 4360
rect 6490 4340 6610 4360
rect 6690 4340 6810 4360
rect 6890 4340 7010 4360
rect 7090 4340 7210 4360
rect 7290 4340 7410 4360
rect 7490 4340 7610 4360
rect 7690 4340 7810 4360
rect 7890 4340 8010 4360
rect 8090 4340 8210 4360
rect 4690 4310 8210 4340
rect 8290 4330 8410 4360
rect 6210 4270 6230 4310
rect 6270 4270 6290 4310
rect 6210 4250 6290 4270
rect 6610 4270 6630 4310
rect 6670 4270 6690 4310
rect 6610 4250 6690 4270
rect 10410 3930 10440 3960
rect 10660 3930 10690 3960
rect 4530 3850 4650 3880
rect 4730 3850 4850 3880
rect 4930 3850 5050 3880
rect 5130 3850 5250 3880
rect 5330 3850 5450 3880
rect 5530 3850 5650 3880
rect 5890 3850 6010 3880
rect 6090 3850 6210 3880
rect 6290 3850 6410 3880
rect 6490 3850 6610 3880
rect 6690 3850 6810 3880
rect 6890 3850 7010 3880
rect 7250 3850 7370 3880
rect 7450 3850 7570 3880
rect 7650 3850 7770 3880
rect 7850 3850 7970 3880
rect 8050 3850 8170 3880
rect 8250 3850 8370 3880
rect 9290 3750 9370 3770
rect 9290 3710 9310 3750
rect 9350 3710 9370 3750
rect 9290 3690 9370 3710
rect 9450 3750 9530 3770
rect 9450 3710 9470 3750
rect 9510 3710 9530 3750
rect 9450 3690 9530 3710
rect 9610 3750 9690 3770
rect 9610 3710 9630 3750
rect 9670 3710 9690 3750
rect 9610 3690 9690 3710
rect 9770 3750 9850 3770
rect 9770 3710 9790 3750
rect 9830 3710 9850 3750
rect 9770 3690 9850 3710
rect 9930 3750 10010 3770
rect 9930 3710 9950 3750
rect 9990 3710 10010 3750
rect 9930 3690 10010 3710
rect 10090 3750 10170 3770
rect 10090 3710 10110 3750
rect 10150 3710 10170 3750
rect 10090 3690 10170 3710
rect 10250 3750 10330 3770
rect 10250 3710 10270 3750
rect 10310 3710 10330 3750
rect 10250 3690 10330 3710
rect 10410 3750 10490 3770
rect 10410 3710 10430 3750
rect 10470 3710 10490 3750
rect 10410 3690 10490 3710
rect 10570 3750 10650 3770
rect 10570 3710 10590 3750
rect 10630 3710 10650 3750
rect 10570 3690 10650 3710
rect 10730 3750 10810 3770
rect 10730 3710 10750 3750
rect 10790 3710 10810 3750
rect 10730 3690 10810 3710
rect 10890 3750 10970 3770
rect 10890 3710 10910 3750
rect 10950 3710 10970 3750
rect 10890 3690 10970 3710
rect 11050 3750 11130 3770
rect 11050 3710 11070 3750
rect 11110 3710 11130 3750
rect 11050 3690 11130 3710
rect 11210 3750 11290 3770
rect 11210 3710 11230 3750
rect 11270 3710 11290 3750
rect 11210 3690 11290 3710
rect 9290 3660 11290 3690
rect 4530 3420 4650 3450
rect 4730 3430 4850 3450
rect 4930 3430 5050 3450
rect 5130 3430 5250 3450
rect 5330 3430 5450 3450
rect 4730 3400 5450 3430
rect 5530 3420 5650 3450
rect 5890 3420 6010 3450
rect 6090 3430 6210 3450
rect 6290 3430 6410 3450
rect 6490 3430 6610 3450
rect 6690 3430 6810 3450
rect 6090 3400 6810 3430
rect 6890 3420 7010 3450
rect 7250 3420 7370 3450
rect 7450 3430 7570 3450
rect 7650 3430 7770 3450
rect 7850 3430 7970 3450
rect 8050 3430 8170 3450
rect 7450 3400 8170 3430
rect 8250 3420 8370 3450
rect 9290 3430 11290 3460
rect 5250 3360 5270 3400
rect 5310 3360 5330 3400
rect 5250 3340 5330 3360
rect 6130 3330 6170 3400
rect 6730 3330 6770 3400
rect 7570 3360 7590 3400
rect 7630 3360 7650 3400
rect 7570 3340 7650 3360
rect 6110 3310 6190 3330
rect 6110 3270 6130 3310
rect 6170 3270 6190 3310
rect 6110 3250 6190 3270
rect 6710 3310 6790 3330
rect 6710 3270 6730 3310
rect 6770 3270 6790 3310
rect 6710 3250 6790 3270
rect 6050 3130 6130 3150
rect 6050 3090 6070 3130
rect 6110 3090 6130 3130
rect 5210 3040 5330 3070
rect 5410 3040 5530 3070
rect 5610 3040 5730 3070
rect 5810 3060 6130 3090
rect 6770 3130 6850 3150
rect 6770 3090 6790 3130
rect 6830 3090 6850 3130
rect 5810 3040 5930 3060
rect 6010 3040 6130 3060
rect 6210 3040 6330 3070
rect 6570 3040 6690 3070
rect 6770 3060 7090 3090
rect 6770 3040 6890 3060
rect 6970 3040 7090 3060
rect 7170 3040 7290 3070
rect 7370 3040 7490 3070
rect 7570 3040 7690 3070
rect 5210 2810 5330 2840
rect 5410 2820 5530 2840
rect 5610 2820 5730 2840
rect 5410 2790 5730 2820
rect 5810 2810 5930 2840
rect 6010 2810 6130 2840
rect 6210 2810 6330 2840
rect 6570 2810 6690 2840
rect 6770 2810 6890 2840
rect 6970 2810 7090 2840
rect 7170 2820 7290 2840
rect 7370 2820 7490 2840
rect 7170 2790 7490 2820
rect 7570 2810 7690 2840
rect 5530 2750 5550 2790
rect 5590 2750 5610 2790
rect 5530 2730 5610 2750
rect 7290 2750 7310 2790
rect 7350 2750 7370 2790
rect 7290 2730 7370 2750
rect 5610 2580 6410 2600
rect 5610 2540 5630 2580
rect 5670 2540 5710 2580
rect 5750 2540 5790 2580
rect 5830 2540 5870 2580
rect 5910 2540 5950 2580
rect 5990 2540 6030 2580
rect 6070 2540 6110 2580
rect 6150 2540 6190 2580
rect 6230 2540 6270 2580
rect 6310 2540 6350 2580
rect 6390 2540 6410 2580
rect 4730 2490 5530 2520
rect 5610 2490 6410 2540
rect 6490 2580 7290 2600
rect 6490 2540 6510 2580
rect 6550 2540 6590 2580
rect 6630 2540 6670 2580
rect 6710 2540 6750 2580
rect 6790 2540 6830 2580
rect 6870 2540 6910 2580
rect 6950 2540 6990 2580
rect 7030 2540 7070 2580
rect 7110 2540 7150 2580
rect 7190 2540 7230 2580
rect 7270 2540 7290 2580
rect 6490 2490 7290 2540
rect 7370 2490 8170 2520
rect 4730 1660 5530 1690
rect 5610 1660 6410 1690
rect 6490 1660 7290 1690
rect 7370 1660 8170 1690
<< polycont >>
rect 10430 4490 10470 4530
rect 10630 4410 10670 4450
rect 6230 4270 6270 4310
rect 6630 4270 6670 4310
rect 9310 3710 9350 3750
rect 9470 3710 9510 3750
rect 9630 3710 9670 3750
rect 9790 3710 9830 3750
rect 9950 3710 9990 3750
rect 10110 3710 10150 3750
rect 10270 3710 10310 3750
rect 10430 3710 10470 3750
rect 10590 3710 10630 3750
rect 10750 3710 10790 3750
rect 10910 3710 10950 3750
rect 11070 3710 11110 3750
rect 11230 3710 11270 3750
rect 5270 3360 5310 3400
rect 7590 3360 7630 3400
rect 6130 3270 6170 3310
rect 6730 3270 6770 3310
rect 6070 3090 6110 3130
rect 6790 3090 6830 3130
rect 5550 2750 5590 2790
rect 7310 2750 7350 2790
rect 5630 2540 5670 2580
rect 5710 2540 5750 2580
rect 5790 2540 5830 2580
rect 5870 2540 5910 2580
rect 5950 2540 5990 2580
rect 6030 2540 6070 2580
rect 6110 2540 6150 2580
rect 6190 2540 6230 2580
rect 6270 2540 6310 2580
rect 6350 2540 6390 2580
rect 6510 2540 6550 2580
rect 6590 2540 6630 2580
rect 6670 2540 6710 2580
rect 6750 2540 6790 2580
rect 6830 2540 6870 2580
rect 6910 2540 6950 2580
rect 6990 2540 7030 2580
rect 7070 2540 7110 2580
rect 7150 2540 7190 2580
rect 7230 2540 7270 2580
<< xpolycontact >>
rect 2010 4680 2450 4750
rect 3790 4680 4230 4750
rect 2010 4560 2450 4630
rect 3790 4560 4230 4630
rect 2010 4440 2450 4510
rect 3790 4440 4230 4510
rect 2010 4320 2450 4390
rect 3790 4320 4230 4390
rect 2010 4200 2450 4270
rect 3790 4200 4230 4270
rect 2010 3680 2450 3750
rect 3790 3680 4230 3750
rect 2010 3560 2450 3630
rect 3790 3560 4230 3630
rect 2010 3440 2450 3510
rect 3790 3440 4230 3510
rect 2010 3320 2450 3390
rect 3790 3320 4230 3390
rect 2010 3200 2450 3270
rect 3790 3200 4230 3270
rect 2010 2730 2450 2800
rect 3150 2730 3590 2800
rect 2010 2610 2450 2680
rect 3790 2610 4230 2680
rect 2010 2490 2450 2560
rect 3790 2490 4230 2560
rect 2010 2370 2450 2440
rect 3790 2370 4230 2440
rect 2010 2250 2450 2320
rect 3790 2250 4230 2320
rect 2010 2130 2450 2200
rect 3790 2130 4230 2200
<< xpolyres >>
rect 2450 4680 3790 4750
rect 2450 4560 3790 4630
rect 2450 4440 3790 4510
rect 2450 4320 3790 4390
rect 2450 4200 3790 4270
rect 2450 3680 3790 3750
rect 2450 3560 3790 3630
rect 2450 3440 3790 3510
rect 2450 3320 3790 3390
rect 2450 3200 3790 3270
rect 2450 2730 3150 2800
rect 2450 2610 3790 2680
rect 2450 2490 3790 2560
rect 2450 2370 3790 2440
rect 2450 2250 3790 2320
rect 2450 2130 3790 2200
<< locali >>
rect 4610 5250 4690 5270
rect 4610 5210 4630 5250
rect 4670 5210 4690 5250
rect 4610 5190 4690 5210
rect 5010 5250 5090 5270
rect 5010 5210 5030 5250
rect 5070 5210 5090 5250
rect 5010 5190 5090 5210
rect 5410 5250 5490 5270
rect 5410 5210 5430 5250
rect 5470 5210 5490 5250
rect 5410 5190 5490 5210
rect 5810 5250 5890 5270
rect 5810 5210 5830 5250
rect 5870 5210 5890 5250
rect 5810 5190 5890 5210
rect 6210 5250 6290 5270
rect 6210 5210 6230 5250
rect 6270 5210 6290 5250
rect 6210 5190 6290 5210
rect 6610 5250 6690 5270
rect 6610 5210 6630 5250
rect 6670 5210 6690 5250
rect 6610 5190 6690 5210
rect 7010 5250 7090 5270
rect 7010 5210 7030 5250
rect 7070 5210 7090 5250
rect 7010 5190 7090 5210
rect 7410 5250 7490 5270
rect 7410 5210 7430 5250
rect 7470 5210 7490 5250
rect 7410 5190 7490 5210
rect 7810 5250 7890 5270
rect 7810 5210 7830 5250
rect 7870 5210 7890 5250
rect 7810 5190 7890 5210
rect 8210 5250 8290 5270
rect 8210 5210 8230 5250
rect 8270 5210 8290 5250
rect 8210 5190 8290 5210
rect 4630 5150 4670 5190
rect 5030 5150 5070 5190
rect 5430 5150 5470 5190
rect 5830 5150 5870 5190
rect 6230 5150 6270 5190
rect 6630 5150 6670 5190
rect 7030 5150 7070 5190
rect 7430 5150 7470 5190
rect 7830 5150 7870 5190
rect 8230 5150 8270 5190
rect 4340 5130 4480 5150
rect 4340 5090 4350 5130
rect 4390 5090 4430 5130
rect 4470 5090 4480 5130
rect 4340 5030 4480 5090
rect 4340 4990 4350 5030
rect 4390 4990 4430 5030
rect 4470 4990 4480 5030
rect 4340 4930 4480 4990
rect 4340 4890 4350 4930
rect 4390 4890 4430 4930
rect 4470 4890 4480 4930
rect 4340 4830 4480 4890
rect 4340 4790 4350 4830
rect 4390 4790 4430 4830
rect 4470 4790 4480 4830
rect 1890 4730 2010 4750
rect 1890 4690 1910 4730
rect 1950 4690 2010 4730
rect 1890 4680 2010 4690
rect 1890 4670 1970 4680
rect 3790 4630 4230 4680
rect 4340 4730 4480 4790
rect 4340 4690 4350 4730
rect 4390 4690 4430 4730
rect 4470 4690 4480 4730
rect 4340 4630 4480 4690
rect 4340 4590 4350 4630
rect 4390 4590 4430 4630
rect 4470 4590 4480 4630
rect 2010 4510 2450 4560
rect 4340 4530 4480 4590
rect 3790 4390 4230 4440
rect 4340 4490 4350 4530
rect 4390 4490 4430 4530
rect 4470 4490 4480 4530
rect 4340 4430 4480 4490
rect 4340 4390 4350 4430
rect 4390 4390 4430 4430
rect 4470 4390 4480 4430
rect 4340 4370 4480 4390
rect 4620 5130 4680 5150
rect 4620 5090 4630 5130
rect 4670 5090 4680 5130
rect 4620 5030 4680 5090
rect 4620 4990 4630 5030
rect 4670 4990 4680 5030
rect 4620 4930 4680 4990
rect 4620 4890 4630 4930
rect 4670 4890 4680 4930
rect 4620 4830 4680 4890
rect 4620 4790 4630 4830
rect 4670 4790 4680 4830
rect 4620 4730 4680 4790
rect 4620 4690 4630 4730
rect 4670 4690 4680 4730
rect 4620 4630 4680 4690
rect 4620 4590 4630 4630
rect 4670 4590 4680 4630
rect 4620 4530 4680 4590
rect 4620 4490 4630 4530
rect 4670 4490 4680 4530
rect 4620 4430 4680 4490
rect 4620 4390 4630 4430
rect 4670 4390 4680 4430
rect 4620 4370 4680 4390
rect 4820 5130 4880 5150
rect 4820 5090 4830 5130
rect 4870 5090 4880 5130
rect 4820 5030 4880 5090
rect 4820 4990 4830 5030
rect 4870 4990 4880 5030
rect 4820 4930 4880 4990
rect 4820 4890 4830 4930
rect 4870 4890 4880 4930
rect 4820 4830 4880 4890
rect 4820 4790 4830 4830
rect 4870 4790 4880 4830
rect 4820 4730 4880 4790
rect 4820 4690 4830 4730
rect 4870 4690 4880 4730
rect 4820 4630 4880 4690
rect 4820 4590 4830 4630
rect 4870 4590 4880 4630
rect 4820 4530 4880 4590
rect 4820 4490 4830 4530
rect 4870 4490 4880 4530
rect 4820 4430 4880 4490
rect 4820 4390 4830 4430
rect 4870 4390 4880 4430
rect 4820 4370 4880 4390
rect 5020 5130 5080 5150
rect 5020 5090 5030 5130
rect 5070 5090 5080 5130
rect 5020 5030 5080 5090
rect 5020 4990 5030 5030
rect 5070 4990 5080 5030
rect 5020 4930 5080 4990
rect 5020 4890 5030 4930
rect 5070 4890 5080 4930
rect 5020 4830 5080 4890
rect 5020 4790 5030 4830
rect 5070 4790 5080 4830
rect 5020 4730 5080 4790
rect 5020 4690 5030 4730
rect 5070 4690 5080 4730
rect 5020 4630 5080 4690
rect 5020 4590 5030 4630
rect 5070 4590 5080 4630
rect 5020 4530 5080 4590
rect 5020 4490 5030 4530
rect 5070 4490 5080 4530
rect 5020 4430 5080 4490
rect 5020 4390 5030 4430
rect 5070 4390 5080 4430
rect 5020 4370 5080 4390
rect 5220 5130 5280 5150
rect 5220 5090 5230 5130
rect 5270 5090 5280 5130
rect 5220 5030 5280 5090
rect 5220 4990 5230 5030
rect 5270 4990 5280 5030
rect 5220 4930 5280 4990
rect 5220 4890 5230 4930
rect 5270 4890 5280 4930
rect 5220 4830 5280 4890
rect 5220 4790 5230 4830
rect 5270 4790 5280 4830
rect 5220 4730 5280 4790
rect 5220 4690 5230 4730
rect 5270 4690 5280 4730
rect 5220 4630 5280 4690
rect 5220 4590 5230 4630
rect 5270 4590 5280 4630
rect 5220 4530 5280 4590
rect 5220 4490 5230 4530
rect 5270 4490 5280 4530
rect 5220 4430 5280 4490
rect 5220 4390 5230 4430
rect 5270 4390 5280 4430
rect 5220 4370 5280 4390
rect 5420 5130 5480 5150
rect 5420 5090 5430 5130
rect 5470 5090 5480 5130
rect 5420 5030 5480 5090
rect 5420 4990 5430 5030
rect 5470 4990 5480 5030
rect 5420 4930 5480 4990
rect 5420 4890 5430 4930
rect 5470 4890 5480 4930
rect 5420 4830 5480 4890
rect 5420 4790 5430 4830
rect 5470 4790 5480 4830
rect 5420 4730 5480 4790
rect 5420 4690 5430 4730
rect 5470 4690 5480 4730
rect 5420 4630 5480 4690
rect 5420 4590 5430 4630
rect 5470 4590 5480 4630
rect 5420 4530 5480 4590
rect 5420 4490 5430 4530
rect 5470 4490 5480 4530
rect 5420 4430 5480 4490
rect 5420 4390 5430 4430
rect 5470 4390 5480 4430
rect 5420 4370 5480 4390
rect 5620 5130 5680 5150
rect 5620 5090 5630 5130
rect 5670 5090 5680 5130
rect 5620 5030 5680 5090
rect 5620 4990 5630 5030
rect 5670 4990 5680 5030
rect 5620 4930 5680 4990
rect 5620 4890 5630 4930
rect 5670 4890 5680 4930
rect 5620 4830 5680 4890
rect 5620 4790 5630 4830
rect 5670 4790 5680 4830
rect 5620 4730 5680 4790
rect 5620 4690 5630 4730
rect 5670 4690 5680 4730
rect 5620 4630 5680 4690
rect 5620 4590 5630 4630
rect 5670 4590 5680 4630
rect 5620 4530 5680 4590
rect 5620 4490 5630 4530
rect 5670 4490 5680 4530
rect 5620 4430 5680 4490
rect 5620 4390 5630 4430
rect 5670 4390 5680 4430
rect 5620 4370 5680 4390
rect 5820 5130 5880 5150
rect 5820 5090 5830 5130
rect 5870 5090 5880 5130
rect 5820 5030 5880 5090
rect 5820 4990 5830 5030
rect 5870 4990 5880 5030
rect 5820 4930 5880 4990
rect 5820 4890 5830 4930
rect 5870 4890 5880 4930
rect 5820 4830 5880 4890
rect 5820 4790 5830 4830
rect 5870 4790 5880 4830
rect 5820 4730 5880 4790
rect 5820 4690 5830 4730
rect 5870 4690 5880 4730
rect 5820 4630 5880 4690
rect 5820 4590 5830 4630
rect 5870 4590 5880 4630
rect 5820 4530 5880 4590
rect 5820 4490 5830 4530
rect 5870 4490 5880 4530
rect 5820 4430 5880 4490
rect 5820 4390 5830 4430
rect 5870 4390 5880 4430
rect 5820 4370 5880 4390
rect 6020 5130 6080 5150
rect 6020 5090 6030 5130
rect 6070 5090 6080 5130
rect 6020 5030 6080 5090
rect 6020 4990 6030 5030
rect 6070 4990 6080 5030
rect 6020 4930 6080 4990
rect 6020 4890 6030 4930
rect 6070 4890 6080 4930
rect 6020 4830 6080 4890
rect 6020 4790 6030 4830
rect 6070 4790 6080 4830
rect 6020 4730 6080 4790
rect 6020 4690 6030 4730
rect 6070 4690 6080 4730
rect 6020 4630 6080 4690
rect 6020 4590 6030 4630
rect 6070 4590 6080 4630
rect 6020 4530 6080 4590
rect 6020 4490 6030 4530
rect 6070 4490 6080 4530
rect 6020 4430 6080 4490
rect 6020 4390 6030 4430
rect 6070 4390 6080 4430
rect 6020 4370 6080 4390
rect 6220 5130 6280 5150
rect 6220 5090 6230 5130
rect 6270 5090 6280 5130
rect 6220 5030 6280 5090
rect 6220 4990 6230 5030
rect 6270 4990 6280 5030
rect 6220 4930 6280 4990
rect 6220 4890 6230 4930
rect 6270 4890 6280 4930
rect 6220 4830 6280 4890
rect 6220 4790 6230 4830
rect 6270 4790 6280 4830
rect 6220 4730 6280 4790
rect 6220 4690 6230 4730
rect 6270 4690 6280 4730
rect 6220 4630 6280 4690
rect 6220 4590 6230 4630
rect 6270 4590 6280 4630
rect 6220 4530 6280 4590
rect 6220 4490 6230 4530
rect 6270 4490 6280 4530
rect 6220 4430 6280 4490
rect 6220 4390 6230 4430
rect 6270 4390 6280 4430
rect 6220 4370 6280 4390
rect 6420 5130 6480 5150
rect 6420 5090 6430 5130
rect 6470 5090 6480 5130
rect 6420 5030 6480 5090
rect 6420 4990 6430 5030
rect 6470 4990 6480 5030
rect 6420 4930 6480 4990
rect 6420 4890 6430 4930
rect 6470 4890 6480 4930
rect 6420 4830 6480 4890
rect 6420 4790 6430 4830
rect 6470 4790 6480 4830
rect 6420 4730 6480 4790
rect 6420 4690 6430 4730
rect 6470 4690 6480 4730
rect 6420 4630 6480 4690
rect 6420 4590 6430 4630
rect 6470 4590 6480 4630
rect 6420 4530 6480 4590
rect 6420 4490 6430 4530
rect 6470 4490 6480 4530
rect 6420 4430 6480 4490
rect 6420 4390 6430 4430
rect 6470 4390 6480 4430
rect 6420 4370 6480 4390
rect 6620 5130 6680 5150
rect 6620 5090 6630 5130
rect 6670 5090 6680 5130
rect 6620 5030 6680 5090
rect 6620 4990 6630 5030
rect 6670 4990 6680 5030
rect 6620 4930 6680 4990
rect 6620 4890 6630 4930
rect 6670 4890 6680 4930
rect 6620 4830 6680 4890
rect 6620 4790 6630 4830
rect 6670 4790 6680 4830
rect 6620 4730 6680 4790
rect 6620 4690 6630 4730
rect 6670 4690 6680 4730
rect 6620 4630 6680 4690
rect 6620 4590 6630 4630
rect 6670 4590 6680 4630
rect 6620 4530 6680 4590
rect 6620 4490 6630 4530
rect 6670 4490 6680 4530
rect 6620 4430 6680 4490
rect 6620 4390 6630 4430
rect 6670 4390 6680 4430
rect 6620 4370 6680 4390
rect 6820 5130 6880 5150
rect 6820 5090 6830 5130
rect 6870 5090 6880 5130
rect 6820 5030 6880 5090
rect 6820 4990 6830 5030
rect 6870 4990 6880 5030
rect 6820 4930 6880 4990
rect 6820 4890 6830 4930
rect 6870 4890 6880 4930
rect 6820 4830 6880 4890
rect 6820 4790 6830 4830
rect 6870 4790 6880 4830
rect 6820 4730 6880 4790
rect 6820 4690 6830 4730
rect 6870 4690 6880 4730
rect 6820 4630 6880 4690
rect 6820 4590 6830 4630
rect 6870 4590 6880 4630
rect 6820 4530 6880 4590
rect 6820 4490 6830 4530
rect 6870 4490 6880 4530
rect 6820 4430 6880 4490
rect 6820 4390 6830 4430
rect 6870 4390 6880 4430
rect 6820 4370 6880 4390
rect 7020 5130 7080 5150
rect 7020 5090 7030 5130
rect 7070 5090 7080 5130
rect 7020 5030 7080 5090
rect 7020 4990 7030 5030
rect 7070 4990 7080 5030
rect 7020 4930 7080 4990
rect 7020 4890 7030 4930
rect 7070 4890 7080 4930
rect 7020 4830 7080 4890
rect 7020 4790 7030 4830
rect 7070 4790 7080 4830
rect 7020 4730 7080 4790
rect 7020 4690 7030 4730
rect 7070 4690 7080 4730
rect 7020 4630 7080 4690
rect 7020 4590 7030 4630
rect 7070 4590 7080 4630
rect 7020 4530 7080 4590
rect 7020 4490 7030 4530
rect 7070 4490 7080 4530
rect 7020 4430 7080 4490
rect 7020 4390 7030 4430
rect 7070 4390 7080 4430
rect 7020 4370 7080 4390
rect 7220 5130 7280 5150
rect 7220 5090 7230 5130
rect 7270 5090 7280 5130
rect 7220 5030 7280 5090
rect 7220 4990 7230 5030
rect 7270 4990 7280 5030
rect 7220 4930 7280 4990
rect 7220 4890 7230 4930
rect 7270 4890 7280 4930
rect 7220 4830 7280 4890
rect 7220 4790 7230 4830
rect 7270 4790 7280 4830
rect 7220 4730 7280 4790
rect 7220 4690 7230 4730
rect 7270 4690 7280 4730
rect 7220 4630 7280 4690
rect 7220 4590 7230 4630
rect 7270 4590 7280 4630
rect 7220 4530 7280 4590
rect 7220 4490 7230 4530
rect 7270 4490 7280 4530
rect 7220 4430 7280 4490
rect 7220 4390 7230 4430
rect 7270 4390 7280 4430
rect 7220 4370 7280 4390
rect 7420 5130 7480 5150
rect 7420 5090 7430 5130
rect 7470 5090 7480 5130
rect 7420 5030 7480 5090
rect 7420 4990 7430 5030
rect 7470 4990 7480 5030
rect 7420 4930 7480 4990
rect 7420 4890 7430 4930
rect 7470 4890 7480 4930
rect 7420 4830 7480 4890
rect 7420 4790 7430 4830
rect 7470 4790 7480 4830
rect 7420 4730 7480 4790
rect 7420 4690 7430 4730
rect 7470 4690 7480 4730
rect 7420 4630 7480 4690
rect 7420 4590 7430 4630
rect 7470 4590 7480 4630
rect 7420 4530 7480 4590
rect 7420 4490 7430 4530
rect 7470 4490 7480 4530
rect 7420 4430 7480 4490
rect 7420 4390 7430 4430
rect 7470 4390 7480 4430
rect 7420 4370 7480 4390
rect 7620 5130 7680 5150
rect 7620 5090 7630 5130
rect 7670 5090 7680 5130
rect 7620 5030 7680 5090
rect 7620 4990 7630 5030
rect 7670 4990 7680 5030
rect 7620 4930 7680 4990
rect 7620 4890 7630 4930
rect 7670 4890 7680 4930
rect 7620 4830 7680 4890
rect 7620 4790 7630 4830
rect 7670 4790 7680 4830
rect 7620 4730 7680 4790
rect 7620 4690 7630 4730
rect 7670 4690 7680 4730
rect 7620 4630 7680 4690
rect 7620 4590 7630 4630
rect 7670 4590 7680 4630
rect 7620 4530 7680 4590
rect 7620 4490 7630 4530
rect 7670 4490 7680 4530
rect 7620 4430 7680 4490
rect 7620 4390 7630 4430
rect 7670 4390 7680 4430
rect 7620 4370 7680 4390
rect 7820 5130 7880 5150
rect 7820 5090 7830 5130
rect 7870 5090 7880 5130
rect 7820 5030 7880 5090
rect 7820 4990 7830 5030
rect 7870 4990 7880 5030
rect 7820 4930 7880 4990
rect 7820 4890 7830 4930
rect 7870 4890 7880 4930
rect 7820 4830 7880 4890
rect 7820 4790 7830 4830
rect 7870 4790 7880 4830
rect 7820 4730 7880 4790
rect 7820 4690 7830 4730
rect 7870 4690 7880 4730
rect 7820 4630 7880 4690
rect 7820 4590 7830 4630
rect 7870 4590 7880 4630
rect 7820 4530 7880 4590
rect 7820 4490 7830 4530
rect 7870 4490 7880 4530
rect 7820 4430 7880 4490
rect 7820 4390 7830 4430
rect 7870 4390 7880 4430
rect 7820 4370 7880 4390
rect 8020 5130 8080 5150
rect 8020 5090 8030 5130
rect 8070 5090 8080 5130
rect 8020 5030 8080 5090
rect 8020 4990 8030 5030
rect 8070 4990 8080 5030
rect 8020 4930 8080 4990
rect 8020 4890 8030 4930
rect 8070 4890 8080 4930
rect 8020 4830 8080 4890
rect 8020 4790 8030 4830
rect 8070 4790 8080 4830
rect 8020 4730 8080 4790
rect 8020 4690 8030 4730
rect 8070 4690 8080 4730
rect 8020 4630 8080 4690
rect 8020 4590 8030 4630
rect 8070 4590 8080 4630
rect 8020 4530 8080 4590
rect 8020 4490 8030 4530
rect 8070 4490 8080 4530
rect 8020 4430 8080 4490
rect 8020 4390 8030 4430
rect 8070 4390 8080 4430
rect 8020 4370 8080 4390
rect 8220 5130 8280 5150
rect 8220 5090 8230 5130
rect 8270 5090 8280 5130
rect 8220 5030 8280 5090
rect 8220 4990 8230 5030
rect 8270 4990 8280 5030
rect 8220 4930 8280 4990
rect 8220 4890 8230 4930
rect 8270 4890 8280 4930
rect 8220 4830 8280 4890
rect 8220 4790 8230 4830
rect 8270 4790 8280 4830
rect 8220 4730 8280 4790
rect 8220 4690 8230 4730
rect 8270 4690 8280 4730
rect 8220 4630 8280 4690
rect 8220 4590 8230 4630
rect 8270 4590 8280 4630
rect 8220 4530 8280 4590
rect 8220 4490 8230 4530
rect 8270 4490 8280 4530
rect 8220 4430 8280 4490
rect 8220 4390 8230 4430
rect 8270 4390 8280 4430
rect 8220 4370 8280 4390
rect 8420 5130 8560 5150
rect 8420 5090 8430 5130
rect 8470 5090 8510 5130
rect 8550 5090 8560 5130
rect 8420 5030 8560 5090
rect 8420 4990 8430 5030
rect 8470 4990 8510 5030
rect 8550 4990 8560 5030
rect 8420 4930 8560 4990
rect 8420 4890 8430 4930
rect 8470 4890 8510 4930
rect 8550 4890 8560 4930
rect 8420 4830 8560 4890
rect 8420 4790 8430 4830
rect 8470 4790 8510 4830
rect 8550 4790 8560 4830
rect 8420 4730 8560 4790
rect 8420 4690 8430 4730
rect 8470 4690 8510 4730
rect 8550 4690 8560 4730
rect 8420 4630 8560 4690
rect 8420 4590 8430 4630
rect 8470 4590 8510 4630
rect 8550 4590 8560 4630
rect 8420 4530 8560 4590
rect 8420 4490 8430 4530
rect 8470 4490 8510 4530
rect 8550 4490 8560 4530
rect 8420 4430 8560 4490
rect 10410 4530 10830 4550
rect 10410 4490 10430 4530
rect 10470 4510 10830 4530
rect 10470 4490 10490 4510
rect 10410 4470 10490 4490
rect 10610 4450 10690 4470
rect 10610 4430 10630 4450
rect 8420 4390 8430 4430
rect 8470 4390 8510 4430
rect 8550 4390 8560 4430
rect 8420 4370 8560 4390
rect 10460 4410 10630 4430
rect 10670 4410 10690 4450
rect 10460 4390 10690 4410
rect 4830 4330 4870 4370
rect 2010 4270 2450 4320
rect 4810 4310 4890 4330
rect 4810 4270 4830 4310
rect 4870 4270 4890 4310
rect 4810 4250 4890 4270
rect 5230 4240 5270 4370
rect 3790 4140 4230 4200
rect 5210 4220 5290 4240
rect 5210 4180 5230 4220
rect 5270 4180 5290 4220
rect 5210 4160 5290 4180
rect 5630 4150 5670 4370
rect 6030 4240 6070 4370
rect 6210 4310 6290 4330
rect 6210 4270 6230 4310
rect 6270 4270 6290 4310
rect 6210 4250 6290 4270
rect 6010 4220 6090 4240
rect 6010 4180 6030 4220
rect 6070 4180 6090 4220
rect 6010 4160 6090 4180
rect 6430 4150 6470 4370
rect 6830 4330 6870 4370
rect 6610 4310 6690 4330
rect 6610 4270 6630 4310
rect 6670 4270 6690 4310
rect 6610 4250 6690 4270
rect 6810 4310 6890 4330
rect 6810 4270 6830 4310
rect 6870 4270 6890 4310
rect 6810 4250 6890 4270
rect 7230 4150 7270 4370
rect 7630 4330 7670 4370
rect 7610 4310 7690 4330
rect 7610 4270 7630 4310
rect 7670 4270 7690 4310
rect 7610 4250 7690 4270
rect 8030 4240 8070 4370
rect 10460 4350 10500 4390
rect 10790 4350 10830 4510
rect 10260 4330 10400 4350
rect 10260 4290 10270 4330
rect 10310 4290 10350 4330
rect 10390 4290 10400 4330
rect 8010 4220 8090 4240
rect 8010 4180 8030 4220
rect 8070 4180 8090 4220
rect 8010 4160 8090 4180
rect 10260 4230 10400 4290
rect 10260 4190 10270 4230
rect 10310 4190 10350 4230
rect 10390 4190 10400 4230
rect 3790 4100 3810 4140
rect 3850 4100 3900 4140
rect 3940 4100 3990 4140
rect 4030 4100 4080 4140
rect 4120 4100 4170 4140
rect 4210 4100 4230 4140
rect 3790 4080 4230 4100
rect 5610 4130 5690 4150
rect 5610 4090 5630 4130
rect 5670 4090 5690 4130
rect 5610 4070 5690 4090
rect 6410 4130 6490 4150
rect 6410 4090 6430 4130
rect 6470 4090 6490 4130
rect 6410 4070 6490 4090
rect 7210 4130 7290 4150
rect 7210 4090 7230 4130
rect 7270 4090 7290 4130
rect 7210 4070 7290 4090
rect 10260 4130 10400 4190
rect 10260 4090 10270 4130
rect 10310 4090 10350 4130
rect 10390 4090 10400 4130
rect 10260 4030 10400 4090
rect 10260 3990 10270 4030
rect 10310 3990 10350 4030
rect 10390 3990 10400 4030
rect 10260 3970 10400 3990
rect 10450 4330 10510 4350
rect 10450 4290 10460 4330
rect 10500 4290 10510 4330
rect 10450 4230 10510 4290
rect 10450 4190 10460 4230
rect 10500 4190 10510 4230
rect 10450 4130 10510 4190
rect 10450 4090 10460 4130
rect 10500 4090 10510 4130
rect 10450 4030 10510 4090
rect 10450 3990 10460 4030
rect 10500 3990 10510 4030
rect 10450 3970 10510 3990
rect 10590 4330 10650 4350
rect 10590 4290 10600 4330
rect 10640 4290 10650 4330
rect 10590 4230 10650 4290
rect 10590 4190 10600 4230
rect 10640 4190 10650 4230
rect 10590 4130 10650 4190
rect 10590 4090 10600 4130
rect 10640 4090 10650 4130
rect 10590 4030 10650 4090
rect 10590 3990 10600 4030
rect 10640 3990 10650 4030
rect 10590 3970 10650 3990
rect 10700 4330 10840 4350
rect 10700 4290 10710 4330
rect 10750 4290 10790 4330
rect 10830 4290 10840 4330
rect 10700 4230 10840 4290
rect 10700 4190 10710 4230
rect 10750 4190 10790 4230
rect 10830 4190 10840 4230
rect 10700 4130 10840 4190
rect 10700 4090 10710 4130
rect 10750 4090 10790 4130
rect 10830 4090 10840 4130
rect 10700 4030 10840 4090
rect 10700 3990 10710 4030
rect 10750 3990 10790 4030
rect 10830 3990 10840 4030
rect 10700 3970 10840 3990
rect 4450 3940 4530 3960
rect 4450 3900 4470 3940
rect 4510 3900 4530 3940
rect 4450 3880 4530 3900
rect 4650 3940 4730 3960
rect 4650 3900 4670 3940
rect 4710 3900 4730 3940
rect 4650 3880 4730 3900
rect 5050 3940 5130 3960
rect 5050 3900 5070 3940
rect 5110 3900 5130 3940
rect 5050 3880 5130 3900
rect 5450 3940 5530 3960
rect 5450 3900 5470 3940
rect 5510 3900 5530 3940
rect 5450 3880 5530 3900
rect 5650 3940 5730 3960
rect 5650 3900 5670 3940
rect 5710 3900 5730 3940
rect 5650 3880 5730 3900
rect 5810 3940 5890 3960
rect 5810 3900 5830 3940
rect 5870 3900 5890 3940
rect 5810 3880 5890 3900
rect 6010 3940 6090 3960
rect 6010 3900 6030 3940
rect 6070 3900 6090 3940
rect 6010 3880 6090 3900
rect 6210 3940 6290 3960
rect 6210 3900 6230 3940
rect 6270 3900 6290 3940
rect 6210 3880 6290 3900
rect 6410 3940 6490 3960
rect 6410 3900 6430 3940
rect 6470 3900 6490 3940
rect 6410 3880 6490 3900
rect 6610 3940 6690 3960
rect 6610 3900 6630 3940
rect 6670 3900 6690 3940
rect 6610 3880 6690 3900
rect 6810 3940 6890 3960
rect 6810 3900 6830 3940
rect 6870 3900 6890 3940
rect 6810 3880 6890 3900
rect 7010 3940 7090 3960
rect 7010 3900 7030 3940
rect 7070 3900 7090 3940
rect 7010 3880 7090 3900
rect 7170 3940 7250 3960
rect 7170 3900 7190 3940
rect 7230 3900 7250 3940
rect 7170 3880 7250 3900
rect 7370 3940 7450 3960
rect 7370 3900 7390 3940
rect 7430 3900 7450 3940
rect 7370 3880 7450 3900
rect 7770 3940 7850 3960
rect 7770 3900 7790 3940
rect 7830 3900 7850 3940
rect 7770 3880 7850 3900
rect 8170 3940 8250 3960
rect 8170 3900 8190 3940
rect 8230 3900 8250 3940
rect 8170 3880 8250 3900
rect 8370 3940 8450 3960
rect 8370 3900 8390 3940
rect 8430 3900 8450 3940
rect 10460 3900 10500 3970
rect 10600 3900 10640 3970
rect 8370 3880 8450 3900
rect 4470 3840 4510 3880
rect 4670 3840 4710 3880
rect 5070 3840 5110 3880
rect 5470 3840 5510 3880
rect 5670 3840 5710 3880
rect 5830 3840 5870 3880
rect 6030 3840 6070 3880
rect 6230 3840 6270 3880
rect 6430 3840 6470 3880
rect 6630 3840 6670 3880
rect 6830 3840 6870 3880
rect 7030 3840 7070 3880
rect 7190 3840 7230 3880
rect 7390 3840 7430 3880
rect 7790 3840 7830 3880
rect 8190 3840 8230 3880
rect 8390 3840 8430 3880
rect 4380 3820 4520 3840
rect 4380 3780 4390 3820
rect 4430 3780 4470 3820
rect 4510 3780 4520 3820
rect 1890 3730 2010 3750
rect 1890 3690 1910 3730
rect 1950 3690 2010 3730
rect 1890 3680 2010 3690
rect 1890 3670 1970 3680
rect 3790 3630 4230 3680
rect 4380 3720 4520 3780
rect 4380 3680 4390 3720
rect 4430 3680 4470 3720
rect 4510 3680 4520 3720
rect 4380 3620 4520 3680
rect 4380 3580 4390 3620
rect 4430 3580 4470 3620
rect 4510 3580 4520 3620
rect 2010 3510 2450 3560
rect 4380 3520 4520 3580
rect 4380 3480 4390 3520
rect 4430 3480 4470 3520
rect 4510 3480 4520 3520
rect 4380 3460 4520 3480
rect 4660 3820 4720 3840
rect 4660 3780 4670 3820
rect 4710 3780 4720 3820
rect 4660 3720 4720 3780
rect 4660 3680 4670 3720
rect 4710 3680 4720 3720
rect 4660 3620 4720 3680
rect 4660 3580 4670 3620
rect 4710 3580 4720 3620
rect 4660 3520 4720 3580
rect 4660 3480 4670 3520
rect 4710 3480 4720 3520
rect 4660 3460 4720 3480
rect 4860 3820 4920 3840
rect 4860 3780 4870 3820
rect 4910 3780 4920 3820
rect 4860 3720 4920 3780
rect 4860 3680 4870 3720
rect 4910 3680 4920 3720
rect 4860 3620 4920 3680
rect 4860 3580 4870 3620
rect 4910 3580 4920 3620
rect 4860 3520 4920 3580
rect 4860 3480 4870 3520
rect 4910 3480 4920 3520
rect 4860 3460 4920 3480
rect 5060 3820 5120 3840
rect 5060 3780 5070 3820
rect 5110 3780 5120 3820
rect 5060 3720 5120 3780
rect 5060 3680 5070 3720
rect 5110 3680 5120 3720
rect 5060 3620 5120 3680
rect 5060 3580 5070 3620
rect 5110 3580 5120 3620
rect 5060 3520 5120 3580
rect 5060 3480 5070 3520
rect 5110 3480 5120 3520
rect 5060 3460 5120 3480
rect 5260 3820 5320 3840
rect 5260 3780 5270 3820
rect 5310 3780 5320 3820
rect 5260 3720 5320 3780
rect 5260 3680 5270 3720
rect 5310 3680 5320 3720
rect 5260 3620 5320 3680
rect 5260 3580 5270 3620
rect 5310 3580 5320 3620
rect 5260 3520 5320 3580
rect 5260 3480 5270 3520
rect 5310 3480 5320 3520
rect 5260 3460 5320 3480
rect 5460 3820 5520 3840
rect 5460 3780 5470 3820
rect 5510 3780 5520 3820
rect 5460 3720 5520 3780
rect 5460 3680 5470 3720
rect 5510 3680 5520 3720
rect 5460 3620 5520 3680
rect 5460 3580 5470 3620
rect 5510 3580 5520 3620
rect 5460 3520 5520 3580
rect 5460 3480 5470 3520
rect 5510 3480 5520 3520
rect 5460 3460 5520 3480
rect 5660 3820 5880 3840
rect 5660 3780 5670 3820
rect 5710 3780 5750 3820
rect 5790 3780 5830 3820
rect 5870 3780 5880 3820
rect 5660 3720 5880 3780
rect 5660 3680 5670 3720
rect 5710 3680 5750 3720
rect 5790 3680 5830 3720
rect 5870 3680 5880 3720
rect 5660 3620 5880 3680
rect 5660 3580 5670 3620
rect 5710 3580 5750 3620
rect 5790 3580 5830 3620
rect 5870 3580 5880 3620
rect 5660 3520 5880 3580
rect 5660 3480 5670 3520
rect 5710 3480 5750 3520
rect 5790 3480 5830 3520
rect 5870 3480 5880 3520
rect 5660 3460 5880 3480
rect 6020 3820 6080 3840
rect 6020 3780 6030 3820
rect 6070 3780 6080 3820
rect 6020 3720 6080 3780
rect 6020 3680 6030 3720
rect 6070 3680 6080 3720
rect 6020 3620 6080 3680
rect 6020 3580 6030 3620
rect 6070 3580 6080 3620
rect 6020 3520 6080 3580
rect 6020 3480 6030 3520
rect 6070 3480 6080 3520
rect 6020 3460 6080 3480
rect 6220 3820 6280 3840
rect 6220 3780 6230 3820
rect 6270 3780 6280 3820
rect 6220 3720 6280 3780
rect 6220 3680 6230 3720
rect 6270 3680 6280 3720
rect 6220 3620 6280 3680
rect 6220 3580 6230 3620
rect 6270 3580 6280 3620
rect 6220 3520 6280 3580
rect 6220 3480 6230 3520
rect 6270 3480 6280 3520
rect 6220 3460 6280 3480
rect 6420 3820 6480 3840
rect 6420 3780 6430 3820
rect 6470 3780 6480 3820
rect 6420 3720 6480 3780
rect 6420 3680 6430 3720
rect 6470 3680 6480 3720
rect 6420 3620 6480 3680
rect 6420 3580 6430 3620
rect 6470 3580 6480 3620
rect 6420 3520 6480 3580
rect 6420 3480 6430 3520
rect 6470 3480 6480 3520
rect 6420 3460 6480 3480
rect 6620 3820 6680 3840
rect 6620 3780 6630 3820
rect 6670 3780 6680 3820
rect 6620 3720 6680 3780
rect 6620 3680 6630 3720
rect 6670 3680 6680 3720
rect 6620 3620 6680 3680
rect 6620 3580 6630 3620
rect 6670 3580 6680 3620
rect 6620 3520 6680 3580
rect 6620 3480 6630 3520
rect 6670 3480 6680 3520
rect 6620 3460 6680 3480
rect 6820 3820 6880 3840
rect 6820 3780 6830 3820
rect 6870 3780 6880 3820
rect 6820 3720 6880 3780
rect 6820 3680 6830 3720
rect 6870 3680 6880 3720
rect 6820 3620 6880 3680
rect 6820 3580 6830 3620
rect 6870 3580 6880 3620
rect 6820 3520 6880 3580
rect 6820 3480 6830 3520
rect 6870 3480 6880 3520
rect 6820 3460 6880 3480
rect 7020 3820 7240 3840
rect 7020 3780 7030 3820
rect 7070 3780 7110 3820
rect 7150 3780 7190 3820
rect 7230 3780 7240 3820
rect 7020 3720 7240 3780
rect 7020 3680 7030 3720
rect 7070 3680 7110 3720
rect 7150 3680 7190 3720
rect 7230 3680 7240 3720
rect 7020 3620 7240 3680
rect 7020 3580 7030 3620
rect 7070 3580 7110 3620
rect 7150 3580 7190 3620
rect 7230 3580 7240 3620
rect 7020 3520 7240 3580
rect 7020 3480 7030 3520
rect 7070 3480 7110 3520
rect 7150 3480 7190 3520
rect 7230 3480 7240 3520
rect 7020 3460 7240 3480
rect 7380 3820 7440 3840
rect 7380 3780 7390 3820
rect 7430 3780 7440 3820
rect 7380 3720 7440 3780
rect 7380 3680 7390 3720
rect 7430 3680 7440 3720
rect 7380 3620 7440 3680
rect 7380 3580 7390 3620
rect 7430 3580 7440 3620
rect 7380 3520 7440 3580
rect 7380 3480 7390 3520
rect 7430 3480 7440 3520
rect 7380 3460 7440 3480
rect 7580 3820 7640 3840
rect 7580 3780 7590 3820
rect 7630 3780 7640 3820
rect 7580 3720 7640 3780
rect 7580 3680 7590 3720
rect 7630 3680 7640 3720
rect 7580 3620 7640 3680
rect 7580 3580 7590 3620
rect 7630 3580 7640 3620
rect 7580 3520 7640 3580
rect 7580 3480 7590 3520
rect 7630 3480 7640 3520
rect 7580 3460 7640 3480
rect 7780 3820 7840 3840
rect 7780 3780 7790 3820
rect 7830 3780 7840 3820
rect 7780 3720 7840 3780
rect 7780 3680 7790 3720
rect 7830 3680 7840 3720
rect 7780 3620 7840 3680
rect 7780 3580 7790 3620
rect 7830 3580 7840 3620
rect 7780 3520 7840 3580
rect 7780 3480 7790 3520
rect 7830 3480 7840 3520
rect 7780 3460 7840 3480
rect 7980 3820 8040 3840
rect 7980 3780 7990 3820
rect 8030 3780 8040 3820
rect 7980 3720 8040 3780
rect 7980 3680 7990 3720
rect 8030 3680 8040 3720
rect 7980 3620 8040 3680
rect 7980 3580 7990 3620
rect 8030 3580 8040 3620
rect 7980 3520 8040 3580
rect 7980 3480 7990 3520
rect 8030 3480 8040 3520
rect 7980 3460 8040 3480
rect 8180 3820 8240 3840
rect 8180 3780 8190 3820
rect 8230 3780 8240 3820
rect 8180 3720 8240 3780
rect 8180 3680 8190 3720
rect 8230 3680 8240 3720
rect 8180 3620 8240 3680
rect 8180 3580 8190 3620
rect 8230 3580 8240 3620
rect 8180 3520 8240 3580
rect 8180 3480 8190 3520
rect 8230 3480 8240 3520
rect 8180 3460 8240 3480
rect 8380 3820 8520 3840
rect 8380 3780 8390 3820
rect 8430 3780 8470 3820
rect 8510 3780 8520 3820
rect 8380 3720 8520 3780
rect 8380 3680 8390 3720
rect 8430 3680 8470 3720
rect 8510 3680 8520 3720
rect 8380 3620 8520 3680
rect 9230 3750 11290 3770
rect 9230 3710 9310 3750
rect 9350 3710 9470 3750
rect 9510 3710 9630 3750
rect 9670 3710 9790 3750
rect 9830 3710 9950 3750
rect 9990 3710 10110 3750
rect 10150 3710 10270 3750
rect 10310 3710 10430 3750
rect 10470 3710 10590 3750
rect 10630 3710 10750 3750
rect 10790 3710 10910 3750
rect 10950 3710 11070 3750
rect 11110 3710 11230 3750
rect 11270 3710 11290 3750
rect 9230 3690 11290 3710
rect 9230 3650 9270 3690
rect 8380 3580 8390 3620
rect 8430 3580 8470 3620
rect 8510 3580 8520 3620
rect 8380 3520 8520 3580
rect 8380 3480 8390 3520
rect 8430 3480 8470 3520
rect 8510 3480 8520 3520
rect 8380 3460 8520 3480
rect 9220 3630 9280 3650
rect 9220 3590 9230 3630
rect 9270 3590 9280 3630
rect 9220 3530 9280 3590
rect 9220 3490 9230 3530
rect 9270 3490 9280 3530
rect 9220 3470 9280 3490
rect 11300 3630 11440 3650
rect 11300 3590 11310 3630
rect 11350 3590 11390 3630
rect 11430 3590 11440 3630
rect 11300 3530 11440 3590
rect 11300 3490 11310 3530
rect 11350 3490 11390 3530
rect 11430 3490 11440 3530
rect 11300 3470 11440 3490
rect 3790 3390 4230 3440
rect 4870 3330 4910 3460
rect 5270 3420 5310 3460
rect 6230 3420 6270 3460
rect 6630 3420 6670 3460
rect 7590 3420 7630 3460
rect 5250 3400 5330 3420
rect 5250 3360 5270 3400
rect 5310 3360 5330 3400
rect 6230 3400 6670 3420
rect 6230 3380 6430 3400
rect 5250 3340 5330 3360
rect 6410 3360 6430 3380
rect 6470 3380 6670 3400
rect 7570 3400 7650 3420
rect 6470 3360 6490 3380
rect 6410 3340 6490 3360
rect 7570 3360 7590 3400
rect 7630 3360 7650 3400
rect 7570 3340 7650 3360
rect 7990 3330 8030 3460
rect 2010 3270 2450 3320
rect 4850 3310 4930 3330
rect 4850 3270 4870 3310
rect 4910 3270 4930 3310
rect 4850 3250 4930 3270
rect 5530 3250 5610 3330
rect 6110 3310 6190 3330
rect 6110 3270 6130 3310
rect 6170 3270 6190 3310
rect 6110 3250 6190 3270
rect 6710 3310 6790 3330
rect 6710 3270 6730 3310
rect 6770 3270 6790 3310
rect 6710 3250 6790 3270
rect 7290 3250 7370 3330
rect 7970 3310 8050 3330
rect 7970 3270 7990 3310
rect 8030 3270 8050 3310
rect 7970 3250 8050 3270
rect 3790 3140 4230 3200
rect 6410 3220 6490 3240
rect 6410 3180 6430 3220
rect 6470 3180 6490 3220
rect 6410 3160 6490 3180
rect 3790 3100 3810 3140
rect 3850 3100 3900 3140
rect 3940 3100 3990 3140
rect 4030 3100 4080 3140
rect 4120 3100 4170 3140
rect 4210 3100 4230 3140
rect 3790 3080 4230 3100
rect 5530 3130 5610 3150
rect 5530 3090 5550 3130
rect 5590 3090 5610 3130
rect 5530 3070 5610 3090
rect 5930 3130 6010 3150
rect 5930 3090 5950 3130
rect 5990 3090 6010 3130
rect 5930 3070 6010 3090
rect 6050 3130 6130 3150
rect 6050 3090 6070 3130
rect 6110 3090 6130 3130
rect 6050 3070 6130 3090
rect 6770 3130 6850 3150
rect 6770 3090 6790 3130
rect 6830 3090 6850 3130
rect 6770 3070 6850 3090
rect 6890 3130 6970 3150
rect 6890 3090 6910 3130
rect 6950 3090 6970 3130
rect 6890 3070 6970 3090
rect 7290 3130 7370 3150
rect 7290 3090 7310 3130
rect 7350 3090 7370 3130
rect 7290 3070 7370 3090
rect 5550 3030 5590 3070
rect 5950 3030 5990 3070
rect 6910 3030 6950 3070
rect 7310 3030 7350 3070
rect 5050 3010 5200 3030
rect 5050 2970 5070 3010
rect 5110 2970 5150 3010
rect 5190 2970 5200 3010
rect 5050 2910 5200 2970
rect 5050 2870 5070 2910
rect 5110 2870 5150 2910
rect 5190 2870 5200 2910
rect 5050 2850 5200 2870
rect 5340 3010 5400 3030
rect 5340 2970 5350 3010
rect 5390 2970 5400 3010
rect 5340 2910 5400 2970
rect 5340 2870 5350 2910
rect 5390 2870 5400 2910
rect 5340 2850 5400 2870
rect 5540 3010 5600 3030
rect 5540 2970 5550 3010
rect 5590 2970 5600 3010
rect 5540 2910 5600 2970
rect 5540 2870 5550 2910
rect 5590 2870 5600 2910
rect 5540 2850 5600 2870
rect 5740 3010 5800 3030
rect 5740 2970 5750 3010
rect 5790 2970 5800 3010
rect 5740 2910 5800 2970
rect 5740 2870 5750 2910
rect 5790 2870 5800 2910
rect 5740 2850 5800 2870
rect 5940 3010 6000 3030
rect 5940 2970 5950 3010
rect 5990 2970 6000 3010
rect 5940 2910 6000 2970
rect 5940 2870 5950 2910
rect 5990 2870 6000 2910
rect 5940 2850 6000 2870
rect 6140 3010 6200 3030
rect 6140 2970 6150 3010
rect 6190 2970 6200 3010
rect 6140 2910 6200 2970
rect 6140 2870 6150 2910
rect 6190 2870 6200 2910
rect 6140 2850 6200 2870
rect 6340 3010 6560 3030
rect 6340 2970 6350 3010
rect 6390 2970 6430 3010
rect 6470 2970 6510 3010
rect 6550 2970 6560 3010
rect 6340 2910 6560 2970
rect 6340 2870 6350 2910
rect 6390 2870 6430 2910
rect 6470 2870 6510 2910
rect 6550 2870 6560 2910
rect 6340 2850 6560 2870
rect 6700 3010 6760 3030
rect 6700 2970 6710 3010
rect 6750 2970 6760 3010
rect 6700 2910 6760 2970
rect 6700 2870 6710 2910
rect 6750 2870 6760 2910
rect 6700 2850 6760 2870
rect 6900 3010 6960 3030
rect 6900 2970 6910 3010
rect 6950 2970 6960 3010
rect 6900 2910 6960 2970
rect 6900 2870 6910 2910
rect 6950 2870 6960 2910
rect 6900 2850 6960 2870
rect 7100 3010 7160 3030
rect 7100 2970 7110 3010
rect 7150 2970 7160 3010
rect 7100 2910 7160 2970
rect 7100 2870 7110 2910
rect 7150 2870 7160 2910
rect 7100 2850 7160 2870
rect 7300 3010 7360 3030
rect 7300 2970 7310 3010
rect 7350 2970 7360 3010
rect 7300 2910 7360 2970
rect 7300 2870 7310 2910
rect 7350 2870 7360 2910
rect 7300 2850 7360 2870
rect 7500 3010 7560 3030
rect 7500 2970 7510 3010
rect 7550 2970 7560 3010
rect 7500 2910 7560 2970
rect 7500 2870 7510 2910
rect 7550 2870 7560 2910
rect 7500 2850 7560 2870
rect 7700 3010 7840 3030
rect 7700 2970 7710 3010
rect 7750 2970 7790 3010
rect 7830 2970 7840 3010
rect 7700 2910 7840 2970
rect 7700 2870 7710 2910
rect 7750 2870 7790 2910
rect 7830 2870 7840 2910
rect 7700 2850 7840 2870
rect 1890 2780 2010 2800
rect 1890 2740 1910 2780
rect 1950 2740 2010 2780
rect 1890 2730 2010 2740
rect 3590 2780 4230 2800
rect 3590 2740 3810 2780
rect 3850 2740 3900 2780
rect 3940 2740 3990 2780
rect 4030 2740 4080 2780
rect 4120 2740 4170 2780
rect 4210 2740 4230 2780
rect 3590 2730 4230 2740
rect 1890 2720 1970 2730
rect 3790 2680 4230 2730
rect 5150 2720 5190 2850
rect 5350 2720 5390 2850
rect 5530 2790 5610 2810
rect 5530 2750 5550 2790
rect 5590 2750 5610 2790
rect 5530 2730 5610 2750
rect 5750 2720 5790 2850
rect 6150 2720 6190 2850
rect 6350 2720 6390 2850
rect 6510 2720 6550 2850
rect 6710 2720 6750 2850
rect 7110 2720 7150 2850
rect 7290 2790 7370 2810
rect 7290 2750 7310 2790
rect 7350 2750 7370 2790
rect 7290 2730 7370 2750
rect 7510 2720 7550 2850
rect 7710 2720 7750 2850
rect 5130 2700 5210 2720
rect 5130 2660 5150 2700
rect 5190 2660 5210 2700
rect 5130 2640 5210 2660
rect 5330 2700 5410 2720
rect 5330 2660 5350 2700
rect 5390 2660 5410 2700
rect 5330 2640 5410 2660
rect 5730 2700 5810 2720
rect 5730 2660 5750 2700
rect 5790 2660 5810 2700
rect 5730 2640 5810 2660
rect 6130 2700 6210 2720
rect 6130 2660 6150 2700
rect 6190 2660 6210 2700
rect 6130 2640 6210 2660
rect 6330 2700 6410 2720
rect 6330 2660 6350 2700
rect 6390 2660 6410 2700
rect 6330 2640 6410 2660
rect 6490 2700 6570 2720
rect 6490 2660 6510 2700
rect 6550 2660 6570 2700
rect 6490 2640 6570 2660
rect 6690 2700 6770 2720
rect 6690 2660 6710 2700
rect 6750 2660 6770 2700
rect 6690 2640 6770 2660
rect 7090 2700 7170 2720
rect 7090 2660 7110 2700
rect 7150 2660 7170 2700
rect 7090 2640 7170 2660
rect 7490 2700 7570 2720
rect 7490 2660 7510 2700
rect 7550 2660 7570 2700
rect 7490 2640 7570 2660
rect 7690 2700 7770 2720
rect 7690 2660 7710 2700
rect 7750 2660 7770 2700
rect 7690 2640 7770 2660
rect 2010 2560 2450 2610
rect 5750 2600 5790 2640
rect 6150 2600 6190 2640
rect 5550 2580 6410 2600
rect 3790 2440 4230 2490
rect 5550 2540 5630 2580
rect 5670 2540 5710 2580
rect 5750 2540 5790 2580
rect 5830 2540 5870 2580
rect 5910 2540 5950 2580
rect 5990 2540 6030 2580
rect 6070 2540 6110 2580
rect 6150 2540 6190 2580
rect 6230 2540 6270 2580
rect 6310 2540 6350 2580
rect 6390 2540 6410 2580
rect 5550 2520 6410 2540
rect 6490 2580 7370 2600
rect 6490 2540 6510 2580
rect 6550 2540 6590 2580
rect 6630 2540 6670 2580
rect 6710 2540 6750 2580
rect 6790 2540 6830 2580
rect 6870 2540 6910 2580
rect 6950 2540 6990 2580
rect 7030 2540 7070 2580
rect 7110 2540 7150 2580
rect 7190 2540 7230 2580
rect 7270 2540 7310 2580
rect 7350 2540 7370 2580
rect 6490 2520 7370 2540
rect 5550 2480 5590 2520
rect 7310 2480 7350 2520
rect 4580 2460 4720 2480
rect 4580 2420 4590 2460
rect 4630 2420 4670 2460
rect 4710 2420 4720 2460
rect 2010 2320 2450 2370
rect 4580 2360 4720 2420
rect 4580 2320 4590 2360
rect 4630 2320 4670 2360
rect 4710 2320 4720 2360
rect 1890 2200 1970 2210
rect 3790 2200 4230 2250
rect 1890 2190 2010 2200
rect 1890 2150 1910 2190
rect 1950 2150 2010 2190
rect 1890 2130 2010 2150
rect 4580 2260 4720 2320
rect 4580 2220 4590 2260
rect 4630 2220 4670 2260
rect 4710 2220 4720 2260
rect 4580 2160 4720 2220
rect 4580 2120 4590 2160
rect 4630 2120 4670 2160
rect 4710 2120 4720 2160
rect 4580 2060 4720 2120
rect 4580 2020 4590 2060
rect 4630 2020 4670 2060
rect 4710 2020 4720 2060
rect 4580 1960 4720 2020
rect 4580 1920 4590 1960
rect 4630 1920 4670 1960
rect 4710 1920 4720 1960
rect 4580 1860 4720 1920
rect 4580 1820 4590 1860
rect 4630 1820 4670 1860
rect 4710 1820 4720 1860
rect 4580 1760 4720 1820
rect 4580 1720 4590 1760
rect 4630 1720 4670 1760
rect 4710 1720 4720 1760
rect 4580 1700 4720 1720
rect 5540 2460 5600 2480
rect 5540 2420 5550 2460
rect 5590 2420 5600 2460
rect 5540 2360 5600 2420
rect 5540 2320 5550 2360
rect 5590 2320 5600 2360
rect 5540 2260 5600 2320
rect 5540 2220 5550 2260
rect 5590 2220 5600 2260
rect 5540 2160 5600 2220
rect 5540 2120 5550 2160
rect 5590 2120 5600 2160
rect 5540 2060 5600 2120
rect 5540 2020 5550 2060
rect 5590 2020 5600 2060
rect 5540 1960 5600 2020
rect 5540 1920 5550 1960
rect 5590 1920 5600 1960
rect 5540 1860 5600 1920
rect 5540 1820 5550 1860
rect 5590 1820 5600 1860
rect 5540 1760 5600 1820
rect 5540 1720 5550 1760
rect 5590 1720 5600 1760
rect 5540 1700 5600 1720
rect 6420 2460 6480 2480
rect 6420 2420 6430 2460
rect 6470 2420 6480 2460
rect 6420 2360 6480 2420
rect 6420 2320 6430 2360
rect 6470 2320 6480 2360
rect 6420 2260 6480 2320
rect 6420 2220 6430 2260
rect 6470 2220 6480 2260
rect 6420 2160 6480 2220
rect 6420 2120 6430 2160
rect 6470 2120 6480 2160
rect 6420 2060 6480 2120
rect 6420 2020 6430 2060
rect 6470 2020 6480 2060
rect 6420 1960 6480 2020
rect 6420 1920 6430 1960
rect 6470 1920 6480 1960
rect 6420 1860 6480 1920
rect 6420 1820 6430 1860
rect 6470 1820 6480 1860
rect 6420 1760 6480 1820
rect 6420 1720 6430 1760
rect 6470 1720 6480 1760
rect 6420 1700 6480 1720
rect 7300 2460 7360 2480
rect 7300 2420 7310 2460
rect 7350 2420 7360 2460
rect 7300 2360 7360 2420
rect 7300 2320 7310 2360
rect 7350 2320 7360 2360
rect 7300 2260 7360 2320
rect 7300 2220 7310 2260
rect 7350 2220 7360 2260
rect 7300 2160 7360 2220
rect 7300 2120 7310 2160
rect 7350 2120 7360 2160
rect 7300 2060 7360 2120
rect 7300 2020 7310 2060
rect 7350 2020 7360 2060
rect 7300 1960 7360 2020
rect 7300 1920 7310 1960
rect 7350 1920 7360 1960
rect 7300 1860 7360 1920
rect 7300 1820 7310 1860
rect 7350 1820 7360 1860
rect 7300 1760 7360 1820
rect 7300 1720 7310 1760
rect 7350 1720 7360 1760
rect 7300 1700 7360 1720
rect 8180 2460 8320 2480
rect 8180 2420 8190 2460
rect 8230 2420 8270 2460
rect 8310 2420 8320 2460
rect 8180 2360 8320 2420
rect 8180 2320 8190 2360
rect 8230 2320 8270 2360
rect 8310 2320 8320 2360
rect 8180 2260 8320 2320
rect 8180 2220 8190 2260
rect 8230 2220 8270 2260
rect 8310 2220 8320 2260
rect 8180 2160 8320 2220
rect 8180 2120 8190 2160
rect 8230 2120 8270 2160
rect 8310 2120 8320 2160
rect 8180 2060 8320 2120
rect 8180 2020 8190 2060
rect 8230 2020 8270 2060
rect 8310 2020 8320 2060
rect 8180 1960 8320 2020
rect 8180 1920 8190 1960
rect 8230 1920 8270 1960
rect 8310 1920 8320 1960
rect 8180 1860 8320 1920
rect 8180 1820 8190 1860
rect 8230 1820 8270 1860
rect 8310 1820 8320 1860
rect 8180 1760 8320 1820
rect 8180 1720 8190 1760
rect 8230 1720 8270 1760
rect 8310 1720 8320 1760
rect 8180 1700 8320 1720
rect 4670 1660 4710 1700
rect 6430 1660 6470 1700
rect 8190 1660 8230 1700
rect 4650 1640 4730 1660
rect 4650 1600 4670 1640
rect 4710 1600 4730 1640
rect 4650 1580 4730 1600
rect 6410 1640 6490 1660
rect 6410 1600 6430 1640
rect 6470 1600 6490 1640
rect 6410 1580 6490 1600
rect 8170 1640 8250 1660
rect 8170 1600 8190 1640
rect 8230 1600 8250 1640
rect 8170 1580 8250 1600
rect 1190 1410 1270 1430
rect 1190 1370 1210 1410
rect 1250 1370 1270 1410
rect 1190 1320 1270 1370
rect 1410 1410 1490 1430
rect 1410 1370 1430 1410
rect 1470 1370 1490 1410
rect 1410 1320 1490 1370
rect 10 1279 9470 1320
rect 10 1256 1506 1279
rect 10 1222 1410 1256
rect 1444 1245 1506 1256
rect 1540 1245 1596 1279
rect 1630 1245 1686 1279
rect 1720 1245 1776 1279
rect 1810 1245 1866 1279
rect 1900 1245 1956 1279
rect 1990 1245 2046 1279
rect 2080 1245 2136 1279
rect 2170 1245 2226 1279
rect 2260 1245 2316 1279
rect 2350 1245 2406 1279
rect 2440 1245 2496 1279
rect 2530 1256 2866 1279
rect 2530 1245 2597 1256
rect 1444 1222 2597 1245
rect 2631 1222 2770 1256
rect 2804 1245 2866 1256
rect 2900 1245 2956 1279
rect 2990 1245 3046 1279
rect 3080 1245 3136 1279
rect 3170 1245 3226 1279
rect 3260 1245 3316 1279
rect 3350 1245 3406 1279
rect 3440 1245 3496 1279
rect 3530 1245 3586 1279
rect 3620 1245 3676 1279
rect 3710 1245 3766 1279
rect 3800 1245 3856 1279
rect 3890 1256 4226 1279
rect 3890 1245 3957 1256
rect 2804 1222 3957 1245
rect 3991 1222 4130 1256
rect 4164 1245 4226 1256
rect 4260 1245 4316 1279
rect 4350 1245 4406 1279
rect 4440 1245 4496 1279
rect 4530 1245 4586 1279
rect 4620 1245 4676 1279
rect 4710 1245 4766 1279
rect 4800 1245 4856 1279
rect 4890 1245 4946 1279
rect 4980 1245 5036 1279
rect 5070 1245 5126 1279
rect 5160 1245 5216 1279
rect 5250 1256 5586 1279
rect 5250 1245 5317 1256
rect 4164 1222 5317 1245
rect 5351 1222 5490 1256
rect 5524 1245 5586 1256
rect 5620 1245 5676 1279
rect 5710 1245 5766 1279
rect 5800 1245 5856 1279
rect 5890 1245 5946 1279
rect 5980 1245 6036 1279
rect 6070 1245 6126 1279
rect 6160 1245 6216 1279
rect 6250 1245 6306 1279
rect 6340 1245 6396 1279
rect 6430 1245 6486 1279
rect 6520 1245 6576 1279
rect 6610 1256 6946 1279
rect 6610 1245 6677 1256
rect 5524 1222 6677 1245
rect 6711 1222 6850 1256
rect 6884 1245 6946 1256
rect 6980 1245 7036 1279
rect 7070 1245 7126 1279
rect 7160 1245 7216 1279
rect 7250 1245 7306 1279
rect 7340 1245 7396 1279
rect 7430 1245 7486 1279
rect 7520 1245 7576 1279
rect 7610 1245 7666 1279
rect 7700 1245 7756 1279
rect 7790 1245 7846 1279
rect 7880 1245 7936 1279
rect 7970 1256 8306 1279
rect 7970 1245 8037 1256
rect 6884 1222 8037 1245
rect 8071 1222 8210 1256
rect 8244 1245 8306 1256
rect 8340 1245 8396 1279
rect 8430 1245 8486 1279
rect 8520 1245 8576 1279
rect 8610 1245 8666 1279
rect 8700 1245 8756 1279
rect 8790 1245 8846 1279
rect 8880 1245 8936 1279
rect 8970 1245 9026 1279
rect 9060 1245 9116 1279
rect 9150 1245 9206 1279
rect 9240 1245 9296 1279
rect 9330 1256 9470 1279
rect 9330 1245 9397 1256
rect 8244 1222 9397 1245
rect 9431 1222 9470 1256
rect 10 1166 9470 1222
rect 10 1132 1410 1166
rect 1444 1132 2597 1166
rect 2631 1132 2770 1166
rect 2804 1132 3957 1166
rect 3991 1132 4130 1166
rect 4164 1132 5317 1166
rect 5351 1132 5490 1166
rect 5524 1132 6677 1166
rect 6711 1132 6850 1166
rect 6884 1132 8037 1166
rect 8071 1132 8210 1166
rect 8244 1132 9397 1166
rect 9431 1132 9470 1166
rect 10 1098 1670 1132
rect 1704 1098 1760 1132
rect 1794 1098 1850 1132
rect 1884 1098 1940 1132
rect 1974 1098 2030 1132
rect 2064 1098 2120 1132
rect 2154 1098 2210 1132
rect 2244 1098 2300 1132
rect 2334 1098 2390 1132
rect 2424 1098 3030 1132
rect 3064 1098 3120 1132
rect 3154 1098 3210 1132
rect 3244 1098 3300 1132
rect 3334 1098 3390 1132
rect 3424 1098 3480 1132
rect 3514 1098 3570 1132
rect 3604 1098 3660 1132
rect 3694 1098 3750 1132
rect 3784 1098 4390 1132
rect 4424 1098 4480 1132
rect 4514 1098 4570 1132
rect 4604 1098 4660 1132
rect 4694 1098 4750 1132
rect 4784 1098 4840 1132
rect 4874 1098 4930 1132
rect 4964 1098 5020 1132
rect 5054 1098 5110 1132
rect 5144 1098 5750 1132
rect 5784 1098 5840 1132
rect 5874 1098 5930 1132
rect 5964 1098 6020 1132
rect 6054 1098 6110 1132
rect 6144 1098 6200 1132
rect 6234 1098 6290 1132
rect 6324 1098 6380 1132
rect 6414 1098 6470 1132
rect 6504 1098 7110 1132
rect 7144 1098 7200 1132
rect 7234 1098 7290 1132
rect 7324 1098 7380 1132
rect 7414 1098 7470 1132
rect 7504 1098 7560 1132
rect 7594 1098 7650 1132
rect 7684 1098 7740 1132
rect 7774 1098 7830 1132
rect 7864 1098 8470 1132
rect 8504 1098 8560 1132
rect 8594 1098 8650 1132
rect 8684 1098 8740 1132
rect 8774 1098 8830 1132
rect 8864 1098 8920 1132
rect 8954 1098 9010 1132
rect 9044 1098 9100 1132
rect 9134 1098 9190 1132
rect 9224 1098 9470 1132
rect 10 1079 9470 1098
rect 10 1076 1620 1079
rect 10 1070 1410 1076
rect 10 270 260 1070
rect 1060 1042 1410 1070
rect 1444 1075 1620 1076
rect 1444 1042 1558 1075
rect 1060 1041 1558 1042
rect 1592 1041 1620 1075
rect 1060 986 1620 1041
rect 2420 1076 2980 1079
rect 2420 1056 2597 1076
rect 2420 1022 2448 1056
rect 2482 1042 2597 1056
rect 2631 1042 2770 1076
rect 2804 1075 2980 1076
rect 2804 1042 2918 1075
rect 2482 1041 2918 1042
rect 2952 1041 2980 1075
rect 2482 1022 2980 1041
rect 1060 952 1410 986
rect 1444 985 1620 986
rect 1444 952 1558 985
rect 1060 951 1558 952
rect 1592 951 1620 985
rect 1060 896 1620 951
rect 1060 862 1410 896
rect 1444 895 1620 896
rect 1444 862 1558 895
rect 1060 861 1558 862
rect 1592 861 1620 895
rect 1060 806 1620 861
rect 1060 772 1410 806
rect 1444 805 1620 806
rect 1444 772 1558 805
rect 1060 771 1558 772
rect 1592 771 1620 805
rect 1060 716 1620 771
rect 1060 682 1410 716
rect 1444 715 1620 716
rect 1444 682 1558 715
rect 1060 681 1558 682
rect 1592 681 1620 715
rect 1060 626 1620 681
rect 1060 592 1410 626
rect 1444 625 1620 626
rect 1444 592 1558 625
rect 1060 591 1558 592
rect 1592 591 1620 625
rect 1060 536 1620 591
rect 1060 502 1410 536
rect 1444 535 1620 536
rect 1444 502 1558 535
rect 1060 501 1558 502
rect 1592 501 1620 535
rect 1060 446 1620 501
rect 1060 412 1410 446
rect 1444 445 1620 446
rect 1444 412 1558 445
rect 1060 411 1558 412
rect 1592 411 1620 445
rect 1060 356 1620 411
rect 1060 322 1410 356
rect 1444 355 1620 356
rect 1444 322 1558 355
rect 1060 321 1558 322
rect 1592 321 1620 355
rect 1673 958 2367 1017
rect 1673 924 1734 958
rect 1768 930 1824 958
rect 1858 930 1914 958
rect 1948 930 2004 958
rect 1780 924 1824 930
rect 1880 924 1914 930
rect 1980 924 2004 930
rect 2038 930 2094 958
rect 2038 924 2046 930
rect 1673 896 1746 924
rect 1780 896 1846 924
rect 1880 896 1946 924
rect 1980 896 2046 924
rect 2080 924 2094 930
rect 2128 930 2184 958
rect 2128 924 2146 930
rect 2080 896 2146 924
rect 2180 924 2184 930
rect 2218 930 2274 958
rect 2218 924 2246 930
rect 2308 924 2367 958
rect 2180 896 2246 924
rect 2280 896 2367 924
rect 1673 868 2367 896
rect 1673 834 1734 868
rect 1768 834 1824 868
rect 1858 834 1914 868
rect 1948 834 2004 868
rect 2038 834 2094 868
rect 2128 834 2184 868
rect 2218 834 2274 868
rect 2308 834 2367 868
rect 1673 830 2367 834
rect 1673 796 1746 830
rect 1780 796 1846 830
rect 1880 796 1946 830
rect 1980 796 2046 830
rect 2080 796 2146 830
rect 2180 796 2246 830
rect 2280 796 2367 830
rect 1673 778 2367 796
rect 1673 744 1734 778
rect 1768 744 1824 778
rect 1858 744 1914 778
rect 1948 744 2004 778
rect 2038 744 2094 778
rect 2128 744 2184 778
rect 2218 744 2274 778
rect 2308 744 2367 778
rect 1673 730 2367 744
rect 1673 696 1746 730
rect 1780 696 1846 730
rect 1880 696 1946 730
rect 1980 696 2046 730
rect 2080 696 2146 730
rect 2180 696 2246 730
rect 2280 696 2367 730
rect 1673 688 2367 696
rect 1673 654 1734 688
rect 1768 654 1824 688
rect 1858 654 1914 688
rect 1948 654 2004 688
rect 2038 654 2094 688
rect 2128 654 2184 688
rect 2218 654 2274 688
rect 2308 654 2367 688
rect 1673 630 2367 654
rect 1673 598 1746 630
rect 1780 598 1846 630
rect 1880 598 1946 630
rect 1980 598 2046 630
rect 1673 564 1734 598
rect 1780 596 1824 598
rect 1880 596 1914 598
rect 1980 596 2004 598
rect 1768 564 1824 596
rect 1858 564 1914 596
rect 1948 564 2004 596
rect 2038 596 2046 598
rect 2080 598 2146 630
rect 2080 596 2094 598
rect 2038 564 2094 596
rect 2128 596 2146 598
rect 2180 598 2246 630
rect 2280 598 2367 630
rect 2180 596 2184 598
rect 2128 564 2184 596
rect 2218 596 2246 598
rect 2218 564 2274 596
rect 2308 564 2367 598
rect 1673 530 2367 564
rect 1673 508 1746 530
rect 1780 508 1846 530
rect 1880 508 1946 530
rect 1980 508 2046 530
rect 1673 474 1734 508
rect 1780 496 1824 508
rect 1880 496 1914 508
rect 1980 496 2004 508
rect 1768 474 1824 496
rect 1858 474 1914 496
rect 1948 474 2004 496
rect 2038 496 2046 508
rect 2080 508 2146 530
rect 2080 496 2094 508
rect 2038 474 2094 496
rect 2128 496 2146 508
rect 2180 508 2246 530
rect 2280 508 2367 530
rect 2180 496 2184 508
rect 2128 474 2184 496
rect 2218 496 2246 508
rect 2218 474 2274 496
rect 2308 474 2367 508
rect 1673 430 2367 474
rect 1673 418 1746 430
rect 1780 418 1846 430
rect 1880 418 1946 430
rect 1980 418 2046 430
rect 1673 384 1734 418
rect 1780 396 1824 418
rect 1880 396 1914 418
rect 1980 396 2004 418
rect 1768 384 1824 396
rect 1858 384 1914 396
rect 1948 384 2004 396
rect 2038 396 2046 418
rect 2080 418 2146 430
rect 2080 396 2094 418
rect 2038 384 2094 396
rect 2128 396 2146 418
rect 2180 418 2246 430
rect 2280 418 2367 430
rect 2180 396 2184 418
rect 2128 384 2184 396
rect 2218 396 2246 418
rect 2218 384 2274 396
rect 2308 384 2367 418
rect 1673 323 2367 384
rect 2420 986 2980 1022
rect 3780 1076 4340 1079
rect 3780 1056 3957 1076
rect 3780 1022 3808 1056
rect 3842 1042 3957 1056
rect 3991 1042 4130 1076
rect 4164 1075 4340 1076
rect 4164 1042 4278 1075
rect 3842 1041 4278 1042
rect 4312 1041 4340 1075
rect 3842 1022 4340 1041
rect 2420 966 2597 986
rect 2420 932 2448 966
rect 2482 952 2597 966
rect 2631 952 2770 986
rect 2804 985 2980 986
rect 2804 952 2918 985
rect 2482 951 2918 952
rect 2952 951 2980 985
rect 2482 932 2980 951
rect 2420 896 2980 932
rect 2420 876 2597 896
rect 2420 842 2448 876
rect 2482 862 2597 876
rect 2631 862 2770 896
rect 2804 895 2980 896
rect 2804 862 2918 895
rect 2482 861 2918 862
rect 2952 861 2980 895
rect 2482 842 2980 861
rect 2420 806 2980 842
rect 2420 786 2597 806
rect 2420 752 2448 786
rect 2482 772 2597 786
rect 2631 772 2770 806
rect 2804 805 2980 806
rect 2804 772 2918 805
rect 2482 771 2918 772
rect 2952 771 2980 805
rect 2482 752 2980 771
rect 2420 716 2980 752
rect 2420 696 2597 716
rect 2420 662 2448 696
rect 2482 682 2597 696
rect 2631 682 2770 716
rect 2804 715 2980 716
rect 2804 682 2918 715
rect 2482 681 2918 682
rect 2952 681 2980 715
rect 2482 662 2980 681
rect 2420 626 2980 662
rect 2420 606 2597 626
rect 2420 572 2448 606
rect 2482 592 2597 606
rect 2631 592 2770 626
rect 2804 625 2980 626
rect 2804 592 2918 625
rect 2482 591 2918 592
rect 2952 591 2980 625
rect 2482 572 2980 591
rect 2420 536 2980 572
rect 2420 516 2597 536
rect 2420 482 2448 516
rect 2482 502 2597 516
rect 2631 502 2770 536
rect 2804 535 2980 536
rect 2804 502 2918 535
rect 2482 501 2918 502
rect 2952 501 2980 535
rect 2482 482 2980 501
rect 2420 446 2980 482
rect 2420 426 2597 446
rect 2420 392 2448 426
rect 2482 412 2597 426
rect 2631 412 2770 446
rect 2804 445 2980 446
rect 2804 412 2918 445
rect 2482 411 2918 412
rect 2952 411 2980 445
rect 2482 392 2980 411
rect 2420 356 2980 392
rect 2420 336 2597 356
rect 1060 270 1620 321
rect 2420 302 2448 336
rect 2482 322 2597 336
rect 2631 322 2770 356
rect 2804 355 2980 356
rect 2804 322 2918 355
rect 2482 321 2918 322
rect 2952 321 2980 355
rect 3033 958 3727 1017
rect 3033 924 3094 958
rect 3128 930 3184 958
rect 3218 930 3274 958
rect 3308 930 3364 958
rect 3140 924 3184 930
rect 3240 924 3274 930
rect 3340 924 3364 930
rect 3398 930 3454 958
rect 3398 924 3406 930
rect 3033 896 3106 924
rect 3140 896 3206 924
rect 3240 896 3306 924
rect 3340 896 3406 924
rect 3440 924 3454 930
rect 3488 930 3544 958
rect 3488 924 3506 930
rect 3440 896 3506 924
rect 3540 924 3544 930
rect 3578 930 3634 958
rect 3578 924 3606 930
rect 3668 924 3727 958
rect 3540 896 3606 924
rect 3640 896 3727 924
rect 3033 868 3727 896
rect 3033 834 3094 868
rect 3128 834 3184 868
rect 3218 834 3274 868
rect 3308 834 3364 868
rect 3398 834 3454 868
rect 3488 834 3544 868
rect 3578 834 3634 868
rect 3668 834 3727 868
rect 3033 830 3727 834
rect 3033 796 3106 830
rect 3140 796 3206 830
rect 3240 796 3306 830
rect 3340 796 3406 830
rect 3440 796 3506 830
rect 3540 796 3606 830
rect 3640 796 3727 830
rect 3033 778 3727 796
rect 3033 744 3094 778
rect 3128 744 3184 778
rect 3218 744 3274 778
rect 3308 744 3364 778
rect 3398 744 3454 778
rect 3488 744 3544 778
rect 3578 744 3634 778
rect 3668 744 3727 778
rect 3033 730 3727 744
rect 3033 696 3106 730
rect 3140 696 3206 730
rect 3240 696 3306 730
rect 3340 696 3406 730
rect 3440 696 3506 730
rect 3540 696 3606 730
rect 3640 696 3727 730
rect 3033 688 3727 696
rect 3033 654 3094 688
rect 3128 654 3184 688
rect 3218 654 3274 688
rect 3308 654 3364 688
rect 3398 654 3454 688
rect 3488 654 3544 688
rect 3578 654 3634 688
rect 3668 654 3727 688
rect 3033 630 3727 654
rect 3033 598 3106 630
rect 3140 598 3206 630
rect 3240 598 3306 630
rect 3340 598 3406 630
rect 3033 564 3094 598
rect 3140 596 3184 598
rect 3240 596 3274 598
rect 3340 596 3364 598
rect 3128 564 3184 596
rect 3218 564 3274 596
rect 3308 564 3364 596
rect 3398 596 3406 598
rect 3440 598 3506 630
rect 3440 596 3454 598
rect 3398 564 3454 596
rect 3488 596 3506 598
rect 3540 598 3606 630
rect 3640 598 3727 630
rect 3540 596 3544 598
rect 3488 564 3544 596
rect 3578 596 3606 598
rect 3578 564 3634 596
rect 3668 564 3727 598
rect 3033 530 3727 564
rect 3033 508 3106 530
rect 3140 508 3206 530
rect 3240 508 3306 530
rect 3340 508 3406 530
rect 3033 474 3094 508
rect 3140 496 3184 508
rect 3240 496 3274 508
rect 3340 496 3364 508
rect 3128 474 3184 496
rect 3218 474 3274 496
rect 3308 474 3364 496
rect 3398 496 3406 508
rect 3440 508 3506 530
rect 3440 496 3454 508
rect 3398 474 3454 496
rect 3488 496 3506 508
rect 3540 508 3606 530
rect 3640 508 3727 530
rect 3540 496 3544 508
rect 3488 474 3544 496
rect 3578 496 3606 508
rect 3578 474 3634 496
rect 3668 474 3727 508
rect 3033 430 3727 474
rect 3033 418 3106 430
rect 3140 418 3206 430
rect 3240 418 3306 430
rect 3340 418 3406 430
rect 3033 384 3094 418
rect 3140 396 3184 418
rect 3240 396 3274 418
rect 3340 396 3364 418
rect 3128 384 3184 396
rect 3218 384 3274 396
rect 3308 384 3364 396
rect 3398 396 3406 418
rect 3440 418 3506 430
rect 3440 396 3454 418
rect 3398 384 3454 396
rect 3488 396 3506 418
rect 3540 418 3606 430
rect 3640 418 3727 430
rect 3540 396 3544 418
rect 3488 384 3544 396
rect 3578 396 3606 418
rect 3578 384 3634 396
rect 3668 384 3727 418
rect 3033 323 3727 384
rect 3780 986 4340 1022
rect 5140 1076 5700 1079
rect 5140 1056 5317 1076
rect 5140 1022 5168 1056
rect 5202 1042 5317 1056
rect 5351 1042 5490 1076
rect 5524 1075 5700 1076
rect 5524 1042 5638 1075
rect 5202 1041 5638 1042
rect 5672 1041 5700 1075
rect 5202 1022 5700 1041
rect 3780 966 3957 986
rect 3780 932 3808 966
rect 3842 952 3957 966
rect 3991 952 4130 986
rect 4164 985 4340 986
rect 4164 952 4278 985
rect 3842 951 4278 952
rect 4312 951 4340 985
rect 3842 932 4340 951
rect 3780 896 4340 932
rect 3780 876 3957 896
rect 3780 842 3808 876
rect 3842 862 3957 876
rect 3991 862 4130 896
rect 4164 895 4340 896
rect 4164 862 4278 895
rect 3842 861 4278 862
rect 4312 861 4340 895
rect 3842 842 4340 861
rect 3780 806 4340 842
rect 3780 786 3957 806
rect 3780 752 3808 786
rect 3842 772 3957 786
rect 3991 772 4130 806
rect 4164 805 4340 806
rect 4164 772 4278 805
rect 3842 771 4278 772
rect 4312 771 4340 805
rect 3842 752 4340 771
rect 3780 716 4340 752
rect 3780 696 3957 716
rect 3780 662 3808 696
rect 3842 682 3957 696
rect 3991 682 4130 716
rect 4164 715 4340 716
rect 4164 682 4278 715
rect 3842 681 4278 682
rect 4312 681 4340 715
rect 3842 662 4340 681
rect 3780 626 4340 662
rect 3780 606 3957 626
rect 3780 572 3808 606
rect 3842 592 3957 606
rect 3991 592 4130 626
rect 4164 625 4340 626
rect 4164 592 4278 625
rect 3842 591 4278 592
rect 4312 591 4340 625
rect 3842 572 4340 591
rect 3780 536 4340 572
rect 3780 516 3957 536
rect 3780 482 3808 516
rect 3842 502 3957 516
rect 3991 502 4130 536
rect 4164 535 4340 536
rect 4164 502 4278 535
rect 3842 501 4278 502
rect 4312 501 4340 535
rect 3842 482 4340 501
rect 3780 446 4340 482
rect 3780 426 3957 446
rect 3780 392 3808 426
rect 3842 412 3957 426
rect 3991 412 4130 446
rect 4164 445 4340 446
rect 4164 412 4278 445
rect 3842 411 4278 412
rect 4312 411 4340 445
rect 3842 392 4340 411
rect 3780 356 4340 392
rect 3780 336 3957 356
rect 2482 302 2980 321
rect 2420 270 2980 302
rect 3780 302 3808 336
rect 3842 322 3957 336
rect 3991 322 4130 356
rect 4164 355 4340 356
rect 4164 322 4278 355
rect 3842 321 4278 322
rect 4312 321 4340 355
rect 4393 958 5087 1017
rect 4393 924 4454 958
rect 4488 930 4544 958
rect 4578 930 4634 958
rect 4668 930 4724 958
rect 4500 924 4544 930
rect 4600 924 4634 930
rect 4700 924 4724 930
rect 4758 930 4814 958
rect 4758 924 4766 930
rect 4393 896 4466 924
rect 4500 896 4566 924
rect 4600 896 4666 924
rect 4700 896 4766 924
rect 4800 924 4814 930
rect 4848 930 4904 958
rect 4848 924 4866 930
rect 4800 896 4866 924
rect 4900 924 4904 930
rect 4938 930 4994 958
rect 4938 924 4966 930
rect 5028 924 5087 958
rect 4900 896 4966 924
rect 5000 896 5087 924
rect 4393 868 5087 896
rect 4393 834 4454 868
rect 4488 834 4544 868
rect 4578 834 4634 868
rect 4668 834 4724 868
rect 4758 834 4814 868
rect 4848 834 4904 868
rect 4938 834 4994 868
rect 5028 834 5087 868
rect 4393 830 5087 834
rect 4393 796 4466 830
rect 4500 796 4566 830
rect 4600 796 4666 830
rect 4700 796 4766 830
rect 4800 796 4866 830
rect 4900 796 4966 830
rect 5000 796 5087 830
rect 4393 778 5087 796
rect 4393 744 4454 778
rect 4488 744 4544 778
rect 4578 744 4634 778
rect 4668 744 4724 778
rect 4758 744 4814 778
rect 4848 744 4904 778
rect 4938 744 4994 778
rect 5028 744 5087 778
rect 4393 730 5087 744
rect 4393 696 4466 730
rect 4500 696 4566 730
rect 4600 696 4666 730
rect 4700 696 4766 730
rect 4800 696 4866 730
rect 4900 696 4966 730
rect 5000 696 5087 730
rect 4393 688 5087 696
rect 4393 654 4454 688
rect 4488 654 4544 688
rect 4578 654 4634 688
rect 4668 654 4724 688
rect 4758 654 4814 688
rect 4848 654 4904 688
rect 4938 654 4994 688
rect 5028 654 5087 688
rect 4393 630 5087 654
rect 4393 598 4466 630
rect 4500 598 4566 630
rect 4600 598 4666 630
rect 4700 598 4766 630
rect 4393 564 4454 598
rect 4500 596 4544 598
rect 4600 596 4634 598
rect 4700 596 4724 598
rect 4488 564 4544 596
rect 4578 564 4634 596
rect 4668 564 4724 596
rect 4758 596 4766 598
rect 4800 598 4866 630
rect 4800 596 4814 598
rect 4758 564 4814 596
rect 4848 596 4866 598
rect 4900 598 4966 630
rect 5000 598 5087 630
rect 4900 596 4904 598
rect 4848 564 4904 596
rect 4938 596 4966 598
rect 4938 564 4994 596
rect 5028 564 5087 598
rect 4393 530 5087 564
rect 4393 508 4466 530
rect 4500 508 4566 530
rect 4600 508 4666 530
rect 4700 508 4766 530
rect 4393 474 4454 508
rect 4500 496 4544 508
rect 4600 496 4634 508
rect 4700 496 4724 508
rect 4488 474 4544 496
rect 4578 474 4634 496
rect 4668 474 4724 496
rect 4758 496 4766 508
rect 4800 508 4866 530
rect 4800 496 4814 508
rect 4758 474 4814 496
rect 4848 496 4866 508
rect 4900 508 4966 530
rect 5000 508 5087 530
rect 4900 496 4904 508
rect 4848 474 4904 496
rect 4938 496 4966 508
rect 4938 474 4994 496
rect 5028 474 5087 508
rect 4393 430 5087 474
rect 4393 418 4466 430
rect 4500 418 4566 430
rect 4600 418 4666 430
rect 4700 418 4766 430
rect 4393 384 4454 418
rect 4500 396 4544 418
rect 4600 396 4634 418
rect 4700 396 4724 418
rect 4488 384 4544 396
rect 4578 384 4634 396
rect 4668 384 4724 396
rect 4758 396 4766 418
rect 4800 418 4866 430
rect 4800 396 4814 418
rect 4758 384 4814 396
rect 4848 396 4866 418
rect 4900 418 4966 430
rect 5000 418 5087 430
rect 4900 396 4904 418
rect 4848 384 4904 396
rect 4938 396 4966 418
rect 4938 384 4994 396
rect 5028 384 5087 418
rect 4393 323 5087 384
rect 5140 986 5700 1022
rect 6500 1076 7060 1079
rect 6500 1056 6677 1076
rect 6500 1022 6528 1056
rect 6562 1042 6677 1056
rect 6711 1042 6850 1076
rect 6884 1075 7060 1076
rect 6884 1042 6998 1075
rect 6562 1041 6998 1042
rect 7032 1041 7060 1075
rect 6562 1022 7060 1041
rect 5140 966 5317 986
rect 5140 932 5168 966
rect 5202 952 5317 966
rect 5351 952 5490 986
rect 5524 985 5700 986
rect 5524 952 5638 985
rect 5202 951 5638 952
rect 5672 951 5700 985
rect 5202 932 5700 951
rect 5140 896 5700 932
rect 5140 876 5317 896
rect 5140 842 5168 876
rect 5202 862 5317 876
rect 5351 862 5490 896
rect 5524 895 5700 896
rect 5524 862 5638 895
rect 5202 861 5638 862
rect 5672 861 5700 895
rect 5202 842 5700 861
rect 5140 806 5700 842
rect 5140 786 5317 806
rect 5140 752 5168 786
rect 5202 772 5317 786
rect 5351 772 5490 806
rect 5524 805 5700 806
rect 5524 772 5638 805
rect 5202 771 5638 772
rect 5672 771 5700 805
rect 5202 752 5700 771
rect 5140 716 5700 752
rect 5140 696 5317 716
rect 5140 662 5168 696
rect 5202 682 5317 696
rect 5351 682 5490 716
rect 5524 715 5700 716
rect 5524 682 5638 715
rect 5202 681 5638 682
rect 5672 681 5700 715
rect 5202 662 5700 681
rect 5140 626 5700 662
rect 5140 606 5317 626
rect 5140 572 5168 606
rect 5202 592 5317 606
rect 5351 592 5490 626
rect 5524 625 5700 626
rect 5524 592 5638 625
rect 5202 591 5638 592
rect 5672 591 5700 625
rect 5202 572 5700 591
rect 5140 536 5700 572
rect 5140 516 5317 536
rect 5140 482 5168 516
rect 5202 502 5317 516
rect 5351 502 5490 536
rect 5524 535 5700 536
rect 5524 502 5638 535
rect 5202 501 5638 502
rect 5672 501 5700 535
rect 5202 482 5700 501
rect 5140 446 5700 482
rect 5140 426 5317 446
rect 5140 392 5168 426
rect 5202 412 5317 426
rect 5351 412 5490 446
rect 5524 445 5700 446
rect 5524 412 5638 445
rect 5202 411 5638 412
rect 5672 411 5700 445
rect 5202 392 5700 411
rect 5140 356 5700 392
rect 5140 336 5317 356
rect 3842 302 4340 321
rect 3780 270 4340 302
rect 5140 302 5168 336
rect 5202 322 5317 336
rect 5351 322 5490 356
rect 5524 355 5700 356
rect 5524 322 5638 355
rect 5202 321 5638 322
rect 5672 321 5700 355
rect 5753 958 6447 1017
rect 5753 924 5814 958
rect 5848 930 5904 958
rect 5938 930 5994 958
rect 6028 930 6084 958
rect 5860 924 5904 930
rect 5960 924 5994 930
rect 6060 924 6084 930
rect 6118 930 6174 958
rect 6118 924 6126 930
rect 5753 896 5826 924
rect 5860 896 5926 924
rect 5960 896 6026 924
rect 6060 896 6126 924
rect 6160 924 6174 930
rect 6208 930 6264 958
rect 6208 924 6226 930
rect 6160 896 6226 924
rect 6260 924 6264 930
rect 6298 930 6354 958
rect 6298 924 6326 930
rect 6388 924 6447 958
rect 6260 896 6326 924
rect 6360 896 6447 924
rect 5753 868 6447 896
rect 5753 834 5814 868
rect 5848 834 5904 868
rect 5938 834 5994 868
rect 6028 834 6084 868
rect 6118 834 6174 868
rect 6208 834 6264 868
rect 6298 834 6354 868
rect 6388 834 6447 868
rect 5753 830 6447 834
rect 5753 796 5826 830
rect 5860 796 5926 830
rect 5960 796 6026 830
rect 6060 796 6126 830
rect 6160 796 6226 830
rect 6260 796 6326 830
rect 6360 796 6447 830
rect 5753 778 6447 796
rect 5753 744 5814 778
rect 5848 744 5904 778
rect 5938 744 5994 778
rect 6028 744 6084 778
rect 6118 744 6174 778
rect 6208 744 6264 778
rect 6298 744 6354 778
rect 6388 744 6447 778
rect 5753 730 6447 744
rect 5753 696 5826 730
rect 5860 696 5926 730
rect 5960 696 6026 730
rect 6060 696 6126 730
rect 6160 696 6226 730
rect 6260 696 6326 730
rect 6360 696 6447 730
rect 5753 688 6447 696
rect 5753 654 5814 688
rect 5848 654 5904 688
rect 5938 654 5994 688
rect 6028 654 6084 688
rect 6118 654 6174 688
rect 6208 654 6264 688
rect 6298 654 6354 688
rect 6388 654 6447 688
rect 5753 630 6447 654
rect 5753 598 5826 630
rect 5860 598 5926 630
rect 5960 598 6026 630
rect 6060 598 6126 630
rect 5753 564 5814 598
rect 5860 596 5904 598
rect 5960 596 5994 598
rect 6060 596 6084 598
rect 5848 564 5904 596
rect 5938 564 5994 596
rect 6028 564 6084 596
rect 6118 596 6126 598
rect 6160 598 6226 630
rect 6160 596 6174 598
rect 6118 564 6174 596
rect 6208 596 6226 598
rect 6260 598 6326 630
rect 6360 598 6447 630
rect 6260 596 6264 598
rect 6208 564 6264 596
rect 6298 596 6326 598
rect 6298 564 6354 596
rect 6388 564 6447 598
rect 5753 530 6447 564
rect 5753 508 5826 530
rect 5860 508 5926 530
rect 5960 508 6026 530
rect 6060 508 6126 530
rect 5753 474 5814 508
rect 5860 496 5904 508
rect 5960 496 5994 508
rect 6060 496 6084 508
rect 5848 474 5904 496
rect 5938 474 5994 496
rect 6028 474 6084 496
rect 6118 496 6126 508
rect 6160 508 6226 530
rect 6160 496 6174 508
rect 6118 474 6174 496
rect 6208 496 6226 508
rect 6260 508 6326 530
rect 6360 508 6447 530
rect 6260 496 6264 508
rect 6208 474 6264 496
rect 6298 496 6326 508
rect 6298 474 6354 496
rect 6388 474 6447 508
rect 5753 430 6447 474
rect 5753 418 5826 430
rect 5860 418 5926 430
rect 5960 418 6026 430
rect 6060 418 6126 430
rect 5753 384 5814 418
rect 5860 396 5904 418
rect 5960 396 5994 418
rect 6060 396 6084 418
rect 5848 384 5904 396
rect 5938 384 5994 396
rect 6028 384 6084 396
rect 6118 396 6126 418
rect 6160 418 6226 430
rect 6160 396 6174 418
rect 6118 384 6174 396
rect 6208 396 6226 418
rect 6260 418 6326 430
rect 6360 418 6447 430
rect 6260 396 6264 418
rect 6208 384 6264 396
rect 6298 396 6326 418
rect 6298 384 6354 396
rect 6388 384 6447 418
rect 5753 323 6447 384
rect 6500 986 7060 1022
rect 7860 1076 8420 1079
rect 7860 1056 8037 1076
rect 7860 1022 7888 1056
rect 7922 1042 8037 1056
rect 8071 1042 8210 1076
rect 8244 1075 8420 1076
rect 8244 1042 8358 1075
rect 7922 1041 8358 1042
rect 8392 1041 8420 1075
rect 7922 1022 8420 1041
rect 6500 966 6677 986
rect 6500 932 6528 966
rect 6562 952 6677 966
rect 6711 952 6850 986
rect 6884 985 7060 986
rect 6884 952 6998 985
rect 6562 951 6998 952
rect 7032 951 7060 985
rect 6562 932 7060 951
rect 6500 896 7060 932
rect 6500 876 6677 896
rect 6500 842 6528 876
rect 6562 862 6677 876
rect 6711 862 6850 896
rect 6884 895 7060 896
rect 6884 862 6998 895
rect 6562 861 6998 862
rect 7032 861 7060 895
rect 6562 842 7060 861
rect 6500 806 7060 842
rect 6500 786 6677 806
rect 6500 752 6528 786
rect 6562 772 6677 786
rect 6711 772 6850 806
rect 6884 805 7060 806
rect 6884 772 6998 805
rect 6562 771 6998 772
rect 7032 771 7060 805
rect 6562 752 7060 771
rect 6500 716 7060 752
rect 6500 696 6677 716
rect 6500 662 6528 696
rect 6562 682 6677 696
rect 6711 682 6850 716
rect 6884 715 7060 716
rect 6884 682 6998 715
rect 6562 681 6998 682
rect 7032 681 7060 715
rect 6562 662 7060 681
rect 6500 626 7060 662
rect 6500 606 6677 626
rect 6500 572 6528 606
rect 6562 592 6677 606
rect 6711 592 6850 626
rect 6884 625 7060 626
rect 6884 592 6998 625
rect 6562 591 6998 592
rect 7032 591 7060 625
rect 6562 572 7060 591
rect 6500 536 7060 572
rect 6500 516 6677 536
rect 6500 482 6528 516
rect 6562 502 6677 516
rect 6711 502 6850 536
rect 6884 535 7060 536
rect 6884 502 6998 535
rect 6562 501 6998 502
rect 7032 501 7060 535
rect 6562 482 7060 501
rect 6500 446 7060 482
rect 6500 426 6677 446
rect 6500 392 6528 426
rect 6562 412 6677 426
rect 6711 412 6850 446
rect 6884 445 7060 446
rect 6884 412 6998 445
rect 6562 411 6998 412
rect 7032 411 7060 445
rect 6562 392 7060 411
rect 6500 356 7060 392
rect 6500 336 6677 356
rect 5202 302 5700 321
rect 5140 270 5700 302
rect 6500 302 6528 336
rect 6562 322 6677 336
rect 6711 322 6850 356
rect 6884 355 7060 356
rect 6884 322 6998 355
rect 6562 321 6998 322
rect 7032 321 7060 355
rect 7113 958 7807 1017
rect 7113 924 7174 958
rect 7208 930 7264 958
rect 7298 930 7354 958
rect 7388 930 7444 958
rect 7220 924 7264 930
rect 7320 924 7354 930
rect 7420 924 7444 930
rect 7478 930 7534 958
rect 7478 924 7486 930
rect 7113 896 7186 924
rect 7220 896 7286 924
rect 7320 896 7386 924
rect 7420 896 7486 924
rect 7520 924 7534 930
rect 7568 930 7624 958
rect 7568 924 7586 930
rect 7520 896 7586 924
rect 7620 924 7624 930
rect 7658 930 7714 958
rect 7658 924 7686 930
rect 7748 924 7807 958
rect 7620 896 7686 924
rect 7720 896 7807 924
rect 7113 868 7807 896
rect 7113 834 7174 868
rect 7208 834 7264 868
rect 7298 834 7354 868
rect 7388 834 7444 868
rect 7478 834 7534 868
rect 7568 834 7624 868
rect 7658 834 7714 868
rect 7748 834 7807 868
rect 7113 830 7807 834
rect 7113 796 7186 830
rect 7220 796 7286 830
rect 7320 796 7386 830
rect 7420 796 7486 830
rect 7520 796 7586 830
rect 7620 796 7686 830
rect 7720 796 7807 830
rect 7113 778 7807 796
rect 7113 744 7174 778
rect 7208 744 7264 778
rect 7298 744 7354 778
rect 7388 744 7444 778
rect 7478 744 7534 778
rect 7568 744 7624 778
rect 7658 744 7714 778
rect 7748 744 7807 778
rect 7113 730 7807 744
rect 7113 696 7186 730
rect 7220 696 7286 730
rect 7320 696 7386 730
rect 7420 696 7486 730
rect 7520 696 7586 730
rect 7620 696 7686 730
rect 7720 696 7807 730
rect 7113 688 7807 696
rect 7113 654 7174 688
rect 7208 654 7264 688
rect 7298 654 7354 688
rect 7388 654 7444 688
rect 7478 654 7534 688
rect 7568 654 7624 688
rect 7658 654 7714 688
rect 7748 654 7807 688
rect 7113 630 7807 654
rect 7113 598 7186 630
rect 7220 598 7286 630
rect 7320 598 7386 630
rect 7420 598 7486 630
rect 7113 564 7174 598
rect 7220 596 7264 598
rect 7320 596 7354 598
rect 7420 596 7444 598
rect 7208 564 7264 596
rect 7298 564 7354 596
rect 7388 564 7444 596
rect 7478 596 7486 598
rect 7520 598 7586 630
rect 7520 596 7534 598
rect 7478 564 7534 596
rect 7568 596 7586 598
rect 7620 598 7686 630
rect 7720 598 7807 630
rect 7620 596 7624 598
rect 7568 564 7624 596
rect 7658 596 7686 598
rect 7658 564 7714 596
rect 7748 564 7807 598
rect 7113 530 7807 564
rect 7113 508 7186 530
rect 7220 508 7286 530
rect 7320 508 7386 530
rect 7420 508 7486 530
rect 7113 474 7174 508
rect 7220 496 7264 508
rect 7320 496 7354 508
rect 7420 496 7444 508
rect 7208 474 7264 496
rect 7298 474 7354 496
rect 7388 474 7444 496
rect 7478 496 7486 508
rect 7520 508 7586 530
rect 7520 496 7534 508
rect 7478 474 7534 496
rect 7568 496 7586 508
rect 7620 508 7686 530
rect 7720 508 7807 530
rect 7620 496 7624 508
rect 7568 474 7624 496
rect 7658 496 7686 508
rect 7658 474 7714 496
rect 7748 474 7807 508
rect 7113 430 7807 474
rect 7113 418 7186 430
rect 7220 418 7286 430
rect 7320 418 7386 430
rect 7420 418 7486 430
rect 7113 384 7174 418
rect 7220 396 7264 418
rect 7320 396 7354 418
rect 7420 396 7444 418
rect 7208 384 7264 396
rect 7298 384 7354 396
rect 7388 384 7444 396
rect 7478 396 7486 418
rect 7520 418 7586 430
rect 7520 396 7534 418
rect 7478 384 7534 396
rect 7568 396 7586 418
rect 7620 418 7686 430
rect 7720 418 7807 430
rect 7620 396 7624 418
rect 7568 384 7624 396
rect 7658 396 7686 418
rect 7658 384 7714 396
rect 7748 384 7807 418
rect 7113 323 7807 384
rect 7860 986 8420 1022
rect 9220 1076 9470 1079
rect 9220 1056 9397 1076
rect 9220 1022 9248 1056
rect 9282 1042 9397 1056
rect 9431 1042 9470 1076
rect 9282 1022 9470 1042
rect 7860 966 8037 986
rect 7860 932 7888 966
rect 7922 952 8037 966
rect 8071 952 8210 986
rect 8244 985 8420 986
rect 8244 952 8358 985
rect 7922 951 8358 952
rect 8392 951 8420 985
rect 7922 932 8420 951
rect 7860 896 8420 932
rect 7860 876 8037 896
rect 7860 842 7888 876
rect 7922 862 8037 876
rect 8071 862 8210 896
rect 8244 895 8420 896
rect 8244 862 8358 895
rect 7922 861 8358 862
rect 8392 861 8420 895
rect 7922 842 8420 861
rect 7860 806 8420 842
rect 7860 786 8037 806
rect 7860 752 7888 786
rect 7922 772 8037 786
rect 8071 772 8210 806
rect 8244 805 8420 806
rect 8244 772 8358 805
rect 7922 771 8358 772
rect 8392 771 8420 805
rect 7922 752 8420 771
rect 7860 716 8420 752
rect 7860 696 8037 716
rect 7860 662 7888 696
rect 7922 682 8037 696
rect 8071 682 8210 716
rect 8244 715 8420 716
rect 8244 682 8358 715
rect 7922 681 8358 682
rect 8392 681 8420 715
rect 7922 662 8420 681
rect 7860 626 8420 662
rect 7860 606 8037 626
rect 7860 572 7888 606
rect 7922 592 8037 606
rect 8071 592 8210 626
rect 8244 625 8420 626
rect 8244 592 8358 625
rect 7922 591 8358 592
rect 8392 591 8420 625
rect 7922 572 8420 591
rect 7860 536 8420 572
rect 7860 516 8037 536
rect 7860 482 7888 516
rect 7922 502 8037 516
rect 8071 502 8210 536
rect 8244 535 8420 536
rect 8244 502 8358 535
rect 7922 501 8358 502
rect 8392 501 8420 535
rect 7922 482 8420 501
rect 7860 446 8420 482
rect 7860 426 8037 446
rect 7860 392 7888 426
rect 7922 412 8037 426
rect 8071 412 8210 446
rect 8244 445 8420 446
rect 8244 412 8358 445
rect 7922 411 8358 412
rect 8392 411 8420 445
rect 7922 392 8420 411
rect 7860 356 8420 392
rect 7860 336 8037 356
rect 6562 302 7060 321
rect 6500 270 7060 302
rect 7860 302 7888 336
rect 7922 322 8037 336
rect 8071 322 8210 356
rect 8244 355 8420 356
rect 8244 322 8358 355
rect 7922 321 8358 322
rect 8392 321 8420 355
rect 8473 958 9167 1017
rect 8473 924 8534 958
rect 8568 930 8624 958
rect 8658 930 8714 958
rect 8748 930 8804 958
rect 8580 924 8624 930
rect 8680 924 8714 930
rect 8780 924 8804 930
rect 8838 930 8894 958
rect 8838 924 8846 930
rect 8473 896 8546 924
rect 8580 896 8646 924
rect 8680 896 8746 924
rect 8780 896 8846 924
rect 8880 924 8894 930
rect 8928 930 8984 958
rect 8928 924 8946 930
rect 8880 896 8946 924
rect 8980 924 8984 930
rect 9018 930 9074 958
rect 9018 924 9046 930
rect 9108 924 9167 958
rect 8980 896 9046 924
rect 9080 896 9167 924
rect 8473 868 9167 896
rect 8473 834 8534 868
rect 8568 834 8624 868
rect 8658 834 8714 868
rect 8748 834 8804 868
rect 8838 834 8894 868
rect 8928 834 8984 868
rect 9018 834 9074 868
rect 9108 834 9167 868
rect 8473 830 9167 834
rect 8473 796 8546 830
rect 8580 796 8646 830
rect 8680 796 8746 830
rect 8780 796 8846 830
rect 8880 796 8946 830
rect 8980 796 9046 830
rect 9080 796 9167 830
rect 8473 778 9167 796
rect 8473 744 8534 778
rect 8568 744 8624 778
rect 8658 744 8714 778
rect 8748 744 8804 778
rect 8838 744 8894 778
rect 8928 744 8984 778
rect 9018 744 9074 778
rect 9108 744 9167 778
rect 8473 730 9167 744
rect 8473 696 8546 730
rect 8580 696 8646 730
rect 8680 696 8746 730
rect 8780 696 8846 730
rect 8880 696 8946 730
rect 8980 696 9046 730
rect 9080 696 9167 730
rect 8473 688 9167 696
rect 8473 654 8534 688
rect 8568 654 8624 688
rect 8658 654 8714 688
rect 8748 654 8804 688
rect 8838 654 8894 688
rect 8928 654 8984 688
rect 9018 654 9074 688
rect 9108 654 9167 688
rect 8473 630 9167 654
rect 8473 598 8546 630
rect 8580 598 8646 630
rect 8680 598 8746 630
rect 8780 598 8846 630
rect 8473 564 8534 598
rect 8580 596 8624 598
rect 8680 596 8714 598
rect 8780 596 8804 598
rect 8568 564 8624 596
rect 8658 564 8714 596
rect 8748 564 8804 596
rect 8838 596 8846 598
rect 8880 598 8946 630
rect 8880 596 8894 598
rect 8838 564 8894 596
rect 8928 596 8946 598
rect 8980 598 9046 630
rect 9080 598 9167 630
rect 8980 596 8984 598
rect 8928 564 8984 596
rect 9018 596 9046 598
rect 9018 564 9074 596
rect 9108 564 9167 598
rect 8473 530 9167 564
rect 8473 508 8546 530
rect 8580 508 8646 530
rect 8680 508 8746 530
rect 8780 508 8846 530
rect 8473 474 8534 508
rect 8580 496 8624 508
rect 8680 496 8714 508
rect 8780 496 8804 508
rect 8568 474 8624 496
rect 8658 474 8714 496
rect 8748 474 8804 496
rect 8838 496 8846 508
rect 8880 508 8946 530
rect 8880 496 8894 508
rect 8838 474 8894 496
rect 8928 496 8946 508
rect 8980 508 9046 530
rect 9080 508 9167 530
rect 8980 496 8984 508
rect 8928 474 8984 496
rect 9018 496 9046 508
rect 9018 474 9074 496
rect 9108 474 9167 508
rect 8473 430 9167 474
rect 8473 418 8546 430
rect 8580 418 8646 430
rect 8680 418 8746 430
rect 8780 418 8846 430
rect 8473 384 8534 418
rect 8580 396 8624 418
rect 8680 396 8714 418
rect 8780 396 8804 418
rect 8568 384 8624 396
rect 8658 384 8714 396
rect 8748 384 8804 396
rect 8838 396 8846 418
rect 8880 418 8946 430
rect 8880 396 8894 418
rect 8838 384 8894 396
rect 8928 396 8946 418
rect 8980 418 9046 430
rect 9080 418 9167 430
rect 8980 396 8984 418
rect 8928 384 8984 396
rect 9018 396 9046 418
rect 9018 384 9074 396
rect 9108 384 9167 418
rect 8473 323 9167 384
rect 9220 986 9470 1022
rect 9220 966 9397 986
rect 9220 932 9248 966
rect 9282 952 9397 966
rect 9431 952 9470 986
rect 9282 932 9470 952
rect 9220 896 9470 932
rect 9220 876 9397 896
rect 9220 842 9248 876
rect 9282 862 9397 876
rect 9431 862 9470 896
rect 9282 842 9470 862
rect 9220 806 9470 842
rect 9220 786 9397 806
rect 9220 752 9248 786
rect 9282 772 9397 786
rect 9431 772 9470 806
rect 9282 752 9470 772
rect 9220 716 9470 752
rect 9220 696 9397 716
rect 9220 662 9248 696
rect 9282 682 9397 696
rect 9431 682 9470 716
rect 9282 662 9470 682
rect 9220 626 9470 662
rect 9220 606 9397 626
rect 9220 572 9248 606
rect 9282 592 9397 606
rect 9431 592 9470 626
rect 9282 572 9470 592
rect 9220 536 9470 572
rect 9220 516 9397 536
rect 9220 482 9248 516
rect 9282 502 9397 516
rect 9431 502 9470 536
rect 9282 482 9470 502
rect 9220 446 9470 482
rect 9220 426 9397 446
rect 9220 392 9248 426
rect 9282 412 9397 426
rect 9431 412 9470 446
rect 9282 392 9470 412
rect 9220 356 9470 392
rect 9220 336 9397 356
rect 7922 302 8420 321
rect 7860 270 8420 302
rect 9220 302 9248 336
rect 9282 322 9397 336
rect 9431 322 9470 356
rect 9282 302 9470 322
rect 9220 270 9470 302
rect 10 266 9470 270
rect 10 232 1410 266
rect 1444 242 2597 266
rect 1444 232 1636 242
rect 10 208 1636 232
rect 1670 208 1726 242
rect 1760 208 1816 242
rect 1850 208 1906 242
rect 1940 208 1996 242
rect 2030 208 2086 242
rect 2120 208 2176 242
rect 2210 208 2266 242
rect 2300 208 2356 242
rect 2390 232 2597 242
rect 2631 232 2770 266
rect 2804 242 3957 266
rect 2804 232 2996 242
rect 2390 208 2996 232
rect 3030 208 3086 242
rect 3120 208 3176 242
rect 3210 208 3266 242
rect 3300 208 3356 242
rect 3390 208 3446 242
rect 3480 208 3536 242
rect 3570 208 3626 242
rect 3660 208 3716 242
rect 3750 232 3957 242
rect 3991 232 4130 266
rect 4164 242 5317 266
rect 4164 232 4356 242
rect 3750 208 4356 232
rect 4390 208 4446 242
rect 4480 208 4536 242
rect 4570 208 4626 242
rect 4660 208 4716 242
rect 4750 208 4806 242
rect 4840 208 4896 242
rect 4930 208 4986 242
rect 5020 208 5076 242
rect 5110 232 5317 242
rect 5351 232 5490 266
rect 5524 242 6677 266
rect 5524 232 5716 242
rect 5110 208 5716 232
rect 5750 208 5806 242
rect 5840 208 5896 242
rect 5930 208 5986 242
rect 6020 208 6076 242
rect 6110 208 6166 242
rect 6200 208 6256 242
rect 6290 208 6346 242
rect 6380 208 6436 242
rect 6470 232 6677 242
rect 6711 232 6850 266
rect 6884 242 8037 266
rect 6884 232 7076 242
rect 6470 208 7076 232
rect 7110 208 7166 242
rect 7200 208 7256 242
rect 7290 208 7346 242
rect 7380 208 7436 242
rect 7470 208 7526 242
rect 7560 208 7616 242
rect 7650 208 7706 242
rect 7740 208 7796 242
rect 7830 232 8037 242
rect 8071 232 8210 266
rect 8244 242 9397 266
rect 8244 232 8436 242
rect 7830 208 8436 232
rect 8470 208 8526 242
rect 8560 208 8616 242
rect 8650 208 8706 242
rect 8740 208 8796 242
rect 8830 208 8886 242
rect 8920 208 8976 242
rect 9010 208 9066 242
rect 9100 208 9156 242
rect 9190 232 9397 242
rect 9431 232 9470 266
rect 9190 208 9470 232
rect 10 176 9470 208
rect 10 142 1410 176
rect 1444 142 2597 176
rect 2631 142 2770 176
rect 2804 142 3957 176
rect 3991 142 4130 176
rect 4164 142 5317 176
rect 5351 142 5490 176
rect 5524 142 6677 176
rect 6711 142 6850 176
rect 6884 142 8037 176
rect 8071 142 8210 176
rect 8244 142 9397 176
rect 9431 142 9470 176
rect 10 92 9470 142
rect 10 58 1506 92
rect 1540 58 1596 92
rect 1630 58 1686 92
rect 1720 58 1776 92
rect 1810 58 1866 92
rect 1900 58 1956 92
rect 1990 58 2046 92
rect 2080 58 2136 92
rect 2170 58 2226 92
rect 2260 58 2316 92
rect 2350 58 2406 92
rect 2440 58 2496 92
rect 2530 58 2866 92
rect 2900 58 2956 92
rect 2990 58 3046 92
rect 3080 58 3136 92
rect 3170 58 3226 92
rect 3260 58 3316 92
rect 3350 58 3406 92
rect 3440 58 3496 92
rect 3530 58 3586 92
rect 3620 58 3676 92
rect 3710 58 3766 92
rect 3800 58 3856 92
rect 3890 58 4226 92
rect 4260 58 4316 92
rect 4350 58 4406 92
rect 4440 58 4496 92
rect 4530 58 4586 92
rect 4620 58 4676 92
rect 4710 58 4766 92
rect 4800 58 4856 92
rect 4890 58 4946 92
rect 4980 58 5036 92
rect 5070 58 5126 92
rect 5160 58 5216 92
rect 5250 58 5586 92
rect 5620 58 5676 92
rect 5710 58 5766 92
rect 5800 58 5856 92
rect 5890 58 5946 92
rect 5980 58 6036 92
rect 6070 58 6126 92
rect 6160 58 6216 92
rect 6250 58 6306 92
rect 6340 58 6396 92
rect 6430 58 6486 92
rect 6520 58 6576 92
rect 6610 58 6946 92
rect 6980 58 7036 92
rect 7070 58 7126 92
rect 7160 58 7216 92
rect 7250 58 7306 92
rect 7340 58 7396 92
rect 7430 58 7486 92
rect 7520 58 7576 92
rect 7610 58 7666 92
rect 7700 58 7756 92
rect 7790 58 7846 92
rect 7880 58 7936 92
rect 7970 58 8306 92
rect 8340 58 8396 92
rect 8430 58 8486 92
rect 8520 58 8576 92
rect 8610 58 8666 92
rect 8700 58 8756 92
rect 8790 58 8846 92
rect 8880 58 8936 92
rect 8970 58 9026 92
rect 9060 58 9116 92
rect 9150 58 9206 92
rect 9240 58 9296 92
rect 9330 58 9470 92
rect 10 20 9470 58
<< viali >>
rect 4630 5210 4670 5250
rect 5030 5210 5070 5250
rect 5430 5210 5470 5250
rect 5830 5210 5870 5250
rect 6230 5210 6270 5250
rect 6630 5210 6670 5250
rect 7030 5210 7070 5250
rect 7430 5210 7470 5250
rect 7830 5210 7870 5250
rect 8230 5210 8270 5250
rect 1910 4690 1950 4730
rect 4830 4270 4870 4310
rect 5230 4180 5270 4220
rect 6230 4270 6270 4310
rect 6030 4180 6070 4220
rect 6630 4270 6670 4310
rect 6830 4270 6870 4310
rect 7630 4270 7670 4310
rect 8030 4180 8070 4220
rect 3810 4100 3850 4140
rect 3900 4100 3940 4140
rect 3990 4100 4030 4140
rect 4080 4100 4120 4140
rect 4170 4100 4210 4140
rect 5630 4090 5670 4130
rect 6430 4090 6470 4130
rect 7230 4090 7270 4130
rect 4470 3900 4510 3940
rect 4670 3900 4710 3940
rect 5070 3900 5110 3940
rect 5470 3900 5510 3940
rect 5670 3900 5710 3940
rect 5830 3900 5870 3940
rect 6030 3900 6070 3940
rect 6230 3900 6270 3940
rect 6430 3900 6470 3940
rect 6630 3900 6670 3940
rect 6830 3900 6870 3940
rect 7030 3900 7070 3940
rect 7190 3900 7230 3940
rect 7390 3900 7430 3940
rect 7790 3900 7830 3940
rect 8190 3900 8230 3940
rect 8390 3900 8430 3940
rect 1910 3690 1950 3730
rect 5270 3360 5310 3400
rect 6430 3360 6470 3400
rect 7590 3360 7630 3400
rect 4870 3270 4910 3310
rect 6130 3270 6170 3310
rect 6730 3270 6770 3310
rect 7990 3270 8030 3310
rect 6430 3180 6470 3220
rect 3810 3100 3850 3140
rect 3900 3100 3940 3140
rect 3990 3100 4030 3140
rect 4080 3100 4120 3140
rect 4170 3100 4210 3140
rect 5550 3090 5590 3130
rect 5950 3090 5990 3130
rect 6070 3090 6110 3130
rect 6790 3090 6830 3130
rect 6910 3090 6950 3130
rect 7310 3090 7350 3130
rect 1910 2740 1950 2780
rect 3810 2740 3850 2780
rect 3900 2740 3940 2780
rect 3990 2740 4030 2780
rect 4080 2740 4120 2780
rect 4170 2740 4210 2780
rect 5550 2750 5590 2790
rect 7310 2750 7350 2790
rect 5150 2660 5190 2700
rect 5350 2660 5390 2700
rect 5750 2660 5790 2700
rect 6150 2660 6190 2700
rect 6350 2660 6390 2700
rect 6510 2660 6550 2700
rect 6710 2660 6750 2700
rect 7110 2660 7150 2700
rect 7510 2660 7550 2700
rect 7710 2660 7750 2700
rect 7310 2540 7350 2580
rect 1910 2150 1950 2190
rect 4670 1600 4710 1640
rect 6430 1600 6470 1640
rect 8190 1600 8230 1640
rect 1210 1370 1250 1410
rect 1430 1370 1470 1410
rect 1746 924 1768 930
rect 1768 924 1780 930
rect 1846 924 1858 930
rect 1858 924 1880 930
rect 1946 924 1948 930
rect 1948 924 1980 930
rect 1746 896 1780 924
rect 1846 896 1880 924
rect 1946 896 1980 924
rect 2046 896 2080 930
rect 2146 896 2180 930
rect 2246 924 2274 930
rect 2274 924 2280 930
rect 2246 896 2280 924
rect 1746 796 1780 830
rect 1846 796 1880 830
rect 1946 796 1980 830
rect 2046 796 2080 830
rect 2146 796 2180 830
rect 2246 796 2280 830
rect 1746 696 1780 730
rect 1846 696 1880 730
rect 1946 696 1980 730
rect 2046 696 2080 730
rect 2146 696 2180 730
rect 2246 696 2280 730
rect 1746 598 1780 630
rect 1846 598 1880 630
rect 1946 598 1980 630
rect 1746 596 1768 598
rect 1768 596 1780 598
rect 1846 596 1858 598
rect 1858 596 1880 598
rect 1946 596 1948 598
rect 1948 596 1980 598
rect 2046 596 2080 630
rect 2146 596 2180 630
rect 2246 598 2280 630
rect 2246 596 2274 598
rect 2274 596 2280 598
rect 1746 508 1780 530
rect 1846 508 1880 530
rect 1946 508 1980 530
rect 1746 496 1768 508
rect 1768 496 1780 508
rect 1846 496 1858 508
rect 1858 496 1880 508
rect 1946 496 1948 508
rect 1948 496 1980 508
rect 2046 496 2080 530
rect 2146 496 2180 530
rect 2246 508 2280 530
rect 2246 496 2274 508
rect 2274 496 2280 508
rect 1746 418 1780 430
rect 1846 418 1880 430
rect 1946 418 1980 430
rect 1746 396 1768 418
rect 1768 396 1780 418
rect 1846 396 1858 418
rect 1858 396 1880 418
rect 1946 396 1948 418
rect 1948 396 1980 418
rect 2046 396 2080 430
rect 2146 396 2180 430
rect 2246 418 2280 430
rect 2246 396 2274 418
rect 2274 396 2280 418
rect 3106 924 3128 930
rect 3128 924 3140 930
rect 3206 924 3218 930
rect 3218 924 3240 930
rect 3306 924 3308 930
rect 3308 924 3340 930
rect 3106 896 3140 924
rect 3206 896 3240 924
rect 3306 896 3340 924
rect 3406 896 3440 930
rect 3506 896 3540 930
rect 3606 924 3634 930
rect 3634 924 3640 930
rect 3606 896 3640 924
rect 3106 796 3140 830
rect 3206 796 3240 830
rect 3306 796 3340 830
rect 3406 796 3440 830
rect 3506 796 3540 830
rect 3606 796 3640 830
rect 3106 696 3140 730
rect 3206 696 3240 730
rect 3306 696 3340 730
rect 3406 696 3440 730
rect 3506 696 3540 730
rect 3606 696 3640 730
rect 3106 598 3140 630
rect 3206 598 3240 630
rect 3306 598 3340 630
rect 3106 596 3128 598
rect 3128 596 3140 598
rect 3206 596 3218 598
rect 3218 596 3240 598
rect 3306 596 3308 598
rect 3308 596 3340 598
rect 3406 596 3440 630
rect 3506 596 3540 630
rect 3606 598 3640 630
rect 3606 596 3634 598
rect 3634 596 3640 598
rect 3106 508 3140 530
rect 3206 508 3240 530
rect 3306 508 3340 530
rect 3106 496 3128 508
rect 3128 496 3140 508
rect 3206 496 3218 508
rect 3218 496 3240 508
rect 3306 496 3308 508
rect 3308 496 3340 508
rect 3406 496 3440 530
rect 3506 496 3540 530
rect 3606 508 3640 530
rect 3606 496 3634 508
rect 3634 496 3640 508
rect 3106 418 3140 430
rect 3206 418 3240 430
rect 3306 418 3340 430
rect 3106 396 3128 418
rect 3128 396 3140 418
rect 3206 396 3218 418
rect 3218 396 3240 418
rect 3306 396 3308 418
rect 3308 396 3340 418
rect 3406 396 3440 430
rect 3506 396 3540 430
rect 3606 418 3640 430
rect 3606 396 3634 418
rect 3634 396 3640 418
rect 4466 924 4488 930
rect 4488 924 4500 930
rect 4566 924 4578 930
rect 4578 924 4600 930
rect 4666 924 4668 930
rect 4668 924 4700 930
rect 4466 896 4500 924
rect 4566 896 4600 924
rect 4666 896 4700 924
rect 4766 896 4800 930
rect 4866 896 4900 930
rect 4966 924 4994 930
rect 4994 924 5000 930
rect 4966 896 5000 924
rect 4466 796 4500 830
rect 4566 796 4600 830
rect 4666 796 4700 830
rect 4766 796 4800 830
rect 4866 796 4900 830
rect 4966 796 5000 830
rect 4466 696 4500 730
rect 4566 696 4600 730
rect 4666 696 4700 730
rect 4766 696 4800 730
rect 4866 696 4900 730
rect 4966 696 5000 730
rect 4466 598 4500 630
rect 4566 598 4600 630
rect 4666 598 4700 630
rect 4466 596 4488 598
rect 4488 596 4500 598
rect 4566 596 4578 598
rect 4578 596 4600 598
rect 4666 596 4668 598
rect 4668 596 4700 598
rect 4766 596 4800 630
rect 4866 596 4900 630
rect 4966 598 5000 630
rect 4966 596 4994 598
rect 4994 596 5000 598
rect 4466 508 4500 530
rect 4566 508 4600 530
rect 4666 508 4700 530
rect 4466 496 4488 508
rect 4488 496 4500 508
rect 4566 496 4578 508
rect 4578 496 4600 508
rect 4666 496 4668 508
rect 4668 496 4700 508
rect 4766 496 4800 530
rect 4866 496 4900 530
rect 4966 508 5000 530
rect 4966 496 4994 508
rect 4994 496 5000 508
rect 4466 418 4500 430
rect 4566 418 4600 430
rect 4666 418 4700 430
rect 4466 396 4488 418
rect 4488 396 4500 418
rect 4566 396 4578 418
rect 4578 396 4600 418
rect 4666 396 4668 418
rect 4668 396 4700 418
rect 4766 396 4800 430
rect 4866 396 4900 430
rect 4966 418 5000 430
rect 4966 396 4994 418
rect 4994 396 5000 418
rect 5826 924 5848 930
rect 5848 924 5860 930
rect 5926 924 5938 930
rect 5938 924 5960 930
rect 6026 924 6028 930
rect 6028 924 6060 930
rect 5826 896 5860 924
rect 5926 896 5960 924
rect 6026 896 6060 924
rect 6126 896 6160 930
rect 6226 896 6260 930
rect 6326 924 6354 930
rect 6354 924 6360 930
rect 6326 896 6360 924
rect 5826 796 5860 830
rect 5926 796 5960 830
rect 6026 796 6060 830
rect 6126 796 6160 830
rect 6226 796 6260 830
rect 6326 796 6360 830
rect 5826 696 5860 730
rect 5926 696 5960 730
rect 6026 696 6060 730
rect 6126 696 6160 730
rect 6226 696 6260 730
rect 6326 696 6360 730
rect 5826 598 5860 630
rect 5926 598 5960 630
rect 6026 598 6060 630
rect 5826 596 5848 598
rect 5848 596 5860 598
rect 5926 596 5938 598
rect 5938 596 5960 598
rect 6026 596 6028 598
rect 6028 596 6060 598
rect 6126 596 6160 630
rect 6226 596 6260 630
rect 6326 598 6360 630
rect 6326 596 6354 598
rect 6354 596 6360 598
rect 5826 508 5860 530
rect 5926 508 5960 530
rect 6026 508 6060 530
rect 5826 496 5848 508
rect 5848 496 5860 508
rect 5926 496 5938 508
rect 5938 496 5960 508
rect 6026 496 6028 508
rect 6028 496 6060 508
rect 6126 496 6160 530
rect 6226 496 6260 530
rect 6326 508 6360 530
rect 6326 496 6354 508
rect 6354 496 6360 508
rect 5826 418 5860 430
rect 5926 418 5960 430
rect 6026 418 6060 430
rect 5826 396 5848 418
rect 5848 396 5860 418
rect 5926 396 5938 418
rect 5938 396 5960 418
rect 6026 396 6028 418
rect 6028 396 6060 418
rect 6126 396 6160 430
rect 6226 396 6260 430
rect 6326 418 6360 430
rect 6326 396 6354 418
rect 6354 396 6360 418
rect 7186 924 7208 930
rect 7208 924 7220 930
rect 7286 924 7298 930
rect 7298 924 7320 930
rect 7386 924 7388 930
rect 7388 924 7420 930
rect 7186 896 7220 924
rect 7286 896 7320 924
rect 7386 896 7420 924
rect 7486 896 7520 930
rect 7586 896 7620 930
rect 7686 924 7714 930
rect 7714 924 7720 930
rect 7686 896 7720 924
rect 7186 796 7220 830
rect 7286 796 7320 830
rect 7386 796 7420 830
rect 7486 796 7520 830
rect 7586 796 7620 830
rect 7686 796 7720 830
rect 7186 696 7220 730
rect 7286 696 7320 730
rect 7386 696 7420 730
rect 7486 696 7520 730
rect 7586 696 7620 730
rect 7686 696 7720 730
rect 7186 598 7220 630
rect 7286 598 7320 630
rect 7386 598 7420 630
rect 7186 596 7208 598
rect 7208 596 7220 598
rect 7286 596 7298 598
rect 7298 596 7320 598
rect 7386 596 7388 598
rect 7388 596 7420 598
rect 7486 596 7520 630
rect 7586 596 7620 630
rect 7686 598 7720 630
rect 7686 596 7714 598
rect 7714 596 7720 598
rect 7186 508 7220 530
rect 7286 508 7320 530
rect 7386 508 7420 530
rect 7186 496 7208 508
rect 7208 496 7220 508
rect 7286 496 7298 508
rect 7298 496 7320 508
rect 7386 496 7388 508
rect 7388 496 7420 508
rect 7486 496 7520 530
rect 7586 496 7620 530
rect 7686 508 7720 530
rect 7686 496 7714 508
rect 7714 496 7720 508
rect 7186 418 7220 430
rect 7286 418 7320 430
rect 7386 418 7420 430
rect 7186 396 7208 418
rect 7208 396 7220 418
rect 7286 396 7298 418
rect 7298 396 7320 418
rect 7386 396 7388 418
rect 7388 396 7420 418
rect 7486 396 7520 430
rect 7586 396 7620 430
rect 7686 418 7720 430
rect 7686 396 7714 418
rect 7714 396 7720 418
rect 8546 924 8568 930
rect 8568 924 8580 930
rect 8646 924 8658 930
rect 8658 924 8680 930
rect 8746 924 8748 930
rect 8748 924 8780 930
rect 8546 896 8580 924
rect 8646 896 8680 924
rect 8746 896 8780 924
rect 8846 896 8880 930
rect 8946 896 8980 930
rect 9046 924 9074 930
rect 9074 924 9080 930
rect 9046 896 9080 924
rect 8546 796 8580 830
rect 8646 796 8680 830
rect 8746 796 8780 830
rect 8846 796 8880 830
rect 8946 796 8980 830
rect 9046 796 9080 830
rect 8546 696 8580 730
rect 8646 696 8680 730
rect 8746 696 8780 730
rect 8846 696 8880 730
rect 8946 696 8980 730
rect 9046 696 9080 730
rect 8546 598 8580 630
rect 8646 598 8680 630
rect 8746 598 8780 630
rect 8546 596 8568 598
rect 8568 596 8580 598
rect 8646 596 8658 598
rect 8658 596 8680 598
rect 8746 596 8748 598
rect 8748 596 8780 598
rect 8846 596 8880 630
rect 8946 596 8980 630
rect 9046 598 9080 630
rect 9046 596 9074 598
rect 9074 596 9080 598
rect 8546 508 8580 530
rect 8646 508 8680 530
rect 8746 508 8780 530
rect 8546 496 8568 508
rect 8568 496 8580 508
rect 8646 496 8658 508
rect 8658 496 8680 508
rect 8746 496 8748 508
rect 8748 496 8780 508
rect 8846 496 8880 530
rect 8946 496 8980 530
rect 9046 508 9080 530
rect 9046 496 9074 508
rect 9074 496 9080 508
rect 8546 418 8580 430
rect 8646 418 8680 430
rect 8746 418 8780 430
rect 8546 396 8568 418
rect 8568 396 8580 418
rect 8646 396 8658 418
rect 8658 396 8680 418
rect 8746 396 8748 418
rect 8748 396 8780 418
rect 8846 396 8880 430
rect 8946 396 8980 430
rect 9046 418 9080 430
rect 9046 396 9074 418
rect 9074 396 9080 418
<< metal1 >>
rect 4610 5260 4690 5270
rect 4610 5200 4620 5260
rect 4680 5200 4690 5260
rect 4610 5190 4690 5200
rect 5010 5260 5090 5270
rect 5010 5200 5020 5260
rect 5080 5200 5090 5260
rect 5010 5190 5090 5200
rect 5410 5260 5490 5270
rect 5410 5200 5420 5260
rect 5480 5200 5490 5260
rect 5410 5190 5490 5200
rect 5810 5260 5890 5270
rect 5810 5200 5820 5260
rect 5880 5200 5890 5260
rect 5810 5190 5890 5200
rect 6210 5260 6290 5270
rect 6210 5200 6220 5260
rect 6280 5200 6290 5260
rect 6210 5190 6290 5200
rect 6610 5260 6690 5270
rect 6610 5200 6620 5260
rect 6680 5200 6690 5260
rect 6610 5190 6690 5200
rect 7010 5260 7090 5270
rect 7010 5200 7020 5260
rect 7080 5200 7090 5260
rect 7010 5190 7090 5200
rect 7410 5260 7490 5270
rect 7410 5200 7420 5260
rect 7480 5200 7490 5260
rect 7410 5190 7490 5200
rect 7810 5260 7890 5270
rect 7810 5200 7820 5260
rect 7880 5200 7890 5260
rect 7810 5190 7890 5200
rect 8210 5260 8290 5270
rect 8210 5200 8220 5260
rect 8280 5200 8290 5260
rect 8210 5190 8290 5200
rect 1190 4740 1270 4750
rect 1190 4680 1200 4740
rect 1260 4680 1270 4740
rect 1190 3740 1270 4680
rect 1890 4740 1970 4750
rect 1890 4680 1900 4740
rect 1960 4680 1970 4740
rect 1890 4670 1970 4680
rect 4810 4320 4890 4330
rect 4810 4260 4820 4320
rect 4880 4260 4890 4320
rect 4810 4250 4890 4260
rect 6210 4310 6290 4330
rect 6210 4270 6230 4310
rect 6270 4270 6290 4310
rect 6210 4250 6290 4270
rect 6610 4310 6690 4330
rect 6610 4270 6630 4310
rect 6670 4270 6690 4310
rect 6610 4250 6690 4270
rect 6810 4320 6890 4330
rect 6810 4260 6820 4320
rect 6880 4260 6890 4320
rect 6810 4250 6890 4260
rect 7610 4320 7690 4330
rect 7610 4260 7620 4320
rect 7680 4260 7690 4320
rect 7610 4250 7690 4260
rect 5210 4230 5290 4240
rect 5210 4170 5220 4230
rect 5280 4170 5290 4230
rect 5210 4160 5290 4170
rect 6010 4230 6090 4240
rect 6010 4170 6020 4230
rect 6080 4170 6090 4230
rect 6010 4160 6090 4170
rect 3790 4150 4230 4160
rect 3790 4090 3800 4150
rect 4220 4090 4230 4150
rect 3790 4080 4230 4090
rect 5610 4140 5690 4150
rect 5610 4080 5620 4140
rect 5680 4080 5690 4140
rect 5610 4070 5690 4080
rect 6230 3960 6270 4250
rect 6410 4140 6490 4150
rect 6410 4080 6420 4140
rect 6480 4080 6490 4140
rect 6410 4070 6490 4080
rect 6630 3960 6670 4250
rect 8010 4230 8090 4240
rect 8010 4170 8020 4230
rect 8080 4170 8090 4230
rect 8010 4160 8090 4170
rect 7210 4140 7290 4150
rect 7210 4080 7220 4140
rect 7280 4080 7290 4140
rect 7210 4070 7290 4080
rect 4450 3950 4530 3960
rect 4450 3890 4460 3950
rect 4520 3890 4530 3950
rect 4450 3880 4530 3890
rect 4650 3950 4730 3960
rect 4650 3890 4660 3950
rect 4720 3890 4730 3950
rect 4650 3880 4730 3890
rect 5050 3950 5130 3960
rect 5050 3890 5060 3950
rect 5120 3890 5130 3950
rect 5050 3880 5130 3890
rect 5450 3950 5530 3960
rect 5450 3890 5460 3950
rect 5520 3890 5530 3950
rect 5450 3880 5530 3890
rect 5650 3950 5730 3960
rect 5650 3890 5660 3950
rect 5720 3890 5730 3950
rect 5650 3880 5730 3890
rect 5810 3950 5890 3960
rect 5810 3890 5820 3950
rect 5880 3890 5890 3950
rect 5810 3880 5890 3890
rect 6010 3950 6090 3960
rect 6010 3890 6020 3950
rect 6080 3890 6090 3950
rect 6010 3880 6090 3890
rect 6210 3940 6290 3960
rect 6210 3900 6230 3940
rect 6270 3900 6290 3940
rect 6210 3880 6290 3900
rect 6410 3950 6490 3960
rect 6410 3890 6420 3950
rect 6480 3890 6490 3950
rect 6410 3880 6490 3890
rect 6610 3940 6690 3960
rect 6610 3900 6630 3940
rect 6670 3900 6690 3940
rect 6610 3880 6690 3900
rect 6810 3950 6890 3960
rect 6810 3890 6820 3950
rect 6880 3890 6890 3950
rect 6810 3880 6890 3890
rect 7010 3950 7090 3960
rect 7010 3890 7020 3950
rect 7080 3890 7090 3950
rect 7010 3880 7090 3890
rect 7170 3950 7250 3960
rect 7170 3890 7180 3950
rect 7240 3890 7250 3950
rect 7170 3880 7250 3890
rect 7370 3950 7450 3960
rect 7370 3890 7380 3950
rect 7440 3890 7450 3950
rect 7370 3880 7450 3890
rect 7770 3950 7850 3960
rect 7770 3890 7780 3950
rect 7840 3890 7850 3950
rect 7770 3880 7850 3890
rect 8170 3950 8250 3960
rect 8170 3890 8180 3950
rect 8240 3890 8250 3950
rect 8170 3880 8250 3890
rect 8370 3950 8450 3960
rect 8370 3890 8380 3950
rect 8440 3890 8450 3950
rect 8370 3880 8450 3890
rect 1190 3680 1200 3740
rect 1260 3680 1270 3740
rect 880 3150 960 3160
rect 880 3090 890 3150
rect 950 3090 960 3150
rect 880 1450 960 3090
rect 360 370 960 1450
rect 1190 1410 1270 3680
rect 1890 3740 1970 3750
rect 1890 3680 1900 3740
rect 1960 3680 1970 3740
rect 1890 3670 1970 3680
rect 5250 3410 5330 3420
rect 5250 3350 5260 3410
rect 5320 3350 5330 3410
rect 5250 3340 5330 3350
rect 5930 3410 6010 3420
rect 5930 3350 5940 3410
rect 6000 3350 6010 3410
rect 5930 3340 6010 3350
rect 6410 3400 6490 3420
rect 6410 3360 6430 3400
rect 6470 3360 6490 3400
rect 6410 3340 6490 3360
rect 6890 3410 6970 3420
rect 6890 3350 6900 3410
rect 6960 3350 6970 3410
rect 6890 3340 6970 3350
rect 7570 3410 7650 3420
rect 7570 3350 7580 3410
rect 7640 3350 7650 3410
rect 7570 3340 7650 3350
rect 4850 3320 4930 3330
rect 4850 3260 4860 3320
rect 4920 3260 4930 3320
rect 4850 3250 4930 3260
rect 5530 3320 5610 3330
rect 5530 3260 5540 3320
rect 5600 3260 5610 3320
rect 5530 3250 5610 3260
rect 3790 3150 4230 3160
rect 5550 3150 5590 3250
rect 5950 3150 5990 3340
rect 6110 3320 6190 3330
rect 6110 3260 6120 3320
rect 6180 3260 6190 3320
rect 6110 3250 6190 3260
rect 6430 3240 6470 3340
rect 6710 3320 6790 3330
rect 6710 3260 6720 3320
rect 6780 3260 6790 3320
rect 6710 3250 6790 3260
rect 6410 3230 6490 3240
rect 6410 3170 6420 3230
rect 6480 3170 6490 3230
rect 6410 3160 6490 3170
rect 6910 3150 6950 3340
rect 7290 3320 7370 3330
rect 7290 3260 7300 3320
rect 7360 3260 7370 3320
rect 7290 3250 7370 3260
rect 7970 3320 8050 3330
rect 7970 3260 7980 3320
rect 8040 3260 8050 3320
rect 7970 3250 8050 3260
rect 7310 3150 7350 3250
rect 7830 3230 7910 3240
rect 7830 3170 7840 3230
rect 7900 3170 7910 3230
rect 7830 3160 7910 3170
rect 3790 3090 3800 3150
rect 4220 3090 4230 3150
rect 3790 3080 4230 3090
rect 5530 3130 5610 3150
rect 5530 3090 5550 3130
rect 5590 3090 5610 3130
rect 5530 3070 5610 3090
rect 5930 3130 6010 3150
rect 5930 3090 5950 3130
rect 5990 3090 6010 3130
rect 5930 3070 6010 3090
rect 6050 3140 6130 3150
rect 6050 3080 6060 3140
rect 6120 3080 6130 3140
rect 6050 3070 6130 3080
rect 6770 3140 6850 3150
rect 6770 3080 6780 3140
rect 6840 3080 6850 3140
rect 6770 3070 6850 3080
rect 6890 3130 6970 3150
rect 6890 3090 6910 3130
rect 6950 3090 6970 3130
rect 6890 3070 6970 3090
rect 7290 3130 7370 3150
rect 7290 3090 7310 3130
rect 7350 3090 7370 3130
rect 7290 3070 7370 3090
rect 5530 2800 5610 2810
rect 1720 2790 1800 2800
rect 1720 2730 1730 2790
rect 1790 2730 1800 2790
rect 1190 1370 1210 1410
rect 1250 1370 1270 1410
rect 1190 1340 1270 1370
rect 1410 2200 1490 2210
rect 1410 2140 1420 2200
rect 1480 2140 1490 2200
rect 1410 1410 1490 2140
rect 1410 1370 1430 1410
rect 1470 1370 1490 1410
rect 1410 1340 1490 1370
rect 1720 1460 1800 2730
rect 1890 2790 1970 2800
rect 1890 2730 1900 2790
rect 1960 2730 1970 2790
rect 1890 2720 1970 2730
rect 3790 2790 4230 2800
rect 3790 2730 3800 2790
rect 4220 2730 4230 2790
rect 5530 2740 5540 2800
rect 5600 2740 5610 2800
rect 5530 2730 5610 2740
rect 7290 2800 7370 2810
rect 7290 2740 7300 2800
rect 7360 2740 7370 2800
rect 7290 2730 7370 2740
rect 3790 2720 4230 2730
rect 5130 2710 5210 2720
rect 5130 2650 5140 2710
rect 5200 2650 5210 2710
rect 5130 2640 5210 2650
rect 5330 2710 5410 2720
rect 5330 2650 5340 2710
rect 5400 2650 5410 2710
rect 5330 2640 5410 2650
rect 5730 2710 5810 2720
rect 5730 2650 5740 2710
rect 5800 2650 5810 2710
rect 5730 2640 5810 2650
rect 6130 2710 6210 2720
rect 6130 2650 6140 2710
rect 6200 2650 6210 2710
rect 6130 2640 6210 2650
rect 6330 2710 6410 2720
rect 6330 2650 6340 2710
rect 6400 2650 6410 2710
rect 6330 2640 6410 2650
rect 6490 2710 6570 2720
rect 6490 2650 6500 2710
rect 6560 2650 6570 2710
rect 6490 2640 6570 2650
rect 6690 2710 6770 2720
rect 6690 2650 6700 2710
rect 6760 2650 6770 2710
rect 6690 2640 6770 2650
rect 7090 2710 7170 2720
rect 7090 2650 7100 2710
rect 7160 2650 7170 2710
rect 7090 2640 7170 2650
rect 7490 2710 7570 2720
rect 7490 2650 7500 2710
rect 7560 2650 7570 2710
rect 7490 2640 7570 2650
rect 7690 2710 7770 2720
rect 7690 2650 7700 2710
rect 7760 2650 7770 2710
rect 7690 2640 7770 2650
rect 7850 2600 7890 3160
rect 7290 2590 7370 2600
rect 7290 2530 7300 2590
rect 7360 2530 7370 2590
rect 7290 2520 7370 2530
rect 7830 2590 7910 2600
rect 7830 2530 7840 2590
rect 7900 2530 7910 2590
rect 7830 2520 7910 2530
rect 1890 2200 1970 2210
rect 1890 2140 1900 2200
rect 1960 2140 1970 2200
rect 1890 2130 1970 2140
rect 4650 1650 4730 1660
rect 4650 1590 4660 1650
rect 4720 1590 4730 1650
rect 4650 1580 4730 1590
rect 6410 1650 6490 1660
rect 6410 1590 6420 1650
rect 6480 1590 6490 1650
rect 6410 1580 6490 1590
rect 8170 1650 8250 1660
rect 8170 1590 8180 1650
rect 8240 1590 8250 1650
rect 8170 1580 8250 1590
rect 1720 1420 9120 1460
rect 1720 975 2320 1420
rect 3080 975 3680 1420
rect 4440 975 5040 1420
rect 5800 975 6400 1420
rect 7160 975 7760 1420
rect 8520 975 9120 1420
rect 1715 930 2325 975
rect 1715 896 1746 930
rect 1780 896 1846 930
rect 1880 896 1946 930
rect 1980 896 2046 930
rect 2080 896 2146 930
rect 2180 896 2246 930
rect 2280 896 2325 930
rect 1715 830 2325 896
rect 1715 796 1746 830
rect 1780 796 1846 830
rect 1880 796 1946 830
rect 1980 796 2046 830
rect 2080 796 2146 830
rect 2180 796 2246 830
rect 2280 796 2325 830
rect 1715 730 2325 796
rect 1715 696 1746 730
rect 1780 696 1846 730
rect 1880 696 1946 730
rect 1980 696 2046 730
rect 2080 696 2146 730
rect 2180 696 2246 730
rect 2280 696 2325 730
rect 1715 630 2325 696
rect 1715 596 1746 630
rect 1780 596 1846 630
rect 1880 596 1946 630
rect 1980 596 2046 630
rect 2080 596 2146 630
rect 2180 596 2246 630
rect 2280 596 2325 630
rect 1715 530 2325 596
rect 1715 496 1746 530
rect 1780 496 1846 530
rect 1880 496 1946 530
rect 1980 496 2046 530
rect 2080 496 2146 530
rect 2180 496 2246 530
rect 2280 496 2325 530
rect 1715 430 2325 496
rect 1715 396 1746 430
rect 1780 396 1846 430
rect 1880 396 1946 430
rect 1980 396 2046 430
rect 2080 396 2146 430
rect 2180 396 2246 430
rect 2280 396 2325 430
rect 1715 365 2325 396
rect 3075 930 3685 975
rect 3075 896 3106 930
rect 3140 896 3206 930
rect 3240 896 3306 930
rect 3340 896 3406 930
rect 3440 896 3506 930
rect 3540 896 3606 930
rect 3640 896 3685 930
rect 3075 830 3685 896
rect 3075 796 3106 830
rect 3140 796 3206 830
rect 3240 796 3306 830
rect 3340 796 3406 830
rect 3440 796 3506 830
rect 3540 796 3606 830
rect 3640 796 3685 830
rect 3075 730 3685 796
rect 3075 696 3106 730
rect 3140 696 3206 730
rect 3240 696 3306 730
rect 3340 696 3406 730
rect 3440 696 3506 730
rect 3540 696 3606 730
rect 3640 696 3685 730
rect 3075 630 3685 696
rect 3075 596 3106 630
rect 3140 596 3206 630
rect 3240 596 3306 630
rect 3340 596 3406 630
rect 3440 596 3506 630
rect 3540 596 3606 630
rect 3640 596 3685 630
rect 3075 530 3685 596
rect 3075 496 3106 530
rect 3140 496 3206 530
rect 3240 496 3306 530
rect 3340 496 3406 530
rect 3440 496 3506 530
rect 3540 496 3606 530
rect 3640 496 3685 530
rect 3075 430 3685 496
rect 3075 396 3106 430
rect 3140 396 3206 430
rect 3240 396 3306 430
rect 3340 396 3406 430
rect 3440 396 3506 430
rect 3540 396 3606 430
rect 3640 396 3685 430
rect 3075 365 3685 396
rect 4435 930 5045 975
rect 4435 896 4466 930
rect 4500 896 4566 930
rect 4600 896 4666 930
rect 4700 896 4766 930
rect 4800 896 4866 930
rect 4900 896 4966 930
rect 5000 896 5045 930
rect 4435 830 5045 896
rect 4435 796 4466 830
rect 4500 796 4566 830
rect 4600 796 4666 830
rect 4700 796 4766 830
rect 4800 796 4866 830
rect 4900 796 4966 830
rect 5000 796 5045 830
rect 4435 730 5045 796
rect 4435 696 4466 730
rect 4500 696 4566 730
rect 4600 696 4666 730
rect 4700 696 4766 730
rect 4800 696 4866 730
rect 4900 696 4966 730
rect 5000 696 5045 730
rect 4435 630 5045 696
rect 4435 596 4466 630
rect 4500 596 4566 630
rect 4600 596 4666 630
rect 4700 596 4766 630
rect 4800 596 4866 630
rect 4900 596 4966 630
rect 5000 596 5045 630
rect 4435 530 5045 596
rect 4435 496 4466 530
rect 4500 496 4566 530
rect 4600 496 4666 530
rect 4700 496 4766 530
rect 4800 496 4866 530
rect 4900 496 4966 530
rect 5000 496 5045 530
rect 4435 430 5045 496
rect 4435 396 4466 430
rect 4500 396 4566 430
rect 4600 396 4666 430
rect 4700 396 4766 430
rect 4800 396 4866 430
rect 4900 396 4966 430
rect 5000 396 5045 430
rect 4435 365 5045 396
rect 5795 930 6405 975
rect 5795 896 5826 930
rect 5860 896 5926 930
rect 5960 896 6026 930
rect 6060 896 6126 930
rect 6160 896 6226 930
rect 6260 896 6326 930
rect 6360 896 6405 930
rect 5795 830 6405 896
rect 5795 796 5826 830
rect 5860 796 5926 830
rect 5960 796 6026 830
rect 6060 796 6126 830
rect 6160 796 6226 830
rect 6260 796 6326 830
rect 6360 796 6405 830
rect 5795 730 6405 796
rect 5795 696 5826 730
rect 5860 696 5926 730
rect 5960 696 6026 730
rect 6060 696 6126 730
rect 6160 696 6226 730
rect 6260 696 6326 730
rect 6360 696 6405 730
rect 5795 630 6405 696
rect 5795 596 5826 630
rect 5860 596 5926 630
rect 5960 596 6026 630
rect 6060 596 6126 630
rect 6160 596 6226 630
rect 6260 596 6326 630
rect 6360 596 6405 630
rect 5795 530 6405 596
rect 5795 496 5826 530
rect 5860 496 5926 530
rect 5960 496 6026 530
rect 6060 496 6126 530
rect 6160 496 6226 530
rect 6260 496 6326 530
rect 6360 496 6405 530
rect 5795 430 6405 496
rect 5795 396 5826 430
rect 5860 396 5926 430
rect 5960 396 6026 430
rect 6060 396 6126 430
rect 6160 396 6226 430
rect 6260 396 6326 430
rect 6360 396 6405 430
rect 5795 365 6405 396
rect 7155 930 7765 975
rect 7155 896 7186 930
rect 7220 896 7286 930
rect 7320 896 7386 930
rect 7420 896 7486 930
rect 7520 896 7586 930
rect 7620 896 7686 930
rect 7720 896 7765 930
rect 7155 830 7765 896
rect 7155 796 7186 830
rect 7220 796 7286 830
rect 7320 796 7386 830
rect 7420 796 7486 830
rect 7520 796 7586 830
rect 7620 796 7686 830
rect 7720 796 7765 830
rect 7155 730 7765 796
rect 7155 696 7186 730
rect 7220 696 7286 730
rect 7320 696 7386 730
rect 7420 696 7486 730
rect 7520 696 7586 730
rect 7620 696 7686 730
rect 7720 696 7765 730
rect 7155 630 7765 696
rect 7155 596 7186 630
rect 7220 596 7286 630
rect 7320 596 7386 630
rect 7420 596 7486 630
rect 7520 596 7586 630
rect 7620 596 7686 630
rect 7720 596 7765 630
rect 7155 530 7765 596
rect 7155 496 7186 530
rect 7220 496 7286 530
rect 7320 496 7386 530
rect 7420 496 7486 530
rect 7520 496 7586 530
rect 7620 496 7686 530
rect 7720 496 7765 530
rect 7155 430 7765 496
rect 7155 396 7186 430
rect 7220 396 7286 430
rect 7320 396 7386 430
rect 7420 396 7486 430
rect 7520 396 7586 430
rect 7620 396 7686 430
rect 7720 396 7765 430
rect 7155 365 7765 396
rect 8515 930 9125 975
rect 8515 896 8546 930
rect 8580 896 8646 930
rect 8680 896 8746 930
rect 8780 896 8846 930
rect 8880 896 8946 930
rect 8980 896 9046 930
rect 9080 896 9125 930
rect 8515 830 9125 896
rect 8515 796 8546 830
rect 8580 796 8646 830
rect 8680 796 8746 830
rect 8780 796 8846 830
rect 8880 796 8946 830
rect 8980 796 9046 830
rect 9080 796 9125 830
rect 8515 730 9125 796
rect 8515 696 8546 730
rect 8580 696 8646 730
rect 8680 696 8746 730
rect 8780 696 8846 730
rect 8880 696 8946 730
rect 8980 696 9046 730
rect 9080 696 9125 730
rect 8515 630 9125 696
rect 8515 596 8546 630
rect 8580 596 8646 630
rect 8680 596 8746 630
rect 8780 596 8846 630
rect 8880 596 8946 630
rect 8980 596 9046 630
rect 9080 596 9125 630
rect 8515 530 9125 596
rect 8515 496 8546 530
rect 8580 496 8646 530
rect 8680 496 8746 530
rect 8780 496 8846 530
rect 8880 496 8946 530
rect 8980 496 9046 530
rect 9080 496 9125 530
rect 8515 430 9125 496
rect 8515 396 8546 430
rect 8580 396 8646 430
rect 8680 396 8746 430
rect 8780 396 8846 430
rect 8880 396 8946 430
rect 8980 396 9046 430
rect 9080 396 9125 430
rect 8515 365 9125 396
<< via1 >>
rect 4620 5250 4680 5260
rect 4620 5210 4630 5250
rect 4630 5210 4670 5250
rect 4670 5210 4680 5250
rect 4620 5200 4680 5210
rect 5020 5250 5080 5260
rect 5020 5210 5030 5250
rect 5030 5210 5070 5250
rect 5070 5210 5080 5250
rect 5020 5200 5080 5210
rect 5420 5250 5480 5260
rect 5420 5210 5430 5250
rect 5430 5210 5470 5250
rect 5470 5210 5480 5250
rect 5420 5200 5480 5210
rect 5820 5250 5880 5260
rect 5820 5210 5830 5250
rect 5830 5210 5870 5250
rect 5870 5210 5880 5250
rect 5820 5200 5880 5210
rect 6220 5250 6280 5260
rect 6220 5210 6230 5250
rect 6230 5210 6270 5250
rect 6270 5210 6280 5250
rect 6220 5200 6280 5210
rect 6620 5250 6680 5260
rect 6620 5210 6630 5250
rect 6630 5210 6670 5250
rect 6670 5210 6680 5250
rect 6620 5200 6680 5210
rect 7020 5250 7080 5260
rect 7020 5210 7030 5250
rect 7030 5210 7070 5250
rect 7070 5210 7080 5250
rect 7020 5200 7080 5210
rect 7420 5250 7480 5260
rect 7420 5210 7430 5250
rect 7430 5210 7470 5250
rect 7470 5210 7480 5250
rect 7420 5200 7480 5210
rect 7820 5250 7880 5260
rect 7820 5210 7830 5250
rect 7830 5210 7870 5250
rect 7870 5210 7880 5250
rect 7820 5200 7880 5210
rect 8220 5250 8280 5260
rect 8220 5210 8230 5250
rect 8230 5210 8270 5250
rect 8270 5210 8280 5250
rect 8220 5200 8280 5210
rect 1200 4680 1260 4740
rect 1900 4730 1960 4740
rect 1900 4690 1910 4730
rect 1910 4690 1950 4730
rect 1950 4690 1960 4730
rect 1900 4680 1960 4690
rect 4820 4310 4880 4320
rect 4820 4270 4830 4310
rect 4830 4270 4870 4310
rect 4870 4270 4880 4310
rect 4820 4260 4880 4270
rect 6820 4310 6880 4320
rect 6820 4270 6830 4310
rect 6830 4270 6870 4310
rect 6870 4270 6880 4310
rect 6820 4260 6880 4270
rect 7620 4310 7680 4320
rect 7620 4270 7630 4310
rect 7630 4270 7670 4310
rect 7670 4270 7680 4310
rect 7620 4260 7680 4270
rect 5220 4220 5280 4230
rect 5220 4180 5230 4220
rect 5230 4180 5270 4220
rect 5270 4180 5280 4220
rect 5220 4170 5280 4180
rect 6020 4220 6080 4230
rect 6020 4180 6030 4220
rect 6030 4180 6070 4220
rect 6070 4180 6080 4220
rect 6020 4170 6080 4180
rect 3800 4140 4220 4150
rect 3800 4100 3810 4140
rect 3810 4100 3850 4140
rect 3850 4100 3900 4140
rect 3900 4100 3940 4140
rect 3940 4100 3990 4140
rect 3990 4100 4030 4140
rect 4030 4100 4080 4140
rect 4080 4100 4120 4140
rect 4120 4100 4170 4140
rect 4170 4100 4210 4140
rect 4210 4100 4220 4140
rect 3800 4090 4220 4100
rect 5620 4130 5680 4140
rect 5620 4090 5630 4130
rect 5630 4090 5670 4130
rect 5670 4090 5680 4130
rect 5620 4080 5680 4090
rect 6420 4130 6480 4140
rect 6420 4090 6430 4130
rect 6430 4090 6470 4130
rect 6470 4090 6480 4130
rect 6420 4080 6480 4090
rect 8020 4220 8080 4230
rect 8020 4180 8030 4220
rect 8030 4180 8070 4220
rect 8070 4180 8080 4220
rect 8020 4170 8080 4180
rect 7220 4130 7280 4140
rect 7220 4090 7230 4130
rect 7230 4090 7270 4130
rect 7270 4090 7280 4130
rect 7220 4080 7280 4090
rect 4460 3940 4520 3950
rect 4460 3900 4470 3940
rect 4470 3900 4510 3940
rect 4510 3900 4520 3940
rect 4460 3890 4520 3900
rect 4660 3940 4720 3950
rect 4660 3900 4670 3940
rect 4670 3900 4710 3940
rect 4710 3900 4720 3940
rect 4660 3890 4720 3900
rect 5060 3940 5120 3950
rect 5060 3900 5070 3940
rect 5070 3900 5110 3940
rect 5110 3900 5120 3940
rect 5060 3890 5120 3900
rect 5460 3940 5520 3950
rect 5460 3900 5470 3940
rect 5470 3900 5510 3940
rect 5510 3900 5520 3940
rect 5460 3890 5520 3900
rect 5660 3940 5720 3950
rect 5660 3900 5670 3940
rect 5670 3900 5710 3940
rect 5710 3900 5720 3940
rect 5660 3890 5720 3900
rect 5820 3940 5880 3950
rect 5820 3900 5830 3940
rect 5830 3900 5870 3940
rect 5870 3900 5880 3940
rect 5820 3890 5880 3900
rect 6020 3940 6080 3950
rect 6020 3900 6030 3940
rect 6030 3900 6070 3940
rect 6070 3900 6080 3940
rect 6020 3890 6080 3900
rect 6420 3940 6480 3950
rect 6420 3900 6430 3940
rect 6430 3900 6470 3940
rect 6470 3900 6480 3940
rect 6420 3890 6480 3900
rect 6820 3940 6880 3950
rect 6820 3900 6830 3940
rect 6830 3900 6870 3940
rect 6870 3900 6880 3940
rect 6820 3890 6880 3900
rect 7020 3940 7080 3950
rect 7020 3900 7030 3940
rect 7030 3900 7070 3940
rect 7070 3900 7080 3940
rect 7020 3890 7080 3900
rect 7180 3940 7240 3950
rect 7180 3900 7190 3940
rect 7190 3900 7230 3940
rect 7230 3900 7240 3940
rect 7180 3890 7240 3900
rect 7380 3940 7440 3950
rect 7380 3900 7390 3940
rect 7390 3900 7430 3940
rect 7430 3900 7440 3940
rect 7380 3890 7440 3900
rect 7780 3940 7840 3950
rect 7780 3900 7790 3940
rect 7790 3900 7830 3940
rect 7830 3900 7840 3940
rect 7780 3890 7840 3900
rect 8180 3940 8240 3950
rect 8180 3900 8190 3940
rect 8190 3900 8230 3940
rect 8230 3900 8240 3940
rect 8180 3890 8240 3900
rect 8380 3940 8440 3950
rect 8380 3900 8390 3940
rect 8390 3900 8430 3940
rect 8430 3900 8440 3940
rect 8380 3890 8440 3900
rect 1200 3680 1260 3740
rect 890 3090 950 3150
rect 1900 3730 1960 3740
rect 1900 3690 1910 3730
rect 1910 3690 1950 3730
rect 1950 3690 1960 3730
rect 1900 3680 1960 3690
rect 5260 3400 5320 3410
rect 5260 3360 5270 3400
rect 5270 3360 5310 3400
rect 5310 3360 5320 3400
rect 5260 3350 5320 3360
rect 5940 3350 6000 3410
rect 6900 3350 6960 3410
rect 7580 3400 7640 3410
rect 7580 3360 7590 3400
rect 7590 3360 7630 3400
rect 7630 3360 7640 3400
rect 7580 3350 7640 3360
rect 4860 3310 4920 3320
rect 4860 3270 4870 3310
rect 4870 3270 4910 3310
rect 4910 3270 4920 3310
rect 4860 3260 4920 3270
rect 5540 3260 5600 3320
rect 6120 3310 6180 3320
rect 6120 3270 6130 3310
rect 6130 3270 6170 3310
rect 6170 3270 6180 3310
rect 6120 3260 6180 3270
rect 6720 3310 6780 3320
rect 6720 3270 6730 3310
rect 6730 3270 6770 3310
rect 6770 3270 6780 3310
rect 6720 3260 6780 3270
rect 6420 3220 6480 3230
rect 6420 3180 6430 3220
rect 6430 3180 6470 3220
rect 6470 3180 6480 3220
rect 6420 3170 6480 3180
rect 7300 3260 7360 3320
rect 7980 3310 8040 3320
rect 7980 3270 7990 3310
rect 7990 3270 8030 3310
rect 8030 3270 8040 3310
rect 7980 3260 8040 3270
rect 7840 3170 7900 3230
rect 3800 3140 4220 3150
rect 3800 3100 3810 3140
rect 3810 3100 3850 3140
rect 3850 3100 3900 3140
rect 3900 3100 3940 3140
rect 3940 3100 3990 3140
rect 3990 3100 4030 3140
rect 4030 3100 4080 3140
rect 4080 3100 4120 3140
rect 4120 3100 4170 3140
rect 4170 3100 4210 3140
rect 4210 3100 4220 3140
rect 3800 3090 4220 3100
rect 6060 3130 6120 3140
rect 6060 3090 6070 3130
rect 6070 3090 6110 3130
rect 6110 3090 6120 3130
rect 6060 3080 6120 3090
rect 6780 3130 6840 3140
rect 6780 3090 6790 3130
rect 6790 3090 6830 3130
rect 6830 3090 6840 3130
rect 6780 3080 6840 3090
rect 1730 2730 1790 2790
rect 1420 2140 1480 2200
rect 1900 2780 1960 2790
rect 1900 2740 1910 2780
rect 1910 2740 1950 2780
rect 1950 2740 1960 2780
rect 1900 2730 1960 2740
rect 3800 2780 4220 2790
rect 3800 2740 3810 2780
rect 3810 2740 3850 2780
rect 3850 2740 3900 2780
rect 3900 2740 3940 2780
rect 3940 2740 3990 2780
rect 3990 2740 4030 2780
rect 4030 2740 4080 2780
rect 4080 2740 4120 2780
rect 4120 2740 4170 2780
rect 4170 2740 4210 2780
rect 4210 2740 4220 2780
rect 3800 2730 4220 2740
rect 5540 2790 5600 2800
rect 5540 2750 5550 2790
rect 5550 2750 5590 2790
rect 5590 2750 5600 2790
rect 5540 2740 5600 2750
rect 7300 2790 7360 2800
rect 7300 2750 7310 2790
rect 7310 2750 7350 2790
rect 7350 2750 7360 2790
rect 7300 2740 7360 2750
rect 5140 2700 5200 2710
rect 5140 2660 5150 2700
rect 5150 2660 5190 2700
rect 5190 2660 5200 2700
rect 5140 2650 5200 2660
rect 5340 2700 5400 2710
rect 5340 2660 5350 2700
rect 5350 2660 5390 2700
rect 5390 2660 5400 2700
rect 5340 2650 5400 2660
rect 5740 2700 5800 2710
rect 5740 2660 5750 2700
rect 5750 2660 5790 2700
rect 5790 2660 5800 2700
rect 5740 2650 5800 2660
rect 6140 2700 6200 2710
rect 6140 2660 6150 2700
rect 6150 2660 6190 2700
rect 6190 2660 6200 2700
rect 6140 2650 6200 2660
rect 6340 2700 6400 2710
rect 6340 2660 6350 2700
rect 6350 2660 6390 2700
rect 6390 2660 6400 2700
rect 6340 2650 6400 2660
rect 6500 2700 6560 2710
rect 6500 2660 6510 2700
rect 6510 2660 6550 2700
rect 6550 2660 6560 2700
rect 6500 2650 6560 2660
rect 6700 2700 6760 2710
rect 6700 2660 6710 2700
rect 6710 2660 6750 2700
rect 6750 2660 6760 2700
rect 6700 2650 6760 2660
rect 7100 2700 7160 2710
rect 7100 2660 7110 2700
rect 7110 2660 7150 2700
rect 7150 2660 7160 2700
rect 7100 2650 7160 2660
rect 7500 2700 7560 2710
rect 7500 2660 7510 2700
rect 7510 2660 7550 2700
rect 7550 2660 7560 2700
rect 7500 2650 7560 2660
rect 7700 2700 7760 2710
rect 7700 2660 7710 2700
rect 7710 2660 7750 2700
rect 7750 2660 7760 2700
rect 7700 2650 7760 2660
rect 7300 2580 7360 2590
rect 7300 2540 7310 2580
rect 7310 2540 7350 2580
rect 7350 2540 7360 2580
rect 7300 2530 7360 2540
rect 7840 2530 7900 2590
rect 1900 2190 1960 2200
rect 1900 2150 1910 2190
rect 1910 2150 1950 2190
rect 1950 2150 1960 2190
rect 1900 2140 1960 2150
rect 4660 1640 4720 1650
rect 4660 1600 4670 1640
rect 4670 1600 4710 1640
rect 4710 1600 4720 1640
rect 4660 1590 4720 1600
rect 6420 1640 6480 1650
rect 6420 1600 6430 1640
rect 6430 1600 6470 1640
rect 6470 1600 6480 1640
rect 6420 1590 6480 1600
rect 8180 1640 8240 1650
rect 8180 1600 8190 1640
rect 8190 1600 8230 1640
rect 8230 1600 8240 1640
rect 8180 1590 8240 1600
<< metal2 >>
rect 4610 5260 4690 5270
rect 4610 5200 4620 5260
rect 4680 5250 4690 5260
rect 5010 5260 5090 5270
rect 5010 5250 5020 5260
rect 4680 5210 5020 5250
rect 4680 5200 4690 5210
rect 4610 5190 4690 5200
rect 5010 5200 5020 5210
rect 5080 5250 5090 5260
rect 5410 5260 5490 5270
rect 5410 5250 5420 5260
rect 5080 5210 5420 5250
rect 5080 5200 5090 5210
rect 5010 5190 5090 5200
rect 5410 5200 5420 5210
rect 5480 5250 5490 5260
rect 5810 5260 5890 5270
rect 5810 5250 5820 5260
rect 5480 5210 5820 5250
rect 5480 5200 5490 5210
rect 5410 5190 5490 5200
rect 5810 5200 5820 5210
rect 5880 5250 5890 5260
rect 6210 5260 6290 5270
rect 6210 5250 6220 5260
rect 5880 5210 6220 5250
rect 5880 5200 5890 5210
rect 5810 5190 5890 5200
rect 6210 5200 6220 5210
rect 6280 5250 6290 5260
rect 6610 5260 6690 5270
rect 6610 5250 6620 5260
rect 6280 5210 6620 5250
rect 6280 5200 6290 5210
rect 6210 5190 6290 5200
rect 6610 5200 6620 5210
rect 6680 5250 6690 5260
rect 7010 5260 7090 5270
rect 7010 5250 7020 5260
rect 6680 5210 7020 5250
rect 6680 5200 6690 5210
rect 6610 5190 6690 5200
rect 7010 5200 7020 5210
rect 7080 5250 7090 5260
rect 7410 5260 7490 5270
rect 7410 5250 7420 5260
rect 7080 5210 7420 5250
rect 7080 5200 7090 5210
rect 7010 5190 7090 5200
rect 7410 5200 7420 5210
rect 7480 5250 7490 5260
rect 7810 5260 7890 5270
rect 7810 5250 7820 5260
rect 7480 5210 7820 5250
rect 7480 5200 7490 5210
rect 7410 5190 7490 5200
rect 7810 5200 7820 5210
rect 7880 5250 7890 5260
rect 8210 5260 8290 5270
rect 8210 5250 8220 5260
rect 7880 5210 8220 5250
rect 7880 5200 7890 5210
rect 7810 5190 7890 5200
rect 8210 5200 8220 5210
rect 8280 5200 8290 5260
rect 8210 5190 8290 5200
rect 1190 4740 1970 4750
rect 1190 4680 1200 4740
rect 1260 4680 1900 4740
rect 1960 4680 1970 4740
rect 1190 4670 1970 4680
rect 4810 4320 4890 4330
rect 4810 4260 4820 4320
rect 4880 4310 4890 4320
rect 6810 4320 6890 4330
rect 6810 4310 6820 4320
rect 4880 4270 6820 4310
rect 4880 4260 4890 4270
rect 4810 4250 4890 4260
rect 6810 4260 6820 4270
rect 6880 4310 6890 4320
rect 7610 4320 7690 4330
rect 7610 4310 7620 4320
rect 6880 4270 7620 4310
rect 6880 4260 6890 4270
rect 6810 4250 6890 4260
rect 7610 4260 7620 4270
rect 7680 4260 7690 4320
rect 7610 4250 7690 4260
rect 5210 4230 5290 4240
rect 5210 4170 5220 4230
rect 5280 4220 5290 4230
rect 6010 4230 6090 4240
rect 6010 4220 6020 4230
rect 5280 4180 6020 4220
rect 5280 4170 5290 4180
rect 5210 4160 5290 4170
rect 6010 4170 6020 4180
rect 6080 4220 6090 4230
rect 8010 4230 8090 4240
rect 8010 4220 8020 4230
rect 6080 4180 8020 4220
rect 6080 4170 6090 4180
rect 6010 4160 6090 4170
rect 8010 4170 8020 4180
rect 8080 4170 8090 4230
rect 8010 4160 8090 4170
rect 3790 4150 4230 4160
rect 3790 4090 3800 4150
rect 4220 4130 4230 4150
rect 5610 4140 5690 4150
rect 5610 4130 5620 4140
rect 4220 4090 5620 4130
rect 3790 4080 4230 4090
rect 5610 4080 5620 4090
rect 5680 4130 5690 4140
rect 6410 4140 6490 4150
rect 6410 4130 6420 4140
rect 5680 4090 6420 4130
rect 5680 4080 5690 4090
rect 5610 4070 5690 4080
rect 6410 4080 6420 4090
rect 6480 4130 6490 4140
rect 7210 4140 7290 4150
rect 7210 4130 7220 4140
rect 6480 4090 7220 4130
rect 6480 4080 6490 4090
rect 6410 4070 6490 4080
rect 7210 4080 7220 4090
rect 7280 4080 7290 4140
rect 7210 4070 7290 4080
rect 4450 3950 4530 3960
rect 4450 3890 4460 3950
rect 4520 3940 4530 3950
rect 4650 3950 4730 3960
rect 4650 3940 4660 3950
rect 4520 3900 4660 3940
rect 4520 3890 4530 3900
rect 4450 3880 4530 3890
rect 4650 3890 4660 3900
rect 4720 3940 4730 3950
rect 5050 3950 5130 3960
rect 5050 3940 5060 3950
rect 4720 3900 5060 3940
rect 4720 3890 4730 3900
rect 4650 3880 4730 3890
rect 5050 3890 5060 3900
rect 5120 3940 5130 3950
rect 5450 3950 5530 3960
rect 5450 3940 5460 3950
rect 5120 3900 5460 3940
rect 5120 3890 5130 3900
rect 5050 3880 5130 3890
rect 5450 3890 5460 3900
rect 5520 3940 5530 3950
rect 5650 3950 5730 3960
rect 5650 3940 5660 3950
rect 5520 3900 5660 3940
rect 5520 3890 5530 3900
rect 5450 3880 5530 3890
rect 5650 3890 5660 3900
rect 5720 3940 5730 3950
rect 5810 3950 5890 3960
rect 5810 3940 5820 3950
rect 5720 3900 5820 3940
rect 5720 3890 5730 3900
rect 5650 3880 5730 3890
rect 5810 3890 5820 3900
rect 5880 3940 5890 3950
rect 6010 3950 6090 3960
rect 6010 3940 6020 3950
rect 5880 3900 6020 3940
rect 5880 3890 5890 3900
rect 5810 3880 5890 3890
rect 6010 3890 6020 3900
rect 6080 3940 6090 3950
rect 6410 3950 6490 3960
rect 6410 3940 6420 3950
rect 6080 3900 6420 3940
rect 6080 3890 6090 3900
rect 6010 3880 6090 3890
rect 6410 3890 6420 3900
rect 6480 3940 6490 3950
rect 6810 3950 6890 3960
rect 6810 3940 6820 3950
rect 6480 3900 6820 3940
rect 6480 3890 6490 3900
rect 6410 3880 6490 3890
rect 6810 3890 6820 3900
rect 6880 3940 6890 3950
rect 7010 3950 7090 3960
rect 7010 3940 7020 3950
rect 6880 3900 7020 3940
rect 6880 3890 6890 3900
rect 6810 3880 6890 3890
rect 7010 3890 7020 3900
rect 7080 3940 7090 3950
rect 7170 3950 7250 3960
rect 7170 3940 7180 3950
rect 7080 3900 7180 3940
rect 7080 3890 7090 3900
rect 7010 3880 7090 3890
rect 7170 3890 7180 3900
rect 7240 3940 7250 3950
rect 7370 3950 7450 3960
rect 7370 3940 7380 3950
rect 7240 3900 7380 3940
rect 7240 3890 7250 3900
rect 7170 3880 7250 3890
rect 7370 3890 7380 3900
rect 7440 3940 7450 3950
rect 7770 3950 7850 3960
rect 7770 3940 7780 3950
rect 7440 3900 7780 3940
rect 7440 3890 7450 3900
rect 7370 3880 7450 3890
rect 7770 3890 7780 3900
rect 7840 3940 7850 3950
rect 8170 3950 8250 3960
rect 8170 3940 8180 3950
rect 7840 3900 8180 3940
rect 7840 3890 7850 3900
rect 7770 3880 7850 3890
rect 8170 3890 8180 3900
rect 8240 3940 8250 3950
rect 8370 3950 8450 3960
rect 8370 3940 8380 3950
rect 8240 3900 8380 3940
rect 8240 3890 8250 3900
rect 8170 3880 8250 3890
rect 8370 3890 8380 3900
rect 8440 3890 8450 3950
rect 8370 3880 8450 3890
rect 1190 3740 1970 3750
rect 1190 3680 1200 3740
rect 1260 3680 1900 3740
rect 1960 3680 1970 3740
rect 1190 3670 1970 3680
rect 5250 3410 5330 3420
rect 5250 3350 5260 3410
rect 5320 3400 5330 3410
rect 5930 3410 6010 3420
rect 5930 3400 5940 3410
rect 5320 3360 5940 3400
rect 5320 3350 5330 3360
rect 5250 3340 5330 3350
rect 5930 3350 5940 3360
rect 6000 3400 6010 3410
rect 6890 3410 6970 3420
rect 6890 3400 6900 3410
rect 6000 3360 6900 3400
rect 6000 3350 6010 3360
rect 5930 3340 6010 3350
rect 6890 3350 6900 3360
rect 6960 3400 6970 3410
rect 7570 3410 7650 3420
rect 7570 3400 7580 3410
rect 6960 3360 7580 3400
rect 6960 3350 6970 3360
rect 6890 3340 6970 3350
rect 7570 3350 7580 3360
rect 7640 3350 7650 3410
rect 7570 3340 7650 3350
rect 4850 3320 4930 3330
rect 4850 3260 4860 3320
rect 4920 3310 4930 3320
rect 5530 3320 5610 3330
rect 5530 3310 5540 3320
rect 4920 3270 5540 3310
rect 4920 3260 4930 3270
rect 4850 3250 4930 3260
rect 5530 3260 5540 3270
rect 5600 3310 5610 3320
rect 6110 3320 6190 3330
rect 6110 3310 6120 3320
rect 5600 3270 6120 3310
rect 5600 3260 5610 3270
rect 5530 3250 5610 3260
rect 6110 3260 6120 3270
rect 6180 3310 6190 3320
rect 6710 3320 6790 3330
rect 6710 3310 6720 3320
rect 6180 3270 6720 3310
rect 6180 3260 6190 3270
rect 6110 3250 6190 3260
rect 6710 3260 6720 3270
rect 6780 3310 6790 3320
rect 7290 3320 7370 3330
rect 7290 3310 7300 3320
rect 6780 3270 7300 3310
rect 6780 3260 6790 3270
rect 6710 3250 6790 3260
rect 7290 3260 7300 3270
rect 7360 3310 7370 3320
rect 7970 3320 8050 3330
rect 7970 3310 7980 3320
rect 7360 3270 7980 3310
rect 7360 3260 7370 3270
rect 7290 3250 7370 3260
rect 7970 3260 7980 3270
rect 8040 3260 8050 3320
rect 7970 3250 8050 3260
rect 6410 3230 6490 3240
rect 6410 3170 6420 3230
rect 6480 3220 6490 3230
rect 7830 3230 7910 3240
rect 7830 3220 7840 3230
rect 6480 3180 7840 3220
rect 6480 3170 6490 3180
rect 6410 3160 6490 3170
rect 7830 3170 7840 3180
rect 7900 3170 7910 3230
rect 7830 3160 7910 3170
rect 880 3150 4230 3160
rect 880 3090 890 3150
rect 950 3090 3800 3150
rect 4220 3130 4230 3150
rect 6050 3140 6130 3150
rect 6050 3130 6060 3140
rect 4220 3090 6060 3130
rect 880 3080 4230 3090
rect 6050 3080 6060 3090
rect 6120 3130 6130 3140
rect 6770 3140 6850 3150
rect 6770 3130 6780 3140
rect 6120 3090 6780 3130
rect 6120 3080 6130 3090
rect 6050 3070 6130 3080
rect 6770 3080 6780 3090
rect 6840 3080 6850 3140
rect 6770 3070 6850 3080
rect 5530 2800 5610 2810
rect 1720 2790 1970 2800
rect 1720 2730 1730 2790
rect 1790 2730 1900 2790
rect 1960 2730 1970 2790
rect 1720 2720 1970 2730
rect 3790 2790 4230 2800
rect 5530 2790 5540 2800
rect 3790 2730 3800 2790
rect 4220 2750 5540 2790
rect 4220 2730 4230 2750
rect 5530 2740 5540 2750
rect 5600 2790 5610 2800
rect 7290 2800 7370 2810
rect 7290 2790 7300 2800
rect 5600 2750 7300 2790
rect 5600 2740 5610 2750
rect 5530 2730 5610 2740
rect 7290 2740 7300 2750
rect 7360 2740 7370 2800
rect 7290 2730 7370 2740
rect 3790 2720 4230 2730
rect 5130 2710 5210 2720
rect 5130 2650 5140 2710
rect 5200 2700 5210 2710
rect 5330 2710 5410 2720
rect 5330 2700 5340 2710
rect 5200 2660 5340 2700
rect 5200 2650 5210 2660
rect 5130 2640 5210 2650
rect 5330 2650 5340 2660
rect 5400 2700 5410 2710
rect 5730 2710 5810 2720
rect 5730 2700 5740 2710
rect 5400 2660 5740 2700
rect 5400 2650 5410 2660
rect 5330 2640 5410 2650
rect 5730 2650 5740 2660
rect 5800 2700 5810 2710
rect 6130 2710 6210 2720
rect 6130 2700 6140 2710
rect 5800 2660 6140 2700
rect 5800 2650 5810 2660
rect 5730 2640 5810 2650
rect 6130 2650 6140 2660
rect 6200 2700 6210 2710
rect 6330 2710 6410 2720
rect 6330 2700 6340 2710
rect 6200 2660 6340 2700
rect 6200 2650 6210 2660
rect 6130 2640 6210 2650
rect 6330 2650 6340 2660
rect 6400 2700 6410 2710
rect 6490 2710 6570 2720
rect 6490 2700 6500 2710
rect 6400 2660 6500 2700
rect 6400 2650 6410 2660
rect 6330 2640 6410 2650
rect 6490 2650 6500 2660
rect 6560 2700 6570 2710
rect 6690 2710 6770 2720
rect 6690 2700 6700 2710
rect 6560 2660 6700 2700
rect 6560 2650 6570 2660
rect 6490 2640 6570 2650
rect 6690 2650 6700 2660
rect 6760 2700 6770 2710
rect 7090 2710 7170 2720
rect 7090 2700 7100 2710
rect 6760 2660 7100 2700
rect 6760 2650 6770 2660
rect 6690 2640 6770 2650
rect 7090 2650 7100 2660
rect 7160 2700 7170 2710
rect 7490 2710 7570 2720
rect 7490 2700 7500 2710
rect 7160 2660 7500 2700
rect 7160 2650 7170 2660
rect 7090 2640 7170 2650
rect 7490 2650 7500 2660
rect 7560 2700 7570 2710
rect 7690 2710 7770 2720
rect 7690 2700 7700 2710
rect 7560 2660 7700 2700
rect 7560 2650 7570 2660
rect 7490 2640 7570 2650
rect 7690 2650 7700 2660
rect 7760 2650 7770 2710
rect 7690 2640 7770 2650
rect 7290 2590 7370 2600
rect 7290 2530 7300 2590
rect 7360 2580 7370 2590
rect 7830 2590 7910 2600
rect 7830 2580 7840 2590
rect 7360 2540 7840 2580
rect 7360 2530 7370 2540
rect 7290 2520 7370 2530
rect 7830 2530 7840 2540
rect 7900 2530 7910 2590
rect 7830 2520 7910 2530
rect 1410 2200 1970 2210
rect 1410 2140 1420 2200
rect 1480 2140 1900 2200
rect 1960 2140 1970 2200
rect 1410 2130 1970 2140
rect 4650 1650 4730 1660
rect 4650 1590 4660 1650
rect 4720 1640 4730 1650
rect 6410 1650 6490 1660
rect 6410 1640 6420 1650
rect 4720 1600 6420 1640
rect 4720 1590 4730 1600
rect 4650 1580 4730 1590
rect 6410 1590 6420 1600
rect 6480 1640 6490 1650
rect 8170 1650 8250 1660
rect 8170 1640 8180 1650
rect 6480 1600 8180 1640
rect 6480 1590 6490 1600
rect 6410 1580 6490 1590
rect 8170 1590 8180 1600
rect 8240 1590 8250 1650
rect 8170 1580 8250 1590
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0 $PDKPATH/libs.ref/sky130_fd_pr/mag
timestamp 1723858470
transform 1 0 -10 0 1 0
box 0 0 1340 1340
<< labels >>
flabel locali s 1940 1102 2058 1142 0 FreeSans 400 0 0 0 Base
port 4 nsew
flabel locali s 1963 1252 2064 1301 0 FreeSans 400 0 0 0 Collector
port 3 nsew
flabel locali s 1904 626 2152 730 0 FreeSans 400 0 0 0 Emitter
port 2 nsew
flabel locali s 3300 1102 3418 1142 0 FreeSans 400 0 0 0 Base
port 4 nsew
flabel locali s 3323 1252 3424 1301 0 FreeSans 400 0 0 0 Collector
port 3 nsew
flabel locali s 3264 626 3512 730 0 FreeSans 400 0 0 0 Emitter
port 2 nsew
flabel locali s 4660 1102 4778 1142 0 FreeSans 400 0 0 0 Base
port 4 nsew
flabel locali s 4683 1252 4784 1301 0 FreeSans 400 0 0 0 Collector
port 3 nsew
flabel locali s 4624 626 4872 730 0 FreeSans 400 0 0 0 Emitter
port 2 nsew
flabel locali s 6020 1102 6138 1142 0 FreeSans 400 0 0 0 Base
port 4 nsew
flabel locali s 6043 1252 6144 1301 0 FreeSans 400 0 0 0 Collector
port 3 nsew
flabel locali s 5984 626 6232 730 0 FreeSans 400 0 0 0 Emitter
port 2 nsew
flabel locali s 7380 1102 7498 1142 0 FreeSans 400 0 0 0 Base
port 4 nsew
flabel locali s 7403 1252 7504 1301 0 FreeSans 400 0 0 0 Collector
port 3 nsew
flabel locali s 7344 626 7592 730 0 FreeSans 400 0 0 0 Emitter
port 2 nsew
flabel locali s 8740 1102 8858 1142 0 FreeSans 400 0 0 0 Base
port 4 nsew
flabel locali s 8763 1252 8864 1301 0 FreeSans 400 0 0 0 Collector
port 3 nsew
flabel locali s 8704 626 8952 730 0 FreeSans 400 0 0 0 Emitter
port 2 nsew
<< end >>
