* PEX produced on Tue Feb 25 01:31:39 PM CET 2025 using /foss/tools/osic-multitool/iic-pex.sh with m=3 and s=1
* NGSPICE file created from full_pll_magic_3.ext - technology: sky130A

.subckt full_pll_magic_2 V_OSC VDDA GNDA F_REF I_IN
X0 GNDA.t187 a_6200_5250.t4 a_6200_5250.t5 GNDA.t186 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X1 a_5970_4630.t6 V_CONT.t8 a_6200_5250.t1 VDDA.t146 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X2 GNDA.t229 GNDA.t227 GNDA.t229 GNDA.t228 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0 ps=0 w=2 l=0.6
X3 a_7630_n1440.t0 VCO_FD_magic_0.div120_2_0.div2.t2 GNDA.t83 GNDA.t82 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X4 a_870_1400.t1 pfd_8_0.QA_b.t3 VDDA.t51 VDDA.t9 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X5 pfd_8_0.DOWN_b.t1 VDDA.t221 pfd_8_0.DOWN_PFD_b.t3 GNDA.t25 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X6 GNDA.t172 VCO_FD_magic_0.div120_2_0.div5_2_0.J.t4 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.t1 GNDA.t171 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X7 VCO_FD_magic_0.div120_2_0.div5_2_0.J.t0 VCO_FD_magic_0.div120_2_0.div24.t3 GNDA.t11 GNDA.t10 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X8 GNDA.t20 VCO_FD_magic_0.div120_2_0.div3_3_0.H.t4 VCO_FD_magic_0.div120_2_0.div3_3_0.I.t0 GNDA.t19 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X9 pfd_8_0.DOWN.t1 pfd_8_0.DOWN_b.t2 VDDA.t12 VDDA.t11 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X10 pfd_8_0.UP_input.t3 pfd_8_0.UP_b.t1 sky130_fd_pr__cap_mim_m3_1 l=6.3 w=5.2
X11 VDDA.t48 VCO_FD_magic_0.vco2_3_0.V1.t3 VCO_FD_magic_0.vco2_3_0.V4.t0 VDDA.t47 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=1.5
X12 VCO_FD_magic_0.div120_2_0.div5_2_0.J.t1 VCO_FD_magic_0.div120_2_0.div5_2_0.G.t3 VDDA.t67 VDDA.t66 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X13 VDDA.t137 pfd_8_0.opamp_out.t10 opamp_cell_4_0.VIN+.t5 VDDA.t136 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X14 opamp_cell_4_0.n_right.t1 opamp_cell_4_0.VIN+.t6 a_6320_5840.t0 GNDA.t87 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X15 opamp_cell_4_0.n_right.t2 opamp_cell_4_0.n_left.t6 VDDA.t46 VDDA.t45 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X16 pfd_8_0.opamp_out.t2 opamp_cell_4_0.n_right.t5 VDDA.t32 VDDA.t31 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X17 GNDA.t90 VCO_FD_magic_0.div120_2_0.div2_4_0.C.t4 VCO_FD_magic_0.div120_2_0.div8.t1 GNDA.t89 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X18 pfd_8_0.opamp_out.t1 a_6490_4630.t5 GNDA.t22 GNDA.t21 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X19 a_2350_1400.t0 pfd_8_0.before_Reset.t3 GNDA.t59 GNDA.t58 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X20 VDDA.t144 GNDA.t270 VCO_FD_magic_0.vco2_3_0.V4.t2 VDDA.t42 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X21 pfd_8_0.DOWN.t0 pfd_8_0.DOWN_b.t3 GNDA.t141 GNDA.t140 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X22 VCO_FD_magic_0.div120_2_0.div2_4_2.B.t0 a_7630_n1440.t3 VCO_FD_magic_0.div120_2_0.div2_4_2.A.t0 GNDA.t168 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X23 VDDA.t39 opamp_cell_4_0.p_bias.t7 opamp_cell_4_0.p_bias.t8 VDDA.t38 sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X24 a_n30_1400.t0 F_REF.t0 VDDA.t218 VDDA.t82 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X25 GNDA.t152 I_IN.t3 I_IN.t4 GNDA.t151 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X26 VDDA.t85 VCO_FD_magic_0.div120_2_0.div4.t2 a_6330_n1440.t2 VDDA.t84 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X27 GNDA.t24 pfd_8_0.QA.t3 pfd_8_0.QA_b.t0 GNDA.t23 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X28 a_6200_5250.t3 a_6200_5250.t2 GNDA.t185 GNDA.t184 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X29 a_6200_5250.t0 V_CONT.t9 a_5970_4630.t5 VDDA.t145 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X30 VDDA.t104 opamp_cell_4_0.p_bias.t9 a_5970_4630.t1 VDDA.t103 sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X31 VDDA.t183 VDDA.t180 VDDA.t182 VDDA.t181 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=0 ps=0 w=2 l=0.6
X32 GNDA.t271 loop_filter_3_0.R1_C1.t1 sky130_fd_pr__cap_mim_m3_1 l=70 w=70
X33 VCO_FD_magic_0.div120_2_0.div2_4_1.C.t2 a_8930_n1440.t3 GNDA.t122 GNDA.t121 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X34 VDDA.t179 VDDA.t177 VDDA.t179 VDDA.t178 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0 ps=0 w=2 l=0.6
X35 pfd_8_0.DOWN_input.t0 pfd_8_0.DOWN_b.t4 I_IN.t0 VDDA.t68 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X36 VDDA.t209 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.t3 VCO_FD_magic_0.div120_2_0.div3_3_0.D.t0 VDDA.t208 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X37 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.t0 VCO_FD_magic_0.div120_2_0.div8.t2 GNDA.t146 GNDA.t145 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X38 VCO_FD_magic_0.div120_2_0.div3_3_0.C.t2 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.t4 GNDA.t118 GNDA.t117 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X39 a_1910_2020.t0 pfd_8_0.QB.t3 GNDA.t15 GNDA.t14 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X40 VDDA.t14 pfd_8_0.UP_input.t4 V_CONT.t0 VDDA.t13 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X41 a_6220_5810.t8 a_6220_5810.t7 GNDA.t75 GNDA.t74 sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0.3125 ps=1.75 w=1.25 l=0.5
X42 GNDA.t92 a_7630_n1440.t4 VCO_FD_magic_0.div120_2_0.div2_4_2.C.t2 GNDA.t91 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X43 pfd_8_0.UP.t1 pfd_8_0.UP_PFD_b.t2 VDDA.t127 VDDA.t126 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X44 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.t2 VCO_FD_magic_0.div120_2_0.div8.t3 VDDA.t217 VDDA.t216 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X45 GNDA.t120 F_VCO.t2 VCO_FD_magic_0.div120_2_0.div5_2_0.I.t2 GNDA.t119 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X46 VCO_FD_magic_0.div120_2_0.div5_2_0.G.t0 VCO_FD_magic_0.div120_2_0.div24.t4 VCO_FD_magic_0.div120_2_0.div5_2_0.H.t0 GNDA.t18 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X47 a_8930_n1440.t0 V_OSC.t2 VDDA.t8 VDDA.t7 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X48 VDDA.t74 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.t2 F_VCO.t0 VDDA.t73 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X49 a_8930_n1440.t1 V_OSC.t3 GNDA.t31 GNDA.t30 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X50 GNDA.t111 VCO_FD_magic_0.div120_2_0.div5_2_0.A.t3 VCO_FD_magic_0.div120_2_0.div5_2_0.C.t1 GNDA.t110 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X51 a_6320_5840.t8 a_6220_5810.t9 GNDA.t174 GNDA.t173 sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0.3125 ps=1.75 w=1.25 l=0.5
X52 pfd_8_0.QA.t2 pfd_8_0.QA_b.t4 GNDA.t55 GNDA.t54 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X53 pfd_8_0.UP_input.t0 pfd_8_0.UP.t2 pfd_8_0.opamp_out.t4 GNDA.t86 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X54 VDDA.t37 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.t3 VCO_FD_magic_0.div120_2_0.div5_2_0.A.t2 VDDA.t36 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X55 a_5970_4630.t3 opamp_cell_4_0.p_bias.t10 VDDA.t125 VDDA.t124 sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X56 a_1390_1400.t1 pfd_8_0.E.t3 pfd_8_0.E_b.t2 VDDA.t58 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X57 pfd_8_0.DOWN_input.t2 pfd_8_0.DOWN.t3 I_IN.t5 GNDA.t41 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X58 a_870_640.t1 pfd_8_0.QB_b.t3 VDDA.t10 VDDA.t9 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X59 I_IN.t2 I_IN.t1 GNDA.t154 GNDA.t153 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X60 VCO_FD_magic_0.div120_2_0.div5_2_0.F.t1 F_VCO.t3 VCO_FD_magic_0.div120_2_0.div5_2_0.G.t2 VDDA.t195 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X61 VDDA.t176 VDDA.t173 VDDA.t175 VDDA.t174 sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0 ps=0 w=1 l=0.15
X62 VDDA.t116 a_2530_190.t2 a_2200_190.t1 VDDA.t115 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=0.15
X63 pfd_8_0.opamp_out.t11 a_9360_3514.t0 sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X64 VCO_FD_magic_0.div120_2_0.div5_2_0.B.t1 VCO_FD_magic_0.div120_2_0.div5_2_0.A.t4 VDDA.t189 VDDA.t188 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X65 GNDA.t226 GNDA.t224 GNDA.t226 GNDA.t225 sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0 ps=0 w=1.25 l=0.5
X66 GNDA.t223 GNDA.t220 GNDA.t222 GNDA.t221 sky130_fd_pr__nfet_01v8 ad=0.25 pd=2 as=0 ps=0 w=0.5 l=0.15
X67 opamp_cell_4_0.p_bias.t6 opamp_cell_4_0.p_bias.t5 VDDA.t4 VDDA.t3 sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X68 VCO_FD_magic_0.vco2_3_0.V1.t2 V_CONT.t10 GNDA.t5 GNDA.t4 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X69 VCO_FD_magic_0.vco2_3_0.V8.t1 VCO_FD_magic_0.vco2_3_0.V9.t2 VCO_FD_magic_0.vco2_3_0.V4.t1 VDDA.t42 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X70 V_CONT.t5 pfd_8_0.UP_input.t5 VDDA.t135 VDDA.t134 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X71 VDDA.t172 VDDA.t170 VDDA.t172 VDDA.t171 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0 ps=0 w=2 l=0.6
X72 V_OSC.t1 VCO_FD_magic_0.vco2_3_0.V8.t2 VCO_FD_magic_0.vco2_3_0.V3.t0 GNDA.t26 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X73 GNDA.t219 GNDA.t216 GNDA.t218 GNDA.t217 sky130_fd_pr__nfet_01v8 ad=1 pd=5 as=0 ps=0 w=2 l=0.6
X74 pfd_8_0.F.t1 pfd_8_0.QB_b.t4 GNDA.t33 GNDA.t32 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X75 GNDA.t77 a_2530_190.t3 a_2200_190.t0 GNDA.t76 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X76 pfd_8_0.DOWN_input.t1 pfd_8_0.DOWN_b.t5 GNDA.t114 GNDA.t113 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X77 GNDA.t47 VCO_FD_magic_0.div120_2_0.div24.t5 VCO_FD_magic_0.div120_2_0.div5_2_0.D.t2 GNDA.t46 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X78 GNDA.t248 VCO_FD_magic_0.div120_2_0.div2_4_2.C.t4 VCO_FD_magic_0.div120_2_0.div4.t1 GNDA.t247 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X79 GNDA.t215 GNDA.t212 GNDA.t214 GNDA.t213 sky130_fd_pr__nfet_01v8 ad=0.625 pd=3.5 as=0 ps=0 w=1.25 l=0.5
X80 VDDA.t57 a_8930_n1440.t4 VCO_FD_magic_0.div120_2_0.div2.t0 VDDA.t56 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X81 VCO_FD_magic_0.div120_2_0.div2_4_1.B.t0 a_8930_n1440.t5 VCO_FD_magic_0.div120_2_0.div2_4_1.A.t0 GNDA.t133 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X82 VCO_FD_magic_0.div120_2_0.div3_3_0.G.t0 VCO_FD_magic_0.div120_2_0.div3_3_0.I.t2 GNDA.t7 GNDA.t6 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X83 GNDA.t1 pfd_8_0.E_b.t3 pfd_8_0.E.t0 GNDA.t0 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X84 pfd_8_0.UP_b.t2 pfd_8_0.UP.t3 GNDA.t52 GNDA.t51 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X85 GNDA.t27 VDDA.t222 VCO_FD_magic_0.vco2_3_0.V3.t2 GNDA.t26 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X86 GNDA.t116 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.t4 VCO_FD_magic_0.div120_2_0.div5_2_0.M.t2 GNDA.t115 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X87 pfd_8_0.opamp_out.t12 a_9360_6440.t0 sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X88 VCO_FD_magic_0.div120_2_0.div2_4_0.A.t1 VCO_FD_magic_0.div120_2_0.div8.t4 VDDA.t94 VDDA.t93 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X89 GNDA.t135 a_6220_5810.t10 a_6320_5840.t7 GNDA.t134 sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0.3125 ps=1.75 w=1.25 l=0.5
X90 a_1390_640.t1 pfd_8_0.F.t3 pfd_8_0.F_b.t1 VDDA.t58 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X91 GNDA.t211 GNDA.t208 GNDA.t210 GNDA.t209 sky130_fd_pr__nfet_01v8 ad=1 pd=5 as=0 ps=0 w=2 l=0.6
X92 GNDA.t259 F_VCO.t4 VCO_FD_magic_0.div120_2_0.div5_2_0.L.t1 GNDA.t258 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X93 VDDA.t16 VCO_FD_magic_0.div120_2_0.div3_3_0.I.t3 VCO_FD_magic_0.div120_2_0.div3_3_0.E.t0 VDDA.t15 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X94 a_2350_1400.t1 pfd_8_0.before_Reset.t4 VDDA.t207 VDDA.t206 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=0.15
X95 VCO_FD_magic_0.div120_2_0.div5_2_0.K.t1 F_VCO.t5 VDDA.t211 VDDA.t210 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X96 GNDA.t240 a_6220_5810.t5 a_6220_5810.t6 GNDA.t239 sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0.3125 ps=1.75 w=1.25 l=0.5
X97 GNDA.t207 GNDA.t204 GNDA.t206 GNDA.t205 sky130_fd_pr__nfet_01v8 ad=1 pd=5 as=0 ps=0 w=2 l=0.6
X98 VDDA.t6 VCO_FD_magic_0.div120_2_0.div2_4_2.A.t2 VCO_FD_magic_0.div120_2_0.div2_4_2.C.t3 VDDA.t5 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X99 GNDA.t203 GNDA.t201 GNDA.t203 GNDA.t202 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0 ps=0 w=0.5 l=0.15
X100 a_5970_4630.t11 a_5970_4630.t10 a_5970_4630.t11 VDDA.t148 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0 ps=0 w=1 l=0.15
X101 VDDA.t65 pfd_8_0.UP_input.t6 V_CONT.t2 VDDA.t64 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X102 pfd_8_0.F_b.t2 pfd_8_0.F.t4 GNDA.t265 GNDA.t264 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X103 VDDA.t79 pfd_8_0.F.t5 a_490_640.t1 VDDA.t49 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X104 VDDA.t169 VDDA.t167 VDDA.t169 VDDA.t168 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0 ps=0 w=1 l=0.15
X105 pfd_8_0.QA_b.t1 pfd_8_0.QA.t4 a_n30_1400.t1 VDDA.t28 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X106 GNDA.t200 GNDA.t198 GNDA.t200 GNDA.t199 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0 ps=0 w=0.5 l=0.15
X107 GNDA.t178 VCO_FD_magic_0.div120_2_0.div8.t5 VCO_FD_magic_0.div120_2_0.div2_4_0.B.t1 GNDA.t177 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X108 GNDA.t132 VCO_FD_magic_0.div120_2_0.div24.t6 VCO_FD_magic_0.div120_2_0.div5_2_0.J.t2 GNDA.t131 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X109 GNDA.t250 pfd_8_0.F.t6 pfd_8_0.QB.t1 GNDA.t249 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X110 GNDA.t244 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.t5 VCO_FD_magic_0.div120_2_0.div3_3_0.H.t3 GNDA.t243 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X111 pfd_8_0.before_Reset.t0 pfd_8_0.QB.t4 VDDA.t18 VDDA.t17 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.805 ps=5 w=2 l=0.15
X112 GNDA.t179 V_CONT.t11 VCO_FD_magic_0.vco2_3_0.V7.t1 GNDA.t45 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X113 GNDA.t49 VDDA.t223 VCO_FD_magic_0.vco2_3_0.V5.t2 GNDA.t48 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X114 VDDA.t185 VCO_FD_magic_0.vco2_3_0.V1.t4 VCO_FD_magic_0.vco2_3_0.V2.t0 VDDA.t184 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=1.5
X115 VDDA.t100 VCO_FD_magic_0.div120_2_0.div24.t7 VCO_FD_magic_0.div120_2_0.div5_2_0.E.t0 VDDA.t99 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X116 VDDA.t1 VCO_FD_magic_0.div120_2_0.div24.t8 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.t0 VDDA.t0 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X117 GNDA.t44 a_6490_4630.t6 pfd_8_0.opamp_out.t3 GNDA.t43 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X118 VDDA.t102 opamp_cell_4_0.n_right.t6 pfd_8_0.opamp_out.t5 VDDA.t101 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X119 opamp_cell_4_0.VIN+.t4 pfd_8_0.opamp_out.t13 VDDA.t72 VDDA.t71 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X120 VDDA.t201 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.t6 VCO_FD_magic_0.div120_2_0.div3_3_0.I.t1 VDDA.t200 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X121 a_490_1400.t0 pfd_8_0.QA_b.t5 pfd_8_0.QA.t1 VDDA.t114 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X122 pfd_8_0.UP_input.t2 pfd_8_0.UP_b.t3 pfd_8_0.opamp_out.t0 VDDA.t68 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X123 V_CONT.t4 pfd_8_0.UP_input.t7 VDDA.t131 VDDA.t130 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X124 VDDA.t143 GNDA.t272 VCO_FD_magic_0.vco2_3_0.V2.t2 VDDA.t2 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X125 GNDA.t79 pfd_8_0.Reset.t2 pfd_8_0.E_b.t0 GNDA.t78 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X126 GNDA.t162 VCO_FD_magic_0.div120_2_0.div2_4_1.C.t4 VCO_FD_magic_0.div120_2_0.div2.t1 GNDA.t161 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X127 GNDA.t255 VCO_FD_magic_0.div120_2_0.div3_3_0.I.t4 VCO_FD_magic_0.div120_2_0.div24.t1 GNDA.t254 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X128 VCO_FD_magic_0.vco2_3_0.V9.t1 V_OSC.t4 VCO_FD_magic_0.vco2_3_0.V7.t0 GNDA.t45 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X129 VCO_FD_magic_0.div120_2_0.div2_4_0.C.t2 a_6330_n1440.t3 GNDA.t242 GNDA.t241 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X130 a_2530_190.t0 a_2350_1400.t2 GNDA.t148 GNDA.t147 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X131 VDDA.t76 opamp_cell_4_0.n_left.t2 opamp_cell_4_0.n_left.t3 VDDA.t75 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X132 VCO_FD_magic_0.div120_2_0.div24.t0 VCO_FD_magic_0.div120_2_0.div3_3_0.I.t5 VDDA.t92 VDDA.t91 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X133 a_6320_5840.t10 V_CONT.t12 opamp_cell_4_0.n_left.t5 GNDA.t112 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X134 a_7630_n1440.t2 VCO_FD_magic_0.div120_2_0.div2.t3 VDDA.t194 VDDA.t193 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X135 VDDA.t215 VCO_FD_magic_0.div120_2_0.div3_3_0.I.t6 VCO_FD_magic_0.div120_2_0.div24.t2 VDDA.t214 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X136 VCO_FD_magic_0.div120_2_0.div3_3_0.C.t1 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.t7 GNDA.t261 GNDA.t260 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X137 GNDA.t170 VCO_FD_magic_0.div120_2_0.div24.t9 VCO_FD_magic_0.div120_2_0.div3_3_0.B.t0 GNDA.t169 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X138 pfd_8_0.E.t1 pfd_8_0.E_b.t4 a_870_1400.t0 VDDA.t33 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X139 pfd_8_0.UP_b.t0 pfd_8_0.UP.t4 VDDA.t19 VDDA.t11 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X140 VCO_FD_magic_0.div120_2_0.div5_2_0.H.t1 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.t5 VCO_FD_magic_0.div120_2_0.div5_2_0.I.t1 GNDA.t253 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X141 pfd_8_0.DOWN_input.t3 pfd_8_0.DOWN.t2 sky130_fd_pr__cap_mim_m3_1 l=3.8 w=2.7
X142 VDDA.t107 V_OSC.t5 a_8930_n1440.t2 VDDA.t106 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X143 VDDA.t133 VCO_FD_magic_0.div120_2_0.div8.t6 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.t1 VDDA.t132 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X144 VCO_FD_magic_0.div120_2_0.div5_2_0.C.t0 VCO_FD_magic_0.div120_2_0.div24.t10 VCO_FD_magic_0.div120_2_0.div5_2_0.B.t0 GNDA.t144 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X145 a_5970_4630.t9 a_5970_4630.t7 a_5970_4630.t8 VDDA.t147 sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0 ps=0 w=1 l=0.15
X146 VCO_FD_magic_0.div120_2_0.div2_4_0.C.t1 a_6330_n1440.t4 GNDA.t128 GNDA.t127 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X147 GNDA.t197 GNDA.t194 GNDA.t196 GNDA.t195 sky130_fd_pr__nfet_01v8 ad=0.25 pd=2 as=0 ps=0 w=0.5 l=0.15
X148 VDDA.t25 a_1870_190.t2 pfd_8_0.Reset.t1 VDDA.t24 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=0.15
X149 pfd_8_0.opamp_out.t6 a_6490_4630.t7 GNDA.t126 GNDA.t125 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X150 pfd_8_0.opamp_out.t7 opamp_cell_4_0.n_right.t7 VDDA.t118 VDDA.t117 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X151 VCO_FD_magic_0.div120_2_0.div5_2_0.G.t1 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.t6 VDDA.t70 VDDA.t69 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X152 GNDA.t103 VCO_FD_magic_0.div120_2_0.div4.t3 VCO_FD_magic_0.div120_2_0.div2_4_2.B.t1 GNDA.t102 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X153 VDDA.t121 VCO_FD_magic_0.div120_2_0.div5_2_0.B.t2 VCO_FD_magic_0.div120_2_0.div5_2_0.D.t3 VDDA.t120 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X154 VDDA.t87 a_7630_n1440.t5 VCO_FD_magic_0.div120_2_0.div4.t0 VDDA.t86 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X155 VCO_FD_magic_0.div120_2_0.div2_4_0.B.t0 a_6330_n1440.t5 VCO_FD_magic_0.div120_2_0.div2_4_0.A.t0 GNDA.t84 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X156 GNDA.t35 a_1870_190.t3 pfd_8_0.Reset.t0 GNDA.t34 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X157 V_OSC.t0 VCO_FD_magic_0.vco2_3_0.V8.t3 VCO_FD_magic_0.vco2_3_0.V2.t1 VDDA.t2 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X158 VCO_FD_magic_0.div120_2_0.div2_4_1.A.t1 VCO_FD_magic_0.div120_2_0.div2.t4 VDDA.t205 VDDA.t204 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X159 VCO_FD_magic_0.div120_2_0.div3_3_0.A.t0 VCO_FD_magic_0.div120_2_0.div24.t11 VDDA.t123 VDDA.t122 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X160 VDDA.t166 VDDA.t163 VDDA.t165 VDDA.t164 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=0 ps=0 w=2 l=0.6
X161 VCO_FD_magic_0.div120_2_0.div5_2_0.D.t1 VCO_FD_magic_0.div120_2_0.div24.t12 GNDA.t17 GNDA.t16 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X162 opamp_cell_4_0.p_bias.t4 opamp_cell_4_0.p_bias.t3 VDDA.t191 VDDA.t190 sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X163 opamp_cell_4_0.p_bias.t0 a_6220_5810.t0 GNDA.t38 sky130_fd_pr__res_xhigh_po_5p73 l=1
X164 VDDA.t44 VCO_FD_magic_0.vco2_3_0.V1.t5 VCO_FD_magic_0.vco2_3_0.V6.t1 VDDA.t43 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=1.5
X165 GNDA.t109 VCO_FD_magic_0.div120_2_0.div3_3_0.C.t4 VCO_FD_magic_0.div120_2_0.div3_3_0.D.t1 GNDA.t108 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X166 VCO_FD_magic_0.div120_2_0.div3_3_0.E.t1 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.t8 VCO_FD_magic_0.div120_2_0.div3_3_0.F.t0 GNDA.t93 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X167 opamp_cell_4_0.n_left.t1 opamp_cell_4_0.n_left.t0 VDDA.t111 VDDA.t110 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X168 GNDA.t65 VCO_FD_magic_0.div120_2_0.div5_2_0.M.t4 F_VCO.t1 GNDA.t64 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X169 GNDA.t273 V_CONT.t6 sky130_fd_pr__cap_mim_m3_1 l=70 w=14
X170 opamp_cell_4_0.n_left.t4 V_CONT.t13 a_6320_5840.t9 GNDA.t175 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X171 VCO_FD_magic_0.div120_2_0.div5_2_0.L.t0 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.t7 VCO_FD_magic_0.div120_2_0.div5_2_0.K.t0 GNDA.t98 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X172 VDDA.t203 VCO_FD_magic_0.div120_2_0.div2_4_0.A.t2 VCO_FD_magic_0.div120_2_0.div2_4_0.C.t3 VDDA.t202 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X173 a_5970_4630.t4 opamp_cell_4_0.p_bias.t11 VDDA.t141 VDDA.t140 sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X174 pfd_8_0.before_Reset.t1 pfd_8_0.QA.t5 a_1910_2020.t1 GNDA.t53 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X175 pfd_8_0.UP_PFD_b.t0 pfd_8_0.QA.t6 GNDA.t40 GNDA.t39 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X176 VDDA.t142 GNDA.t274 VCO_FD_magic_0.vco2_3_0.V6.t2 VDDA.t119 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X177 VCO_FD_magic_0.div120_2_0.div2_4_2.C.t1 a_7630_n1440.t6 GNDA.t234 GNDA.t233 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X178 GNDA.t130 pfd_8_0.E.t4 pfd_8_0.QA.t0 GNDA.t129 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X179 VDDA.t60 VCO_FD_magic_0.div120_2_0.div5_2_0.K.t2 VCO_FD_magic_0.div120_2_0.div5_2_0.M.t3 VDDA.t59 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X180 a_9360_6440.t1 a_6490_4630.t4 GNDA.t176 sky130_fd_pr__res_xhigh_po_0p35 l=0.86
X181 VDDA.t162 VDDA.t160 VDDA.t162 VDDA.t161 sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0 ps=0 w=2.5 l=0.5
X182 VDDA.t63 pfd_8_0.Reset.t3 a_1390_1400.t0 VDDA.t61 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X183 pfd_8_0.F.t0 pfd_8_0.F_b.t3 a_870_640.t0 VDDA.t33 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X184 a_2530_190.t1 a_2350_1400.t3 VDDA.t197 VDDA.t196 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=0.15
X185 GNDA.t193 GNDA.t191 GNDA.t193 GNDA.t192 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0 ps=0 w=2 l=0.6
X186 GNDA.t95 a_6220_5810.t3 a_6220_5810.t4 GNDA.t94 sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0.3125 ps=1.75 w=1.25 l=0.5
X187 GNDA.t167 a_6490_4630.t8 pfd_8_0.opamp_out.t8 GNDA.t166 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X188 VDDA.t139 opamp_cell_4_0.n_right.t8 pfd_8_0.opamp_out.t9 VDDA.t138 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X189 VDDA.t159 VDDA.t156 VDDA.t158 VDDA.t157 sky130_fd_pr__pfet_01v8 ad=1.25 pd=6 as=0 ps=0 w=2.5 l=0.5
X190 GNDA.t156 a_8930_n1440.t6 VCO_FD_magic_0.div120_2_0.div2_4_1.C.t1 GNDA.t155 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X191 GNDA.t164 pfd_8_0.F_b.t4 pfd_8_0.F.t2 GNDA.t163 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X192 VCO_FD_magic_0.div120_2_0.div5_2_0.J.t3 VCO_FD_magic_0.div120_2_0.div24.t13 GNDA.t143 GNDA.t142 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X193 GNDA.t263 a_6220_5810.t11 a_6320_5840.t12 GNDA.t262 sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0.3125 ps=1.75 w=1.25 l=0.5
X194 pfd_8_0.QB_b.t1 pfd_8_0.QB.t5 a_n30_640.t0 VDDA.t28 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X195 VCO_FD_magic_0.div120_2_0.div2_4_2.C.t0 a_7630_n1440.t7 GNDA.t9 GNDA.t8 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X196 GNDA.t183 a_6200_5250.t6 a_6490_4630.t3 GNDA.t182 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X197 a_5970_4630.t0 opamp_cell_4_0.VIN+.t7 a_6490_4630.t1 VDDA.t90 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X198 VDDA.t113 opamp_cell_4_0.p_bias.t12 a_5970_4630.t2 VDDA.t112 sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X199 VCO_FD_magic_0.div120_2_0.div3_3_0.H.t2 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.t9 GNDA.t107 GNDA.t106 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X200 GNDA.t124 VCO_FD_magic_0.div120_2_0.div2.t5 VCO_FD_magic_0.div120_2_0.div2_4_1.B.t1 GNDA.t123 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X201 VDDA.t62 pfd_8_0.Reset.t4 a_1390_640.t0 VDDA.t61 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X202 VDDA.t81 opamp_cell_4_0.p_bias.t1 opamp_cell_4_0.p_bias.t2 VDDA.t80 sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X203 opamp_cell_4_0.n_right.t4 a_9360_3514.t1 GNDA.t176 sky130_fd_pr__res_xhigh_po_0p35 l=1.14
X204 pfd_8_0.UP_input.t1 pfd_8_0.UP.t5 VDDA.t96 VDDA.t95 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X205 VDDA.t155 VDDA.t152 VDDA.t154 VDDA.t153 sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0 ps=0 w=1 l=0.15
X206 a_6320_5840.t6 a_6320_5840.t4 a_6320_5840.t5 GNDA.t88 sky130_fd_pr__nfet_01v8 ad=0.25 pd=2 as=0 ps=0 w=0.5 l=0.15
X207 GNDA.t73 pfd_8_0.QB.t6 pfd_8_0.QB_b.t0 GNDA.t72 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X208 a_6320_5840.t11 a_6220_5810.t12 GNDA.t246 GNDA.t245 sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0.3125 ps=1.75 w=1.25 l=0.5
X209 GNDA.t252 pfd_8_0.Reset.t5 pfd_8_0.F_b.t0 GNDA.t251 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X210 a_6330_n1440.t1 VCO_FD_magic_0.div120_2_0.div4.t4 VDDA.t187 VDDA.t186 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X211 VCO_FD_magic_0.vco2_3_0.V9.t0 V_OSC.t6 VCO_FD_magic_0.vco2_3_0.V6.t0 VDDA.t119 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X212 GNDA.t71 pfd_8_0.DOWN_input.t4 V_CONT.t1 GNDA.t70 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X213 a_6320_5840.t3 a_6320_5840.t2 a_6320_5840.t3 GNDA.t99 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0 ps=0 w=0.5 l=0.15
X214 VDDA.t151 VDDA.t149 VDDA.t151 VDDA.t150 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0 ps=0 w=1 l=0.15
X215 a_6220_5810.t2 a_6220_5810.t1 GNDA.t257 GNDA.t256 sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0.3125 ps=1.75 w=1.25 l=0.5
X216 GNDA.t67 V_CONT.t14 VCO_FD_magic_0.vco2_3_0.V3.t1 GNDA.t26 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X217 VDDA.t213 VCO_FD_magic_0.div120_2_0.div2.t6 a_7630_n1440.t1 VDDA.t212 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X218 pfd_8_0.E.t2 pfd_8_0.QA_b.t6 GNDA.t139 GNDA.t138 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X219 GNDA.t160 I_IN.t6 opamp_cell_4_0.VIN+.t1 GNDA.t159 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X220 GNDA.t238 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.t10 VCO_FD_magic_0.div120_2_0.div3_3_0.C.t0 GNDA.t237 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X221 a_6330_n1440.t0 VCO_FD_magic_0.div120_2_0.div4.t5 GNDA.t150 GNDA.t149 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X222 VCO_FD_magic_0.div120_2_0.div3_3_0.B.t1 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.t11 VCO_FD_magic_0.div120_2_0.div3_3_0.A.t1 GNDA.t230 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X223 GNDA.t236 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.t8 VCO_FD_magic_0.div120_2_0.div5_2_0.A.t0 GNDA.t235 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X224 VDDA.t199 pfd_8_0.QA.t7 pfd_8_0.before_Reset.t2 VDDA.t198 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X225 pfd_8_0.UP_PFD_b.t1 pfd_8_0.QA.t8 VDDA.t78 VDDA.t77 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X226 a_n30_640.t1 F_VCO.t6 VDDA.t83 VDDA.t82 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X227 GNDA.t50 VDDA.t224 VCO_FD_magic_0.vco2_3_0.V7.t2 GNDA.t45 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X228 VCO_FD_magic_0.div120_2_0.div5_2_0.I.t0 VCO_FD_magic_0.div120_2_0.div5_2_0.E.t2 GNDA.t37 GNDA.t36 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X229 a_6490_4630.t2 a_6200_5250.t7 GNDA.t181 GNDA.t180 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X230 a_6490_4630.t0 opamp_cell_4_0.VIN+.t8 a_5970_4630.t12 VDDA.t192 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X231 VDDA.t23 a_6330_n1440.t6 VCO_FD_magic_0.div120_2_0.div8.t0 VDDA.t22 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X232 VCO_FD_magic_0.div120_2_0.div5_2_0.A.t1 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.t9 VDDA.t35 VDDA.t34 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X233 VDDA.t50 pfd_8_0.E.t5 a_490_1400.t1 VDDA.t49 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X234 VCO_FD_magic_0.div120_2_0.div2_4_2.A.t1 VCO_FD_magic_0.div120_2_0.div4.t6 VDDA.t55 VDDA.t54 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X235 VDDA.t220 a_2200_190.t2 a_1870_190.t1 VDDA.t219 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=0.15
X236 V_CONT.t3 loop_filter_3_0.R1_C1.t0 GNDA.t165 sky130_fd_pr__res_xhigh_po_0p35 l=6.8
X237 VDDA.t21 VCO_FD_magic_0.div120_2_0.div5_2_0.E.t3 VCO_FD_magic_0.div120_2_0.div5_2_0.F.t0 VDDA.t20 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X238 pfd_8_0.QA_b.t2 F_REF.t1 GNDA.t101 GNDA.t100 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X239 VDDA.t89 pfd_8_0.opamp_out.t14 opamp_cell_4_0.VIN+.t3 VDDA.t88 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X240 a_490_640.t0 pfd_8_0.QB_b.t5 pfd_8_0.QB.t0 VDDA.t114 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X241 V_CONT.t7 pfd_8_0.DOWN_input.t5 GNDA.t267 GNDA.t266 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X242 pfd_8_0.QB_b.t2 F_VCO.t7 GNDA.t97 GNDA.t96 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X243 VCO_FD_magic_0.div120_2_0.div5_2_0.M.t1 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.t10 GNDA.t69 GNDA.t68 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X244 VCO_FD_magic_0.div120_2_0.div2_4_1.C.t0 a_8930_n1440.t7 GNDA.t232 GNDA.t231 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X245 VDDA.t98 VCO_FD_magic_0.div120_2_0.div2_4_1.A.t2 VCO_FD_magic_0.div120_2_0.div2_4_1.C.t3 VDDA.t97 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X246 VDDA.t129 VCO_FD_magic_0.div120_2_0.div3_3_0.A.t2 VCO_FD_magic_0.div120_2_0.div3_3_0.C.t3 VDDA.t128 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X247 VCO_FD_magic_0.vco2_3_0.V8.t0 VCO_FD_magic_0.vco2_3_0.V9.t3 VCO_FD_magic_0.vco2_3_0.V5.t0 GNDA.t48 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X248 GNDA.t63 a_2200_190.t3 a_1870_190.t0 GNDA.t62 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X249 GNDA.t3 VCO_FD_magic_0.div120_2_0.div5_2_0.D.t4 VCO_FD_magic_0.div120_2_0.div5_2_0.E.t1 GNDA.t2 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X250 VCO_FD_magic_0.div120_2_0.div5_2_0.D.t0 VCO_FD_magic_0.div120_2_0.div24.t14 GNDA.t81 GNDA.t80 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X251 opamp_cell_4_0.VIN+.t0 I_IN.t7 GNDA.t158 GNDA.t157 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X252 a_6320_5840.t1 opamp_cell_4_0.VIN+.t9 opamp_cell_4_0.n_right.t0 GNDA.t42 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X253 VDDA.t109 opamp_cell_4_0.n_left.t7 opamp_cell_4_0.n_right.t3 VDDA.t108 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X254 pfd_8_0.DOWN_PFD_b.t1 pfd_8_0.QB.t7 VDDA.t105 VDDA.t77 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X255 pfd_8_0.QB.t2 pfd_8_0.QB_b.t6 GNDA.t269 GNDA.t268 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X256 GNDA.t66 V_CONT.t15 VCO_FD_magic_0.vco2_3_0.V5.t1 GNDA.t48 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X257 VCO_FD_magic_0.div120_2_0.div3_3_0.F.t1 VCO_FD_magic_0.div120_2_0.div3_3_0.D.t2 VCO_FD_magic_0.div120_2_0.div3_3_0.G.t1 GNDA.t85 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X258 VCO_FD_magic_0.div120_2_0.div3_3_0.H.t0 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.t12 GNDA.t13 GNDA.t12 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X259 VCO_FD_magic_0.div120_2_0.div5_2_0.M.t0 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.t11 GNDA.t57 GNDA.t56 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X260 pfd_8_0.UP.t0 pfd_8_0.UP_PFD_b.t3 GNDA.t29 GNDA.t28 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X261 VCO_FD_magic_0.div120_2_0.div3_3_0.E.t2 VCO_FD_magic_0.div120_2_0.div3_3_0.D.t3 VDDA.t41 VDDA.t40 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X262 VCO_FD_magic_0.div120_2_0.div3_3_0.H.t1 VCO_FD_magic_0.div120_2_0.div3_3_0.E.t3 VDDA.t27 VDDA.t26 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X263 GNDA.t190 GNDA.t188 GNDA.t190 GNDA.t189 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0 ps=0 w=2 l=0.6
X264 pfd_8_0.E_b.t1 pfd_8_0.E.t6 GNDA.t137 GNDA.t136 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X265 pfd_8_0.DOWN_PFD_b.t0 pfd_8_0.QB.t8 GNDA.t61 GNDA.t60 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X266 VCO_FD_magic_0.vco2_3_0.V1.t1 VCO_FD_magic_0.vco2_3_0.V1.t0 VDDA.t30 VDDA.t29 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=1.5
X267 opamp_cell_4_0.VIN+.t2 pfd_8_0.opamp_out.t15 VDDA.t53 VDDA.t52 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X268 pfd_8_0.DOWN_b.t0 GNDA.t275 pfd_8_0.DOWN_PFD_b.t2 VDDA.t126 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X269 GNDA.t105 a_6330_n1440.t7 VCO_FD_magic_0.div120_2_0.div2_4_0.C.t0 GNDA.t104 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
R0 a_6200_5250.n4 a_6200_5250.n0 427.647
R1 a_6200_5250.n1 a_6200_5250.t6 321.334
R2 a_6200_5250.n5 a_6200_5250.n4 210.601
R3 a_6200_5250.n2 a_6200_5250.n1 208.868
R4 a_6200_5250.n3 a_6200_5250.t2 174.056
R5 a_6200_5250.n4 a_6200_5250.n3 152
R6 a_6200_5250.n1 a_6200_5250.t7 112.468
R7 a_6200_5250.n2 a_6200_5250.t4 112.468
R8 a_6200_5250.n3 a_6200_5250.n2 61.5894
R9 a_6200_5250.t5 a_6200_5250.n5 60.0005
R10 a_6200_5250.n5 a_6200_5250.t3 60.0005
R11 a_6200_5250.n0 a_6200_5250.t1 49.2505
R12 a_6200_5250.n0 a_6200_5250.t0 49.2505
R13 GNDA.n725 GNDA.n724 337993
R14 GNDA.n724 GNDA.n723 309276
R15 GNDA.n207 GNDA.n24 204624
R16 GNDA.n725 GNDA.n23 164874
R17 GNDA.n495 GNDA.n494 36300
R18 GNDA.n493 GNDA.t86 10524.4
R19 GNDA.n131 GNDA.t165 1824.86
R20 GNDA.n558 GNDA.n60 1204.13
R21 GNDA.n533 GNDA.n532 1204.13
R22 GNDA.n426 GNDA.n425 1204.13
R23 GNDA.n253 GNDA.n252 1186
R24 GNDA.n206 GNDA.n205 1186
R25 GNDA.n199 GNDA.n198 1186
R26 GNDA.n260 GNDA.n259 1186
R27 GNDA.n689 GNDA.n688 1182.8
R28 GNDA.n50 GNDA.n25 1182.8
R29 GNDA.n498 GNDA.n497 1173.78
R30 GNDA.n169 GNDA.n112 1173.78
R31 GNDA.n123 GNDA.n122 1173.78
R32 GNDA.n132 GNDA.n131 1170
R33 GNDA.t235 GNDA.t25 800
R34 GNDA.n299 GNDA.t100 783.001
R35 GNDA.t119 GNDA.t10 776.471
R36 GNDA.n123 GNDA.t272 728.524
R37 GNDA.n497 GNDA.t274 728.524
R38 GNDA.n112 GNDA.t270 728.524
R39 GNDA.n131 GNDA.n23 726.415
R40 GNDA.n126 GNDA.n120 686.717
R41 GNDA.n500 GNDA.n499 686.717
R42 GNDA.n168 GNDA.n167 686.717
R43 GNDA.n168 GNDA.n114 686.717
R44 GNDA.n499 GNDA.n111 686.717
R45 GNDA.n125 GNDA.n120 686.717
R46 GNDA.n530 GNDA.n529 669.307
R47 GNDA.n527 GNDA.n73 669.307
R48 GNDA.n464 GNDA.n463 669.307
R49 GNDA.n467 GNDA.n466 669.307
R50 GNDA.n491 GNDA.n490 669.307
R51 GNDA.n485 GNDA.n369 669.307
R52 GNDA.t108 GNDA.t93 613.048
R53 GNDA.t0 GNDA.t136 601.333
R54 GNDA.t23 GNDA.t54 601.333
R55 GNDA.n728 GNDA.n727 585.003
R56 GNDA.n298 GNDA.n297 585.003
R57 GNDA.n295 GNDA.n294 585.001
R58 GNDA.n293 GNDA.n279 585.001
R59 GNDA.n292 GNDA.n276 585.001
R60 GNDA.n273 GNDA.n272 585.001
R61 GNDA.n251 GNDA.n250 585.001
R62 GNDA.n208 GNDA.n207 585.001
R63 GNDA.n368 GNDA.n367 585.001
R64 GNDA.n270 GNDA.n264 585.001
R65 GNDA.n271 GNDA.n267 585.001
R66 GNDA.n722 GNDA.n721 585.001
R67 GNDA.n36 GNDA.n31 585.001
R68 GNDA.n691 GNDA.n690 585.001
R69 GNDA.n733 GNDA.n732 585.001
R70 GNDA.n731 GNDA.n19 585.001
R71 GNDA.n730 GNDA.n16 585.001
R72 GNDA.n729 GNDA.n13 585.001
R73 GNDA.n726 GNDA.n2 585.001
R74 GNDA.n489 GNDA.n427 585
R75 GNDA.n487 GNDA.n486 585
R76 GNDA.n442 GNDA.n438 585
R77 GNDA.n440 GNDA.n437 585
R78 GNDA.n77 GNDA.n74 585
R79 GNDA.n80 GNDA.n79 585
R80 GNDA.n99 GNDA.n98 585
R81 GNDA.n100 GNDA.n99 585
R82 GNDA.n97 GNDA.n95 585
R83 GNDA.n93 GNDA.n91 585
R84 GNDA.n102 GNDA.n101 585
R85 GNDA.n101 GNDA.n100 585
R86 GNDA.n704 GNDA.t275 566.966
R87 GNDA.n100 GNDA.t260 522.179
R88 GNDA.t34 GNDA.t18 517.648
R89 GNDA.t254 GNDA.n36 482.353
R90 GNDA.t64 GNDA.n725 482.353
R91 GNDA.t76 GNDA.n731 458.825
R92 GNDA.t86 GNDA.t51 425.334
R93 GNDA.t147 GNDA.n271 418
R94 GNDA.n690 GNDA.t60 388.236
R95 GNDA.t217 GNDA.t266 376.654
R96 GNDA.t98 GNDA.t72 376.471
R97 GNDA.t209 GNDA.n531 359.534
R98 GNDA.n368 GNDA.t28 344.668
R99 GNDA.t39 GNDA.n270 344.668
R100 GNDA.n75 GNDA.t227 336.329
R101 GNDA.n75 GNDA.t208 336.329
R102 GNDA.n439 GNDA.t188 336.329
R103 GNDA.n439 GNDA.t216 336.329
R104 GNDA.t268 GNDA.t258 329.413
R105 GNDA.n103 GNDA.t204 320.7
R106 GNDA.n484 GNDA.t191 320.7
R107 GNDA.n689 GNDA.t110 317.647
R108 GNDA.t82 GNDA.t192 316.733
R109 GNDA.t159 GNDA.t149 316.733
R110 GNDA.t145 GNDA.t153 316.733
R111 GNDA.n532 GNDA.t189 308.171
R112 GNDA.t151 GNDA.n60 308.171
R113 GNDA.t2 GNDA.t34 305.882
R114 GNDA.n170 GNDA.t198 304.634
R115 GNDA.n254 GNDA.t220 304.634
R116 GNDA.n204 GNDA.t194 304.634
R117 GNDA.n200 GNDA.t201 304.634
R118 GNDA.n635 GNDA.t259 295.933
R119 GNDA.n607 GNDA.t236 295.933
R120 GNDA.n42 GNDA.t255 295.933
R121 GNDA.n249 GNDA.t224 292.584
R122 GNDA.n209 GNDA.t212 292.584
R123 GNDA.n492 GNDA.n426 291.051
R124 GNDA.t53 GNDA.n292 286
R125 GNDA.t41 GNDA.n25 270.589
R126 GNDA.n126 GNDA.t67 260
R127 GNDA.t67 GNDA.n125 260
R128 GNDA.t85 GNDA.t6 258.825
R129 GNDA.n722 GNDA.n25 258.825
R130 GNDA.t243 GNDA.t12 258.825
R131 GNDA.t19 GNDA.t106 258.825
R132 GNDA.t80 GNDA.t46 258.825
R133 GNDA.t249 GNDA.t268 258.825
R134 GNDA.t258 GNDA.t98 258.825
R135 GNDA.t56 GNDA.t64 258.825
R136 GNDA.n640 GNDA.n637 256.207
R137 GNDA.n492 GNDA.n491 250.349
R138 GNDA.n492 GNDA.n369 250.349
R139 GNDA.n465 GNDA.n464 250.349
R140 GNDA.n466 GNDA.n465 250.349
R141 GNDA.n531 GNDA.n530 250.349
R142 GNDA.n531 GNDA.n73 250.349
R143 GNDA.n100 GNDA.n94 250.349
R144 GNDA.n639 GNDA.n638 247.934
R145 GNDA.n631 GNDA.n630 247.934
R146 GNDA.n656 GNDA.n629 247.934
R147 GNDA.n663 GNDA.n626 247.934
R148 GNDA.n675 GNDA.n621 247.934
R149 GNDA.n619 GNDA.n618 247.934
R150 GNDA.n45 GNDA.n44 247.934
R151 GNDA.n595 GNDA.n47 247.934
R152 GNDA.n576 GNDA.n575 247.934
R153 GNDA.n573 GNDA.n55 247.934
R154 GNDA.t16 GNDA.n730 247.06
R155 GNDA.n561 GNDA.n560 246.714
R156 GNDA.n259 GNDA.t200 245
R157 GNDA.n253 GNDA.t223 245
R158 GNDA.n205 GNDA.t197 245
R159 GNDA.n199 GNDA.t203 245
R160 GNDA.n169 GNDA.n168 241.643
R161 GNDA.n499 GNDA.n498 241.643
R162 GNDA.n122 GNDA.n120 241.643
R163 GNDA.t140 GNDA.t243 235.294
R164 GNDA.n690 GNDA.n689 235.294
R165 GNDA.n124 GNDA.t27 233
R166 GNDA.n688 GNDA.t111 233
R167 GNDA.n50 GNDA.t7 233
R168 GNDA.n496 GNDA.t50 233
R169 GNDA.n113 GNDA.t49 233
R170 GNDA.t51 GNDA.n368 227.333
R171 GNDA.n270 GNDA.t28 227.333
R172 GNDA.n271 GNDA.t39 227.333
R173 GNDA.n552 GNDA.n63 219.133
R174 GNDA.n65 GNDA.n64 219.133
R175 GNDA.n540 GNDA.n69 219.133
R176 GNDA.n405 GNDA.n404 219.133
R177 GNDA.n411 GNDA.n402 219.133
R178 GNDA.n419 GNDA.n399 219.133
R179 GNDA.n393 GNDA.n373 219.133
R180 GNDA.n387 GNDA.n386 219.133
R181 GNDA.n379 GNDA.n378 219.133
R182 GNDA.t62 GNDA.t16 211.766
R183 GNDA.t171 GNDA.t249 211.766
R184 GNDA.t72 GNDA.t68 211.766
R185 GNDA.t96 GNDA.t115 211.766
R186 GNDA.n295 GNDA.n293 205.333
R187 GNDA.n256 GNDA.n172 204.201
R188 GNDA.n202 GNDA.n196 204.201
R189 GNDA.n203 GNDA.n195 204.201
R190 GNDA.n201 GNDA.n197 204.201
R191 GNDA.n255 GNDA.n173 204.201
R192 GNDA.n258 GNDA.n257 204.201
R193 GNDA.n732 GNDA.t144 200
R194 GNDA.n3 GNDA.t73 198.058
R195 GNDA.n774 GNDA.t269 198.058
R196 GNDA.n762 GNDA.t164 198.058
R197 GNDA.n11 GNDA.t265 198.058
R198 GNDA.n324 GNDA.t137 198.058
R199 GNDA.n319 GNDA.t1 198.058
R200 GNDA.n289 GNDA.t55 198.058
R201 GNDA.n305 GNDA.t24 198.058
R202 GNDA.n272 GNDA.t147 198
R203 GNDA.n292 GNDA.t58 198
R204 GNDA.n293 GNDA.t14 198
R205 GNDA.t78 GNDA.n295 198
R206 GNDA.n298 GNDA.t138 198
R207 GNDA.t129 GNDA.n298 198
R208 GNDA.n79 GNDA.n74 197
R209 GNDA.n438 GNDA.n437 197
R210 GNDA.n486 GNDA.n427 197
R211 GNDA.n99 GNDA.n95 197
R212 GNDA.n101 GNDA.n93 197
R213 GNDA.t4 GNDA.n23 189.173
R214 GNDA.t168 GNDA.t102 188.327
R215 GNDA.t91 GNDA.t233 188.327
R216 GNDA.t8 GNDA.t247 188.327
R217 GNDA.t177 GNDA.t84 188.327
R218 GNDA.t241 GNDA.t104 188.327
R219 GNDA.t127 GNDA.t89 188.327
R220 GNDA.t230 GNDA.t169 188.327
R221 GNDA.t237 GNDA.t117 188.327
R222 GNDA.t117 GNDA.t108 188.327
R223 GNDA.t93 GNDA.t113 188.236
R224 GNDA.t12 GNDA.t41 188.236
R225 GNDA.n529 GNDA.n528 185
R226 GNDA.n528 GNDA.n527 185
R227 GNDA.n463 GNDA.n436 185
R228 GNDA.n467 GNDA.n436 185
R229 GNDA.n490 GNDA.n428 185
R230 GNDA.n485 GNDA.n428 185
R231 GNDA.n98 GNDA.n92 185
R232 GNDA.n102 GNDA.n92 185
R233 GNDA.n529 GNDA.n75 166.63
R234 GNDA.n463 GNDA.n439 166.63
R235 GNDA.t253 GNDA.t251 164.707
R236 GNDA.t36 GNDA.t264 164.707
R237 GNDA.t163 GNDA.t131 164.707
R238 GNDA.t32 GNDA.t142 164.707
R239 GNDA.t228 GNDA.t127 162.647
R240 GNDA.t14 GNDA.t53 161.333
R241 GNDA.t136 GNDA.t78 161.333
R242 GNDA.t138 GNDA.t0 161.333
R243 GNDA.t54 GNDA.t129 161.333
R244 GNDA.t100 GNDA.t23 161.333
R245 GNDA.n729 GNDA.t253 152.941
R246 GNDA.t142 GNDA.n728 152.941
R247 GNDA.n726 GNDA.t56 152.941
R248 GNDA.n465 GNDA.t8 145.525
R249 GNDA.n531 GNDA.t241 145.525
R250 GNDA.n723 GNDA.t260 145.525
R251 GNDA.n134 GNDA.n133 142.694
R252 GNDA.n724 GNDA.t58 139.333
R253 GNDA.n250 GNDA.t226 134.501
R254 GNDA.n208 GNDA.t215 134.501
R255 GNDA.n7 GNDA.t250 130.713
R256 GNDA.n169 GNDA.t26 130.319
R257 GNDA.n498 GNDA.t48 130.319
R258 GNDA.n2 GNDA.t97 130.001
R259 GNDA.n13 GNDA.t252 130.001
R260 GNDA.n16 GNDA.t35 130.001
R261 GNDA.n19 GNDA.t63 130.001
R262 GNDA.n733 GNDA.t77 130.001
R263 GNDA.n299 GNDA.t101 130.001
R264 GNDA.n294 GNDA.t79 130.001
R265 GNDA.n279 GNDA.t15 130.001
R266 GNDA.n276 GNDA.t59 130.001
R267 GNDA.n273 GNDA.t148 130.001
R268 GNDA.n8 GNDA.t33 130.001
R269 GNDA.n296 GNDA.t139 130.001
R270 GNDA.n288 GNDA.t130 130.001
R271 GNDA.t45 GNDA.t30 128.917
R272 GNDA.n121 GNDA.t5 128.562
R273 GNDA.t102 GNDA.t70 128.405
R274 GNDA.t233 GNDA.t217 128.405
R275 GNDA.t157 GNDA.t177 128.405
R276 GNDA.t169 GNDA.t205 128.405
R277 GNDA.n166 GNDA.t66 127.754
R278 GNDA.n110 GNDA.t179 127.754
R279 GNDA.n691 GNDA.t61 122.501
R280 GNDA.n31 GNDA.t141 122.501
R281 GNDA.n721 GNDA.t114 122.501
R282 GNDA.n267 GNDA.t40 122.501
R283 GNDA.n264 GNDA.t29 122.501
R284 GNDA.n367 GNDA.t52 122.501
R285 GNDA.t60 GNDA.t235 117.647
R286 GNDA.t144 GNDA.t76 117.647
R287 GNDA.n493 GNDA.t161 111.284
R288 GNDA.n36 GNDA.t19 105.882
R289 GNDA.t18 GNDA.n729 105.882
R290 GNDA.n728 GNDA.t171 105.882
R291 GNDA.t115 GNDA.n726 105.882
R292 GNDA.t121 GNDA.t155 100.001
R293 GNDA.t155 GNDA.t231 100.001
R294 GNDA.n177 GNDA.n176 97.8707
R295 GNDA.n181 GNDA.n180 97.8707
R296 GNDA.n185 GNDA.n184 97.8707
R297 GNDA.n189 GNDA.n188 97.8707
R298 GNDA.n194 GNDA.n193 97.8707
R299 GNDA.t251 GNDA.t36 94.1181
R300 GNDA.t264 GNDA.t119 94.1181
R301 GNDA.t10 GNDA.t163 94.1181
R302 GNDA.t131 GNDA.t32 94.1181
R303 GNDA.n474 GNDA.n473 92.2612
R304 GNDA.n482 GNDA.n481 92.2612
R305 GNDA.n460 GNDA.n459 92.2612
R306 GNDA.n453 GNDA.n448 92.2612
R307 GNDA.n521 GNDA.n87 92.2612
R308 GNDA.n515 GNDA.n90 92.2612
R309 GNDA.n528 GNDA.n78 91.3721
R310 GNDA.n86 GNDA.n76 91.3721
R311 GNDA.n86 GNDA.n81 91.3721
R312 GNDA.n441 GNDA.n436 91.3721
R313 GNDA.n462 GNDA.n461 91.3721
R314 GNDA.n461 GNDA.n435 91.3721
R315 GNDA.n488 GNDA.n428 90.7567
R316 GNDA.n96 GNDA.n92 90.7567
R317 GNDA.n251 GNDA.t99 89.0971
R318 GNDA.n491 GNDA.n427 84.306
R319 GNDA.n486 GNDA.n369 84.306
R320 GNDA.n464 GNDA.n438 84.306
R321 GNDA.n466 GNDA.n437 84.306
R322 GNDA.n530 GNDA.n74 84.306
R323 GNDA.n79 GNDA.n73 84.306
R324 GNDA.n95 GNDA.n94 84.306
R325 GNDA.n94 GNDA.n93 84.306
R326 GNDA.n202 GNDA.n201 83.2005
R327 GNDA.n203 GNDA.n202 83.2005
R328 GNDA.n132 GNDA.t271 82.8829
R329 GNDA.n133 GNDA.t273 81.6029
R330 GNDA.n724 GNDA.n24 80.6672
R331 GNDA.n198 GNDA.t74 77.6744
R332 GNDA.n252 GNDA.t221 75.3899
R333 GNDA.n260 GNDA.t199 75.2337
R334 GNDA.t74 GNDA.t88 70.8209
R335 GNDA.t113 GNDA.t85 70.5887
R336 GNDA.n206 GNDA.t213 68.5363
R337 GNDA.t192 GNDA.n426 68.483
R338 GNDA.n532 GNDA.t159 68.483
R339 GNDA.t153 GNDA.n60 68.483
R340 GNDA.n257 GNDA.n256 66.5605
R341 GNDA.n256 GNDA.n255 66.5605
R342 GNDA.n272 GNDA.n24 66.0005
R343 GNDA.n256 GNDA.n171 65.9634
R344 GNDA.t239 GNDA.t202 61.6827
R345 GNDA.n734 GNDA.n733 60.29
R346 GNDA.n741 GNDA.n19 60.29
R347 GNDA.n747 GNDA.n16 60.29
R348 GNDA.n754 GNDA.n13 60.29
R349 GNDA.n782 GNDA.n2 60.29
R350 GNDA.n300 GNDA.n299 60.29
R351 GNDA.n294 GNDA.n282 60.29
R352 GNDA.n332 GNDA.n279 60.29
R353 GNDA.n339 GNDA.n276 60.29
R354 GNDA.n345 GNDA.n273 60.29
R355 GNDA.n172 GNDA.t126 60.0005
R356 GNDA.n172 GNDA.t167 60.0005
R357 GNDA.n196 GNDA.t181 60.0005
R358 GNDA.n196 GNDA.t187 60.0005
R359 GNDA.n195 GNDA.t185 60.0005
R360 GNDA.n195 GNDA.t196 60.0005
R361 GNDA.t203 GNDA.n197 60.0005
R362 GNDA.n197 GNDA.t183 60.0005
R363 GNDA.n173 GNDA.t22 60.0005
R364 GNDA.n173 GNDA.t222 60.0005
R365 GNDA.t200 GNDA.n258 60.0005
R366 GNDA.n258 GNDA.t44 60.0005
R367 GNDA.t70 GNDA.t82 59.9227
R368 GNDA.t266 GNDA.t168 59.9227
R369 GNDA.t149 GNDA.t157 59.9227
R370 GNDA.t84 GNDA.t209 59.9227
R371 GNDA.t205 GNDA.t145 59.9227
R372 GNDA.n353 GNDA.n267 59.5478
R373 GNDA.n360 GNDA.n264 59.5478
R374 GNDA.n367 GNDA.n366 59.5478
R375 GNDA.n252 GNDA.n251 59.3982
R376 GNDA.t112 GNDA.t87 59.3982
R377 GNDA.t182 GNDA.t180 59.3982
R378 GNDA.t184 GNDA.t195 59.3982
R379 GNDA.t221 GNDA.t21 59.3367
R380 GNDA.t43 GNDA.t199 59.2751
R381 GNDA.t125 GNDA.t43 59.2751
R382 GNDA.t166 GNDA.t125 59.2751
R383 GNDA.t21 GNDA.t166 59.2751
R384 GNDA.n494 GNDA.t121 59.0914
R385 GNDA.n709 GNDA.n31 58.9809
R386 GNDA.n692 GNDA.n691 58.9809
R387 GNDA.n721 GNDA.n720 58.9809
R388 GNDA.t6 GNDA.n722 58.824
R389 GNDA.n732 GNDA.t110 58.824
R390 GNDA.t42 GNDA.t225 57.1137
R391 GNDA.t134 GNDA.t186 57.1137
R392 GNDA.n767 GNDA.n8 54.4005
R393 GNDA.n769 GNDA.n7 54.4005
R394 GNDA.n688 GNDA.n687 54.4005
R395 GNDA.n589 GNDA.n50 54.4005
R396 GNDA.n313 GNDA.n288 54.4005
R397 GNDA.n296 GNDA.n287 54.4005
R398 GNDA.t175 GNDA.t173 52.5446
R399 GNDA.n637 GNDA.t57 48.0005
R400 GNDA.n637 GNDA.t65 48.0005
R401 GNDA.n638 GNDA.t69 48.0005
R402 GNDA.n638 GNDA.t116 48.0005
R403 GNDA.n630 GNDA.t143 48.0005
R404 GNDA.n630 GNDA.t172 48.0005
R405 GNDA.n629 GNDA.t11 48.0005
R406 GNDA.n629 GNDA.t132 48.0005
R407 GNDA.n626 GNDA.t37 48.0005
R408 GNDA.n626 GNDA.t120 48.0005
R409 GNDA.n621 GNDA.t17 48.0005
R410 GNDA.n621 GNDA.t3 48.0005
R411 GNDA.n618 GNDA.t81 48.0005
R412 GNDA.n618 GNDA.t47 48.0005
R413 GNDA.n44 GNDA.t107 48.0005
R414 GNDA.n44 GNDA.t20 48.0005
R415 GNDA.n47 GNDA.t13 48.0005
R416 GNDA.n47 GNDA.t244 48.0005
R417 GNDA.n575 GNDA.t118 48.0005
R418 GNDA.n575 GNDA.t109 48.0005
R419 GNDA.n55 GNDA.t261 48.0005
R420 GNDA.n55 GNDA.t238 48.0005
R421 GNDA.n560 GNDA.t146 48.0005
R422 GNDA.n560 GNDA.t170 48.0005
R423 GNDA.n63 GNDA.t128 48.0005
R424 GNDA.n63 GNDA.t90 48.0005
R425 GNDA.n64 GNDA.t242 48.0005
R426 GNDA.n64 GNDA.t105 48.0005
R427 GNDA.n69 GNDA.t150 48.0005
R428 GNDA.n69 GNDA.t178 48.0005
R429 GNDA.n404 GNDA.t9 48.0005
R430 GNDA.n404 GNDA.t248 48.0005
R431 GNDA.n402 GNDA.t234 48.0005
R432 GNDA.n402 GNDA.t92 48.0005
R433 GNDA.n399 GNDA.t83 48.0005
R434 GNDA.n399 GNDA.t103 48.0005
R435 GNDA.n373 GNDA.t232 48.0005
R436 GNDA.n373 GNDA.t162 48.0005
R437 GNDA.n386 GNDA.t122 48.0005
R438 GNDA.n386 GNDA.t156 48.0005
R439 GNDA.n378 GNDA.t31 48.0005
R440 GNDA.n378 GNDA.t124 48.0005
R441 GNDA.t25 GNDA.t254 47.0593
R442 GNDA.t46 GNDA.t62 47.0593
R443 GNDA.t68 GNDA.t96 47.0593
R444 GNDA.t161 GNDA.n492 42.8021
R445 GNDA.n465 GNDA.t91 42.8021
R446 GNDA.n100 GNDA.t230 42.8021
R447 GNDA.n723 GNDA.t237 42.8021
R448 GNDA.n202 GNDA.n191 41.6005
R449 GNDA.n510 GNDA.n509 41.3005
R450 GNDA.n494 GNDA.n260 41.0368
R451 GNDA.t231 GNDA.n493 40.9096
R452 GNDA.n135 GNDA.n134 39.4989
R453 GNDA.n246 GNDA.n171 39.4985
R454 GNDA.t133 GNDA.t176 39.2362
R455 GNDA.t94 GNDA.t175 38.8375
R456 GNDA.n122 GNDA.t4 37.8349
R457 GNDA.n122 GNDA.t26 37.8349
R458 GNDA.t48 GNDA.n169 37.8349
R459 GNDA.n498 GNDA.t45 37.8349
R460 GNDA.n496 GNDA.n111 35.6576
R461 GNDA.n501 GNDA.n500 35.6576
R462 GNDA.n167 GNDA.n165 35.6576
R463 GNDA.n114 GNDA.n113 35.6576
R464 GNDA.t176 GNDA.n494 35.0323
R465 GNDA.n125 GNDA.n124 34.3278
R466 GNDA.n147 GNDA.n126 34.3278
R467 GNDA.t262 GNDA.t42 34.2684
R468 GNDA.t186 GNDA.t245 34.2684
R469 GNDA.n783 GNDA.n782 33.0991
R470 GNDA.n300 GNDA.n0 33.0991
R471 GNDA.n474 GNDA.n472 32.0005
R472 GNDA.n472 GNDA.n432 32.0005
R473 GNDA.n480 GNDA.n479 32.0005
R474 GNDA.n479 GNDA.n430 32.0005
R475 GNDA.n475 GNDA.n430 32.0005
R476 GNDA.n443 GNDA.n434 32.0005
R477 GNDA.n458 GNDA.n446 32.0005
R478 GNDA.n454 GNDA.n446 32.0005
R479 GNDA.n454 GNDA.n453 32.0005
R480 GNDA.n452 GNDA.n449 32.0005
R481 GNDA.n449 GNDA.n82 32.0005
R482 GNDA.n526 GNDA.n83 32.0005
R483 GNDA.n522 GNDA.n83 32.0005
R484 GNDA.n520 GNDA.n88 32.0005
R485 GNDA.n516 GNDA.n88 32.0005
R486 GNDA.n514 GNDA.n104 32.0005
R487 GNDA.n719 GNDA.n27 32.0005
R488 GNDA.n715 GNDA.n27 32.0005
R489 GNDA.n715 GNDA.n714 32.0005
R490 GNDA.n714 GNDA.n713 32.0005
R491 GNDA.n713 GNDA.n29 32.0005
R492 GNDA.n709 GNDA.n29 32.0005
R493 GNDA.n709 GNDA.n708 32.0005
R494 GNDA.n708 GNDA.n707 32.0005
R495 GNDA.n707 GNDA.n32 32.0005
R496 GNDA.n702 GNDA.n32 32.0005
R497 GNDA.n702 GNDA.n701 32.0005
R498 GNDA.n701 GNDA.n700 32.0005
R499 GNDA.n700 GNDA.n34 32.0005
R500 GNDA.n696 GNDA.n695 32.0005
R501 GNDA.n695 GNDA.n694 32.0005
R502 GNDA.n694 GNDA.n22 32.0005
R503 GNDA.n735 GNDA.n22 32.0005
R504 GNDA.n739 GNDA.n20 32.0005
R505 GNDA.n740 GNDA.n739 32.0005
R506 GNDA.n742 GNDA.n17 32.0005
R507 GNDA.n746 GNDA.n17 32.0005
R508 GNDA.n749 GNDA.n748 32.0005
R509 GNDA.n749 GNDA.n14 32.0005
R510 GNDA.n753 GNDA.n14 32.0005
R511 GNDA.n756 GNDA.n755 32.0005
R512 GNDA.n756 GNDA.n11 32.0005
R513 GNDA.n760 GNDA.n11 32.0005
R514 GNDA.n761 GNDA.n760 32.0005
R515 GNDA.n762 GNDA.n761 32.0005
R516 GNDA.n762 GNDA.n9 32.0005
R517 GNDA.n766 GNDA.n9 32.0005
R518 GNDA.n770 GNDA.n5 32.0005
R519 GNDA.n774 GNDA.n5 32.0005
R520 GNDA.n775 GNDA.n774 32.0005
R521 GNDA.n776 GNDA.n775 32.0005
R522 GNDA.n776 GNDA.n3 32.0005
R523 GNDA.n780 GNDA.n3 32.0005
R524 GNDA.n781 GNDA.n780 32.0005
R525 GNDA.n148 GNDA.n118 32.0005
R526 GNDA.n152 GNDA.n118 32.0005
R527 GNDA.n153 GNDA.n152 32.0005
R528 GNDA.n154 GNDA.n153 32.0005
R529 GNDA.n154 GNDA.n115 32.0005
R530 GNDA.n380 GNDA.n376 32.0005
R531 GNDA.n384 GNDA.n376 32.0005
R532 GNDA.n385 GNDA.n384 32.0005
R533 GNDA.n388 GNDA.n385 32.0005
R534 GNDA.n392 GNDA.n374 32.0005
R535 GNDA.n395 GNDA.n394 32.0005
R536 GNDA.n395 GNDA.n370 32.0005
R537 GNDA.n424 GNDA.n371 32.0005
R538 GNDA.n420 GNDA.n371 32.0005
R539 GNDA.n418 GNDA.n417 32.0005
R540 GNDA.n417 GNDA.n400 32.0005
R541 GNDA.n413 GNDA.n400 32.0005
R542 GNDA.n413 GNDA.n412 32.0005
R543 GNDA.n410 GNDA.n403 32.0005
R544 GNDA.n406 GNDA.n72 32.0005
R545 GNDA.n534 GNDA.n72 32.0005
R546 GNDA.n538 GNDA.n70 32.0005
R547 GNDA.n539 GNDA.n538 32.0005
R548 GNDA.n541 GNDA.n67 32.0005
R549 GNDA.n545 GNDA.n67 32.0005
R550 GNDA.n546 GNDA.n545 32.0005
R551 GNDA.n547 GNDA.n546 32.0005
R552 GNDA.n551 GNDA.n550 32.0005
R553 GNDA.n553 GNDA.n61 32.0005
R554 GNDA.n557 GNDA.n61 32.0005
R555 GNDA.n562 GNDA.n559 32.0005
R556 GNDA.n566 GNDA.n58 32.0005
R557 GNDA.n567 GNDA.n566 32.0005
R558 GNDA.n568 GNDA.n567 32.0005
R559 GNDA.n568 GNDA.n56 32.0005
R560 GNDA.n572 GNDA.n56 32.0005
R561 GNDA.n577 GNDA.n574 32.0005
R562 GNDA.n581 GNDA.n53 32.0005
R563 GNDA.n582 GNDA.n581 32.0005
R564 GNDA.n583 GNDA.n582 32.0005
R565 GNDA.n583 GNDA.n51 32.0005
R566 GNDA.n587 GNDA.n51 32.0005
R567 GNDA.n588 GNDA.n587 32.0005
R568 GNDA.n590 GNDA.n48 32.0005
R569 GNDA.n594 GNDA.n48 32.0005
R570 GNDA.n597 GNDA.n596 32.0005
R571 GNDA.n601 GNDA.n600 32.0005
R572 GNDA.n602 GNDA.n601 32.0005
R573 GNDA.n606 GNDA.n605 32.0005
R574 GNDA.n608 GNDA.n606 32.0005
R575 GNDA.n612 GNDA.n40 32.0005
R576 GNDA.n613 GNDA.n612 32.0005
R577 GNDA.n614 GNDA.n613 32.0005
R578 GNDA.n614 GNDA.n37 32.0005
R579 GNDA.n686 GNDA.n38 32.0005
R580 GNDA.n682 GNDA.n38 32.0005
R581 GNDA.n682 GNDA.n681 32.0005
R582 GNDA.n681 GNDA.n680 32.0005
R583 GNDA.n677 GNDA.n676 32.0005
R584 GNDA.n674 GNDA.n622 32.0005
R585 GNDA.n670 GNDA.n622 32.0005
R586 GNDA.n670 GNDA.n669 32.0005
R587 GNDA.n669 GNDA.n668 32.0005
R588 GNDA.n668 GNDA.n624 32.0005
R589 GNDA.n664 GNDA.n624 32.0005
R590 GNDA.n662 GNDA.n661 32.0005
R591 GNDA.n661 GNDA.n627 32.0005
R592 GNDA.n657 GNDA.n627 32.0005
R593 GNDA.n655 GNDA.n654 32.0005
R594 GNDA.n651 GNDA.n650 32.0005
R595 GNDA.n650 GNDA.n649 32.0005
R596 GNDA.n649 GNDA.n633 32.0005
R597 GNDA.n645 GNDA.n644 32.0005
R598 GNDA.n644 GNDA.n643 32.0005
R599 GNDA.n643 GNDA.n636 32.0005
R600 GNDA.n165 GNDA.n116 32.0005
R601 GNDA.n161 GNDA.n116 32.0005
R602 GNDA.n161 GNDA.n160 32.0005
R603 GNDA.n160 GNDA.n159 32.0005
R604 GNDA.n159 GNDA.n109 32.0005
R605 GNDA.n501 GNDA.n107 32.0005
R606 GNDA.n505 GNDA.n107 32.0005
R607 GNDA.n366 GNDA.n365 32.0005
R608 GNDA.n365 GNDA.n262 32.0005
R609 GNDA.n361 GNDA.n262 32.0005
R610 GNDA.n359 GNDA.n358 32.0005
R611 GNDA.n358 GNDA.n265 32.0005
R612 GNDA.n354 GNDA.n265 32.0005
R613 GNDA.n352 GNDA.n351 32.0005
R614 GNDA.n351 GNDA.n268 32.0005
R615 GNDA.n347 GNDA.n268 32.0005
R616 GNDA.n347 GNDA.n346 32.0005
R617 GNDA.n344 GNDA.n274 32.0005
R618 GNDA.n340 GNDA.n274 32.0005
R619 GNDA.n338 GNDA.n337 32.0005
R620 GNDA.n337 GNDA.n277 32.0005
R621 GNDA.n333 GNDA.n277 32.0005
R622 GNDA.n331 GNDA.n330 32.0005
R623 GNDA.n330 GNDA.n280 32.0005
R624 GNDA.n326 GNDA.n325 32.0005
R625 GNDA.n325 GNDA.n324 32.0005
R626 GNDA.n324 GNDA.n283 32.0005
R627 GNDA.n320 GNDA.n283 32.0005
R628 GNDA.n320 GNDA.n319 32.0005
R629 GNDA.n319 GNDA.n318 32.0005
R630 GNDA.n318 GNDA.n285 32.0005
R631 GNDA.n312 GNDA.n311 32.0005
R632 GNDA.n311 GNDA.n289 32.0005
R633 GNDA.n307 GNDA.n289 32.0005
R634 GNDA.n307 GNDA.n306 32.0005
R635 GNDA.n306 GNDA.n305 32.0005
R636 GNDA.n305 GNDA.n291 32.0005
R637 GNDA.n301 GNDA.n291 32.0005
R638 GNDA.n246 GNDA.n245 32.0005
R639 GNDA.n245 GNDA.n244 32.0005
R640 GNDA.n244 GNDA.n175 32.0005
R641 GNDA.n240 GNDA.n175 32.0005
R642 GNDA.n240 GNDA.n239 32.0005
R643 GNDA.n239 GNDA.n238 32.0005
R644 GNDA.n238 GNDA.n179 32.0005
R645 GNDA.n234 GNDA.n179 32.0005
R646 GNDA.n234 GNDA.n233 32.0005
R647 GNDA.n233 GNDA.n232 32.0005
R648 GNDA.n232 GNDA.n183 32.0005
R649 GNDA.n228 GNDA.n183 32.0005
R650 GNDA.n228 GNDA.n227 32.0005
R651 GNDA.n227 GNDA.n226 32.0005
R652 GNDA.n226 GNDA.n187 32.0005
R653 GNDA.n222 GNDA.n221 32.0005
R654 GNDA.n221 GNDA.n220 32.0005
R655 GNDA.n220 GNDA.n192 32.0005
R656 GNDA.n215 GNDA.n192 32.0005
R657 GNDA.n215 GNDA.n214 32.0005
R658 GNDA.n214 GNDA.n213 32.0005
R659 GNDA.n136 GNDA.n135 32.0005
R660 GNDA.n136 GNDA.n129 32.0005
R661 GNDA.n140 GNDA.n129 32.0005
R662 GNDA.n141 GNDA.n140 32.0005
R663 GNDA.n142 GNDA.n141 32.0005
R664 GNDA.n142 GNDA.n127 32.0005
R665 GNDA.n146 GNDA.n127 32.0005
R666 GNDA.t123 GNDA.t133 30.8285
R667 GNDA.t202 GNDA.t256 29.6994
R668 GNDA.t256 GNDA.t182 29.6994
R669 GNDA.n506 GNDA.n505 29.4625
R670 GNDA.n527 GNDA.n526 29.0291
R671 GNDA.n468 GNDA.n467 29.0291
R672 GNDA.n380 GNDA.n379 28.8005
R673 GNDA.n419 GNDA.n418 28.8005
R674 GNDA.n541 GNDA.n540 28.8005
R675 GNDA.n562 GNDA.n561 28.8005
R676 GNDA.n597 GNDA.n45 28.8005
R677 GNDA.n608 GNDA.n607 28.8005
R678 GNDA.n639 GNDA.n636 28.8005
R679 GNDA.n361 GNDA.n360 28.8005
R680 GNDA.n345 GNDA.n344 28.8005
R681 GNDA.n254 GNDA.n253 27.2005
R682 GNDA.n259 GNDA.n170 27.2005
R683 GNDA.t247 GNDA.t189 25.6814
R684 GNDA.t104 GNDA.t228 25.6814
R685 GNDA.t89 GNDA.t151 25.6814
R686 GNDA.n468 GNDA.n434 25.6005
R687 GNDA.n521 GNDA.n520 25.6005
R688 GNDA.n516 GNDA.n515 25.6005
R689 GNDA.n720 GNDA.n719 25.6005
R690 GNDA.n692 GNDA.n34 25.6005
R691 GNDA.n734 GNDA.n20 25.6005
R692 GNDA.n747 GNDA.n746 25.6005
R693 GNDA.n754 GNDA.n753 25.6005
R694 GNDA.n768 GNDA.n767 25.6005
R695 GNDA.n148 GNDA.n147 25.6005
R696 GNDA.n393 GNDA.n392 25.6005
R697 GNDA.n405 GNDA.n403 25.6005
R698 GNDA.n552 GNDA.n551 25.6005
R699 GNDA.n577 GNDA.n576 25.6005
R700 GNDA.n677 GNDA.n619 25.6005
R701 GNDA.n663 GNDA.n662 25.6005
R702 GNDA.n654 GNDA.n631 25.6005
R703 GNDA.n645 GNDA.n635 25.6005
R704 GNDA.n354 GNDA.n353 25.6005
R705 GNDA.n333 GNDA.n332 25.6005
R706 GNDA.n282 GNDA.n280 25.6005
R707 GNDA.n314 GNDA.n287 25.6005
R708 GNDA.n314 GNDA.n313 25.6005
R709 GNDA.n205 GNDA.n204 25.6005
R710 GNDA.n200 GNDA.n199 25.6005
R711 GNDA.n222 GNDA.n191 25.6005
R712 GNDA.n213 GNDA 25.6005
R713 GNDA.t87 GNDA.t262 25.1303
R714 GNDA.n250 GNDA.n249 24.8279
R715 GNDA.n209 GNDA.n208 24.8279
R716 GNDA.n176 GNDA.t226 24.0005
R717 GNDA.n176 GNDA.t263 24.0005
R718 GNDA.n180 GNDA.t174 24.0005
R719 GNDA.n180 GNDA.t95 24.0005
R720 GNDA.n184 GNDA.t75 24.0005
R721 GNDA.n184 GNDA.t240 24.0005
R722 GNDA.n188 GNDA.t257 24.0005
R723 GNDA.n188 GNDA.t135 24.0005
R724 GNDA.n193 GNDA.t246 24.0005
R725 GNDA.n193 GNDA.t214 24.0005
R726 GNDA.t106 GNDA.t140 23.5299
R727 GNDA.n377 GNDA.n106 23.1831
R728 GNDA.n207 GNDA.n206 22.8458
R729 GNDA.t30 GNDA.n495 22.4209
R730 GNDA.n769 GNDA.n768 22.4005
R731 GNDA.n425 GNDA.n424 22.4005
R732 GNDA.n533 GNDA.n70 22.4005
R733 GNDA.n559 GNDA.n558 22.4005
R734 GNDA.n595 GNDA.n594 22.4005
R735 GNDA.n484 GNDA.n483 20.9665
R736 GNDA.t88 GNDA.t94 20.5612
R737 GNDA.n507 GNDA.n506 19.4202
R738 GNDA.n459 GNDA.n443 19.2005
R739 GNDA.n459 GNDA.n458 19.2005
R740 GNDA.n388 GNDA.n387 19.2005
R741 GNDA.n412 GNDA.n411 19.2005
R742 GNDA.n547 GNDA.n65 19.2005
R743 GNDA.n573 GNDA.n572 19.2005
R744 GNDA.n590 GNDA.n589 19.2005
R745 GNDA.n605 GNDA.n42 19.2005
R746 GNDA.n675 GNDA.n674 19.2005
R747 GNDA.n657 GNDA.n656 19.2005
R748 GNDA.n339 GNDA.n338 19.2005
R749 GNDA.n147 GNDA.n146 19.2005
R750 GNDA.n741 GNDA.n740 16.0005
R751 GNDA.n742 GNDA.n741 16.0005
R752 GNDA.n687 GNDA.n37 16.0005
R753 GNDA.n687 GNDA.n686 16.0005
R754 GNDA.n211 GNDA 15.7005
R755 GNDA.n485 GNDA.n484 15.6449
R756 GNDA.n103 GNDA.n102 15.6449
R757 GNDA.n473 GNDA.t267 15.0005
R758 GNDA.n473 GNDA.t218 15.0005
R759 GNDA.n481 GNDA.t193 15.0005
R760 GNDA.n481 GNDA.t71 15.0005
R761 GNDA.t190 GNDA.n460 15.0005
R762 GNDA.n460 GNDA.t160 15.0005
R763 GNDA.n448 GNDA.t158 15.0005
R764 GNDA.n448 GNDA.t210 15.0005
R765 GNDA.n87 GNDA.t229 15.0005
R766 GNDA.n87 GNDA.t152 15.0005
R767 GNDA.n90 GNDA.t154 15.0005
R768 GNDA.n90 GNDA.t206 15.0005
R769 GNDA.t229 GNDA.n86 15.0005
R770 GNDA.n528 GNDA.t211 15.0005
R771 GNDA.n461 GNDA.t190 15.0005
R772 GNDA.n436 GNDA.t219 15.0005
R773 GNDA.t193 GNDA.n428 15.0005
R774 GNDA.n92 GNDA.t207 15.0005
R775 GNDA.n104 GNDA.n103 14.4005
R776 GNDA.t38 GNDA.t184 14.1646
R777 GNDA.n255 GNDA.n254 14.0805
R778 GNDA.n257 GNDA.n170 14.0805
R779 GNDA.n720 GNDA.n26 13.9181
R780 GNDA.n198 GNDA.t239 13.7077
R781 GNDA.n211 GNDA.n105 13.1958
R782 GNDA.n261 GNDA.n105 12.8163
R783 GNDA.n468 GNDA.n432 12.8005
R784 GNDA.n482 GNDA.n480 12.8005
R785 GNDA.n522 GNDA.n521 12.8005
R786 GNDA.n515 GNDA.n514 12.8005
R787 GNDA.n165 GNDA.n115 12.8005
R788 GNDA.n387 GNDA.n374 12.8005
R789 GNDA.n411 GNDA.n410 12.8005
R790 GNDA.n550 GNDA.n65 12.8005
R791 GNDA.n574 GNDA.n573 12.8005
R792 GNDA.n589 GNDA.n588 12.8005
R793 GNDA.n602 GNDA.n42 12.8005
R794 GNDA.n676 GNDA.n675 12.8005
R795 GNDA.n656 GNDA.n655 12.8005
R796 GNDA.n501 GNDA.n109 12.8005
R797 GNDA.n340 GNDA.n339 12.8005
R798 GNDA.n204 GNDA.n203 12.8005
R799 GNDA.n201 GNDA.n200 12.8005
R800 GNDA GNDA.n0 12.7806
R801 GNDA GNDA.n783 11.8829
R802 GNDA.n731 GNDA.t80 11.7652
R803 GNDA.n730 GNDA.t2 11.7652
R804 GNDA.n507 GNDA.n26 11.7212
R805 GNDA.n509 GNDA.n508 11.6542
R806 GNDA.t245 GNDA.t38 10.9662
R807 GNDA.n379 GNDA.n377 10.7016
R808 GNDA.n640 GNDA.n639 10.4505
R809 GNDA.n770 GNDA.n769 9.6005
R810 GNDA.n425 GNDA.n370 9.6005
R811 GNDA.n534 GNDA.n533 9.6005
R812 GNDA.n558 GNDA.n557 9.6005
R813 GNDA.n596 GNDA.n595 9.6005
R814 GNDA.n249 GNDA.n248 9.58175
R815 GNDA.n217 GNDA.n209 9.58175
R816 GNDA.n641 GNDA.n636 9.3005
R817 GNDA.n643 GNDA.n642 9.3005
R818 GNDA.n644 GNDA.n634 9.3005
R819 GNDA.n646 GNDA.n645 9.3005
R820 GNDA.n647 GNDA.n633 9.3005
R821 GNDA.n649 GNDA.n648 9.3005
R822 GNDA.n650 GNDA.n632 9.3005
R823 GNDA.n652 GNDA.n651 9.3005
R824 GNDA.n654 GNDA.n653 9.3005
R825 GNDA.n655 GNDA.n628 9.3005
R826 GNDA.n658 GNDA.n657 9.3005
R827 GNDA.n659 GNDA.n627 9.3005
R828 GNDA.n661 GNDA.n660 9.3005
R829 GNDA.n662 GNDA.n625 9.3005
R830 GNDA.n665 GNDA.n664 9.3005
R831 GNDA.n666 GNDA.n624 9.3005
R832 GNDA.n668 GNDA.n667 9.3005
R833 GNDA.n669 GNDA.n623 9.3005
R834 GNDA.n671 GNDA.n670 9.3005
R835 GNDA.n672 GNDA.n622 9.3005
R836 GNDA.n674 GNDA.n673 9.3005
R837 GNDA.n676 GNDA.n620 9.3005
R838 GNDA.n678 GNDA.n677 9.3005
R839 GNDA.n680 GNDA.n679 9.3005
R840 GNDA.n681 GNDA.n617 9.3005
R841 GNDA.n683 GNDA.n682 9.3005
R842 GNDA.n684 GNDA.n38 9.3005
R843 GNDA.n686 GNDA.n685 9.3005
R844 GNDA.n616 GNDA.n37 9.3005
R845 GNDA.n615 GNDA.n614 9.3005
R846 GNDA.n613 GNDA.n39 9.3005
R847 GNDA.n612 GNDA.n611 9.3005
R848 GNDA.n610 GNDA.n40 9.3005
R849 GNDA.n609 GNDA.n608 9.3005
R850 GNDA.n606 GNDA.n41 9.3005
R851 GNDA.n605 GNDA.n604 9.3005
R852 GNDA.n603 GNDA.n602 9.3005
R853 GNDA.n601 GNDA.n43 9.3005
R854 GNDA.n600 GNDA.n599 9.3005
R855 GNDA.n598 GNDA.n597 9.3005
R856 GNDA.n596 GNDA.n46 9.3005
R857 GNDA.n594 GNDA.n593 9.3005
R858 GNDA.n592 GNDA.n48 9.3005
R859 GNDA.n591 GNDA.n590 9.3005
R860 GNDA.n588 GNDA.n49 9.3005
R861 GNDA.n587 GNDA.n586 9.3005
R862 GNDA.n585 GNDA.n51 9.3005
R863 GNDA.n584 GNDA.n583 9.3005
R864 GNDA.n582 GNDA.n52 9.3005
R865 GNDA.n581 GNDA.n580 9.3005
R866 GNDA.n579 GNDA.n53 9.3005
R867 GNDA.n578 GNDA.n577 9.3005
R868 GNDA.n574 GNDA.n54 9.3005
R869 GNDA.n572 GNDA.n571 9.3005
R870 GNDA.n570 GNDA.n56 9.3005
R871 GNDA.n569 GNDA.n568 9.3005
R872 GNDA.n567 GNDA.n57 9.3005
R873 GNDA.n566 GNDA.n565 9.3005
R874 GNDA.n564 GNDA.n58 9.3005
R875 GNDA.n563 GNDA.n562 9.3005
R876 GNDA.n559 GNDA.n59 9.3005
R877 GNDA.n557 GNDA.n556 9.3005
R878 GNDA.n555 GNDA.n61 9.3005
R879 GNDA.n554 GNDA.n553 9.3005
R880 GNDA.n551 GNDA.n62 9.3005
R881 GNDA.n550 GNDA.n549 9.3005
R882 GNDA.n548 GNDA.n547 9.3005
R883 GNDA.n546 GNDA.n66 9.3005
R884 GNDA.n545 GNDA.n544 9.3005
R885 GNDA.n543 GNDA.n67 9.3005
R886 GNDA.n542 GNDA.n541 9.3005
R887 GNDA.n539 GNDA.n68 9.3005
R888 GNDA.n538 GNDA.n537 9.3005
R889 GNDA.n536 GNDA.n70 9.3005
R890 GNDA.n535 GNDA.n534 9.3005
R891 GNDA.n72 GNDA.n71 9.3005
R892 GNDA.n407 GNDA.n406 9.3005
R893 GNDA.n408 GNDA.n403 9.3005
R894 GNDA.n410 GNDA.n409 9.3005
R895 GNDA.n412 GNDA.n401 9.3005
R896 GNDA.n414 GNDA.n413 9.3005
R897 GNDA.n415 GNDA.n400 9.3005
R898 GNDA.n417 GNDA.n416 9.3005
R899 GNDA.n418 GNDA.n398 9.3005
R900 GNDA.n421 GNDA.n420 9.3005
R901 GNDA.n422 GNDA.n371 9.3005
R902 GNDA.n424 GNDA.n423 9.3005
R903 GNDA.n397 GNDA.n370 9.3005
R904 GNDA.n396 GNDA.n395 9.3005
R905 GNDA.n394 GNDA.n372 9.3005
R906 GNDA.n392 GNDA.n391 9.3005
R907 GNDA.n390 GNDA.n374 9.3005
R908 GNDA.n389 GNDA.n388 9.3005
R909 GNDA.n385 GNDA.n375 9.3005
R910 GNDA.n384 GNDA.n383 9.3005
R911 GNDA.n382 GNDA.n376 9.3005
R912 GNDA.n381 GNDA.n380 9.3005
R913 GNDA.n149 GNDA.n148 9.3005
R914 GNDA.n150 GNDA.n118 9.3005
R915 GNDA.n152 GNDA.n151 9.3005
R916 GNDA.n153 GNDA.n117 9.3005
R917 GNDA.n155 GNDA.n154 9.3005
R918 GNDA.n156 GNDA.n115 9.3005
R919 GNDA.n163 GNDA.n116 9.3005
R920 GNDA.n162 GNDA.n161 9.3005
R921 GNDA.n160 GNDA.n157 9.3005
R922 GNDA.n159 GNDA.n158 9.3005
R923 GNDA.n109 GNDA.n108 9.3005
R924 GNDA.n505 GNDA.n504 9.3005
R925 GNDA.n503 GNDA.n107 9.3005
R926 GNDA.n502 GNDA.n501 9.3005
R927 GNDA.n165 GNDA.n164 9.3005
R928 GNDA.n315 GNDA.n314 9.3005
R929 GNDA.n302 GNDA.n301 9.3005
R930 GNDA.n303 GNDA.n291 9.3005
R931 GNDA.n305 GNDA.n304 9.3005
R932 GNDA.n306 GNDA.n290 9.3005
R933 GNDA.n308 GNDA.n307 9.3005
R934 GNDA.n309 GNDA.n289 9.3005
R935 GNDA.n311 GNDA.n310 9.3005
R936 GNDA.n312 GNDA.n286 9.3005
R937 GNDA.n316 GNDA.n285 9.3005
R938 GNDA.n318 GNDA.n317 9.3005
R939 GNDA.n319 GNDA.n284 9.3005
R940 GNDA.n321 GNDA.n320 9.3005
R941 GNDA.n322 GNDA.n283 9.3005
R942 GNDA.n324 GNDA.n323 9.3005
R943 GNDA.n325 GNDA.n281 9.3005
R944 GNDA.n327 GNDA.n326 9.3005
R945 GNDA.n328 GNDA.n280 9.3005
R946 GNDA.n330 GNDA.n329 9.3005
R947 GNDA.n331 GNDA.n278 9.3005
R948 GNDA.n334 GNDA.n333 9.3005
R949 GNDA.n335 GNDA.n277 9.3005
R950 GNDA.n337 GNDA.n336 9.3005
R951 GNDA.n338 GNDA.n275 9.3005
R952 GNDA.n341 GNDA.n340 9.3005
R953 GNDA.n342 GNDA.n274 9.3005
R954 GNDA.n344 GNDA.n343 9.3005
R955 GNDA.n346 GNDA.n269 9.3005
R956 GNDA.n348 GNDA.n347 9.3005
R957 GNDA.n349 GNDA.n268 9.3005
R958 GNDA.n351 GNDA.n350 9.3005
R959 GNDA.n352 GNDA.n266 9.3005
R960 GNDA.n355 GNDA.n354 9.3005
R961 GNDA.n356 GNDA.n265 9.3005
R962 GNDA.n358 GNDA.n357 9.3005
R963 GNDA.n359 GNDA.n263 9.3005
R964 GNDA.n362 GNDA.n361 9.3005
R965 GNDA.n363 GNDA.n262 9.3005
R966 GNDA.n365 GNDA.n364 9.3005
R967 GNDA.n247 GNDA.n246 9.3005
R968 GNDA.n245 GNDA.n174 9.3005
R969 GNDA.n244 GNDA.n243 9.3005
R970 GNDA.n242 GNDA.n175 9.3005
R971 GNDA.n241 GNDA.n240 9.3005
R972 GNDA.n239 GNDA.n178 9.3005
R973 GNDA.n238 GNDA.n237 9.3005
R974 GNDA.n236 GNDA.n179 9.3005
R975 GNDA.n235 GNDA.n234 9.3005
R976 GNDA.n233 GNDA.n182 9.3005
R977 GNDA.n232 GNDA.n231 9.3005
R978 GNDA.n230 GNDA.n183 9.3005
R979 GNDA.n229 GNDA.n228 9.3005
R980 GNDA.n227 GNDA.n186 9.3005
R981 GNDA.n226 GNDA.n225 9.3005
R982 GNDA.n224 GNDA.n187 9.3005
R983 GNDA.n223 GNDA.n222 9.3005
R984 GNDA.n221 GNDA.n190 9.3005
R985 GNDA.n220 GNDA.n219 9.3005
R986 GNDA.n218 GNDA.n192 9.3005
R987 GNDA.n216 GNDA.n215 9.3005
R988 GNDA.n214 GNDA.n210 9.3005
R989 GNDA.n213 GNDA.n212 9.3005
R990 GNDA.n147 GNDA.n119 9.3005
R991 GNDA.n135 GNDA.n130 9.3005
R992 GNDA.n137 GNDA.n136 9.3005
R993 GNDA.n138 GNDA.n129 9.3005
R994 GNDA.n140 GNDA.n139 9.3005
R995 GNDA.n141 GNDA.n128 9.3005
R996 GNDA.n143 GNDA.n142 9.3005
R997 GNDA.n144 GNDA.n127 9.3005
R998 GNDA.n146 GNDA.n145 9.3005
R999 GNDA.n511 GNDA.n510 9.3005
R1000 GNDA.n512 GNDA.n104 9.3005
R1001 GNDA.n514 GNDA.n513 9.3005
R1002 GNDA.n515 GNDA.n89 9.3005
R1003 GNDA.n517 GNDA.n516 9.3005
R1004 GNDA.n518 GNDA.n88 9.3005
R1005 GNDA.n520 GNDA.n519 9.3005
R1006 GNDA.n521 GNDA.n85 9.3005
R1007 GNDA.n523 GNDA.n522 9.3005
R1008 GNDA.n524 GNDA.n83 9.3005
R1009 GNDA.n526 GNDA.n525 9.3005
R1010 GNDA.n480 GNDA.n429 9.3005
R1011 GNDA.n479 GNDA.n478 9.3005
R1012 GNDA.n477 GNDA.n430 9.3005
R1013 GNDA.n476 GNDA.n475 9.3005
R1014 GNDA.n474 GNDA.n431 9.3005
R1015 GNDA.n472 GNDA.n471 9.3005
R1016 GNDA.n470 GNDA.n432 9.3005
R1017 GNDA.n469 GNDA.n468 9.3005
R1018 GNDA.n434 GNDA.n433 9.3005
R1019 GNDA.n444 GNDA.n443 9.3005
R1020 GNDA.n459 GNDA.n445 9.3005
R1021 GNDA.n458 GNDA.n457 9.3005
R1022 GNDA.n456 GNDA.n446 9.3005
R1023 GNDA.n455 GNDA.n454 9.3005
R1024 GNDA.n453 GNDA.n447 9.3005
R1025 GNDA.n452 GNDA.n451 9.3005
R1026 GNDA.n450 GNDA.n449 9.3005
R1027 GNDA.n84 GNDA.n82 9.3005
R1028 GNDA.n719 GNDA.n718 9.3005
R1029 GNDA.n717 GNDA.n27 9.3005
R1030 GNDA.n716 GNDA.n715 9.3005
R1031 GNDA.n714 GNDA.n28 9.3005
R1032 GNDA.n713 GNDA.n712 9.3005
R1033 GNDA.n711 GNDA.n29 9.3005
R1034 GNDA.n710 GNDA.n709 9.3005
R1035 GNDA.n708 GNDA.n30 9.3005
R1036 GNDA.n707 GNDA.n706 9.3005
R1037 GNDA.n705 GNDA.n32 9.3005
R1038 GNDA.n703 GNDA.n702 9.3005
R1039 GNDA.n701 GNDA.n33 9.3005
R1040 GNDA.n700 GNDA.n699 9.3005
R1041 GNDA.n698 GNDA.n34 9.3005
R1042 GNDA.n697 GNDA.n696 9.3005
R1043 GNDA.n695 GNDA.n35 9.3005
R1044 GNDA.n694 GNDA.n693 9.3005
R1045 GNDA.n22 GNDA.n21 9.3005
R1046 GNDA.n736 GNDA.n735 9.3005
R1047 GNDA.n737 GNDA.n20 9.3005
R1048 GNDA.n739 GNDA.n738 9.3005
R1049 GNDA.n740 GNDA.n18 9.3005
R1050 GNDA.n743 GNDA.n742 9.3005
R1051 GNDA.n744 GNDA.n17 9.3005
R1052 GNDA.n746 GNDA.n745 9.3005
R1053 GNDA.n748 GNDA.n15 9.3005
R1054 GNDA.n750 GNDA.n749 9.3005
R1055 GNDA.n751 GNDA.n14 9.3005
R1056 GNDA.n753 GNDA.n752 9.3005
R1057 GNDA.n755 GNDA.n12 9.3005
R1058 GNDA.n757 GNDA.n756 9.3005
R1059 GNDA.n758 GNDA.n11 9.3005
R1060 GNDA.n760 GNDA.n759 9.3005
R1061 GNDA.n761 GNDA.n10 9.3005
R1062 GNDA.n763 GNDA.n762 9.3005
R1063 GNDA.n764 GNDA.n9 9.3005
R1064 GNDA.n766 GNDA.n765 9.3005
R1065 GNDA.n768 GNDA.n6 9.3005
R1066 GNDA.n771 GNDA.n770 9.3005
R1067 GNDA.n772 GNDA.n5 9.3005
R1068 GNDA.n774 GNDA.n773 9.3005
R1069 GNDA.n775 GNDA.n4 9.3005
R1070 GNDA.n777 GNDA.n776 9.3005
R1071 GNDA.n778 GNDA.n3 9.3005
R1072 GNDA.n780 GNDA.n779 9.3005
R1073 GNDA.n781 GNDA.n1 9.3005
R1074 GNDA.n495 GNDA.t123 8.40814
R1075 GNDA.n366 GNDA.n261 7.49888
R1076 GNDA.n490 GNDA.n489 7.11161
R1077 GNDA.n487 GNDA.n485 7.11161
R1078 GNDA.n98 GNDA.n97 7.11161
R1079 GNDA.n102 GNDA.n91 7.11161
R1080 GNDA.t173 GNDA.t112 6.85408
R1081 GNDA.t195 GNDA.t213 6.85408
R1082 GNDA.n483 GNDA.n482 6.69883
R1083 GNDA.n475 GNDA.n474 6.4005
R1084 GNDA.n453 GNDA.n452 6.4005
R1085 GNDA.n526 GNDA.n82 6.4005
R1086 GNDA.n696 GNDA.n692 6.4005
R1087 GNDA.n735 GNDA.n734 6.4005
R1088 GNDA.n748 GNDA.n747 6.4005
R1089 GNDA.n755 GNDA.n754 6.4005
R1090 GNDA.n767 GNDA.n766 6.4005
R1091 GNDA.n782 GNDA.n781 6.4005
R1092 GNDA.n394 GNDA.n393 6.4005
R1093 GNDA.n406 GNDA.n405 6.4005
R1094 GNDA.n553 GNDA.n552 6.4005
R1095 GNDA.n576 GNDA.n53 6.4005
R1096 GNDA.n680 GNDA.n619 6.4005
R1097 GNDA.n664 GNDA.n663 6.4005
R1098 GNDA.n651 GNDA.n631 6.4005
R1099 GNDA.n635 GNDA.n633 6.4005
R1100 GNDA.n353 GNDA.n352 6.4005
R1101 GNDA.n332 GNDA.n331 6.4005
R1102 GNDA.n326 GNDA.n282 6.4005
R1103 GNDA.n287 GNDA.n285 6.4005
R1104 GNDA.n313 GNDA.n312 6.4005
R1105 GNDA.n301 GNDA.n300 6.4005
R1106 GNDA.n191 GNDA.n187 6.4005
R1107 GNDA.n510 GNDA.n104 6.4005
R1108 GNDA.n727 GNDA.n8 5.68939
R1109 GNDA.n297 GNDA.n296 5.68939
R1110 GNDA.n297 GNDA.n288 5.68939
R1111 GNDA.n727 GNDA.n7 4.97828
R1112 GNDA.n166 GNDA.n114 4.49344
R1113 GNDA.n111 GNDA.n110 4.49344
R1114 GNDA.n500 GNDA.n110 4.49344
R1115 GNDA.n167 GNDA.n166 4.49344
R1116 GNDA.n133 GNDA.n132 4.4805
R1117 GNDA.n497 GNDA.n496 3.8278
R1118 GNDA.n113 GNDA.n112 3.8278
R1119 GNDA.n124 GNDA.n123 3.8278
R1120 GNDA.n489 GNDA.n488 3.48951
R1121 GNDA.n488 GNDA.n487 3.48951
R1122 GNDA.n97 GNDA.n96 3.48951
R1123 GNDA.n96 GNDA.n91 3.48951
R1124 GNDA.n420 GNDA.n419 3.2005
R1125 GNDA.n540 GNDA.n539 3.2005
R1126 GNDA.n561 GNDA.n58 3.2005
R1127 GNDA.n600 GNDA.n45 3.2005
R1128 GNDA.n607 GNDA.n40 3.2005
R1129 GNDA.n360 GNDA.n359 3.2005
R1130 GNDA.n346 GNDA.n345 3.2005
R1131 GNDA.n125 GNDA.n121 2.8779
R1132 GNDA.n126 GNDA.n121 2.8779
R1133 GNDA.t225 GNDA.t99 2.28503
R1134 GNDA.t180 GNDA.t134 2.28503
R1135 GNDA.n77 GNDA.n76 2.25882
R1136 GNDA.n78 GNDA.n77 2.25882
R1137 GNDA.n527 GNDA.n81 2.25882
R1138 GNDA.n80 GNDA.n78 2.25882
R1139 GNDA.n529 GNDA.n76 2.25882
R1140 GNDA.n81 GNDA.n80 2.25882
R1141 GNDA.n462 GNDA.n442 2.25882
R1142 GNDA.n442 GNDA.n441 2.25882
R1143 GNDA.n467 GNDA.n435 2.25882
R1144 GNDA.n441 GNDA.n440 2.25882
R1145 GNDA.n463 GNDA.n462 2.25882
R1146 GNDA.n440 GNDA.n435 2.25882
R1147 GNDA.n508 GNDA.n105 0.9875
R1148 GNDA.n483 GNDA.n429 0.703977
R1149 GNDA.n641 GNDA.n640 0.442364
R1150 GNDA.n364 GNDA.n261 0.193977
R1151 GNDA.n302 GNDA.n0 0.193881
R1152 GNDA.n783 GNDA.n1 0.193881
R1153 GNDA.n718 GNDA.n26 0.193695
R1154 GNDA.n381 GNDA.n377 0.193477
R1155 GNDA.n212 GNDA.n211 0.188
R1156 GNDA.n134 GNDA 0.162727
R1157 GNDA.n382 GNDA.n381 0.15675
R1158 GNDA.n383 GNDA.n382 0.15675
R1159 GNDA.n383 GNDA.n375 0.15675
R1160 GNDA.n389 GNDA.n375 0.15675
R1161 GNDA.n390 GNDA.n389 0.15675
R1162 GNDA.n391 GNDA.n390 0.15675
R1163 GNDA.n391 GNDA.n372 0.15675
R1164 GNDA.n396 GNDA.n372 0.15675
R1165 GNDA.n397 GNDA.n396 0.15675
R1166 GNDA.n423 GNDA.n397 0.15675
R1167 GNDA.n423 GNDA.n422 0.15675
R1168 GNDA.n422 GNDA.n421 0.15675
R1169 GNDA.n421 GNDA.n398 0.15675
R1170 GNDA.n416 GNDA.n398 0.15675
R1171 GNDA.n416 GNDA.n415 0.15675
R1172 GNDA.n415 GNDA.n414 0.15675
R1173 GNDA.n414 GNDA.n401 0.15675
R1174 GNDA.n409 GNDA.n401 0.15675
R1175 GNDA.n409 GNDA.n408 0.15675
R1176 GNDA.n408 GNDA.n407 0.15675
R1177 GNDA.n407 GNDA.n71 0.15675
R1178 GNDA.n535 GNDA.n71 0.15675
R1179 GNDA.n536 GNDA.n535 0.15675
R1180 GNDA.n537 GNDA.n536 0.15675
R1181 GNDA.n537 GNDA.n68 0.15675
R1182 GNDA.n542 GNDA.n68 0.15675
R1183 GNDA.n543 GNDA.n542 0.15675
R1184 GNDA.n544 GNDA.n543 0.15675
R1185 GNDA.n544 GNDA.n66 0.15675
R1186 GNDA.n548 GNDA.n66 0.15675
R1187 GNDA.n549 GNDA.n548 0.15675
R1188 GNDA.n549 GNDA.n62 0.15675
R1189 GNDA.n554 GNDA.n62 0.15675
R1190 GNDA.n555 GNDA.n554 0.15675
R1191 GNDA.n556 GNDA.n555 0.15675
R1192 GNDA.n556 GNDA.n59 0.15675
R1193 GNDA.n563 GNDA.n59 0.15675
R1194 GNDA.n564 GNDA.n563 0.15675
R1195 GNDA.n565 GNDA.n564 0.15675
R1196 GNDA.n565 GNDA.n57 0.15675
R1197 GNDA.n569 GNDA.n57 0.15675
R1198 GNDA.n570 GNDA.n569 0.15675
R1199 GNDA.n571 GNDA.n570 0.15675
R1200 GNDA.n571 GNDA.n54 0.15675
R1201 GNDA.n578 GNDA.n54 0.15675
R1202 GNDA.n579 GNDA.n578 0.15675
R1203 GNDA.n580 GNDA.n579 0.15675
R1204 GNDA.n580 GNDA.n52 0.15675
R1205 GNDA.n584 GNDA.n52 0.15675
R1206 GNDA.n585 GNDA.n584 0.15675
R1207 GNDA.n586 GNDA.n585 0.15675
R1208 GNDA.n586 GNDA.n49 0.15675
R1209 GNDA.n591 GNDA.n49 0.15675
R1210 GNDA.n592 GNDA.n591 0.15675
R1211 GNDA.n593 GNDA.n592 0.15675
R1212 GNDA.n593 GNDA.n46 0.15675
R1213 GNDA.n598 GNDA.n46 0.15675
R1214 GNDA.n599 GNDA.n598 0.15675
R1215 GNDA.n599 GNDA.n43 0.15675
R1216 GNDA.n603 GNDA.n43 0.15675
R1217 GNDA.n604 GNDA.n603 0.15675
R1218 GNDA.n604 GNDA.n41 0.15675
R1219 GNDA.n609 GNDA.n41 0.15675
R1220 GNDA.n610 GNDA.n609 0.15675
R1221 GNDA.n611 GNDA.n610 0.15675
R1222 GNDA.n611 GNDA.n39 0.15675
R1223 GNDA.n615 GNDA.n39 0.15675
R1224 GNDA.n616 GNDA.n615 0.15675
R1225 GNDA.n685 GNDA.n616 0.15675
R1226 GNDA.n685 GNDA.n684 0.15675
R1227 GNDA.n684 GNDA.n683 0.15675
R1228 GNDA.n683 GNDA.n617 0.15675
R1229 GNDA.n679 GNDA.n617 0.15675
R1230 GNDA.n679 GNDA.n678 0.15675
R1231 GNDA.n678 GNDA.n620 0.15675
R1232 GNDA.n673 GNDA.n620 0.15675
R1233 GNDA.n673 GNDA.n672 0.15675
R1234 GNDA.n672 GNDA.n671 0.15675
R1235 GNDA.n671 GNDA.n623 0.15675
R1236 GNDA.n667 GNDA.n623 0.15675
R1237 GNDA.n667 GNDA.n666 0.15675
R1238 GNDA.n666 GNDA.n665 0.15675
R1239 GNDA.n665 GNDA.n625 0.15675
R1240 GNDA.n660 GNDA.n625 0.15675
R1241 GNDA.n660 GNDA.n659 0.15675
R1242 GNDA.n659 GNDA.n658 0.15675
R1243 GNDA.n658 GNDA.n628 0.15675
R1244 GNDA.n653 GNDA.n628 0.15675
R1245 GNDA.n653 GNDA.n652 0.15675
R1246 GNDA.n652 GNDA.n632 0.15675
R1247 GNDA.n648 GNDA.n632 0.15675
R1248 GNDA.n648 GNDA.n647 0.15675
R1249 GNDA.n647 GNDA.n646 0.15675
R1250 GNDA.n646 GNDA.n634 0.15675
R1251 GNDA.n642 GNDA.n634 0.15675
R1252 GNDA.n642 GNDA.n641 0.15675
R1253 GNDA.n137 GNDA.n130 0.15675
R1254 GNDA.n138 GNDA.n137 0.15675
R1255 GNDA.n139 GNDA.n138 0.15675
R1256 GNDA.n139 GNDA.n128 0.15675
R1257 GNDA.n143 GNDA.n128 0.15675
R1258 GNDA.n144 GNDA.n143 0.15675
R1259 GNDA.n145 GNDA.n144 0.15675
R1260 GNDA.n145 GNDA.n119 0.15675
R1261 GNDA.n149 GNDA.n119 0.15675
R1262 GNDA.n150 GNDA.n149 0.15675
R1263 GNDA.n151 GNDA.n150 0.15675
R1264 GNDA.n151 GNDA.n117 0.15675
R1265 GNDA.n155 GNDA.n117 0.15675
R1266 GNDA.n156 GNDA.n155 0.15675
R1267 GNDA.n164 GNDA.n156 0.15675
R1268 GNDA.n164 GNDA.n163 0.15675
R1269 GNDA.n163 GNDA.n162 0.15675
R1270 GNDA.n162 GNDA.n157 0.15675
R1271 GNDA.n158 GNDA.n157 0.15675
R1272 GNDA.n158 GNDA.n108 0.15675
R1273 GNDA.n502 GNDA.n108 0.15675
R1274 GNDA.n503 GNDA.n502 0.15675
R1275 GNDA.n504 GNDA.n503 0.15675
R1276 GNDA.n364 GNDA.n363 0.15675
R1277 GNDA.n363 GNDA.n362 0.15675
R1278 GNDA.n362 GNDA.n263 0.15675
R1279 GNDA.n357 GNDA.n263 0.15675
R1280 GNDA.n357 GNDA.n356 0.15675
R1281 GNDA.n356 GNDA.n355 0.15675
R1282 GNDA.n355 GNDA.n266 0.15675
R1283 GNDA.n350 GNDA.n266 0.15675
R1284 GNDA.n350 GNDA.n349 0.15675
R1285 GNDA.n349 GNDA.n348 0.15675
R1286 GNDA.n348 GNDA.n269 0.15675
R1287 GNDA.n343 GNDA.n269 0.15675
R1288 GNDA.n343 GNDA.n342 0.15675
R1289 GNDA.n342 GNDA.n341 0.15675
R1290 GNDA.n341 GNDA.n275 0.15675
R1291 GNDA.n336 GNDA.n275 0.15675
R1292 GNDA.n336 GNDA.n335 0.15675
R1293 GNDA.n335 GNDA.n334 0.15675
R1294 GNDA.n334 GNDA.n278 0.15675
R1295 GNDA.n329 GNDA.n278 0.15675
R1296 GNDA.n329 GNDA.n328 0.15675
R1297 GNDA.n328 GNDA.n327 0.15675
R1298 GNDA.n327 GNDA.n281 0.15675
R1299 GNDA.n323 GNDA.n281 0.15675
R1300 GNDA.n323 GNDA.n322 0.15675
R1301 GNDA.n322 GNDA.n321 0.15675
R1302 GNDA.n321 GNDA.n284 0.15675
R1303 GNDA.n317 GNDA.n284 0.15675
R1304 GNDA.n317 GNDA.n316 0.15675
R1305 GNDA.n316 GNDA.n315 0.15675
R1306 GNDA.n315 GNDA.n286 0.15675
R1307 GNDA.n310 GNDA.n286 0.15675
R1308 GNDA.n310 GNDA.n309 0.15675
R1309 GNDA.n309 GNDA.n308 0.15675
R1310 GNDA.n308 GNDA.n290 0.15675
R1311 GNDA.n304 GNDA.n290 0.15675
R1312 GNDA.n304 GNDA.n303 0.15675
R1313 GNDA.n303 GNDA.n302 0.15675
R1314 GNDA.n247 GNDA.n174 0.15675
R1315 GNDA.n243 GNDA.n242 0.15675
R1316 GNDA.n242 GNDA.n241 0.15675
R1317 GNDA.n241 GNDA.n178 0.15675
R1318 GNDA.n237 GNDA.n236 0.15675
R1319 GNDA.n236 GNDA.n235 0.15675
R1320 GNDA.n235 GNDA.n182 0.15675
R1321 GNDA.n231 GNDA.n230 0.15675
R1322 GNDA.n230 GNDA.n229 0.15675
R1323 GNDA.n229 GNDA.n186 0.15675
R1324 GNDA.n225 GNDA.n224 0.15675
R1325 GNDA.n224 GNDA.n223 0.15675
R1326 GNDA.n223 GNDA.n190 0.15675
R1327 GNDA.n219 GNDA.n218 0.15675
R1328 GNDA.n216 GNDA.n210 0.15675
R1329 GNDA.n212 GNDA.n210 0.15675
R1330 GNDA.n478 GNDA.n429 0.15675
R1331 GNDA.n478 GNDA.n477 0.15675
R1332 GNDA.n477 GNDA.n476 0.15675
R1333 GNDA.n476 GNDA.n431 0.15675
R1334 GNDA.n471 GNDA.n431 0.15675
R1335 GNDA.n471 GNDA.n470 0.15675
R1336 GNDA.n470 GNDA.n469 0.15675
R1337 GNDA.n469 GNDA.n433 0.15675
R1338 GNDA.n444 GNDA.n433 0.15675
R1339 GNDA.n445 GNDA.n444 0.15675
R1340 GNDA.n457 GNDA.n445 0.15675
R1341 GNDA.n457 GNDA.n456 0.15675
R1342 GNDA.n456 GNDA.n455 0.15675
R1343 GNDA.n455 GNDA.n447 0.15675
R1344 GNDA.n451 GNDA.n447 0.15675
R1345 GNDA.n451 GNDA.n450 0.15675
R1346 GNDA.n450 GNDA.n84 0.15675
R1347 GNDA.n525 GNDA.n84 0.15675
R1348 GNDA.n525 GNDA.n524 0.15675
R1349 GNDA.n524 GNDA.n523 0.15675
R1350 GNDA.n523 GNDA.n85 0.15675
R1351 GNDA.n519 GNDA.n85 0.15675
R1352 GNDA.n519 GNDA.n518 0.15675
R1353 GNDA.n518 GNDA.n517 0.15675
R1354 GNDA.n517 GNDA.n89 0.15675
R1355 GNDA.n513 GNDA.n89 0.15675
R1356 GNDA.n513 GNDA.n512 0.15675
R1357 GNDA.n512 GNDA.n511 0.15675
R1358 GNDA.n718 GNDA.n717 0.15675
R1359 GNDA.n717 GNDA.n716 0.15675
R1360 GNDA.n716 GNDA.n28 0.15675
R1361 GNDA.n712 GNDA.n28 0.15675
R1362 GNDA.n712 GNDA.n711 0.15675
R1363 GNDA.n711 GNDA.n710 0.15675
R1364 GNDA.n710 GNDA.n30 0.15675
R1365 GNDA.n706 GNDA.n30 0.15675
R1366 GNDA.n706 GNDA.n705 0.15675
R1367 GNDA.n703 GNDA.n33 0.15675
R1368 GNDA.n699 GNDA.n33 0.15675
R1369 GNDA.n699 GNDA.n698 0.15675
R1370 GNDA.n698 GNDA.n697 0.15675
R1371 GNDA.n697 GNDA.n35 0.15675
R1372 GNDA.n693 GNDA.n35 0.15675
R1373 GNDA.n693 GNDA.n21 0.15675
R1374 GNDA.n736 GNDA.n21 0.15675
R1375 GNDA.n737 GNDA.n736 0.15675
R1376 GNDA.n738 GNDA.n737 0.15675
R1377 GNDA.n738 GNDA.n18 0.15675
R1378 GNDA.n743 GNDA.n18 0.15675
R1379 GNDA.n744 GNDA.n743 0.15675
R1380 GNDA.n745 GNDA.n744 0.15675
R1381 GNDA.n745 GNDA.n15 0.15675
R1382 GNDA.n750 GNDA.n15 0.15675
R1383 GNDA.n751 GNDA.n750 0.15675
R1384 GNDA.n752 GNDA.n751 0.15675
R1385 GNDA.n752 GNDA.n12 0.15675
R1386 GNDA.n757 GNDA.n12 0.15675
R1387 GNDA.n758 GNDA.n757 0.15675
R1388 GNDA.n759 GNDA.n758 0.15675
R1389 GNDA.n759 GNDA.n10 0.15675
R1390 GNDA.n763 GNDA.n10 0.15675
R1391 GNDA.n764 GNDA.n763 0.15675
R1392 GNDA.n765 GNDA.n764 0.15675
R1393 GNDA.n765 GNDA.n6 0.15675
R1394 GNDA.n771 GNDA.n6 0.15675
R1395 GNDA.n772 GNDA.n771 0.15675
R1396 GNDA.n773 GNDA.n772 0.15675
R1397 GNDA.n773 GNDA.n4 0.15675
R1398 GNDA.n777 GNDA.n4 0.15675
R1399 GNDA.n778 GNDA.n777 0.15675
R1400 GNDA.n779 GNDA.n778 0.15675
R1401 GNDA.n779 GNDA.n1 0.15675
R1402 GNDA.n504 GNDA.n106 0.141125
R1403 GNDA.n508 GNDA.n507 0.1321
R1404 GNDA.n248 GNDA.n171 0.131895
R1405 GNDA.n511 GNDA 0.1255
R1406 GNDA.n705 GNDA.n704 0.109875
R1407 GNDA.n177 GNDA.n174 0.09425
R1408 GNDA.n181 GNDA.n178 0.09425
R1409 GNDA.n185 GNDA.n182 0.09425
R1410 GNDA.n189 GNDA.n186 0.09425
R1411 GNDA.n194 GNDA.n190 0.09425
R1412 GNDA.n218 GNDA.n217 0.09425
R1413 GNDA.n248 GNDA.n247 0.063
R1414 GNDA.n243 GNDA.n177 0.063
R1415 GNDA.n237 GNDA.n181 0.063
R1416 GNDA.n231 GNDA.n185 0.063
R1417 GNDA.n225 GNDA.n189 0.063
R1418 GNDA.n219 GNDA.n194 0.063
R1419 GNDA.n217 GNDA.n216 0.063
R1420 GNDA.n509 GNDA 0.063
R1421 GNDA.n704 GNDA.n703 0.047375
R1422 GNDA.n506 GNDA.n106 0.0430057
R1423 GNDA GNDA.n130 0.03175
R1424 V_CONT.n10 V_CONT.t11 1156.8
R1425 V_CONT.n11 V_CONT.n10 964
R1426 VCO_FD_magic_0.V_CONT V_CONT.n12 562.333
R1427 V_CONT.n12 V_CONT.n11 433.8
R1428 V_CONT.n1 V_CONT.t8 377.567
R1429 V_CONT.n0 V_CONT.t12 297.233
R1430 V_CONT.n5 V_CONT.n4 242.903
R1431 V_CONT.n2 V_CONT.n0 237.851
R1432 V_CONT.n2 V_CONT.n1 232.809
R1433 V_CONT.n1 V_CONT.t9 216.9
R1434 V_CONT.n12 V_CONT.t10 192.8
R1435 V_CONT.n11 V_CONT.t14 192.8
R1436 V_CONT.n10 V_CONT.t15 192.8
R1437 V_CONT.n5 V_CONT.n3 172.502
R1438 V_CONT.n13 VCO_FD_magic_0.V_CONT 168.037
R1439 V_CONT.n8 V_CONT.t3 164.457
R1440 V_CONT.n0 V_CONT.t13 136.567
R1441 V_CONT.n15 V_CONT.n7 118.35
R1442 V_CONT.n7 V_CONT.n6 106.662
R1443 opamp_cell_4_0.VIN- V_CONT.n15 50.938
R1444 V_CONT.n3 V_CONT.t2 24.6255
R1445 V_CONT.n3 V_CONT.t4 24.6255
R1446 V_CONT.n4 V_CONT.t0 24.6255
R1447 V_CONT.n4 V_CONT.t5 24.6255
R1448 V_CONT.n7 V_CONT.n5 22.4005
R1449 V_CONT.n6 V_CONT.t1 15.0005
R1450 V_CONT.n6 V_CONT.t7 15.0005
R1451 V_CONT.n15 V_CONT.n14 9.45883
R1452 V_CONT.n14 V_CONT.n13 4.5005
R1453 V_CONT.n9 V_CONT.n8 4.5005
R1454 V_CONT.n9 V_CONT.t6 3.76103
R1455 opamp_cell_4_0.VIN- V_CONT.n2 1.39633
R1456 V_CONT.n13 V_CONT.n9 0.172375
R1457 V_CONT.n14 V_CONT.n8 0.172375
R1458 a_5970_4630.n8 a_5970_4630.n6 522.322
R1459 a_5970_4630.n3 a_5970_4630.t7 384.967
R1460 a_5970_4630.n0 a_5970_4630.t10 384.967
R1461 a_5970_4630.n3 a_5970_4630.t9 379.166
R1462 a_5970_4630.t11 a_5970_4630.n0 376.56
R1463 a_5970_4630.n5 a_5970_4630.n1 315.647
R1464 a_5970_4630.n4 a_5970_4630.n2 315.647
R1465 a_5970_4630.n11 a_5970_4630.n10 314.502
R1466 a_5970_4630.n8 a_5970_4630.n7 160.721
R1467 a_5970_4630.n5 a_5970_4630.n4 83.2005
R1468 a_5970_4630.n1 a_5970_4630.t12 49.2505
R1469 a_5970_4630.n1 a_5970_4630.t6 49.2505
R1470 a_5970_4630.n2 a_5970_4630.t5 49.2505
R1471 a_5970_4630.n2 a_5970_4630.t8 49.2505
R1472 a_5970_4630.t11 a_5970_4630.n11 49.2505
R1473 a_5970_4630.n11 a_5970_4630.t0 49.2505
R1474 a_5970_4630.n10 a_5970_4630.n9 42.6672
R1475 a_5970_4630.n9 a_5970_4630.n8 37.763
R1476 a_5970_4630.n9 a_5970_4630.n5 23.4672
R1477 a_5970_4630.n6 a_5970_4630.t1 19.7005
R1478 a_5970_4630.n6 a_5970_4630.t4 19.7005
R1479 a_5970_4630.n7 a_5970_4630.t2 19.7005
R1480 a_5970_4630.n7 a_5970_4630.t3 19.7005
R1481 a_5970_4630.n4 a_5970_4630.n3 16.0005
R1482 a_5970_4630.n10 a_5970_4630.n0 16.0005
R1483 VDDA.t99 VDDA.t69 2804.76
R1484 VDDA.t0 VDDA.t210 2533.33
R1485 VDDA.t208 VDDA.t40 2307.14
R1486 VDDA.t56 VDDA.t193 2216.67
R1487 VDDA.t86 VDDA.t186 2216.67
R1488 VDDA.t22 VDDA.t216 2216.67
R1489 VDDA.t200 VDDA.t214 2126.19
R1490 VDDA.t36 VDDA.t188 1538.1
R1491 VDDA.t15 VDDA.t26 1492.86
R1492 VDDA.t195 VDDA.t66 1492.86
R1493 VDDA.t119 VDDA.t7 1317.78
R1494 VDDA.t120 VDDA.n91 1289.29
R1495 VDDA.t59 VDDA.n90 1289.29
R1496 VDDA.t106 VDDA.t204 1130.95
R1497 VDDA.t212 VDDA.t54 1130.95
R1498 VDDA.t84 VDDA.t93 1130.95
R1499 VDDA.t132 VDDA.t122 1130.95
R1500 VDDA.t91 VDDA.t34 1130.95
R1501 VDDA.t97 VDDA.n97 927.381
R1502 VDDA.t5 VDDA.n95 927.381
R1503 VDDA.t202 VDDA.n94 927.381
R1504 VDDA.t128 VDDA.n92 927.381
R1505 VDDA.n86 VDDA.n75 831.25
R1506 VDDA.n80 VDDA.n78 831.25
R1507 VDDA.n768 VDDA.n760 831.25
R1508 VDDA.n763 VDDA.n762 831.25
R1509 VDDA.n757 VDDA.n749 831.25
R1510 VDDA.n752 VDDA.n751 831.25
R1511 VDDA.n236 VDDA.t215 726.734
R1512 VDDA.n238 VDDA.t92 726.734
R1513 VDDA.n96 VDDA.t57 663.801
R1514 VDDA.n53 VDDA.t87 663.801
R1515 VDDA.n93 VDDA.t23 663.801
R1516 VDDA.n35 VDDA.t209 663.801
R1517 VDDA.n17 VDDA.t100 663.801
R1518 VDDA.n89 VDDA.t74 663.801
R1519 VDDA.n67 VDDA.n66 647.933
R1520 VDDA.n134 VDDA.n133 647.933
R1521 VDDA.n152 VDDA.n59 647.933
R1522 VDDA.n158 VDDA.n56 647.933
R1523 VDDA.n49 VDDA.n48 647.933
R1524 VDDA.n179 VDDA.n178 647.933
R1525 VDDA.n197 VDDA.n41 647.933
R1526 VDDA.n203 VDDA.n38 647.933
R1527 VDDA.n219 VDDA.n218 647.933
R1528 VDDA.n29 VDDA.n28 647.933
R1529 VDDA.n245 VDDA.n23 647.933
R1530 VDDA.n252 VDDA.n20 647.933
R1531 VDDA.n8 VDDA.n7 647.933
R1532 VDDA.n291 VDDA.n290 647.933
R1533 VDDA.n271 VDDA.n12 646.715
R1534 VDDA.n97 VDDA.t56 610.715
R1535 VDDA.n95 VDDA.t86 610.715
R1536 VDDA.n94 VDDA.t22 610.715
R1537 VDDA.n92 VDDA.t208 610.715
R1538 VDDA.n91 VDDA.t99 610.715
R1539 VDDA.n90 VDDA.t73 610.715
R1540 VDDA.n83 VDDA.n75 585
R1541 VDDA.n82 VDDA.n78 585
R1542 VDDA.n761 VDDA.n760 585
R1543 VDDA.n765 VDDA.n763 585
R1544 VDDA.n661 VDDA.n655 585
R1545 VDDA.n656 VDDA.n655 585
R1546 VDDA.n667 VDDA.n344 585
R1547 VDDA.n671 VDDA.n344 585
R1548 VDDA.n612 VDDA.n350 585
R1549 VDDA.n607 VDDA.n350 585
R1550 VDDA.n588 VDDA.n583 585
R1551 VDDA.n592 VDDA.n583 585
R1552 VDDA.n750 VDDA.n749 585
R1553 VDDA.n754 VDDA.n752 585
R1554 VDDA.n652 VDDA.n646 585
R1555 VDDA.n647 VDDA.n646 585
R1556 VDDA.n358 VDDA.n351 585
R1557 VDDA.n353 VDDA.n351 585
R1558 VDDA.n423 VDDA.n416 585
R1559 VDDA.n405 VDDA.n397 585
R1560 VDDA.n571 VDDA.n475 585
R1561 VDDA.n564 VDDA.n475 585
R1562 VDDA.n561 VDDA.n560 585
R1563 VDDA.n560 VDDA.n559 585
R1564 VDDA.n530 VDDA.n529 585
R1565 VDDA.n530 VDDA.n519 585
R1566 VDDA.n99 VDDA.t224 537.492
R1567 VDDA.n110 VDDA.t223 537.491
R1568 VDDA.n87 VDDA.t222 537.491
R1569 VDDA.t7 VDDA.t106 497.62
R1570 VDDA.t204 VDDA.t97 497.62
R1571 VDDA.t193 VDDA.t212 497.62
R1572 VDDA.t54 VDDA.t5 497.62
R1573 VDDA.t186 VDDA.t84 497.62
R1574 VDDA.t93 VDDA.t202 497.62
R1575 VDDA.t216 VDDA.t132 497.62
R1576 VDDA.t122 VDDA.t128 497.62
R1577 VDDA.t40 VDDA.t15 497.62
R1578 VDDA.t26 VDDA.t200 497.62
R1579 VDDA.t214 VDDA.t91 497.62
R1580 VDDA.t34 VDDA.t36 497.62
R1581 VDDA.t188 VDDA.t120 497.62
R1582 VDDA.t69 VDDA.t20 497.62
R1583 VDDA.t20 VDDA.t195 497.62
R1584 VDDA.t66 VDDA.t0 497.62
R1585 VDDA.t210 VDDA.t59 497.62
R1586 VDDA.t30 VDDA.n76 465.079
R1587 VDDA.n81 VDDA.t30 465.079
R1588 VDDA.n767 VDDA.t51 465.079
R1589 VDDA.t51 VDDA.n766 465.079
R1590 VDDA.n756 VDDA.t10 465.079
R1591 VDDA.t10 VDDA.n755 465.079
R1592 VDDA.n105 VDDA.t44 464.281
R1593 VDDA.n102 VDDA.t44 464.281
R1594 VDDA.n113 VDDA.t48 464.281
R1595 VDDA.t48 VDDA.n72 464.281
R1596 VDDA.t116 VDDA.n636 464.281
R1597 VDDA.n638 VDDA.t116 464.281
R1598 VDDA.n744 VDDA.t218 464.281
R1599 VDDA.t218 VDDA.n743 464.281
R1600 VDDA.n781 VDDA.t63 464.281
R1601 VDDA.t63 VDDA.n780 464.281
R1602 VDDA.n725 VDDA.t18 464.281
R1603 VDDA.t18 VDDA.n724 464.281
R1604 VDDA.n703 VDDA.t207 464.281
R1605 VDDA.t207 VDDA.n702 464.281
R1606 VDDA.n633 VDDA.t197 464.281
R1607 VDDA.t197 VDDA.n632 464.281
R1608 VDDA.t83 VDDA.n733 464.281
R1609 VDDA.n734 VDDA.t83 464.281
R1610 VDDA.t62 VDDA.n317 464.281
R1611 VDDA.n771 VDDA.t62 464.281
R1612 VDDA.t25 VDDA.n325 464.281
R1613 VDDA.n706 VDDA.t25 464.281
R1614 VDDA.t220 VDDA.n621 464.281
R1615 VDDA.n622 VDDA.t220 464.281
R1616 VDDA.n341 VDDA.t221 415.336
R1617 VDDA.n386 VDDA.t167 384.967
R1618 VDDA.n428 VDDA.t173 384.967
R1619 VDDA.n391 VDDA.t152 384.967
R1620 VDDA.n411 VDDA.t149 384.967
R1621 VDDA.n95 VDDA.n53 382.8
R1622 VDDA.n94 VDDA.n93 382.8
R1623 VDDA.n92 VDDA.n35 382.8
R1624 VDDA.n91 VDDA.n17 382.8
R1625 VDDA.n90 VDDA.n89 382.8
R1626 VDDA.n97 VDDA.n96 382.8
R1627 VDDA.n423 VDDA.t160 374.878
R1628 VDDA.t171 VDDA.t64 360.346
R1629 VDDA.t64 VDDA.t130 360.346
R1630 VDDA.t130 VDDA.t13 360.346
R1631 VDDA.t13 VDDA.t134 360.346
R1632 VDDA.t134 VDDA.t164 360.346
R1633 VDDA.t88 VDDA.t178 360.346
R1634 VDDA.t52 VDDA.t88 360.346
R1635 VDDA.t136 VDDA.t52 360.346
R1636 VDDA.t71 VDDA.t136 360.346
R1637 VDDA.t181 VDDA.t71 360.346
R1638 VDDA.n110 VDDA.t144 359.752
R1639 VDDA.n87 VDDA.t143 359.752
R1640 VDDA.n99 VDDA.t142 359.752
R1641 VDDA.n396 VDDA.t156 352.834
R1642 VDDA.n525 VDDA.t171 343.966
R1643 VDDA.n563 VDDA.t164 343.966
R1644 VDDA.t178 VDDA.n563 343.966
R1645 VDDA.n569 VDDA.t181 343.966
R1646 VDDA.n412 VDDA.t151 341.752
R1647 VDDA.n427 VDDA.t176 341.752
R1648 VDDA.n387 VDDA.t169 341.752
R1649 VDDA.n392 VDDA.t155 341.752
R1650 VDDA.n558 VDDA.t177 336.329
R1651 VDDA.n558 VDDA.t163 336.329
R1652 VDDA.n520 VDDA.t170 320.7
R1653 VDDA.n572 VDDA.t180 320.7
R1654 VDDA.n385 VDDA.n383 315.647
R1655 VDDA.n379 VDDA.n378 315.647
R1656 VDDA.n410 VDDA.n409 315.647
R1657 VDDA.n390 VDDA.n389 315.647
R1658 VDDA.n430 VDDA.n382 315.647
R1659 VDDA.n429 VDDA.n384 315.647
R1660 VDDA.n324 VDDA.t199 315.25
R1661 VDDA.t58 VDDA.t33 314.113
R1662 VDDA.t114 VDDA.t28 314.113
R1663 VDDA.t168 VDDA.n387 304.659
R1664 VDDA.n560 VDDA.n483 291.363
R1665 VDDA.n556 VDDA.n481 291.363
R1666 VDDA.n557 VDDA.n556 291.363
R1667 VDDA.n659 VDDA.n655 290.733
R1668 VDDA.n665 VDDA.n344 290.733
R1669 VDDA.n610 VDDA.n350 290.733
R1670 VDDA.n586 VDDA.n583 290.733
R1671 VDDA.n650 VDDA.n646 290.733
R1672 VDDA.n352 VDDA.n351 290.733
R1673 VDDA.n421 VDDA.n416 290.733
R1674 VDDA.n417 VDDA.n416 290.733
R1675 VDDA.n403 VDDA.n397 290.733
R1676 VDDA.n398 VDDA.n397 290.733
R1677 VDDA.n565 VDDA.n475 290.733
R1678 VDDA.n530 VDDA.n518 290.733
R1679 VDDA.n745 VDDA.n744 243.698
R1680 VDDA.n782 VDDA.n781 243.698
R1681 VDDA.n726 VDDA.n725 243.698
R1682 VDDA.n704 VDDA.n703 243.698
R1683 VDDA.n634 VDDA.n633 243.698
R1684 VDDA.n734 VDDA.n731 243.698
R1685 VDDA.n775 VDDA.n771 243.698
R1686 VDDA.n710 VDDA.n706 243.698
R1687 VDDA.n622 VDDA.n619 243.698
R1688 VDDA.n107 VDDA.n106 238.367
R1689 VDDA.n101 VDDA.n88 238.367
R1690 VDDA.n115 VDDA.n114 238.367
R1691 VDDA.n118 VDDA.n117 238.367
R1692 VDDA.n86 VDDA.n85 238.367
R1693 VDDA.n80 VDDA.n79 238.367
R1694 VDDA.n730 VDDA.n301 238.367
R1695 VDDA.n769 VDDA.n768 238.367
R1696 VDDA.n762 VDDA.n729 238.367
R1697 VDDA.n728 VDDA.n316 238.367
R1698 VDDA.n721 VDDA.n319 238.367
R1699 VDDA.n699 VDDA.n327 238.367
R1700 VDDA.n618 VDDA.n335 238.367
R1701 VDDA.n738 VDDA.n302 238.367
R1702 VDDA.n758 VDDA.n757 238.367
R1703 VDDA.n785 VDDA.n784 238.367
R1704 VDDA.n713 VDDA.n712 238.367
R1705 VDDA.n626 VDDA.n331 238.367
R1706 VDDA.n751 VDDA.n747 238.367
R1707 VDDA.n417 VDDA.n388 233.841
R1708 VDDA.n398 VDDA.n394 233.841
R1709 VDDA.n662 VDDA.n661 230.308
R1710 VDDA.n656 VDDA.n615 230.308
R1711 VDDA.n668 VDDA.n667 230.308
R1712 VDDA.n671 VDDA.n670 230.308
R1713 VDDA.n613 VDDA.n612 230.308
R1714 VDDA.n607 VDDA.n346 230.308
R1715 VDDA.n589 VDDA.n588 230.308
R1716 VDDA.n592 VDDA.n591 230.308
R1717 VDDA.n653 VDDA.n652 230.308
R1718 VDDA.n358 VDDA.n348 230.308
R1719 VDDA.n353 VDDA.n347 230.308
R1720 VDDA.n647 VDDA.n644 230.308
R1721 VDDA.n424 VDDA.n423 230.308
R1722 VDDA.n571 VDDA.n570 230.308
R1723 VDDA.n568 VDDA.n564 230.308
R1724 VDDA.n562 VDDA.n561 230.308
R1725 VDDA.n559 VDDA.n478 230.308
R1726 VDDA.t68 VDDA.t11 222.178
R1727 VDDA.n74 VDDA.t29 219.232
R1728 VDDA.t184 VDDA.n74 219.232
R1729 VDDA.n116 VDDA.t47 219.232
R1730 VDDA.n108 VDDA.t43 219.232
R1731 VDDA.n663 VDDA.n643 199.195
R1732 VDDA.n492 VDDA.n491 196.502
R1733 VDDA.n489 VDDA.n488 196.502
R1734 VDDA.n555 VDDA.n554 196.502
R1735 VDDA.n546 VDDA.n511 196.502
R1736 VDDA.n539 VDDA.n514 196.502
R1737 VDDA.n532 VDDA.n531 196.502
R1738 VDDA.n638 VDDA.n617 190.333
R1739 VDDA.n110 VDDA.t47 185.002
R1740 VDDA.t184 VDDA.n87 185.002
R1741 VDDA.n99 VDDA.t43 185.002
R1742 VDDA.n427 VDDA.n426 185.001
R1743 VDDA.n413 VDDA.n412 185.001
R1744 VDDA.n408 VDDA.n392 185.001
R1745 VDDA.n84 VDDA.n83 185
R1746 VDDA.n82 VDDA.n77 185
R1747 VDDA.n112 VDDA.n109 185
R1748 VDDA.n111 VDDA.n73 185
R1749 VDDA.n104 VDDA.n98 185
R1750 VDDA.n103 VDDA.n100 185
R1751 VDDA.n357 VDDA.n356 185
R1752 VDDA.n355 VDDA.n354 185
R1753 VDDA.n651 VDDA.n645 185
R1754 VDDA.n649 VDDA.n648 185
R1755 VDDA.n625 VDDA.n624 185
R1756 VDDA.n623 VDDA.n620 185
R1757 VDDA.n707 VDDA.n326 185
R1758 VDDA.n709 VDDA.n708 185
R1759 VDDA.n772 VDDA.n318 185
R1760 VDDA.n774 VDDA.n773 185
R1761 VDDA.n750 VDDA.n748 185
R1762 VDDA.n754 VDDA.n753 185
R1763 VDDA.n737 VDDA.n736 185
R1764 VDDA.n735 VDDA.n732 185
R1765 VDDA.n587 VDDA.n585 185
R1766 VDDA.n584 VDDA.n582 185
R1767 VDDA.n611 VDDA.n349 185
R1768 VDDA.n609 VDDA.n608 185
R1769 VDDA.n666 VDDA.n664 185
R1770 VDDA.n345 VDDA.n343 185
R1771 VDDA.n660 VDDA.n654 185
R1772 VDDA.n658 VDDA.n657 185
R1773 VDDA.n629 VDDA.n628 185
R1774 VDDA.n631 VDDA.n630 185
R1775 VDDA.n329 VDDA.n328 185
R1776 VDDA.n701 VDDA.n700 185
R1777 VDDA.n321 VDDA.n320 185
R1778 VDDA.n723 VDDA.n722 185
R1779 VDDA.n777 VDDA.n776 185
R1780 VDDA.n779 VDDA.n778 185
R1781 VDDA.n761 VDDA.n759 185
R1782 VDDA.n765 VDDA.n764 185
R1783 VDDA.n740 VDDA.n739 185
R1784 VDDA.n742 VDDA.n741 185
R1785 VDDA.n642 VDDA.n334 185
R1786 VDDA.n643 VDDA.n642 185
R1787 VDDA.n641 VDDA.n640 185
R1788 VDDA.n639 VDDA.n637 185
R1789 VDDA.n643 VDDA.n617 185
R1790 VDDA.n422 VDDA.n415 185
R1791 VDDA.n420 VDDA.n414 185
R1792 VDDA.n425 VDDA.n414 185
R1793 VDDA.n419 VDDA.n418 185
R1794 VDDA.n406 VDDA.n405 185
R1795 VDDA.n407 VDDA.n406 185
R1796 VDDA.n404 VDDA.n395 185
R1797 VDDA.n402 VDDA.n401 185
R1798 VDDA.n400 VDDA.n399 185
R1799 VDDA.n482 VDDA.n479 185
R1800 VDDA.n485 VDDA.n484 185
R1801 VDDA.n477 VDDA.n476 185
R1802 VDDA.n567 VDDA.n566 185
R1803 VDDA.n529 VDDA.n521 185
R1804 VDDA.n525 VDDA.n521 185
R1805 VDDA.n528 VDDA.n527 185
R1806 VDDA.n523 VDDA.n522 185
R1807 VDDA.n524 VDDA.n519 185
R1808 VDDA.n525 VDDA.n524 185
R1809 VDDA.n590 VDDA.t68 172.38
R1810 VDDA.t126 VDDA.n614 172.38
R1811 VDDA.n669 VDDA.t77 172.38
R1812 VDDA.n559 VDDA.n558 166.63
R1813 VDDA.n116 VDDA.t2 158.333
R1814 VDDA.t42 VDDA.n108 158.333
R1815 VDDA.n100 VDDA.n98 150
R1816 VDDA.n109 VDDA.n73 150
R1817 VDDA.n84 VDDA.n77 150
R1818 VDDA.n741 VDDA.n739 150
R1819 VDDA.n764 VDDA.n759 150
R1820 VDDA.n778 VDDA.n776 150
R1821 VDDA.n722 VDDA.n320 150
R1822 VDDA.n700 VDDA.n328 150
R1823 VDDA.n630 VDDA.n628 150
R1824 VDDA.n737 VDDA.n732 150
R1825 VDDA.n753 VDDA.n748 150
R1826 VDDA.n774 VDDA.n318 150
R1827 VDDA.n709 VDDA.n326 150
R1828 VDDA.n625 VDDA.n620 150
R1829 VDDA.n642 VDDA.n641 150
R1830 VDDA.n637 VDDA.n617 150
R1831 VDDA.t80 VDDA.t3 145.038
R1832 VDDA.n635 VDDA.n627 137.904
R1833 VDDA.n711 VDDA.n705 137.904
R1834 VDDA.n590 VDDA.t95 126.412
R1835 VDDA.n614 VDDA.t11 126.412
R1836 VDDA.n669 VDDA.t126 126.412
R1837 VDDA.t77 VDDA.n663 126.412
R1838 VDDA.t185 VDDA.n75 123.126
R1839 VDDA.n78 VDDA.t185 123.126
R1840 VDDA.t50 VDDA.n760 123.126
R1841 VDDA.n763 VDDA.t50 123.126
R1842 VDDA.t79 VDDA.n749 123.126
R1843 VDDA.n752 VDDA.t79 123.126
R1844 VDDA.n657 VDDA.n654 120.001
R1845 VDDA.n664 VDDA.n345 120.001
R1846 VDDA.n608 VDDA.n349 120.001
R1847 VDDA.n585 VDDA.n584 120.001
R1848 VDDA.n648 VDDA.n645 120.001
R1849 VDDA.n356 VDDA.n355 120.001
R1850 VDDA.n415 VDDA.n414 120.001
R1851 VDDA.n418 VDDA.n414 120.001
R1852 VDDA.n406 VDDA.n395 120.001
R1853 VDDA.n401 VDDA.n400 120.001
R1854 VDDA.n567 VDDA.n477 120.001
R1855 VDDA.n484 VDDA.n479 120.001
R1856 VDDA.n527 VDDA.n521 120.001
R1857 VDDA.n524 VDDA.n523 120.001
R1858 VDDA.n461 VDDA.n367 119.737
R1859 VDDA.n454 VDDA.n370 119.737
R1860 VDDA.n447 VDDA.n373 119.737
R1861 VDDA.n440 VDDA.n376 119.737
R1862 VDDA.n432 VDDA.n381 119.737
R1863 VDDA.n426 VDDA.t174 119.656
R1864 VDDA.t2 VDDA.t184 109.615
R1865 VDDA.t47 VDDA.t42 109.615
R1866 VDDA.t43 VDDA.t119 109.615
R1867 VDDA.n425 VDDA.n413 108.779
R1868 VDDA.n783 VDDA.n727 107.258
R1869 VDDA.n783 VDDA.t61 103.427
R1870 VDDA.t9 VDDA.n770 103.427
R1871 VDDA.n770 VDDA.t49 103.427
R1872 VDDA.t82 VDDA.n746 103.427
R1873 VDDA.n727 VDDA.t24 95.7666
R1874 VDDA.t101 VDDA.t168 94.2753
R1875 VDDA.t117 VDDA.t101 94.2753
R1876 VDDA.t138 VDDA.t117 94.2753
R1877 VDDA.t31 VDDA.t138 94.2753
R1878 VDDA.t174 VDDA.t31 94.2753
R1879 VDDA.t108 VDDA.t45 94.2753
R1880 VDDA.t110 VDDA.t153 94.2753
R1881 VDDA.t190 VDDA.n408 94.2753
R1882 VDDA.t148 VDDA.t90 94.2753
R1883 VDDA.t146 VDDA.t145 94.2753
R1884 VDDA.t196 VDDA.t115 91.936
R1885 VDDA.t206 VDDA.t219 91.936
R1886 VDDA.n87 VDDA.n86 90.5056
R1887 VDDA.t198 VDDA.t17 84.2747
R1888 VDDA.t61 VDDA.t58 84.2747
R1889 VDDA.t33 VDDA.t9 84.2747
R1890 VDDA.t49 VDDA.t114 84.2747
R1891 VDDA.t28 VDDA.t82 84.2747
R1892 VDDA.t161 VDDA.t150 83.3974
R1893 VDDA.t112 VDDA.t192 83.3974
R1894 VDDA.n410 VDDA.n379 83.2005
R1895 VDDA.n390 VDDA.n379 83.2005
R1896 VDDA.n430 VDDA.n383 83.2005
R1897 VDDA.n430 VDDA.n429 83.2005
R1898 VDDA.n66 VDDA.t8 78.8005
R1899 VDDA.n66 VDDA.t107 78.8005
R1900 VDDA.n133 VDDA.t205 78.8005
R1901 VDDA.n133 VDDA.t98 78.8005
R1902 VDDA.n59 VDDA.t194 78.8005
R1903 VDDA.n59 VDDA.t213 78.8005
R1904 VDDA.n56 VDDA.t55 78.8005
R1905 VDDA.n56 VDDA.t6 78.8005
R1906 VDDA.n48 VDDA.t187 78.8005
R1907 VDDA.n48 VDDA.t85 78.8005
R1908 VDDA.n178 VDDA.t94 78.8005
R1909 VDDA.n178 VDDA.t203 78.8005
R1910 VDDA.n41 VDDA.t217 78.8005
R1911 VDDA.n41 VDDA.t133 78.8005
R1912 VDDA.n38 VDDA.t123 78.8005
R1913 VDDA.n38 VDDA.t129 78.8005
R1914 VDDA.n218 VDDA.t41 78.8005
R1915 VDDA.n218 VDDA.t16 78.8005
R1916 VDDA.n28 VDDA.t27 78.8005
R1917 VDDA.n28 VDDA.t201 78.8005
R1918 VDDA.n23 VDDA.t35 78.8005
R1919 VDDA.n23 VDDA.t37 78.8005
R1920 VDDA.n20 VDDA.t189 78.8005
R1921 VDDA.n20 VDDA.t121 78.8005
R1922 VDDA.n12 VDDA.t70 78.8005
R1923 VDDA.n12 VDDA.t21 78.8005
R1924 VDDA.n7 VDDA.t67 78.8005
R1925 VDDA.n7 VDDA.t1 78.8005
R1926 VDDA.n290 VDDA.t211 78.8005
R1927 VDDA.n290 VDDA.t60 78.8005
R1928 VDDA.t140 VDDA.t75 76.1455
R1929 VDDA.t157 VDDA.t147 76.1455
R1930 VDDA.n114 VDDA.n110 74.7688
R1931 VDDA.n106 VDDA.n99 74.7688
R1932 VDDA.n614 VDDA.n348 69.8479
R1933 VDDA.n614 VDDA.n347 69.8479
R1934 VDDA.n663 VDDA.n653 69.8479
R1935 VDDA.n663 VDDA.n644 69.8479
R1936 VDDA.n590 VDDA.n589 69.8479
R1937 VDDA.n591 VDDA.n590 69.8479
R1938 VDDA.n614 VDDA.n613 69.8479
R1939 VDDA.n614 VDDA.n346 69.8479
R1940 VDDA.n669 VDDA.n668 69.8479
R1941 VDDA.n670 VDDA.n669 69.8479
R1942 VDDA.n663 VDDA.n662 69.8479
R1943 VDDA.n663 VDDA.n615 69.8479
R1944 VDDA.n425 VDDA.n424 69.8479
R1945 VDDA.n425 VDDA.n388 69.8479
R1946 VDDA.n407 VDDA.n393 69.8479
R1947 VDDA.n407 VDDA.n394 69.8479
R1948 VDDA.n563 VDDA.n562 69.8479
R1949 VDDA.n563 VDDA.n478 69.8479
R1950 VDDA.n570 VDDA.n569 69.8479
R1951 VDDA.n569 VDDA.n568 69.8479
R1952 VDDA.n526 VDDA.n525 69.8479
R1953 VDDA.n431 VDDA.n430 69.3203
R1954 VDDA.t75 VDDA.t38 68.8936
R1955 VDDA.t147 VDDA.n407 68.8936
R1956 VDDA.n85 VDDA.n74 65.8183
R1957 VDDA.n79 VDDA.n74 65.8183
R1958 VDDA.n116 VDDA.n115 65.8183
R1959 VDDA.n117 VDDA.n116 65.8183
R1960 VDDA.n108 VDDA.n107 65.8183
R1961 VDDA.n108 VDDA.n88 65.8183
R1962 VDDA.n627 VDDA.n626 65.8183
R1963 VDDA.n627 VDDA.n619 65.8183
R1964 VDDA.n712 VDDA.n711 65.8183
R1965 VDDA.n711 VDDA.n710 65.8183
R1966 VDDA.n784 VDDA.n783 65.8183
R1967 VDDA.n783 VDDA.n775 65.8183
R1968 VDDA.n770 VDDA.n758 65.8183
R1969 VDDA.n770 VDDA.n747 65.8183
R1970 VDDA.n746 VDDA.n738 65.8183
R1971 VDDA.n746 VDDA.n731 65.8183
R1972 VDDA.n635 VDDA.n634 65.8183
R1973 VDDA.n635 VDDA.n618 65.8183
R1974 VDDA.n705 VDDA.n704 65.8183
R1975 VDDA.n705 VDDA.n327 65.8183
R1976 VDDA.n727 VDDA.n726 65.8183
R1977 VDDA.n727 VDDA.n319 65.8183
R1978 VDDA.n783 VDDA.n782 65.8183
R1979 VDDA.n783 VDDA.n728 65.8183
R1980 VDDA.n770 VDDA.n769 65.8183
R1981 VDDA.n770 VDDA.n729 65.8183
R1982 VDDA.n746 VDDA.n745 65.8183
R1983 VDDA.n746 VDDA.n730 65.8183
R1984 VDDA.n643 VDDA.n616 65.8183
R1985 VDDA.t150 VDDA.t103 61.6417
R1986 VDDA.t192 VDDA.t124 61.6417
R1987 VDDA.n816 VDDA.n301 58.0576
R1988 VDDA.n786 VDDA.n316 58.0576
R1989 VDDA.n721 VDDA.n720 58.0576
R1990 VDDA.n699 VDDA.n698 58.0576
R1991 VDDA.n689 VDDA.n335 58.0576
R1992 VDDA.n816 VDDA.n302 58.0576
R1993 VDDA.n786 VDDA.n785 58.0576
R1994 VDDA.n714 VDDA.n713 58.0576
R1995 VDDA.n697 VDDA.n331 58.0576
R1996 VDDA.n690 VDDA.n334 58.0576
R1997 VDDA.n656 VDDA.n338 57.2449
R1998 VDDA.n672 VDDA.n671 57.2449
R1999 VDDA.n607 VDDA.n606 57.2449
R2000 VDDA.n593 VDDA.n592 57.2449
R2001 VDDA.n652 VDDA.n338 57.2449
R2002 VDDA.n606 VDDA.n358 57.2449
R2003 VDDA.n165 VDDA.n53 54.4005
R2004 VDDA.n93 VDDA.n44 54.4005
R2005 VDDA.n210 VDDA.n35 54.4005
R2006 VDDA.n259 VDDA.n17 54.4005
R2007 VDDA.n89 VDDA.n1 54.4005
R2008 VDDA.n96 VDDA.n62 54.4005
R2009 VDDA.n803 VDDA.n307 54.4005
R2010 VDDA.n309 VDDA.n307 54.4005
R2011 VDDA.n309 VDDA.n308 54.4005
R2012 VDDA.n803 VDDA.n308 54.4005
R2013 VDDA.n85 VDDA.n84 53.3664
R2014 VDDA.n79 VDDA.n77 53.3664
R2015 VDDA.n115 VDDA.n109 53.3664
R2016 VDDA.n117 VDDA.n73 53.3664
R2017 VDDA.n107 VDDA.n98 53.3664
R2018 VDDA.n100 VDDA.n88 53.3664
R2019 VDDA.n732 VDDA.n731 53.3664
R2020 VDDA.n753 VDDA.n747 53.3664
R2021 VDDA.n775 VDDA.n774 53.3664
R2022 VDDA.n626 VDDA.n625 53.3664
R2023 VDDA.n620 VDDA.n619 53.3664
R2024 VDDA.n712 VDDA.n326 53.3664
R2025 VDDA.n710 VDDA.n709 53.3664
R2026 VDDA.n784 VDDA.n318 53.3664
R2027 VDDA.n758 VDDA.n748 53.3664
R2028 VDDA.n738 VDDA.n737 53.3664
R2029 VDDA.n634 VDDA.n628 53.3664
R2030 VDDA.n630 VDDA.n618 53.3664
R2031 VDDA.n704 VDDA.n328 53.3664
R2032 VDDA.n700 VDDA.n327 53.3664
R2033 VDDA.n726 VDDA.n320 53.3664
R2034 VDDA.n722 VDDA.n319 53.3664
R2035 VDDA.n782 VDDA.n776 53.3664
R2036 VDDA.n778 VDDA.n728 53.3664
R2037 VDDA.n769 VDDA.n759 53.3664
R2038 VDDA.n764 VDDA.n729 53.3664
R2039 VDDA.n745 VDDA.n739 53.3664
R2040 VDDA.n741 VDDA.n730 53.3664
R2041 VDDA.n641 VDDA.n616 53.3664
R2042 VDDA.n637 VDDA.n616 53.3664
R2043 VDDA.n408 VDDA.t80 50.7639
R2044 VDDA.t169 VDDA.n385 49.2505
R2045 VDDA.n385 VDDA.t102 49.2505
R2046 VDDA.n378 VDDA.t46 49.2505
R2047 VDDA.n378 VDDA.t76 49.2505
R2048 VDDA.n409 VDDA.t151 49.2505
R2049 VDDA.n409 VDDA.t109 49.2505
R2050 VDDA.n389 VDDA.t111 49.2505
R2051 VDDA.n389 VDDA.t154 49.2505
R2052 VDDA.n382 VDDA.t118 49.2505
R2053 VDDA.n382 VDDA.t139 49.2505
R2054 VDDA.n384 VDDA.t32 49.2505
R2055 VDDA.n384 VDDA.t175 49.2505
R2056 VDDA.n818 VDDA.n817 47.7005
R2057 VDDA.n648 VDDA.n644 45.3071
R2058 VDDA.n355 VDDA.n347 45.3071
R2059 VDDA.n356 VDDA.n348 45.3071
R2060 VDDA.n653 VDDA.n645 45.3071
R2061 VDDA.n589 VDDA.n585 45.3071
R2062 VDDA.n591 VDDA.n584 45.3071
R2063 VDDA.n613 VDDA.n349 45.3071
R2064 VDDA.n608 VDDA.n346 45.3071
R2065 VDDA.n668 VDDA.n664 45.3071
R2066 VDDA.n670 VDDA.n345 45.3071
R2067 VDDA.n662 VDDA.n654 45.3071
R2068 VDDA.n657 VDDA.n615 45.3071
R2069 VDDA.n418 VDDA.n388 45.3071
R2070 VDDA.n424 VDDA.n415 45.3071
R2071 VDDA.n395 VDDA.n393 45.3071
R2072 VDDA.n400 VDDA.n394 45.3071
R2073 VDDA.n401 VDDA.n393 45.3071
R2074 VDDA.n562 VDDA.n479 45.3071
R2075 VDDA.n484 VDDA.n478 45.3071
R2076 VDDA.n570 VDDA.n477 45.3071
R2077 VDDA.n568 VDDA.n567 45.3071
R2078 VDDA.n527 VDDA.n526 45.3071
R2079 VDDA.n526 VDDA.n523 45.3071
R2080 VDDA.n437 VDDA.n379 41.6005
R2081 VDDA.t3 VDDA.t148 39.886
R2082 VDDA.n431 VDDA.n380 39.4988
R2083 VDDA.n579 VDDA.n578 38.1005
R2084 VDDA.n413 VDDA.t161 36.26
R2085 VDDA.t103 VDDA.t108 32.6341
R2086 VDDA.t124 VDDA.t146 32.6341
R2087 VDDA.n561 VDDA.n480 32.2291
R2088 VDDA.n120 VDDA.n70 32.0005
R2089 VDDA.n124 VDDA.n70 32.0005
R2090 VDDA.n125 VDDA.n124 32.0005
R2091 VDDA.n126 VDDA.n125 32.0005
R2092 VDDA.n132 VDDA.n131 32.0005
R2093 VDDA.n135 VDDA.n132 32.0005
R2094 VDDA.n139 VDDA.n64 32.0005
R2095 VDDA.n140 VDDA.n139 32.0005
R2096 VDDA.n141 VDDA.n140 32.0005
R2097 VDDA.n145 VDDA.n144 32.0005
R2098 VDDA.n146 VDDA.n145 32.0005
R2099 VDDA.n146 VDDA.n60 32.0005
R2100 VDDA.n150 VDDA.n60 32.0005
R2101 VDDA.n151 VDDA.n150 32.0005
R2102 VDDA.n153 VDDA.n57 32.0005
R2103 VDDA.n157 VDDA.n57 32.0005
R2104 VDDA.n160 VDDA.n159 32.0005
R2105 VDDA.n160 VDDA.n54 32.0005
R2106 VDDA.n164 VDDA.n54 32.0005
R2107 VDDA.n167 VDDA.n166 32.0005
R2108 VDDA.n167 VDDA.n51 32.0005
R2109 VDDA.n171 VDDA.n51 32.0005
R2110 VDDA.n172 VDDA.n171 32.0005
R2111 VDDA.n173 VDDA.n172 32.0005
R2112 VDDA.n177 VDDA.n176 32.0005
R2113 VDDA.n180 VDDA.n177 32.0005
R2114 VDDA.n184 VDDA.n46 32.0005
R2115 VDDA.n185 VDDA.n184 32.0005
R2116 VDDA.n186 VDDA.n185 32.0005
R2117 VDDA.n190 VDDA.n189 32.0005
R2118 VDDA.n191 VDDA.n190 32.0005
R2119 VDDA.n191 VDDA.n42 32.0005
R2120 VDDA.n195 VDDA.n42 32.0005
R2121 VDDA.n196 VDDA.n195 32.0005
R2122 VDDA.n198 VDDA.n39 32.0005
R2123 VDDA.n202 VDDA.n39 32.0005
R2124 VDDA.n205 VDDA.n204 32.0005
R2125 VDDA.n205 VDDA.n36 32.0005
R2126 VDDA.n209 VDDA.n36 32.0005
R2127 VDDA.n212 VDDA.n211 32.0005
R2128 VDDA.n212 VDDA.n33 32.0005
R2129 VDDA.n216 VDDA.n33 32.0005
R2130 VDDA.n217 VDDA.n216 32.0005
R2131 VDDA.n220 VDDA.n217 32.0005
R2132 VDDA.n224 VDDA.n31 32.0005
R2133 VDDA.n225 VDDA.n224 32.0005
R2134 VDDA.n226 VDDA.n225 32.0005
R2135 VDDA.n230 VDDA.n229 32.0005
R2136 VDDA.n231 VDDA.n230 32.0005
R2137 VDDA.n231 VDDA.n26 32.0005
R2138 VDDA.n235 VDDA.n26 32.0005
R2139 VDDA.n239 VDDA.n237 32.0005
R2140 VDDA.n243 VDDA.n24 32.0005
R2141 VDDA.n244 VDDA.n243 32.0005
R2142 VDDA.n246 VDDA.n21 32.0005
R2143 VDDA.n250 VDDA.n21 32.0005
R2144 VDDA.n251 VDDA.n250 32.0005
R2145 VDDA.n253 VDDA.n18 32.0005
R2146 VDDA.n257 VDDA.n18 32.0005
R2147 VDDA.n258 VDDA.n257 32.0005
R2148 VDDA.n260 VDDA.n15 32.0005
R2149 VDDA.n264 VDDA.n15 32.0005
R2150 VDDA.n265 VDDA.n264 32.0005
R2151 VDDA.n266 VDDA.n265 32.0005
R2152 VDDA.n266 VDDA.n13 32.0005
R2153 VDDA.n270 VDDA.n13 32.0005
R2154 VDDA.n273 VDDA.n272 32.0005
R2155 VDDA.n273 VDDA.n10 32.0005
R2156 VDDA.n277 VDDA.n10 32.0005
R2157 VDDA.n278 VDDA.n277 32.0005
R2158 VDDA.n279 VDDA.n278 32.0005
R2159 VDDA.n283 VDDA.n282 32.0005
R2160 VDDA.n284 VDDA.n283 32.0005
R2161 VDDA.n284 VDDA.n5 32.0005
R2162 VDDA.n288 VDDA.n5 32.0005
R2163 VDDA.n289 VDDA.n288 32.0005
R2164 VDDA.n292 VDDA.n289 32.0005
R2165 VDDA.n296 VDDA.n3 32.0005
R2166 VDDA.n297 VDDA.n296 32.0005
R2167 VDDA.n298 VDDA.n297 32.0005
R2168 VDDA.n594 VDDA.n362 32.0005
R2169 VDDA.n598 VDDA.n362 32.0005
R2170 VDDA.n599 VDDA.n598 32.0005
R2171 VDDA.n600 VDDA.n599 32.0005
R2172 VDDA.n600 VDDA.n359 32.0005
R2173 VDDA.n606 VDDA.n359 32.0005
R2174 VDDA.n606 VDDA.n360 32.0005
R2175 VDDA.n360 VDDA.n342 32.0005
R2176 VDDA.n673 VDDA.n342 32.0005
R2177 VDDA.n677 VDDA.n340 32.0005
R2178 VDDA.n678 VDDA.n677 32.0005
R2179 VDDA.n679 VDDA.n678 32.0005
R2180 VDDA.n683 VDDA.n682 32.0005
R2181 VDDA.n684 VDDA.n683 32.0005
R2182 VDDA.n684 VDDA.n336 32.0005
R2183 VDDA.n688 VDDA.n336 32.0005
R2184 VDDA.n692 VDDA.n691 32.0005
R2185 VDDA.n692 VDDA.n330 32.0005
R2186 VDDA.n696 VDDA.n332 32.0005
R2187 VDDA.n719 VDDA.n322 32.0005
R2188 VDDA.n787 VDDA.n315 32.0005
R2189 VDDA.n791 VDDA.n313 32.0005
R2190 VDDA.n792 VDDA.n791 32.0005
R2191 VDDA.n793 VDDA.n792 32.0005
R2192 VDDA.n793 VDDA.n311 32.0005
R2193 VDDA.n797 VDDA.n311 32.0005
R2194 VDDA.n798 VDDA.n797 32.0005
R2195 VDDA.n799 VDDA.n798 32.0005
R2196 VDDA.n805 VDDA.n804 32.0005
R2197 VDDA.n805 VDDA.n305 32.0005
R2198 VDDA.n809 VDDA.n305 32.0005
R2199 VDDA.n810 VDDA.n809 32.0005
R2200 VDDA.n811 VDDA.n810 32.0005
R2201 VDDA.n811 VDDA.n303 32.0005
R2202 VDDA.n815 VDDA.n303 32.0005
R2203 VDDA.n435 VDDA.n380 32.0005
R2204 VDDA.n436 VDDA.n435 32.0005
R2205 VDDA.n438 VDDA.n375 32.0005
R2206 VDDA.n443 VDDA.n375 32.0005
R2207 VDDA.n444 VDDA.n443 32.0005
R2208 VDDA.n445 VDDA.n444 32.0005
R2209 VDDA.n445 VDDA.n372 32.0005
R2210 VDDA.n450 VDDA.n372 32.0005
R2211 VDDA.n451 VDDA.n450 32.0005
R2212 VDDA.n452 VDDA.n451 32.0005
R2213 VDDA.n452 VDDA.n369 32.0005
R2214 VDDA.n457 VDDA.n369 32.0005
R2215 VDDA.n458 VDDA.n457 32.0005
R2216 VDDA.n459 VDDA.n458 32.0005
R2217 VDDA.n459 VDDA.n366 32.0005
R2218 VDDA.n464 VDDA.n366 32.0005
R2219 VDDA.n465 VDDA.n464 32.0005
R2220 VDDA.n465 VDDA.n364 32.0005
R2221 VDDA.n469 VDDA.n364 32.0005
R2222 VDDA.n470 VDDA.n469 32.0005
R2223 VDDA.n574 VDDA.n472 32.0005
R2224 VDDA.n578 VDDA.n472 32.0005
R2225 VDDA.n498 VDDA.n497 32.0005
R2226 VDDA.n497 VDDA.n496 32.0005
R2227 VDDA.n504 VDDA.n486 32.0005
R2228 VDDA.n504 VDDA.n503 32.0005
R2229 VDDA.n503 VDDA.n502 32.0005
R2230 VDDA.n553 VDDA.n508 32.0005
R2231 VDDA.n548 VDDA.n547 32.0005
R2232 VDDA.n541 VDDA.n540 32.0005
R2233 VDDA.n541 VDDA.n512 32.0005
R2234 VDDA.n545 VDDA.n512 32.0005
R2235 VDDA.n534 VDDA.n533 32.0005
R2236 VDDA.n534 VDDA.n515 32.0005
R2237 VDDA.n538 VDDA.n515 32.0005
R2238 VDDA.n428 VDDA.n427 30.754
R2239 VDDA.n392 VDDA.n391 30.754
R2240 VDDA.n80 VDDA.n71 30.2632
R2241 VDDA.n412 VDDA.n411 30.186
R2242 VDDA.n387 VDDA.n386 30.186
R2243 VDDA.n131 VDDA.n67 28.8005
R2244 VDDA.n144 VDDA.n62 28.8005
R2245 VDDA.n153 VDDA.n152 28.8005
R2246 VDDA.n166 VDDA.n165 28.8005
R2247 VDDA.n176 VDDA.n49 28.8005
R2248 VDDA.n189 VDDA.n44 28.8005
R2249 VDDA.n198 VDDA.n197 28.8005
R2250 VDDA.n211 VDDA.n210 28.8005
R2251 VDDA.n246 VDDA.n245 28.8005
R2252 VDDA.n271 VDDA.n270 28.8005
R2253 VDDA.n673 VDDA.n672 28.8005
R2254 VDDA.n573 VDDA.n474 28.8005
R2255 VDDA.n498 VDDA.n489 28.8005
R2256 VDDA.n554 VDDA.n553 28.8005
R2257 VDDA.n259 VDDA.n258 25.6005
R2258 VDDA.n594 VDDA.n593 25.6005
R2259 VDDA.n679 VDDA.n338 25.6005
R2260 VDDA.n691 VDDA.n690 25.6005
R2261 VDDA.n715 VDDA.n714 25.6005
R2262 VDDA.n720 VDDA.n315 25.6005
R2263 VDDA.n787 VDDA.n786 25.6005
R2264 VDDA.n802 VDDA.n309 25.6005
R2265 VDDA.n803 VDDA.n802 25.6005
R2266 VDDA.n817 VDDA.n816 25.6005
R2267 VDDA.n437 VDDA.n436 25.6005
R2268 VDDA VDDA.n470 25.6005
R2269 VDDA.t38 VDDA.t110 25.3822
R2270 VDDA.t153 VDDA.t190 25.3822
R2271 VDDA.n119 VDDA.n118 24.991
R2272 VDDA.n101 VDDA.n68 24.991
R2273 VDDA.n818 VDDA.n300 24.8806
R2274 VDDA.n655 VDDA.t78 24.6255
R2275 VDDA.n344 VDDA.t127 24.6255
R2276 VDDA.n350 VDDA.t19 24.6255
R2277 VDDA.n583 VDDA.t96 24.6255
R2278 VDDA.n646 VDDA.t105 24.6255
R2279 VDDA.n351 VDDA.t12 24.6255
R2280 VDDA.n491 VDDA.t72 24.6255
R2281 VDDA.n491 VDDA.t182 24.6255
R2282 VDDA.n488 VDDA.t53 24.6255
R2283 VDDA.n488 VDDA.t137 24.6255
R2284 VDDA.t179 VDDA.n555 24.6255
R2285 VDDA.n555 VDDA.t89 24.6255
R2286 VDDA.n511 VDDA.t135 24.6255
R2287 VDDA.n511 VDDA.t165 24.6255
R2288 VDDA.n514 VDDA.t131 24.6255
R2289 VDDA.n514 VDDA.t14 24.6255
R2290 VDDA.n531 VDDA.t172 24.6255
R2291 VDDA.n531 VDDA.t65 24.6255
R2292 VDDA.t172 VDDA.n530 24.6255
R2293 VDDA.n475 VDDA.t183 24.6255
R2294 VDDA.n556 VDDA.t179 24.6255
R2295 VDDA.n560 VDDA.t166 24.6255
R2296 VDDA.n520 VDDA.n517 24.361
R2297 VDDA.n129 VDDA.n128 24.1919
R2298 VDDA.n300 VDDA.n1 23.4989
R2299 VDDA.n120 VDDA.n119 22.4005
R2300 VDDA.n126 VDDA.n68 22.4005
R2301 VDDA.n135 VDDA.n134 22.4005
R2302 VDDA.n158 VDDA.n157 22.4005
R2303 VDDA.n180 VDDA.n179 22.4005
R2304 VDDA.n203 VDDA.n202 22.4005
R2305 VDDA.n219 VDDA.n31 22.4005
R2306 VDDA.n226 VDDA.n29 22.4005
R2307 VDDA.n291 VDDA.n3 22.4005
R2308 VDDA.n496 VDDA.n492 22.4005
R2309 VDDA.n547 VDDA.n546 22.4005
R2310 VDDA.n548 VDDA.n480 22.4005
R2311 VDDA.n405 VDDA.n396 22.0449
R2312 VDDA.n416 VDDA.t162 19.7005
R2313 VDDA.n397 VDDA.t159 19.7005
R2314 VDDA.n367 VDDA.t125 19.7005
R2315 VDDA.n367 VDDA.t158 19.7005
R2316 VDDA.n370 VDDA.t4 19.7005
R2317 VDDA.n370 VDDA.t113 19.7005
R2318 VDDA.n373 VDDA.t191 19.7005
R2319 VDDA.n373 VDDA.t81 19.7005
R2320 VDDA.n376 VDDA.t141 19.7005
R2321 VDDA.n376 VDDA.t39 19.7005
R2322 VDDA.t162 VDDA.n381 19.7005
R2323 VDDA.n381 VDDA.t104 19.7005
R2324 VDDA.n237 VDDA.n236 19.2005
R2325 VDDA.n239 VDDA.n238 19.2005
R2326 VDDA.n279 VDDA.n8 19.2005
R2327 VDDA.n332 VDDA.n324 19.2005
R2328 VDDA.t45 VDDA.t140 18.1303
R2329 VDDA.t145 VDDA.t157 18.1303
R2330 VDDA.n573 VDDA.n572 17.6005
R2331 VDDA.n252 VDDA.n251 16.0005
R2332 VDDA.n253 VDDA.n252 16.0005
R2333 VDDA.n298 VDDA.n1 16.0005
R2334 VDDA.n697 VDDA.n696 16.0005
R2335 VDDA.n429 VDDA.n428 16.0005
R2336 VDDA.n391 VDDA.n390 16.0005
R2337 VDDA.n411 VDDA.n410 16.0005
R2338 VDDA.n386 VDDA.n383 16.0005
R2339 VDDA.n492 VDDA.n474 16.0005
R2340 VDDA.n508 VDDA.n480 16.0005
R2341 VDDA.n546 VDDA.n545 16.0005
R2342 VDDA.n533 VDDA.n532 16.0005
R2343 VDDA.n471 VDDA 15.7005
R2344 VDDA.n572 VDDA.n571 15.6449
R2345 VDDA.n529 VDDA.n520 15.6449
R2346 VDDA.n593 VDDA.n581 13.8989
R2347 VDDA.n236 VDDA.n235 12.8005
R2348 VDDA.n238 VDDA.n24 12.8005
R2349 VDDA.n282 VDDA.n8 12.8005
R2350 VDDA.n698 VDDA.n330 12.8005
R2351 VDDA.n715 VDDA.n324 12.8005
R2352 VDDA.n580 VDDA.n471 12.7493
R2353 VDDA.n581 VDDA.n580 12.3383
R2354 VDDA.n580 VDDA.n579 11.579
R2355 VDDA.n643 VDDA.t196 11.4924
R2356 VDDA.t115 VDDA.n635 11.4924
R2357 VDDA.n627 VDDA.t206 11.4924
R2358 VDDA.n705 VDDA.t219 11.4924
R2359 VDDA.n711 VDDA.t198 11.4924
R2360 VDDA.t90 VDDA.t112 10.8784
R2361 VDDA.n129 VDDA.n67 10.7016
R2362 VDDA.n396 VDDA.n365 9.613
R2363 VDDA.n134 VDDA.n64 9.6005
R2364 VDDA.n159 VDDA.n158 9.6005
R2365 VDDA.n179 VDDA.n46 9.6005
R2366 VDDA.n204 VDDA.n203 9.6005
R2367 VDDA.n220 VDDA.n219 9.6005
R2368 VDDA.n229 VDDA.n29 9.6005
R2369 VDDA.n292 VDDA.n291 9.6005
R2370 VDDA.n574 VDDA.n573 9.6005
R2371 VDDA.n554 VDDA.n486 9.6005
R2372 VDDA.n502 VDDA.n489 9.6005
R2373 VDDA.n121 VDDA.n120 9.3005
R2374 VDDA.n122 VDDA.n70 9.3005
R2375 VDDA.n124 VDDA.n123 9.3005
R2376 VDDA.n125 VDDA.n69 9.3005
R2377 VDDA.n127 VDDA.n126 9.3005
R2378 VDDA.n131 VDDA.n130 9.3005
R2379 VDDA.n132 VDDA.n65 9.3005
R2380 VDDA.n136 VDDA.n135 9.3005
R2381 VDDA.n137 VDDA.n64 9.3005
R2382 VDDA.n139 VDDA.n138 9.3005
R2383 VDDA.n140 VDDA.n63 9.3005
R2384 VDDA.n142 VDDA.n141 9.3005
R2385 VDDA.n144 VDDA.n143 9.3005
R2386 VDDA.n145 VDDA.n61 9.3005
R2387 VDDA.n147 VDDA.n146 9.3005
R2388 VDDA.n148 VDDA.n60 9.3005
R2389 VDDA.n150 VDDA.n149 9.3005
R2390 VDDA.n151 VDDA.n58 9.3005
R2391 VDDA.n154 VDDA.n153 9.3005
R2392 VDDA.n155 VDDA.n57 9.3005
R2393 VDDA.n157 VDDA.n156 9.3005
R2394 VDDA.n159 VDDA.n55 9.3005
R2395 VDDA.n161 VDDA.n160 9.3005
R2396 VDDA.n162 VDDA.n54 9.3005
R2397 VDDA.n164 VDDA.n163 9.3005
R2398 VDDA.n166 VDDA.n52 9.3005
R2399 VDDA.n168 VDDA.n167 9.3005
R2400 VDDA.n169 VDDA.n51 9.3005
R2401 VDDA.n171 VDDA.n170 9.3005
R2402 VDDA.n172 VDDA.n50 9.3005
R2403 VDDA.n174 VDDA.n173 9.3005
R2404 VDDA.n176 VDDA.n175 9.3005
R2405 VDDA.n177 VDDA.n47 9.3005
R2406 VDDA.n181 VDDA.n180 9.3005
R2407 VDDA.n182 VDDA.n46 9.3005
R2408 VDDA.n184 VDDA.n183 9.3005
R2409 VDDA.n185 VDDA.n45 9.3005
R2410 VDDA.n187 VDDA.n186 9.3005
R2411 VDDA.n189 VDDA.n188 9.3005
R2412 VDDA.n190 VDDA.n43 9.3005
R2413 VDDA.n192 VDDA.n191 9.3005
R2414 VDDA.n193 VDDA.n42 9.3005
R2415 VDDA.n195 VDDA.n194 9.3005
R2416 VDDA.n196 VDDA.n40 9.3005
R2417 VDDA.n199 VDDA.n198 9.3005
R2418 VDDA.n200 VDDA.n39 9.3005
R2419 VDDA.n202 VDDA.n201 9.3005
R2420 VDDA.n204 VDDA.n37 9.3005
R2421 VDDA.n206 VDDA.n205 9.3005
R2422 VDDA.n207 VDDA.n36 9.3005
R2423 VDDA.n209 VDDA.n208 9.3005
R2424 VDDA.n211 VDDA.n34 9.3005
R2425 VDDA.n213 VDDA.n212 9.3005
R2426 VDDA.n214 VDDA.n33 9.3005
R2427 VDDA.n216 VDDA.n215 9.3005
R2428 VDDA.n217 VDDA.n32 9.3005
R2429 VDDA.n221 VDDA.n220 9.3005
R2430 VDDA.n222 VDDA.n31 9.3005
R2431 VDDA.n224 VDDA.n223 9.3005
R2432 VDDA.n225 VDDA.n30 9.3005
R2433 VDDA.n227 VDDA.n226 9.3005
R2434 VDDA.n229 VDDA.n228 9.3005
R2435 VDDA.n230 VDDA.n27 9.3005
R2436 VDDA.n232 VDDA.n231 9.3005
R2437 VDDA.n233 VDDA.n26 9.3005
R2438 VDDA.n235 VDDA.n234 9.3005
R2439 VDDA.n237 VDDA.n25 9.3005
R2440 VDDA.n240 VDDA.n239 9.3005
R2441 VDDA.n241 VDDA.n24 9.3005
R2442 VDDA.n243 VDDA.n242 9.3005
R2443 VDDA.n244 VDDA.n22 9.3005
R2444 VDDA.n247 VDDA.n246 9.3005
R2445 VDDA.n248 VDDA.n21 9.3005
R2446 VDDA.n250 VDDA.n249 9.3005
R2447 VDDA.n251 VDDA.n19 9.3005
R2448 VDDA.n254 VDDA.n253 9.3005
R2449 VDDA.n255 VDDA.n18 9.3005
R2450 VDDA.n257 VDDA.n256 9.3005
R2451 VDDA.n258 VDDA.n16 9.3005
R2452 VDDA.n261 VDDA.n260 9.3005
R2453 VDDA.n262 VDDA.n15 9.3005
R2454 VDDA.n264 VDDA.n263 9.3005
R2455 VDDA.n265 VDDA.n14 9.3005
R2456 VDDA.n267 VDDA.n266 9.3005
R2457 VDDA.n268 VDDA.n13 9.3005
R2458 VDDA.n270 VDDA.n269 9.3005
R2459 VDDA.n272 VDDA.n11 9.3005
R2460 VDDA.n274 VDDA.n273 9.3005
R2461 VDDA.n275 VDDA.n10 9.3005
R2462 VDDA.n277 VDDA.n276 9.3005
R2463 VDDA.n278 VDDA.n9 9.3005
R2464 VDDA.n280 VDDA.n279 9.3005
R2465 VDDA.n282 VDDA.n281 9.3005
R2466 VDDA.n283 VDDA.n6 9.3005
R2467 VDDA.n285 VDDA.n284 9.3005
R2468 VDDA.n286 VDDA.n5 9.3005
R2469 VDDA.n288 VDDA.n287 9.3005
R2470 VDDA.n289 VDDA.n4 9.3005
R2471 VDDA.n293 VDDA.n292 9.3005
R2472 VDDA.n294 VDDA.n3 9.3005
R2473 VDDA.n296 VDDA.n295 9.3005
R2474 VDDA.n297 VDDA.n2 9.3005
R2475 VDDA.n299 VDDA.n298 9.3005
R2476 VDDA.n470 VDDA.n363 9.3005
R2477 VDDA.n469 VDDA.n468 9.3005
R2478 VDDA.n467 VDDA.n364 9.3005
R2479 VDDA.n466 VDDA.n465 9.3005
R2480 VDDA.n464 VDDA.n463 9.3005
R2481 VDDA.n462 VDDA.n366 9.3005
R2482 VDDA.n460 VDDA.n459 9.3005
R2483 VDDA.n458 VDDA.n368 9.3005
R2484 VDDA.n457 VDDA.n456 9.3005
R2485 VDDA.n455 VDDA.n369 9.3005
R2486 VDDA.n453 VDDA.n452 9.3005
R2487 VDDA.n451 VDDA.n371 9.3005
R2488 VDDA.n450 VDDA.n449 9.3005
R2489 VDDA.n448 VDDA.n372 9.3005
R2490 VDDA.n446 VDDA.n445 9.3005
R2491 VDDA.n444 VDDA.n374 9.3005
R2492 VDDA.n443 VDDA.n442 9.3005
R2493 VDDA.n441 VDDA.n375 9.3005
R2494 VDDA.n439 VDDA.n438 9.3005
R2495 VDDA.n433 VDDA.n380 9.3005
R2496 VDDA.n435 VDDA.n434 9.3005
R2497 VDDA.n436 VDDA.n377 9.3005
R2498 VDDA.n533 VDDA.n516 9.3005
R2499 VDDA.n535 VDDA.n534 9.3005
R2500 VDDA.n536 VDDA.n515 9.3005
R2501 VDDA.n538 VDDA.n537 9.3005
R2502 VDDA.n540 VDDA.n513 9.3005
R2503 VDDA.n542 VDDA.n541 9.3005
R2504 VDDA.n543 VDDA.n512 9.3005
R2505 VDDA.n545 VDDA.n544 9.3005
R2506 VDDA.n546 VDDA.n510 9.3005
R2507 VDDA.n547 VDDA.n509 9.3005
R2508 VDDA.n549 VDDA.n548 9.3005
R2509 VDDA.n550 VDDA.n480 9.3005
R2510 VDDA.n551 VDDA.n508 9.3005
R2511 VDDA.n553 VDDA.n552 9.3005
R2512 VDDA.n554 VDDA.n507 9.3005
R2513 VDDA.n506 VDDA.n486 9.3005
R2514 VDDA.n505 VDDA.n504 9.3005
R2515 VDDA.n503 VDDA.n487 9.3005
R2516 VDDA.n502 VDDA.n501 9.3005
R2517 VDDA.n500 VDDA.n489 9.3005
R2518 VDDA.n499 VDDA.n498 9.3005
R2519 VDDA.n497 VDDA.n490 9.3005
R2520 VDDA.n496 VDDA.n495 9.3005
R2521 VDDA.n494 VDDA.n492 9.3005
R2522 VDDA.n493 VDDA.n474 9.3005
R2523 VDDA.n573 VDDA.n473 9.3005
R2524 VDDA.n575 VDDA.n574 9.3005
R2525 VDDA.n576 VDDA.n472 9.3005
R2526 VDDA.n578 VDDA.n577 9.3005
R2527 VDDA.n817 VDDA.n0 9.3005
R2528 VDDA.n595 VDDA.n594 9.3005
R2529 VDDA.n596 VDDA.n362 9.3005
R2530 VDDA.n598 VDDA.n597 9.3005
R2531 VDDA.n599 VDDA.n361 9.3005
R2532 VDDA.n601 VDDA.n600 9.3005
R2533 VDDA.n602 VDDA.n359 9.3005
R2534 VDDA.n606 VDDA.n605 9.3005
R2535 VDDA.n604 VDDA.n360 9.3005
R2536 VDDA.n603 VDDA.n342 9.3005
R2537 VDDA.n674 VDDA.n673 9.3005
R2538 VDDA.n675 VDDA.n340 9.3005
R2539 VDDA.n677 VDDA.n676 9.3005
R2540 VDDA.n678 VDDA.n339 9.3005
R2541 VDDA.n680 VDDA.n679 9.3005
R2542 VDDA.n682 VDDA.n681 9.3005
R2543 VDDA.n683 VDDA.n337 9.3005
R2544 VDDA.n685 VDDA.n684 9.3005
R2545 VDDA.n686 VDDA.n336 9.3005
R2546 VDDA.n688 VDDA.n687 9.3005
R2547 VDDA.n691 VDDA.n333 9.3005
R2548 VDDA.n693 VDDA.n692 9.3005
R2549 VDDA.n694 VDDA.n330 9.3005
R2550 VDDA.n696 VDDA.n695 9.3005
R2551 VDDA.n332 VDDA.n323 9.3005
R2552 VDDA.n716 VDDA.n715 9.3005
R2553 VDDA.n717 VDDA.n322 9.3005
R2554 VDDA.n719 VDDA.n718 9.3005
R2555 VDDA.n315 VDDA.n314 9.3005
R2556 VDDA.n788 VDDA.n787 9.3005
R2557 VDDA.n789 VDDA.n313 9.3005
R2558 VDDA.n791 VDDA.n790 9.3005
R2559 VDDA.n792 VDDA.n312 9.3005
R2560 VDDA.n794 VDDA.n793 9.3005
R2561 VDDA.n795 VDDA.n311 9.3005
R2562 VDDA.n797 VDDA.n796 9.3005
R2563 VDDA.n798 VDDA.n310 9.3005
R2564 VDDA.n800 VDDA.n799 9.3005
R2565 VDDA.n802 VDDA.n801 9.3005
R2566 VDDA.n804 VDDA.n306 9.3005
R2567 VDDA.n806 VDDA.n805 9.3005
R2568 VDDA.n807 VDDA.n305 9.3005
R2569 VDDA.n809 VDDA.n808 9.3005
R2570 VDDA.n810 VDDA.n304 9.3005
R2571 VDDA.n812 VDDA.n811 9.3005
R2572 VDDA.n813 VDDA.n303 9.3005
R2573 VDDA.n815 VDDA.n814 9.3005
R2574 VDDA.n112 VDDA.n111 9.14336
R2575 VDDA.n104 VDDA.n103 9.14336
R2576 VDDA.n742 VDDA.n740 9.14336
R2577 VDDA.n779 VDDA.n777 9.14336
R2578 VDDA.n723 VDDA.n321 9.14336
R2579 VDDA.n701 VDDA.n329 9.14336
R2580 VDDA.n631 VDDA.n629 9.14336
R2581 VDDA.n736 VDDA.n735 9.14336
R2582 VDDA.n773 VDDA.n772 9.14336
R2583 VDDA.n708 VDDA.n707 9.14336
R2584 VDDA.n624 VDDA.n623 9.14336
R2585 VDDA.n640 VDDA.n639 9.14336
R2586 VDDA.t17 VDDA.t24 7.66179
R2587 VDDA.n426 VDDA.n425 7.25241
R2588 VDDA.n661 VDDA.n660 7.11161
R2589 VDDA.n658 VDDA.n656 7.11161
R2590 VDDA.n667 VDDA.n666 7.11161
R2591 VDDA.n671 VDDA.n343 7.11161
R2592 VDDA.n612 VDDA.n611 7.11161
R2593 VDDA.n609 VDDA.n607 7.11161
R2594 VDDA.n588 VDDA.n587 7.11161
R2595 VDDA.n592 VDDA.n582 7.11161
R2596 VDDA.n652 VDDA.n651 7.11161
R2597 VDDA.n649 VDDA.n647 7.11161
R2598 VDDA.n358 VDDA.n357 7.11161
R2599 VDDA.n354 VDDA.n353 7.11161
R2600 VDDA.n423 VDDA.n422 7.11161
R2601 VDDA.n420 VDDA.n419 7.11161
R2602 VDDA.n405 VDDA.n404 7.11161
R2603 VDDA.n402 VDDA.n399 7.11161
R2604 VDDA.n571 VDDA.n476 7.11161
R2605 VDDA.n566 VDDA.n564 7.11161
R2606 VDDA.n529 VDDA.n528 7.11161
R2607 VDDA.n522 VDDA.n519 7.11161
R2608 VDDA.n128 VDDA.n68 7.05969
R2609 VDDA.n119 VDDA.n71 7.05957
R2610 VDDA.n532 VDDA.n517 6.54033
R2611 VDDA.n260 VDDA.n259 6.4005
R2612 VDDA.n682 VDDA.n338 6.4005
R2613 VDDA.n714 VDDA.n322 6.4005
R2614 VDDA.n720 VDDA.n719 6.4005
R2615 VDDA.n786 VDDA.n313 6.4005
R2616 VDDA.n799 VDDA.n309 6.4005
R2617 VDDA.n804 VDDA.n803 6.4005
R2618 VDDA.n816 VDDA.n815 6.4005
R2619 VDDA.n438 VDDA.n437 6.4005
R2620 VDDA.n83 VDDA.n82 5.81868
R2621 VDDA.n765 VDDA.n761 5.81868
R2622 VDDA.n754 VDDA.n750 5.81868
R2623 VDDA.n106 VDDA.n105 5.33286
R2624 VDDA.n114 VDDA.n113 5.33286
R2625 VDDA.n118 VDDA.n72 5.33286
R2626 VDDA.n102 VDDA.n101 5.33286
R2627 VDDA.n636 VDDA.n334 5.33286
R2628 VDDA.n743 VDDA.n301 5.33286
R2629 VDDA.n780 VDDA.n316 5.33286
R2630 VDDA.n724 VDDA.n721 5.33286
R2631 VDDA.n702 VDDA.n699 5.33286
R2632 VDDA.n632 VDDA.n335 5.33286
R2633 VDDA.n733 VDDA.n302 5.33286
R2634 VDDA.n785 VDDA.n317 5.33286
R2635 VDDA.n713 VDDA.n325 5.33286
R2636 VDDA.n621 VDDA.n331 5.33286
R2637 VDDA.n113 VDDA.n112 3.75335
R2638 VDDA.n111 VDDA.n72 3.75335
R2639 VDDA.n105 VDDA.n104 3.75335
R2640 VDDA.n103 VDDA.n102 3.75335
R2641 VDDA.n744 VDDA.n740 3.75335
R2642 VDDA.n743 VDDA.n742 3.75335
R2643 VDDA.n781 VDDA.n777 3.75335
R2644 VDDA.n780 VDDA.n779 3.75335
R2645 VDDA.n725 VDDA.n321 3.75335
R2646 VDDA.n724 VDDA.n723 3.75335
R2647 VDDA.n703 VDDA.n329 3.75335
R2648 VDDA.n702 VDDA.n701 3.75335
R2649 VDDA.n633 VDDA.n629 3.75335
R2650 VDDA.n632 VDDA.n631 3.75335
R2651 VDDA.n736 VDDA.n733 3.75335
R2652 VDDA.n735 VDDA.n734 3.75335
R2653 VDDA.n772 VDDA.n317 3.75335
R2654 VDDA.n773 VDDA.n771 3.75335
R2655 VDDA.n707 VDDA.n325 3.75335
R2656 VDDA.n708 VDDA.n706 3.75335
R2657 VDDA.n624 VDDA.n621 3.75335
R2658 VDDA.n623 VDDA.n622 3.75335
R2659 VDDA.n640 VDDA.n636 3.75335
R2660 VDDA.n639 VDDA.n638 3.75335
R2661 VDDA.n660 VDDA.n659 3.53508
R2662 VDDA.n659 VDDA.n658 3.53508
R2663 VDDA.n666 VDDA.n665 3.53508
R2664 VDDA.n665 VDDA.n343 3.53508
R2665 VDDA.n611 VDDA.n610 3.53508
R2666 VDDA.n610 VDDA.n609 3.53508
R2667 VDDA.n587 VDDA.n586 3.53508
R2668 VDDA.n586 VDDA.n582 3.53508
R2669 VDDA.n651 VDDA.n650 3.53508
R2670 VDDA.n650 VDDA.n649 3.53508
R2671 VDDA.n357 VDDA.n352 3.53508
R2672 VDDA.n354 VDDA.n352 3.53508
R2673 VDDA.n422 VDDA.n421 3.53508
R2674 VDDA.n419 VDDA.n417 3.53508
R2675 VDDA.n421 VDDA.n420 3.53508
R2676 VDDA.n404 VDDA.n403 3.53508
R2677 VDDA.n399 VDDA.n398 3.53508
R2678 VDDA.n403 VDDA.n402 3.53508
R2679 VDDA.n565 VDDA.n476 3.53508
R2680 VDDA.n566 VDDA.n565 3.53508
R2681 VDDA.n528 VDDA.n518 3.53508
R2682 VDDA.n522 VDDA.n518 3.53508
R2683 VDDA.n86 VDDA.n76 3.40194
R2684 VDDA.n81 VDDA.n80 3.40194
R2685 VDDA.n768 VDDA.n767 3.40194
R2686 VDDA.n766 VDDA.n762 3.40194
R2687 VDDA.n757 VDDA.n756 3.40194
R2688 VDDA.n755 VDDA.n751 3.40194
R2689 VDDA.n141 VDDA.n62 3.2005
R2690 VDDA.n152 VDDA.n151 3.2005
R2691 VDDA.n165 VDDA.n164 3.2005
R2692 VDDA.n173 VDDA.n49 3.2005
R2693 VDDA.n186 VDDA.n44 3.2005
R2694 VDDA.n197 VDDA.n196 3.2005
R2695 VDDA.n210 VDDA.n209 3.2005
R2696 VDDA.n245 VDDA.n244 3.2005
R2697 VDDA.n272 VDDA.n271 3.2005
R2698 VDDA.n672 VDDA.n340 3.2005
R2699 VDDA.n689 VDDA.n688 3.2005
R2700 VDDA.n690 VDDA.n689 3.2005
R2701 VDDA.n698 VDDA.n697 3.2005
R2702 VDDA.n540 VDDA.n539 3.2005
R2703 VDDA.n539 VDDA.n538 3.2005
R2704 VDDA.n83 VDDA.n76 2.39444
R2705 VDDA.n82 VDDA.n81 2.39444
R2706 VDDA.n767 VDDA.n761 2.39444
R2707 VDDA.n766 VDDA.n765 2.39444
R2708 VDDA.n756 VDDA.n750 2.39444
R2709 VDDA.n755 VDDA.n754 2.39444
R2710 VDDA.n762 VDDA.n307 2.32777
R2711 VDDA.n757 VDDA.n308 2.32777
R2712 VDDA.n482 VDDA.n481 2.27782
R2713 VDDA.n483 VDDA.n482 2.27782
R2714 VDDA.n559 VDDA.n557 2.27782
R2715 VDDA.n485 VDDA.n483 2.27782
R2716 VDDA.n561 VDDA.n481 2.27782
R2717 VDDA.n557 VDDA.n485 2.27782
R2718 VDDA.n517 VDDA.n516 0.703395
R2719 VDDA.n121 VDDA.n71 0.203053
R2720 VDDA.n128 VDDA.n127 0.202927
R2721 VDDA.n595 VDDA.n581 0.193961
R2722 VDDA.n300 VDDA.n299 0.193958
R2723 VDDA.n130 VDDA.n129 0.193477
R2724 VDDA.n471 VDDA.n363 0.188
R2725 VDDA.n122 VDDA.n121 0.15675
R2726 VDDA.n123 VDDA.n122 0.15675
R2727 VDDA.n123 VDDA.n69 0.15675
R2728 VDDA.n127 VDDA.n69 0.15675
R2729 VDDA.n130 VDDA.n65 0.15675
R2730 VDDA.n136 VDDA.n65 0.15675
R2731 VDDA.n137 VDDA.n136 0.15675
R2732 VDDA.n138 VDDA.n137 0.15675
R2733 VDDA.n138 VDDA.n63 0.15675
R2734 VDDA.n142 VDDA.n63 0.15675
R2735 VDDA.n143 VDDA.n142 0.15675
R2736 VDDA.n143 VDDA.n61 0.15675
R2737 VDDA.n147 VDDA.n61 0.15675
R2738 VDDA.n148 VDDA.n147 0.15675
R2739 VDDA.n149 VDDA.n148 0.15675
R2740 VDDA.n149 VDDA.n58 0.15675
R2741 VDDA.n154 VDDA.n58 0.15675
R2742 VDDA.n155 VDDA.n154 0.15675
R2743 VDDA.n156 VDDA.n155 0.15675
R2744 VDDA.n156 VDDA.n55 0.15675
R2745 VDDA.n161 VDDA.n55 0.15675
R2746 VDDA.n162 VDDA.n161 0.15675
R2747 VDDA.n163 VDDA.n162 0.15675
R2748 VDDA.n163 VDDA.n52 0.15675
R2749 VDDA.n168 VDDA.n52 0.15675
R2750 VDDA.n169 VDDA.n168 0.15675
R2751 VDDA.n170 VDDA.n169 0.15675
R2752 VDDA.n170 VDDA.n50 0.15675
R2753 VDDA.n174 VDDA.n50 0.15675
R2754 VDDA.n175 VDDA.n174 0.15675
R2755 VDDA.n175 VDDA.n47 0.15675
R2756 VDDA.n181 VDDA.n47 0.15675
R2757 VDDA.n182 VDDA.n181 0.15675
R2758 VDDA.n183 VDDA.n182 0.15675
R2759 VDDA.n183 VDDA.n45 0.15675
R2760 VDDA.n187 VDDA.n45 0.15675
R2761 VDDA.n188 VDDA.n187 0.15675
R2762 VDDA.n188 VDDA.n43 0.15675
R2763 VDDA.n192 VDDA.n43 0.15675
R2764 VDDA.n193 VDDA.n192 0.15675
R2765 VDDA.n194 VDDA.n193 0.15675
R2766 VDDA.n194 VDDA.n40 0.15675
R2767 VDDA.n199 VDDA.n40 0.15675
R2768 VDDA.n200 VDDA.n199 0.15675
R2769 VDDA.n201 VDDA.n200 0.15675
R2770 VDDA.n201 VDDA.n37 0.15675
R2771 VDDA.n206 VDDA.n37 0.15675
R2772 VDDA.n207 VDDA.n206 0.15675
R2773 VDDA.n208 VDDA.n207 0.15675
R2774 VDDA.n208 VDDA.n34 0.15675
R2775 VDDA.n213 VDDA.n34 0.15675
R2776 VDDA.n214 VDDA.n213 0.15675
R2777 VDDA.n215 VDDA.n214 0.15675
R2778 VDDA.n215 VDDA.n32 0.15675
R2779 VDDA.n221 VDDA.n32 0.15675
R2780 VDDA.n222 VDDA.n221 0.15675
R2781 VDDA.n223 VDDA.n222 0.15675
R2782 VDDA.n223 VDDA.n30 0.15675
R2783 VDDA.n227 VDDA.n30 0.15675
R2784 VDDA.n228 VDDA.n227 0.15675
R2785 VDDA.n228 VDDA.n27 0.15675
R2786 VDDA.n232 VDDA.n27 0.15675
R2787 VDDA.n233 VDDA.n232 0.15675
R2788 VDDA.n234 VDDA.n233 0.15675
R2789 VDDA.n234 VDDA.n25 0.15675
R2790 VDDA.n240 VDDA.n25 0.15675
R2791 VDDA.n241 VDDA.n240 0.15675
R2792 VDDA.n242 VDDA.n241 0.15675
R2793 VDDA.n242 VDDA.n22 0.15675
R2794 VDDA.n247 VDDA.n22 0.15675
R2795 VDDA.n248 VDDA.n247 0.15675
R2796 VDDA.n249 VDDA.n248 0.15675
R2797 VDDA.n249 VDDA.n19 0.15675
R2798 VDDA.n254 VDDA.n19 0.15675
R2799 VDDA.n255 VDDA.n254 0.15675
R2800 VDDA.n256 VDDA.n255 0.15675
R2801 VDDA.n256 VDDA.n16 0.15675
R2802 VDDA.n261 VDDA.n16 0.15675
R2803 VDDA.n262 VDDA.n261 0.15675
R2804 VDDA.n263 VDDA.n262 0.15675
R2805 VDDA.n263 VDDA.n14 0.15675
R2806 VDDA.n267 VDDA.n14 0.15675
R2807 VDDA.n268 VDDA.n267 0.15675
R2808 VDDA.n269 VDDA.n268 0.15675
R2809 VDDA.n269 VDDA.n11 0.15675
R2810 VDDA.n274 VDDA.n11 0.15675
R2811 VDDA.n275 VDDA.n274 0.15675
R2812 VDDA.n276 VDDA.n275 0.15675
R2813 VDDA.n276 VDDA.n9 0.15675
R2814 VDDA.n280 VDDA.n9 0.15675
R2815 VDDA.n281 VDDA.n280 0.15675
R2816 VDDA.n281 VDDA.n6 0.15675
R2817 VDDA.n285 VDDA.n6 0.15675
R2818 VDDA.n286 VDDA.n285 0.15675
R2819 VDDA.n287 VDDA.n286 0.15675
R2820 VDDA.n287 VDDA.n4 0.15675
R2821 VDDA.n293 VDDA.n4 0.15675
R2822 VDDA.n294 VDDA.n293 0.15675
R2823 VDDA.n295 VDDA.n294 0.15675
R2824 VDDA.n295 VDDA.n2 0.15675
R2825 VDDA.n299 VDDA.n2 0.15675
R2826 VDDA.n434 VDDA.n433 0.15675
R2827 VDDA.n434 VDDA.n377 0.15675
R2828 VDDA.n439 VDDA.n377 0.15675
R2829 VDDA.n442 VDDA.n441 0.15675
R2830 VDDA.n442 VDDA.n374 0.15675
R2831 VDDA.n446 VDDA.n374 0.15675
R2832 VDDA.n449 VDDA.n448 0.15675
R2833 VDDA.n449 VDDA.n371 0.15675
R2834 VDDA.n453 VDDA.n371 0.15675
R2835 VDDA.n456 VDDA.n455 0.15675
R2836 VDDA.n456 VDDA.n368 0.15675
R2837 VDDA.n460 VDDA.n368 0.15675
R2838 VDDA.n463 VDDA.n462 0.15675
R2839 VDDA.n467 VDDA.n466 0.15675
R2840 VDDA.n468 VDDA.n467 0.15675
R2841 VDDA.n468 VDDA.n363 0.15675
R2842 VDDA.n535 VDDA.n516 0.15675
R2843 VDDA.n536 VDDA.n535 0.15675
R2844 VDDA.n537 VDDA.n536 0.15675
R2845 VDDA.n537 VDDA.n513 0.15675
R2846 VDDA.n542 VDDA.n513 0.15675
R2847 VDDA.n543 VDDA.n542 0.15675
R2848 VDDA.n544 VDDA.n543 0.15675
R2849 VDDA.n544 VDDA.n510 0.15675
R2850 VDDA.n510 VDDA.n509 0.15675
R2851 VDDA.n549 VDDA.n509 0.15675
R2852 VDDA.n550 VDDA.n549 0.15675
R2853 VDDA.n551 VDDA.n550 0.15675
R2854 VDDA.n552 VDDA.n551 0.15675
R2855 VDDA.n552 VDDA.n507 0.15675
R2856 VDDA.n507 VDDA.n506 0.15675
R2857 VDDA.n506 VDDA.n505 0.15675
R2858 VDDA.n505 VDDA.n487 0.15675
R2859 VDDA.n501 VDDA.n487 0.15675
R2860 VDDA.n501 VDDA.n500 0.15675
R2861 VDDA.n500 VDDA.n499 0.15675
R2862 VDDA.n499 VDDA.n490 0.15675
R2863 VDDA.n495 VDDA.n490 0.15675
R2864 VDDA.n495 VDDA.n494 0.15675
R2865 VDDA.n494 VDDA.n493 0.15675
R2866 VDDA.n493 VDDA.n473 0.15675
R2867 VDDA.n575 VDDA.n473 0.15675
R2868 VDDA.n576 VDDA.n575 0.15675
R2869 VDDA.n577 VDDA.n576 0.15675
R2870 VDDA.n596 VDDA.n595 0.15675
R2871 VDDA.n597 VDDA.n596 0.15675
R2872 VDDA.n597 VDDA.n361 0.15675
R2873 VDDA.n601 VDDA.n361 0.15675
R2874 VDDA.n602 VDDA.n601 0.15675
R2875 VDDA.n605 VDDA.n602 0.15675
R2876 VDDA.n605 VDDA.n604 0.15675
R2877 VDDA.n604 VDDA.n603 0.15675
R2878 VDDA.n675 VDDA.n674 0.15675
R2879 VDDA.n676 VDDA.n675 0.15675
R2880 VDDA.n676 VDDA.n339 0.15675
R2881 VDDA.n680 VDDA.n339 0.15675
R2882 VDDA.n681 VDDA.n680 0.15675
R2883 VDDA.n681 VDDA.n337 0.15675
R2884 VDDA.n685 VDDA.n337 0.15675
R2885 VDDA.n686 VDDA.n685 0.15675
R2886 VDDA.n687 VDDA.n686 0.15675
R2887 VDDA.n687 VDDA.n333 0.15675
R2888 VDDA.n693 VDDA.n333 0.15675
R2889 VDDA.n694 VDDA.n693 0.15675
R2890 VDDA.n695 VDDA.n694 0.15675
R2891 VDDA.n695 VDDA.n323 0.15675
R2892 VDDA.n716 VDDA.n323 0.15675
R2893 VDDA.n717 VDDA.n716 0.15675
R2894 VDDA.n718 VDDA.n717 0.15675
R2895 VDDA.n718 VDDA.n314 0.15675
R2896 VDDA.n788 VDDA.n314 0.15675
R2897 VDDA.n789 VDDA.n788 0.15675
R2898 VDDA.n790 VDDA.n789 0.15675
R2899 VDDA.n790 VDDA.n312 0.15675
R2900 VDDA.n794 VDDA.n312 0.15675
R2901 VDDA.n795 VDDA.n794 0.15675
R2902 VDDA.n796 VDDA.n795 0.15675
R2903 VDDA.n796 VDDA.n310 0.15675
R2904 VDDA.n800 VDDA.n310 0.15675
R2905 VDDA.n801 VDDA.n800 0.15675
R2906 VDDA.n801 VDDA.n306 0.15675
R2907 VDDA.n806 VDDA.n306 0.15675
R2908 VDDA.n807 VDDA.n806 0.15675
R2909 VDDA.n808 VDDA.n807 0.15675
R2910 VDDA.n808 VDDA.n304 0.15675
R2911 VDDA.n812 VDDA.n304 0.15675
R2912 VDDA.n813 VDDA.n812 0.15675
R2913 VDDA.n814 VDDA.n813 0.15675
R2914 VDDA.n814 VDDA.n0 0.15675
R2915 VDDA VDDA.n0 0.1255
R2916 VDDA.n577 VDDA 0.122375
R2917 VDDA.n432 VDDA.n431 0.100307
R2918 VDDA.n433 VDDA.n432 0.09425
R2919 VDDA.n441 VDDA.n440 0.09425
R2920 VDDA.n448 VDDA.n447 0.09425
R2921 VDDA.n455 VDDA.n454 0.09425
R2922 VDDA.n462 VDDA.n461 0.09425
R2923 VDDA.n466 VDDA.n365 0.09425
R2924 VDDA.n603 VDDA.n341 0.078625
R2925 VDDA.n674 VDDA.n341 0.078625
R2926 VDDA VDDA.n818 0.063
R2927 VDDA.n440 VDDA.n439 0.063
R2928 VDDA.n447 VDDA.n446 0.063
R2929 VDDA.n454 VDDA.n453 0.063
R2930 VDDA.n461 VDDA.n460 0.063
R2931 VDDA.n463 VDDA.n365 0.063
R2932 VDDA.n579 VDDA 0.0505
R2933 VCO_FD_magic_0.div120_2_0.div2.t4 VCO_FD_magic_0.div120_2_0.div2.t5 1012.2
R2934 VCO_FD_magic_0.div120_2_0.div2.n0 VCO_FD_magic_0.div120_2_0.div2.t0 663.801
R2935 VCO_FD_magic_0.div120_2_0.div2.n2 VCO_FD_magic_0.div120_2_0.div2.n1 431.401
R2936 VCO_FD_magic_0.div120_2_0.div2.t3 VCO_FD_magic_0.div120_2_0.div2.t6 401.668
R2937 VCO_FD_magic_0.div120_2_0.div2.n0 VCO_FD_magic_0.div120_2_0.div2.t4 361.692
R2938 VCO_FD_magic_0.div120_2_0.div2.n1 VCO_FD_magic_0.div120_2_0.div2.t2 353.467
R2939 VCO_FD_magic_0.div120_2_0.div2.t1 VCO_FD_magic_0.div120_2_0.div2.n2 298.921
R2940 VCO_FD_magic_0.div120_2_0.div2.n1 VCO_FD_magic_0.div120_2_0.div2.t3 257.067
R2941 VCO_FD_magic_0.div120_2_0.div2.n2 VCO_FD_magic_0.div120_2_0.div2.n0 67.2005
R2942 a_7630_n1440.n4 a_7630_n1440.t1 752.333
R2943 a_7630_n1440.t2 a_7630_n1440.n5 752.333
R2944 a_7630_n1440.n0 a_7630_n1440.t5 514.134
R2945 a_7630_n1440.n3 a_7630_n1440.n2 366.856
R2946 a_7630_n1440.n5 a_7630_n1440.t0 254.333
R2947 a_7630_n1440.n3 a_7630_n1440.t3 190.123
R2948 a_7630_n1440.n4 a_7630_n1440.n3 187.201
R2949 a_7630_n1440.n2 a_7630_n1440.n1 176.733
R2950 a_7630_n1440.n1 a_7630_n1440.n0 176.733
R2951 a_7630_n1440.n2 a_7630_n1440.t6 112.468
R2952 a_7630_n1440.n1 a_7630_n1440.t4 112.468
R2953 a_7630_n1440.n0 a_7630_n1440.t7 112.468
R2954 a_7630_n1440.n5 a_7630_n1440.n4 70.4005
R2955 pfd_8_0.QA_b.t4 pfd_8_0.QA_b.t6 1188.93
R2956 pfd_8_0.QA_b pfd_8_0.QA_b.n2 837.38
R2957 pfd_8_0.QA_b.t6 pfd_8_0.QA_b.t3 835.467
R2958 pfd_8_0.QA_b.n0 pfd_8_0.QA_b.t5 562.333
R2959 pfd_8_0.QA_b pfd_8_0.QA_b.n0 482
R2960 pfd_8_0.QA_b.n2 pfd_8_0.QA_b.n1 247.917
R2961 pfd_8_0.QA_b.n0 pfd_8_0.QA_b.t4 224.934
R2962 pfd_8_0.QA_b.n2 pfd_8_0.QA_b.t1 221.411
R2963 pfd_8_0.QA_b.n1 pfd_8_0.QA_b.t0 24.0005
R2964 pfd_8_0.QA_b.n1 pfd_8_0.QA_b.t2 24.0005
R2965 a_870_1400.t0 a_870_1400.t1 39.4005
R2966 pfd_8_0.DOWN_PFD_b.t1 pfd_8_0.DOWN_PFD_b.n1 203.528
R2967 pfd_8_0.DOWN_PFD_b.n0 pfd_8_0.DOWN_PFD_b.t2 203.528
R2968 pfd_8_0.DOWN_PFD_b.n1 pfd_8_0.DOWN_PFD_b.t0 183.935
R2969 pfd_8_0.DOWN_PFD_b.n0 pfd_8_0.DOWN_PFD_b.t3 183.935
R2970 pfd_8_0.DOWN_PFD_b.n1 pfd_8_0.DOWN_PFD_b.n0 83.2005
R2971 pfd_8_0.DOWN_b.n0 pfd_8_0.DOWN_b.t5 1028.27
R2972 pfd_8_0.DOWN_b.n2 pfd_8_0.DOWN_b.n1 569.734
R2973 pfd_8_0.DOWN_b.n1 pfd_8_0.DOWN_b.n0 465.933
R2974 pfd_8_0.DOWN_b.n1 pfd_8_0.DOWN_b.t3 401.668
R2975 pfd_8_0.DOWN_b.n0 pfd_8_0.DOWN_b.t4 385.601
R2976 pfd_8_0.DOWN_b.n1 pfd_8_0.DOWN_b.t2 385.601
R2977 pfd_8_0.DOWN_b.t0 pfd_8_0.DOWN_b.n2 211.847
R2978 pfd_8_0.DOWN_b.n2 pfd_8_0.DOWN_b.t1 173.055
R2979 VCO_FD_magic_0.div120_2_0.div5_2_0.J VCO_FD_magic_0.div120_2_0.div5_2_0.J.t1 710.734
R2980 VCO_FD_magic_0.div120_2_0.div5_2_0.J.n1 VCO_FD_magic_0.div120_2_0.div5_2_0.J.t4 553.534
R2981 VCO_FD_magic_0.div120_2_0.div5_2_0.J.n2 VCO_FD_magic_0.div120_2_0.div5_2_0.J.t0 254.333
R2982 VCO_FD_magic_0.div120_2_0.div5_2_0.J.n1 VCO_FD_magic_0.div120_2_0.div5_2_0.J.n0 206.333
R2983 VCO_FD_magic_0.div120_2_0.div5_2_0.J.n2 VCO_FD_magic_0.div120_2_0.div5_2_0.J.n1 70.4005
R2984 VCO_FD_magic_0.div120_2_0.div5_2_0.J.n0 VCO_FD_magic_0.div120_2_0.div5_2_0.J.t2 48.0005
R2985 VCO_FD_magic_0.div120_2_0.div5_2_0.J.n0 VCO_FD_magic_0.div120_2_0.div5_2_0.J.t3 48.0005
R2986 VCO_FD_magic_0.div120_2_0.div5_2_0.J VCO_FD_magic_0.div120_2_0.div5_2_0.J.n2 12.8005
R2987 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.n6 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.t0 777.4
R2988 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.t5 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.t6 514.134
R2989 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.n5 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.n4 364.178
R2990 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.t8 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.n0 353.467
R2991 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.n2 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.t2 353.467
R2992 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.n1 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.t8 318.702
R2993 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.n1 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.t5 307.909
R2994 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.n0 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.t3 289.2
R2995 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.n6 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.n5 257.079
R2996 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.t1 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.n7 233
R2997 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.n2 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.t11 192.8
R2998 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.n4 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.n3 176.733
R2999 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.n0 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.t9 112.468
R3000 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.n4 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.t10 112.468
R3001 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.n3 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.t4 112.468
R3002 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.n5 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.t7 112.468
R3003 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.n3 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.n2 96.4005
R3004 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.n7 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.n1 38.2642
R3005 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.n7 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.n6 21.3338
R3006 VCO_FD_magic_0.div120_2_0.div24.n3 VCO_FD_magic_0.div120_2_0.div24.n2 919.244
R3007 VCO_FD_magic_0.div120_2_0.div24 VCO_FD_magic_0.div120_2_0.div24.n7 912.303
R3008 VCO_FD_magic_0.div120_2_0.div24.t9 VCO_FD_magic_0.div120_2_0.div24.t11 819.4
R3009 VCO_FD_magic_0.div120_2_0.div24.n9 VCO_FD_magic_0.div120_2_0.div24.n8 628.734
R3010 VCO_FD_magic_0.div120_2_0.div24.n2 VCO_FD_magic_0.div120_2_0.div24.n1 520.361
R3011 VCO_FD_magic_0.div120_2_0.div24.n7 VCO_FD_magic_0.div120_2_0.div24.n6 364.178
R3012 VCO_FD_magic_0.div120_2_0.div24.n0 VCO_FD_magic_0.div120_2_0.div24.t8 337.401
R3013 VCO_FD_magic_0.div120_2_0.div24.n10 VCO_FD_magic_0.div120_2_0.div24.t9 336.25
R3014 VCO_FD_magic_0.div120_2_0.div24.n0 VCO_FD_magic_0.div120_2_0.div24.t13 305.267
R3015 VCO_FD_magic_0.div120_2_0.div24.n9 VCO_FD_magic_0.div120_2_0.div24.t1 257.534
R3016 VCO_FD_magic_0.div120_2_0.div24.n4 VCO_FD_magic_0.div120_2_0.div24.t12 192.8
R3017 VCO_FD_magic_0.div120_2_0.div24.n1 VCO_FD_magic_0.div120_2_0.div24.n0 176.733
R3018 VCO_FD_magic_0.div120_2_0.div24.n6 VCO_FD_magic_0.div120_2_0.div24.n5 176.733
R3019 VCO_FD_magic_0.div120_2_0.div24.n4 VCO_FD_magic_0.div120_2_0.div24.n3 160.667
R3020 VCO_FD_magic_0.div120_2_0.div24.n3 VCO_FD_magic_0.div120_2_0.div24.t7 144.601
R3021 VCO_FD_magic_0.div120_2_0.div24.n2 VCO_FD_magic_0.div120_2_0.div24.t4 131.976
R3022 VCO_FD_magic_0.div120_2_0.div24.n1 VCO_FD_magic_0.div120_2_0.div24.t3 128.534
R3023 VCO_FD_magic_0.div120_2_0.div24.n0 VCO_FD_magic_0.div120_2_0.div24.t6 128.534
R3024 VCO_FD_magic_0.div120_2_0.div24.n6 VCO_FD_magic_0.div120_2_0.div24.t14 112.468
R3025 VCO_FD_magic_0.div120_2_0.div24.n5 VCO_FD_magic_0.div120_2_0.div24.t5 112.468
R3026 VCO_FD_magic_0.div120_2_0.div24.n7 VCO_FD_magic_0.div120_2_0.div24.t10 112.468
R3027 VCO_FD_magic_0.div120_2_0.div24.n5 VCO_FD_magic_0.div120_2_0.div24.n4 96.4005
R3028 VCO_FD_magic_0.div120_2_0.div24.n8 VCO_FD_magic_0.div120_2_0.div24.t2 78.8005
R3029 VCO_FD_magic_0.div120_2_0.div24.n8 VCO_FD_magic_0.div120_2_0.div24.t0 78.8005
R3030 VCO_FD_magic_0.div120_2_0.div24.n10 VCO_FD_magic_0.div120_2_0.div24.n9 11.2005
R3031 VCO_FD_magic_0.div120_2_0.div24 VCO_FD_magic_0.div120_2_0.div24.n10 6.4005
R3032 VCO_FD_magic_0.div120_2_0.div3_3_0.H VCO_FD_magic_0.div120_2_0.div3_3_0.H.t1 710.734
R3033 VCO_FD_magic_0.div120_2_0.div3_3_0.H.n1 VCO_FD_magic_0.div120_2_0.div3_3_0.H.t4 553.534
R3034 VCO_FD_magic_0.div120_2_0.div3_3_0.H.n2 VCO_FD_magic_0.div120_2_0.div3_3_0.H.t0 254.333
R3035 VCO_FD_magic_0.div120_2_0.div3_3_0.H.n1 VCO_FD_magic_0.div120_2_0.div3_3_0.H.n0 206.333
R3036 VCO_FD_magic_0.div120_2_0.div3_3_0.H.n2 VCO_FD_magic_0.div120_2_0.div3_3_0.H.n1 70.4005
R3037 VCO_FD_magic_0.div120_2_0.div3_3_0.H.n0 VCO_FD_magic_0.div120_2_0.div3_3_0.H.t3 48.0005
R3038 VCO_FD_magic_0.div120_2_0.div3_3_0.H.n0 VCO_FD_magic_0.div120_2_0.div3_3_0.H.t2 48.0005
R3039 VCO_FD_magic_0.div120_2_0.div3_3_0.H VCO_FD_magic_0.div120_2_0.div3_3_0.H.n2 12.8005
R3040 VCO_FD_magic_0.div120_2_0.div3_3_0.I.n0 VCO_FD_magic_0.div120_2_0.div3_3_0.I.t1 663.801
R3041 VCO_FD_magic_0.div120_2_0.div3_3_0.I.t3 VCO_FD_magic_0.div120_2_0.div3_3_0.I.t2 514.134
R3042 VCO_FD_magic_0.div120_2_0.div3_3_0.I.n0 VCO_FD_magic_0.div120_2_0.div3_3_0.I.t3 479.284
R3043 VCO_FD_magic_0.div120_2_0.div3_3_0.I.n3 VCO_FD_magic_0.div120_2_0.div3_3_0.I.n2 344.8
R3044 VCO_FD_magic_0.div120_2_0.div3_3_0.I.n1 VCO_FD_magic_0.div120_2_0.div3_3_0.I.t5 289.2
R3045 VCO_FD_magic_0.div120_2_0.div3_3_0.I.t0 VCO_FD_magic_0.div120_2_0.div3_3_0.I.n3 275.454
R3046 VCO_FD_magic_0.div120_2_0.div3_3_0.I.n2 VCO_FD_magic_0.div120_2_0.div3_3_0.I.t4 241
R3047 VCO_FD_magic_0.div120_2_0.div3_3_0.I.n1 VCO_FD_magic_0.div120_2_0.div3_3_0.I.t6 112.468
R3048 VCO_FD_magic_0.div120_2_0.div3_3_0.I.n3 VCO_FD_magic_0.div120_2_0.div3_3_0.I.n0 97.9205
R3049 VCO_FD_magic_0.div120_2_0.div3_3_0.I.n2 VCO_FD_magic_0.div120_2_0.div3_3_0.I.n1 64.2672
R3050 pfd_8_0.DOWN.t3 pfd_8_0.DOWN.n0 605.311
R3051 charge_pump_cell_6_0.DOWN pfd_8_0.DOWN.t3 399.497
R3052 pfd_8_0.DOWN.n0 pfd_8_0.DOWN.t1 240.327
R3053 pfd_8_0.DOWN.n0 pfd_8_0.DOWN.t0 148.736
R3054 charge_pump_cell_6_0.DOWN pfd_8_0.DOWN.t2 24.487
R3055 pfd_8_0.UP_input.n2 pfd_8_0.UP_input.t3 326.658
R3056 pfd_8_0.UP_input.n4 pfd_8_0.UP_input.t6 297.233
R3057 pfd_8_0.UP_input.t5 pfd_8_0.UP_input.n5 297.233
R3058 pfd_8_0.UP_input.n3 pfd_8_0.UP_input.n1 257.067
R3059 pfd_8_0.UP_input.n7 pfd_8_0.UP_input.n6 246.275
R3060 pfd_8_0.UP_input.n0 pfd_8_0.UP_input.t2 241.928
R3061 pfd_8_0.UP_input.n6 pfd_8_0.UP_input.n1 226.942
R3062 pfd_8_0.UP_input.n3 pfd_8_0.UP_input.n2 226.942
R3063 pfd_8_0.UP_input.n5 pfd_8_0.UP_input.n4 216.9
R3064 pfd_8_0.UP_input.t1 pfd_8_0.UP_input.n7 209.928
R3065 pfd_8_0.UP_input.n0 pfd_8_0.UP_input.t0 145.536
R3066 pfd_8_0.UP_input.n7 pfd_8_0.UP_input.n0 144
R3067 pfd_8_0.UP_input.n2 pfd_8_0.UP_input.t6 92.3838
R3068 pfd_8_0.UP_input.n6 pfd_8_0.UP_input.t5 92.3838
R3069 pfd_8_0.UP_input.n4 pfd_8_0.UP_input.t7 80.3338
R3070 pfd_8_0.UP_input.t7 pfd_8_0.UP_input.n3 80.3338
R3071 pfd_8_0.UP_input.n5 pfd_8_0.UP_input.t4 80.3338
R3072 pfd_8_0.UP_input.t4 pfd_8_0.UP_input.n1 80.3338
R3073 charge_pump_cell_6_0.UP_b pfd_8_0.UP_b.n1 507.072
R3074 pfd_8_0.UP_b.n1 pfd_8_0.UP_b.n0 409.067
R3075 pfd_8_0.UP_b.n1 pfd_8_0.UP_b.t3 369.534
R3076 pfd_8_0.UP_b.n0 pfd_8_0.UP_b.t0 209.928
R3077 pfd_8_0.UP_b.n0 pfd_8_0.UP_b.t2 177.536
R3078 charge_pump_cell_6_0.UP_b pfd_8_0.UP_b.t1 24.0223
R3079 VCO_FD_magic_0.vco2_3_0.V1.n1 VCO_FD_magic_0.vco2_3_0.V1.t5 600.206
R3080 VCO_FD_magic_0.vco2_3_0.V1.t2 VCO_FD_magic_0.vco2_3_0.V1.n5 576.192
R3081 VCO_FD_magic_0.vco2_3_0.V1.n2 VCO_FD_magic_0.vco2_3_0.V1.n1 568.072
R3082 VCO_FD_magic_0.vco2_3_0.V1.n4 VCO_FD_magic_0.vco2_3_0.V1.n2 392.486
R3083 VCO_FD_magic_0.vco2_3_0.V1.n0 VCO_FD_magic_0.vco2_3_0.V1.t1 289.791
R3084 VCO_FD_magic_0.vco2_3_0.V1.n5 VCO_FD_magic_0.vco2_3_0.V1.n4 168.067
R3085 VCO_FD_magic_0.vco2_3_0.V1.n3 VCO_FD_magic_0.vco2_3_0.V1.n0 97.9242
R3086 VCO_FD_magic_0.vco2_3_0.V1.n4 VCO_FD_magic_0.vco2_3_0.V1.n3 37.7572
R3087 VCO_FD_magic_0.vco2_3_0.V1.n1 VCO_FD_magic_0.vco2_3_0.V1.t3 32.1338
R3088 VCO_FD_magic_0.vco2_3_0.V1.n2 VCO_FD_magic_0.vco2_3_0.V1.t4 32.1338
R3089 VCO_FD_magic_0.vco2_3_0.V1.n3 VCO_FD_magic_0.vco2_3_0.V1.t0 32.1338
R3090 VCO_FD_magic_0.vco2_3_0.V1.n5 VCO_FD_magic_0.vco2_3_0.V1.n0 28.3357
R3091 VCO_FD_magic_0.vco2_3_0.V4.n0 VCO_FD_magic_0.vco2_3_0.V4.t1 421.027
R3092 VCO_FD_magic_0.vco2_3_0.V4.n0 VCO_FD_magic_0.vco2_3_0.V4.t2 348.81
R3093 VCO_FD_magic_0.vco2_3_0.V4 VCO_FD_magic_0.vco2_3_0.V4.t0 280.05
R3094 VCO_FD_magic_0.vco2_3_0.V4 VCO_FD_magic_0.vco2_3_0.V4.n0 36.1094
R3095 VCO_FD_magic_0.div120_2_0.div5_2_0.G.n0 VCO_FD_magic_0.div120_2_0.div5_2_0.G.t1 685.134
R3096 VCO_FD_magic_0.div120_2_0.div5_2_0.G VCO_FD_magic_0.div120_2_0.div5_2_0.G.t2 663.801
R3097 VCO_FD_magic_0.div120_2_0.div5_2_0.G.n1 VCO_FD_magic_0.div120_2_0.div5_2_0.G.t3 534.268
R3098 VCO_FD_magic_0.div120_2_0.div5_2_0.G.n0 VCO_FD_magic_0.div120_2_0.div5_2_0.G.t0 340.521
R3099 VCO_FD_magic_0.div120_2_0.div5_2_0.G.n1 VCO_FD_magic_0.div120_2_0.div5_2_0.G.n0 105.6
R3100 VCO_FD_magic_0.div120_2_0.div5_2_0.G VCO_FD_magic_0.div120_2_0.div5_2_0.G.n1 21.3338
R3101 pfd_8_0.opamp_out.n6 pfd_8_0.opamp_out.n5 424.447
R3102 pfd_8_0.opamp_out.n6 pfd_8_0.opamp_out.n4 354.048
R3103 pfd_8_0.opamp_out.n2 pfd_8_0.opamp_out.n1 313
R3104 pfd_8_0.opamp_out.n9 pfd_8_0.opamp_out.t14 297.233
R3105 pfd_8_0.opamp_out.n10 pfd_8_0.opamp_out.t14 297.233
R3106 pfd_8_0.opamp_out.t13 pfd_8_0.opamp_out.n11 297.233
R3107 pfd_8_0.opamp_out.n13 pfd_8_0.opamp_out.t0 281.596
R3108 pfd_8_0.opamp_out.n2 pfd_8_0.opamp_out.n0 242.601
R3109 pfd_8_0.opamp_out.n3 pfd_8_0.opamp_out.n2 220.8
R3110 pfd_8_0.opamp_out.n7 pfd_8_0.opamp_out.n6 220.8
R3111 pfd_8_0.opamp_out.n11 pfd_8_0.opamp_out.n10 216.9
R3112 pfd_8_0.opamp_out.n9 pfd_8_0.opamp_out.n8 216.9
R3113 pfd_8_0.opamp_out.n14 pfd_8_0.opamp_out.n12 215.107
R3114 pfd_8_0.opamp_out.n12 pfd_8_0.opamp_out.n8 184.768
R3115 pfd_8_0.opamp_out.n13 pfd_8_0.opamp_out.t4 118.666
R3116 pfd_8_0.opamp_out.n10 pfd_8_0.opamp_out.t15 80.3338
R3117 pfd_8_0.opamp_out.t15 pfd_8_0.opamp_out.n9 80.3338
R3118 pfd_8_0.opamp_out.n11 pfd_8_0.opamp_out.t10 80.3338
R3119 pfd_8_0.opamp_out.t10 pfd_8_0.opamp_out.n8 80.3338
R3120 pfd_8_0.opamp_out.n12 pfd_8_0.opamp_out.t13 80.3338
R3121 pfd_8_0.opamp_out.n15 pfd_8_0.opamp_out.n14 78.9255
R3122 pfd_8_0.opamp_out.n3 pfd_8_0.opamp_out.t12 70.0829
R3123 pfd_8_0.opamp_out.n7 pfd_8_0.opamp_out.t11 63.6829
R3124 opamp_cell_4_0.VOUT pfd_8_0.opamp_out.n3 62.4005
R3125 pfd_8_0.opamp_out.n15 pfd_8_0.opamp_out.n7 60.8005
R3126 pfd_8_0.opamp_out.n14 pfd_8_0.opamp_out.n13 60.2361
R3127 pfd_8_0.opamp_out.n0 pfd_8_0.opamp_out.t3 60.0005
R3128 pfd_8_0.opamp_out.n0 pfd_8_0.opamp_out.t6 60.0005
R3129 pfd_8_0.opamp_out.n1 pfd_8_0.opamp_out.t8 60.0005
R3130 pfd_8_0.opamp_out.n1 pfd_8_0.opamp_out.t1 60.0005
R3131 pfd_8_0.opamp_out.n5 pfd_8_0.opamp_out.t9 49.2505
R3132 pfd_8_0.opamp_out.n5 pfd_8_0.opamp_out.t2 49.2505
R3133 pfd_8_0.opamp_out.n4 pfd_8_0.opamp_out.t5 49.2505
R3134 pfd_8_0.opamp_out.n4 pfd_8_0.opamp_out.t7 49.2505
R3135 opamp_cell_4_0.VOUT pfd_8_0.opamp_out.n15 1.6005
R3136 opamp_cell_4_0.VIN+.n1 opamp_cell_4_0.VIN+.t8 377.567
R3137 opamp_cell_4_0.VIN+.n0 opamp_cell_4_0.VIN+.t6 321.334
R3138 opamp_cell_4_0.VIN+.n2 opamp_cell_4_0.VIN+.n1 233.476
R3139 opamp_cell_4_0.VIN+.n1 opamp_cell_4_0.VIN+.t7 216.9
R3140 opamp_cell_4_0.VIN+.n5 opamp_cell_4_0.VIN+.n4 199.462
R3141 opamp_cell_4_0.VIN+.n2 opamp_cell_4_0.VIN+.n0 189.898
R3142 opamp_cell_4_0.VIN+.n5 opamp_cell_4_0.VIN+.n3 172.502
R3143 opamp_cell_4_0.VIN+.n7 opamp_cell_4_0.VIN+.n6 172.5
R3144 opamp_cell_4_0.VIN+.n0 opamp_cell_4_0.VIN+.t9 112.468
R3145 opamp_cell_4_0.VIN+.n7 opamp_cell_4_0.VIN+.n5 70.4005
R3146 opamp_cell_4_0.VIN+ opamp_cell_4_0.VIN+.n7 50.088
R3147 opamp_cell_4_0.VIN+.n3 opamp_cell_4_0.VIN+.t3 24.6255
R3148 opamp_cell_4_0.VIN+.n3 opamp_cell_4_0.VIN+.t2 24.6255
R3149 opamp_cell_4_0.VIN+.n6 opamp_cell_4_0.VIN+.t5 24.6255
R3150 opamp_cell_4_0.VIN+.n6 opamp_cell_4_0.VIN+.t4 24.6255
R3151 opamp_cell_4_0.VIN+.n4 opamp_cell_4_0.VIN+.t1 15.0005
R3152 opamp_cell_4_0.VIN+.n4 opamp_cell_4_0.VIN+.t0 15.0005
R3153 opamp_cell_4_0.VIN+ opamp_cell_4_0.VIN+.n2 3.313
R3154 a_6320_5840.n7 a_6320_5840.n5 482.582
R3155 a_6320_5840.n10 a_6320_5840.t4 304.634
R3156 a_6320_5840.n3 a_6320_5840.t2 304.634
R3157 a_6320_5840.t6 a_6320_5840.n10 277.914
R3158 a_6320_5840.n3 a_6320_5840.t3 276.289
R3159 a_6320_5840.n8 a_6320_5840.n1 204.201
R3160 a_6320_5840.n4 a_6320_5840.n2 204.201
R3161 a_6320_5840.n9 a_6320_5840.n0 204.201
R3162 a_6320_5840.n7 a_6320_5840.n6 120.981
R3163 a_6320_5840.n8 a_6320_5840.n4 74.6672
R3164 a_6320_5840.n9 a_6320_5840.n8 74.6672
R3165 a_6320_5840.n1 a_6320_5840.t0 60.0005
R3166 a_6320_5840.n1 a_6320_5840.t10 60.0005
R3167 a_6320_5840.t3 a_6320_5840.n2 60.0005
R3168 a_6320_5840.n2 a_6320_5840.t1 60.0005
R3169 a_6320_5840.n0 a_6320_5840.t9 60.0005
R3170 a_6320_5840.n0 a_6320_5840.t5 60.0005
R3171 a_6320_5840.n8 a_6320_5840.n7 37.763
R3172 a_6320_5840.n5 a_6320_5840.t7 24.0005
R3173 a_6320_5840.n5 a_6320_5840.t11 24.0005
R3174 a_6320_5840.n6 a_6320_5840.t12 24.0005
R3175 a_6320_5840.n6 a_6320_5840.t8 24.0005
R3176 a_6320_5840.n4 a_6320_5840.n3 16.0005
R3177 a_6320_5840.n10 a_6320_5840.n9 16.0005
R3178 opamp_cell_4_0.n_right.t4 opamp_cell_4_0.n_right.n6 1010.36
R3179 opamp_cell_4_0.n_right.n3 opamp_cell_4_0.n_right.n2 404.8
R3180 opamp_cell_4_0.n_right.n2 opamp_cell_4_0.n_right.n1 322.048
R3181 opamp_cell_4_0.n_right.n2 opamp_cell_4_0.n_right.n0 316.2
R3182 opamp_cell_4_0.n_right.n4 opamp_cell_4_0.n_right.t8 289.2
R3183 opamp_cell_4_0.n_right.n5 opamp_cell_4_0.n_right.t7 289.2
R3184 opamp_cell_4_0.n_right.n6 opamp_cell_4_0.n_right.t6 289.2
R3185 opamp_cell_4_0.n_right.n3 opamp_cell_4_0.n_right.t5 232.968
R3186 opamp_cell_4_0.n_right.n6 opamp_cell_4_0.n_right.n5 208.868
R3187 opamp_cell_4_0.n_right.n5 opamp_cell_4_0.n_right.n4 208.868
R3188 opamp_cell_4_0.n_right.n4 opamp_cell_4_0.n_right.n3 199.829
R3189 opamp_cell_4_0.n_right.n0 opamp_cell_4_0.n_right.t0 60.0005
R3190 opamp_cell_4_0.n_right.n0 opamp_cell_4_0.n_right.t1 60.0005
R3191 opamp_cell_4_0.n_right.n1 opamp_cell_4_0.n_right.t3 49.2505
R3192 opamp_cell_4_0.n_right.n1 opamp_cell_4_0.n_right.t2 49.2505
R3193 opamp_cell_4_0.n_left.n1 opamp_cell_4_0.n_left.t7 359.894
R3194 opamp_cell_4_0.n_left.n5 opamp_cell_4_0.n_left.n4 325.248
R3195 opamp_cell_4_0.n_left.n4 opamp_cell_4_0.n_left.n0 313
R3196 opamp_cell_4_0.n_left.n3 opamp_cell_4_0.n_left.t0 252.248
R3197 opamp_cell_4_0.n_left.n2 opamp_cell_4_0.n_left.n1 208.868
R3198 opamp_cell_4_0.n_left.n2 opamp_cell_4_0.n_left.t2 192.8
R3199 opamp_cell_4_0.n_left.n1 opamp_cell_4_0.n_left.t6 192.8
R3200 opamp_cell_4_0.n_left.n4 opamp_cell_4_0.n_left.n3 152
R3201 opamp_cell_4_0.n_left.n0 opamp_cell_4_0.n_left.t5 60.0005
R3202 opamp_cell_4_0.n_left.n0 opamp_cell_4_0.n_left.t4 60.0005
R3203 opamp_cell_4_0.n_left.n3 opamp_cell_4_0.n_left.n2 59.4472
R3204 opamp_cell_4_0.n_left.t3 opamp_cell_4_0.n_left.n5 49.2505
R3205 opamp_cell_4_0.n_left.n5 opamp_cell_4_0.n_left.t1 49.2505
R3206 VCO_FD_magic_0.div120_2_0.div2_4_0.C VCO_FD_magic_0.div120_2_0.div2_4_0.C.t3 702.201
R3207 VCO_FD_magic_0.div120_2_0.div2_4_0.C.n1 VCO_FD_magic_0.div120_2_0.div2_4_0.C.t4 349.433
R3208 VCO_FD_magic_0.div120_2_0.div2_4_0.C.n2 VCO_FD_magic_0.div120_2_0.div2_4_0.C.t2 276.733
R3209 VCO_FD_magic_0.div120_2_0.div2_4_0.C.n1 VCO_FD_magic_0.div120_2_0.div2_4_0.C.n0 206.333
R3210 VCO_FD_magic_0.div120_2_0.div2_4_0.C VCO_FD_magic_0.div120_2_0.div2_4_0.C.n2 48.0005
R3211 VCO_FD_magic_0.div120_2_0.div2_4_0.C.n2 VCO_FD_magic_0.div120_2_0.div2_4_0.C.n1 48.0005
R3212 VCO_FD_magic_0.div120_2_0.div2_4_0.C.n0 VCO_FD_magic_0.div120_2_0.div2_4_0.C.t0 48.0005
R3213 VCO_FD_magic_0.div120_2_0.div2_4_0.C.n0 VCO_FD_magic_0.div120_2_0.div2_4_0.C.t1 48.0005
R3214 VCO_FD_magic_0.div120_2_0.div8.t4 VCO_FD_magic_0.div120_2_0.div8.t5 1012.2
R3215 VCO_FD_magic_0.div120_2_0.div8.n0 VCO_FD_magic_0.div120_2_0.div8.t0 663.801
R3216 VCO_FD_magic_0.div120_2_0.div8.n2 VCO_FD_magic_0.div120_2_0.div8.n1 431.401
R3217 VCO_FD_magic_0.div120_2_0.div8.t3 VCO_FD_magic_0.div120_2_0.div8.t6 401.668
R3218 VCO_FD_magic_0.div120_2_0.div8.n0 VCO_FD_magic_0.div120_2_0.div8.t4 361.692
R3219 VCO_FD_magic_0.div120_2_0.div8.t1 VCO_FD_magic_0.div120_2_0.div8.n2 298.921
R3220 VCO_FD_magic_0.div120_2_0.div8.n1 VCO_FD_magic_0.div120_2_0.div8.t3 257.067
R3221 VCO_FD_magic_0.div120_2_0.div8.n1 VCO_FD_magic_0.div120_2_0.div8.t2 208.868
R3222 VCO_FD_magic_0.div120_2_0.div8.n2 VCO_FD_magic_0.div120_2_0.div8.n0 67.2005
R3223 a_6490_4630.t4 a_6490_4630.n6 1112.76
R3224 a_6490_4630.n3 a_6490_4630.n2 441.433
R3225 a_6490_4630.n2 a_6490_4630.n1 379.647
R3226 a_6490_4630.n2 a_6490_4630.n0 258.601
R3227 a_6490_4630.n6 a_6490_4630.t6 208.868
R3228 a_6490_4630.n5 a_6490_4630.t7 208.868
R3229 a_6490_4630.n4 a_6490_4630.t8 208.868
R3230 a_6490_4630.n3 a_6490_4630.t5 208.868
R3231 a_6490_4630.n6 a_6490_4630.n5 208.868
R3232 a_6490_4630.n5 a_6490_4630.n4 208.868
R3233 a_6490_4630.n4 a_6490_4630.n3 208.868
R3234 a_6490_4630.n0 a_6490_4630.t3 60.0005
R3235 a_6490_4630.n0 a_6490_4630.t2 60.0005
R3236 a_6490_4630.n1 a_6490_4630.t1 49.2505
R3237 a_6490_4630.n1 a_6490_4630.t0 49.2505
R3238 pfd_8_0.before_Reset.n1 pfd_8_0.before_Reset.n0 481.334
R3239 pfd_8_0.before_Reset.n0 pfd_8_0.before_Reset.t4 465.933
R3240 pfd_8_0.before_Reset.n0 pfd_8_0.before_Reset.t3 321.334
R3241 pfd_8_0.before_Reset.n2 pfd_8_0.before_Reset.n1 226.889
R3242 pfd_8_0.before_Reset.n1 pfd_8_0.before_Reset.t1 172.458
R3243 pfd_8_0.before_Reset.n2 pfd_8_0.before_Reset.t2 19.7005
R3244 pfd_8_0.before_Reset.t0 pfd_8_0.before_Reset.n2 19.7005
R3245 a_2350_1400.t1 a_2350_1400.n2 500.086
R3246 a_2350_1400.n1 a_2350_1400.n0 473.334
R3247 a_2350_1400.n0 a_2350_1400.t3 465.933
R3248 a_2350_1400.t1 a_2350_1400.n2 461.389
R3249 a_2350_1400.n0 a_2350_1400.t2 321.334
R3250 a_2350_1400.n1 a_2350_1400.t0 177.577
R3251 a_2350_1400.n2 a_2350_1400.n1 48.3899
R3252 VCO_FD_magic_0.div120_2_0.div2_4_2.A.n0 VCO_FD_magic_0.div120_2_0.div2_4_2.A.t1 713.933
R3253 VCO_FD_magic_0.div120_2_0.div2_4_2.A VCO_FD_magic_0.div120_2_0.div2_4_2.A.t0 327.401
R3254 VCO_FD_magic_0.div120_2_0.div2_4_2.A.n0 VCO_FD_magic_0.div120_2_0.div2_4_2.A.t2 314.233
R3255 VCO_FD_magic_0.div120_2_0.div2_4_2.A VCO_FD_magic_0.div120_2_0.div2_4_2.A.n0 9.6005
R3256 VCO_FD_magic_0.div120_2_0.div2_4_2.B.t0 VCO_FD_magic_0.div120_2_0.div2_4_2.B.t1 96.0005
R3257 opamp_cell_4_0.p_bias opamp_cell_4_0.p_bias.t0 918.318
R3258 opamp_cell_4_0.p_bias opamp_cell_4_0.p_bias.n11 540.801
R3259 opamp_cell_4_0.p_bias.n8 opamp_cell_4_0.p_bias.t10 377.567
R3260 opamp_cell_4_0.p_bias.n3 opamp_cell_4_0.p_bias.t9 377.567
R3261 opamp_cell_4_0.p_bias.n9 opamp_cell_4_0.p_bias.n8 257.067
R3262 opamp_cell_4_0.p_bias.n7 opamp_cell_4_0.p_bias.n6 257.067
R3263 opamp_cell_4_0.p_bias.n4 opamp_cell_4_0.p_bias.n3 257.067
R3264 opamp_cell_4_0.p_bias.n11 opamp_cell_4_0.p_bias.n0 154.321
R3265 opamp_cell_4_0.p_bias.n2 opamp_cell_4_0.p_bias.n1 154.321
R3266 opamp_cell_4_0.p_bias.n5 opamp_cell_4_0.p_bias.n2 152
R3267 opamp_cell_4_0.p_bias.n11 opamp_cell_4_0.p_bias.n10 152
R3268 opamp_cell_4_0.p_bias.n8 opamp_cell_4_0.p_bias.t12 120.501
R3269 opamp_cell_4_0.p_bias.n9 opamp_cell_4_0.p_bias.t5 120.501
R3270 opamp_cell_4_0.p_bias.n7 opamp_cell_4_0.p_bias.t1 120.501
R3271 opamp_cell_4_0.p_bias.n6 opamp_cell_4_0.p_bias.t3 120.501
R3272 opamp_cell_4_0.p_bias.n3 opamp_cell_4_0.p_bias.t11 120.501
R3273 opamp_cell_4_0.p_bias.n4 opamp_cell_4_0.p_bias.t7 120.501
R3274 opamp_cell_4_0.p_bias.n11 opamp_cell_4_0.p_bias.n2 115.201
R3275 opamp_cell_4_0.p_bias.n10 opamp_cell_4_0.p_bias.n9 85.6894
R3276 opamp_cell_4_0.p_bias.n10 opamp_cell_4_0.p_bias.n7 85.6894
R3277 opamp_cell_4_0.p_bias.n6 opamp_cell_4_0.p_bias.n5 85.6894
R3278 opamp_cell_4_0.p_bias.n5 opamp_cell_4_0.p_bias.n4 85.6894
R3279 opamp_cell_4_0.p_bias.n0 opamp_cell_4_0.p_bias.t2 19.7005
R3280 opamp_cell_4_0.p_bias.n0 opamp_cell_4_0.p_bias.t6 19.7005
R3281 opamp_cell_4_0.p_bias.n1 opamp_cell_4_0.p_bias.t8 19.7005
R3282 opamp_cell_4_0.p_bias.n1 opamp_cell_4_0.p_bias.t4 19.7005
R3283 F_REF.n0 F_REF.t0 514.134
R3284 F_REF.n0 F_REF.t1 273.134
R3285 F_REF F_REF.n0 216.9
R3286 a_n30_1400.t0 a_n30_1400.t1 39.4005
R3287 I_IN.n1 I_IN.n0 1269.42
R3288 I_IN.n1 I_IN.t1 275.325
R3289 I_IN.n6 I_IN.n2 248.4
R3290 I_IN.n4 I_IN.t5 238.892
R3291 I_IN.n4 I_IN.t0 161.371
R3292 I_IN.n0 I_IN.t6 151.792
R3293 I_IN.n5 I_IN.n4 151.34
R3294 I_IN.n2 I_IN.t3 140.583
R3295 I_IN.n2 I_IN.t1 140.583
R3296 I_IN.n6 I_IN.n3 98.6614
R3297 I_IN.t3 I_IN.n1 80.3338
R3298 I_IN.n0 I_IN.t7 44.2902
R3299 I_IN.n3 I_IN.t4 15.0005
R3300 I_IN.n3 I_IN.t2 15.0005
R3301 I_IN.n6 I_IN.n5 9.3005
R3302 I_IN I_IN.n6 3.2005
R3303 I_IN.n5 I_IN 0.063
R3304 VCO_FD_magic_0.div120_2_0.div4.t6 VCO_FD_magic_0.div120_2_0.div4.t3 1012.2
R3305 VCO_FD_magic_0.div120_2_0.div4.n0 VCO_FD_magic_0.div120_2_0.div4.t0 663.801
R3306 VCO_FD_magic_0.div120_2_0.div4.n2 VCO_FD_magic_0.div120_2_0.div4.n1 431.401
R3307 VCO_FD_magic_0.div120_2_0.div4.t4 VCO_FD_magic_0.div120_2_0.div4.t2 401.668
R3308 VCO_FD_magic_0.div120_2_0.div4.n0 VCO_FD_magic_0.div120_2_0.div4.t6 361.692
R3309 VCO_FD_magic_0.div120_2_0.div4.n1 VCO_FD_magic_0.div120_2_0.div4.t5 353.467
R3310 VCO_FD_magic_0.div120_2_0.div4.t1 VCO_FD_magic_0.div120_2_0.div4.n2 298.921
R3311 VCO_FD_magic_0.div120_2_0.div4.n1 VCO_FD_magic_0.div120_2_0.div4.t4 257.067
R3312 VCO_FD_magic_0.div120_2_0.div4.n2 VCO_FD_magic_0.div120_2_0.div4.n0 67.2005
R3313 a_6330_n1440.n0 a_6330_n1440.t1 752.333
R3314 a_6330_n1440.t2 a_6330_n1440.n5 752.333
R3315 a_6330_n1440.n1 a_6330_n1440.t6 514.134
R3316 a_6330_n1440.n4 a_6330_n1440.n3 366.856
R3317 a_6330_n1440.n0 a_6330_n1440.t0 254.333
R3318 a_6330_n1440.n4 a_6330_n1440.t5 190.123
R3319 a_6330_n1440.n5 a_6330_n1440.n4 187.201
R3320 a_6330_n1440.n3 a_6330_n1440.n2 176.733
R3321 a_6330_n1440.n2 a_6330_n1440.n1 176.733
R3322 a_6330_n1440.n3 a_6330_n1440.t3 112.468
R3323 a_6330_n1440.n2 a_6330_n1440.t7 112.468
R3324 a_6330_n1440.n1 a_6330_n1440.t4 112.468
R3325 a_6330_n1440.n5 a_6330_n1440.n0 70.4005
R3326 pfd_8_0.QA.t5 pfd_8_0.QA.t7 835.467
R3327 pfd_8_0.QA.n2 pfd_8_0.QA.t4 517.347
R3328 pfd_8_0.QA.n0 pfd_8_0.QA.t8 465.933
R3329 pfd_8_0.QA.n1 pfd_8_0.QA.n0 454.031
R3330 pfd_8_0.QA.n1 pfd_8_0.QA.t5 394.267
R3331 pfd_8_0.QA.n0 pfd_8_0.QA.t6 321.334
R3332 pfd_8_0.QA.n4 pfd_8_0.QA.n3 244.715
R3333 pfd_8_0.QA.n2 pfd_8_0.QA.t3 228.148
R3334 pfd_8_0.QA.n4 pfd_8_0.QA.t1 221.411
R3335 pfd_8_0.QA.n5 pfd_8_0.QA.n2 216
R3336 pfd_8_0.QA.n5 pfd_8_0.QA.n4 201.573
R3337 pfd_8_0.QA pfd_8_0.QA.n5 60.8005
R3338 pfd_8_0.QA pfd_8_0.QA.n1 56.1505
R3339 pfd_8_0.QA.n3 pfd_8_0.QA.t0 24.0005
R3340 pfd_8_0.QA.n3 pfd_8_0.QA.t2 24.0005
R3341 loop_filter_3_0.R1_C1.t0 loop_filter_3_0.R1_C1.t1 167.486
R3342 a_8930_n1440.n5 a_8930_n1440.t0 752.333
R3343 a_8930_n1440.n4 a_8930_n1440.t2 752.333
R3344 a_8930_n1440.n0 a_8930_n1440.t4 514.134
R3345 a_8930_n1440.n3 a_8930_n1440.n2 366.856
R3346 a_8930_n1440.t1 a_8930_n1440.n5 254.333
R3347 a_8930_n1440.n3 a_8930_n1440.t5 190.123
R3348 a_8930_n1440.n4 a_8930_n1440.n3 187.201
R3349 a_8930_n1440.n2 a_8930_n1440.n1 176.733
R3350 a_8930_n1440.n1 a_8930_n1440.n0 176.733
R3351 a_8930_n1440.n2 a_8930_n1440.t3 112.468
R3352 a_8930_n1440.n1 a_8930_n1440.t6 112.468
R3353 a_8930_n1440.n0 a_8930_n1440.t7 112.468
R3354 a_8930_n1440.n5 a_8930_n1440.n4 70.4005
R3355 VCO_FD_magic_0.div120_2_0.div2_4_1.C VCO_FD_magic_0.div120_2_0.div2_4_1.C.t3 702.201
R3356 VCO_FD_magic_0.div120_2_0.div2_4_1.C.n1 VCO_FD_magic_0.div120_2_0.div2_4_1.C.t4 349.433
R3357 VCO_FD_magic_0.div120_2_0.div2_4_1.C.n2 VCO_FD_magic_0.div120_2_0.div2_4_1.C.t2 276.733
R3358 VCO_FD_magic_0.div120_2_0.div2_4_1.C.n1 VCO_FD_magic_0.div120_2_0.div2_4_1.C.n0 206.333
R3359 VCO_FD_magic_0.div120_2_0.div2_4_1.C.n0 VCO_FD_magic_0.div120_2_0.div2_4_1.C.t1 48.0005
R3360 VCO_FD_magic_0.div120_2_0.div2_4_1.C.n0 VCO_FD_magic_0.div120_2_0.div2_4_1.C.t0 48.0005
R3361 VCO_FD_magic_0.div120_2_0.div2_4_1.C VCO_FD_magic_0.div120_2_0.div2_4_1.C.n2 48.0005
R3362 VCO_FD_magic_0.div120_2_0.div2_4_1.C.n2 VCO_FD_magic_0.div120_2_0.div2_4_1.C.n1 48.0005
R3363 pfd_8_0.DOWN_input.t5 pfd_8_0.DOWN_input.t4 377.567
R3364 pfd_8_0.DOWN_input.n2 pfd_8_0.DOWN_input.t3 326.658
R3365 pfd_8_0.DOWN_input pfd_8_0.DOWN_input.n3 237.65
R3366 pfd_8_0.DOWN_input.n0 pfd_8_0.DOWN_input.t0 229.127
R3367 pfd_8_0.DOWN_input.n3 pfd_8_0.DOWN_input.n2 196.817
R3368 pfd_8_0.DOWN_input.n0 pfd_8_0.DOWN_input.t2 158.335
R3369 pfd_8_0.DOWN_input.n1 pfd_8_0.DOWN_input.t1 158.335
R3370 pfd_8_0.DOWN_input.n1 pfd_8_0.DOWN_input.n0 121.6
R3371 pfd_8_0.DOWN_input.t4 pfd_8_0.DOWN_input.n2 92.3838
R3372 pfd_8_0.DOWN_input.n3 pfd_8_0.DOWN_input.t5 92.3838
R3373 pfd_8_0.DOWN_input pfd_8_0.DOWN_input.n1 3.2005
R3374 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.n3 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.n2 742.51
R3375 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.n8 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.t1 723.534
R3376 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.t2 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.n9 723.534
R3377 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.n2 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.n1 684.806
R3378 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.n7 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.n6 366.856
R3379 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.n0 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.t6 337.401
R3380 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.n0 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.t9 305.267
R3381 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.n9 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.t0 254.333
R3382 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.n4 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.n3 224.934
R3383 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.n7 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.t11 190.123
R3384 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.n8 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.n7 187.201
R3385 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.n1 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.n0 176.733
R3386 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.n6 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.n5 176.733
R3387 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.n5 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.n4 176.733
R3388 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.n3 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.t3 144.601
R3389 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.n2 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.t8 131.976
R3390 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.n1 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.t12 128.534
R3391 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.n0 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.t5 128.534
R3392 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.n6 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.t7 112.468
R3393 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.n5 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.t10 112.468
R3394 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.n4 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.t4 112.468
R3395 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.n9 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.n8 70.4005
R3396 VCO_FD_magic_0.div120_2_0.div3_3_0.D.n1 VCO_FD_magic_0.div120_2_0.div3_3_0.D.n0 701.467
R3397 VCO_FD_magic_0.div120_2_0.div3_3_0.D.n1 VCO_FD_magic_0.div120_2_0.div3_3_0.D.t0 694.201
R3398 VCO_FD_magic_0.div120_2_0.div3_3_0.D.n0 VCO_FD_magic_0.div120_2_0.div3_3_0.D.t2 321.334
R3399 VCO_FD_magic_0.div120_2_0.div3_3_0.D VCO_FD_magic_0.div120_2_0.div3_3_0.D.t1 260.521
R3400 VCO_FD_magic_0.div120_2_0.div3_3_0.D.n0 VCO_FD_magic_0.div120_2_0.div3_3_0.D.t3 144.601
R3401 VCO_FD_magic_0.div120_2_0.div3_3_0.D VCO_FD_magic_0.div120_2_0.div3_3_0.D.n1 54.4005
R3402 VCO_FD_magic_0.div120_2_0.div3_3_0.C VCO_FD_magic_0.div120_2_0.div3_3_0.C.t3 702.201
R3403 VCO_FD_magic_0.div120_2_0.div3_3_0.C.n1 VCO_FD_magic_0.div120_2_0.div3_3_0.C.t4 350.349
R3404 VCO_FD_magic_0.div120_2_0.div3_3_0.C.n2 VCO_FD_magic_0.div120_2_0.div3_3_0.C.t1 276.733
R3405 VCO_FD_magic_0.div120_2_0.div3_3_0.C.n1 VCO_FD_magic_0.div120_2_0.div3_3_0.C.n0 206.333
R3406 VCO_FD_magic_0.div120_2_0.div3_3_0.C.n2 VCO_FD_magic_0.div120_2_0.div3_3_0.C.n1 48.0005
R3407 VCO_FD_magic_0.div120_2_0.div3_3_0.C.n0 VCO_FD_magic_0.div120_2_0.div3_3_0.C.t0 48.0005
R3408 VCO_FD_magic_0.div120_2_0.div3_3_0.C.n0 VCO_FD_magic_0.div120_2_0.div3_3_0.C.t2 48.0005
R3409 VCO_FD_magic_0.div120_2_0.div3_3_0.C VCO_FD_magic_0.div120_2_0.div3_3_0.C.n2 19.2005
R3410 pfd_8_0.QB.t4 pfd_8_0.QB.t3 835.467
R3411 pfd_8_0.QB.n1 pfd_8_0.QB.t4 564.496
R3412 pfd_8_0.QB.n2 pfd_8_0.QB.t5 517.347
R3413 pfd_8_0.QB.n0 pfd_8_0.QB.t7 514.134
R3414 pfd_8_0.QB.n1 pfd_8_0.QB.n0 455.219
R3415 pfd_8_0.QB.n5 pfd_8_0.QB.n2 363.2
R3416 pfd_8_0.QB.n0 pfd_8_0.QB.t8 273.134
R3417 pfd_8_0.QB.n4 pfd_8_0.QB.n3 244.716
R3418 pfd_8_0.QB.n2 pfd_8_0.QB.t6 228.148
R3419 pfd_8_0.QB.n4 pfd_8_0.QB.t0 221.411
R3420 pfd_8_0.QB.n5 pfd_8_0.QB.n4 54.3734
R3421 pfd_8_0.QB pfd_8_0.QB.n1 26.7568
R3422 pfd_8_0.QB.n3 pfd_8_0.QB.t1 24.0005
R3423 pfd_8_0.QB.n3 pfd_8_0.QB.t2 24.0005
R3424 pfd_8_0.QB pfd_8_0.QB.n5 6.4005
R3425 a_1910_2020.t0 a_1910_2020.t1 48.0005
R3426 a_6220_5810.n4 a_6220_5810.t12 317.317
R3427 a_6220_5810.n2 a_6220_5810.t11 317.317
R3428 a_6220_5810.n5 a_6220_5810.n4 257.067
R3429 a_6220_5810.n3 a_6220_5810.n2 257.067
R3430 a_6220_5810.n10 a_6220_5810.n9 257.067
R3431 a_6220_5810.t0 a_6220_5810.n12 194.478
R3432 a_6220_5810.n8 a_6220_5810.n7 152
R3433 a_6220_5810.n12 a_6220_5810.n11 152
R3434 a_6220_5810.n1 a_6220_5810.n0 120.981
R3435 a_6220_5810.n7 a_6220_5810.n6 117.781
R3436 a_6220_5810.n7 a_6220_5810.n1 108.8
R3437 a_6220_5810.n8 a_6220_5810.n5 85.6894
R3438 a_6220_5810.n11 a_6220_5810.n3 85.6894
R3439 a_6220_5810.n11 a_6220_5810.n10 85.6894
R3440 a_6220_5810.n9 a_6220_5810.n8 85.6894
R3441 a_6220_5810.n4 a_6220_5810.t10 60.2505
R3442 a_6220_5810.n5 a_6220_5810.t1 60.2505
R3443 a_6220_5810.n2 a_6220_5810.t9 60.2505
R3444 a_6220_5810.n3 a_6220_5810.t3 60.2505
R3445 a_6220_5810.n10 a_6220_5810.t7 60.2505
R3446 a_6220_5810.n9 a_6220_5810.t5 60.2505
R3447 a_6220_5810.n6 a_6220_5810.t6 24.0005
R3448 a_6220_5810.n6 a_6220_5810.t2 24.0005
R3449 a_6220_5810.n0 a_6220_5810.t4 24.0005
R3450 a_6220_5810.n0 a_6220_5810.t8 24.0005
R3451 a_6220_5810.n12 a_6220_5810.n1 3.2005
R3452 VCO_FD_magic_0.div120_2_0.div2_4_2.C VCO_FD_magic_0.div120_2_0.div2_4_2.C.t3 702.201
R3453 VCO_FD_magic_0.div120_2_0.div2_4_2.C.n1 VCO_FD_magic_0.div120_2_0.div2_4_2.C.t4 349.433
R3454 VCO_FD_magic_0.div120_2_0.div2_4_2.C.n2 VCO_FD_magic_0.div120_2_0.div2_4_2.C.t1 276.733
R3455 VCO_FD_magic_0.div120_2_0.div2_4_2.C.n1 VCO_FD_magic_0.div120_2_0.div2_4_2.C.n0 206.333
R3456 VCO_FD_magic_0.div120_2_0.div2_4_2.C VCO_FD_magic_0.div120_2_0.div2_4_2.C.n2 48.0005
R3457 VCO_FD_magic_0.div120_2_0.div2_4_2.C.n2 VCO_FD_magic_0.div120_2_0.div2_4_2.C.n1 48.0005
R3458 VCO_FD_magic_0.div120_2_0.div2_4_2.C.n0 VCO_FD_magic_0.div120_2_0.div2_4_2.C.t2 48.0005
R3459 VCO_FD_magic_0.div120_2_0.div2_4_2.C.n0 VCO_FD_magic_0.div120_2_0.div2_4_2.C.t0 48.0005
R3460 pfd_8_0.UP_PFD_b.n0 pfd_8_0.UP_PFD_b.t2 441.834
R3461 pfd_8_0.UP_PFD_b.n0 pfd_8_0.UP_PFD_b.t3 313.3
R3462 pfd_8_0.UP_PFD_b.n1 pfd_8_0.UP_PFD_b.n0 235.201
R3463 pfd_8_0.UP_PFD_b.t1 pfd_8_0.UP_PFD_b.n1 219.528
R3464 pfd_8_0.UP_PFD_b.n1 pfd_8_0.UP_PFD_b.t0 167.935
R3465 pfd_8_0.UP.n0 pfd_8_0.UP.t5 1205
R3466 pfd_8_0.UP.n2 pfd_8_0.UP.t4 522.168
R3467 pfd_8_0.UP.n1 pfd_8_0.UP.n0 441.834
R3468 pfd_8_0.UP.n3 pfd_8_0.UP.n2 235.201
R3469 pfd_8_0.UP.t1 pfd_8_0.UP.n3 229.127
R3470 pfd_8_0.UP.n1 pfd_8_0.UP.t3 217.905
R3471 pfd_8_0.UP.n0 pfd_8_0.UP.t2 208.868
R3472 pfd_8_0.UP.n3 pfd_8_0.UP.t0 158.335
R3473 pfd_8_0.UP.n2 pfd_8_0.UP.n1 15.063
R3474 F_VCO.n3 F_VCO.t3 772.196
R3475 F_VCO.n5 F_VCO.t0 751.801
R3476 F_VCO.n4 F_VCO.n3 607.465
R3477 F_VCO.t3 F_VCO.t2 514.134
R3478 F_VCO.n0 F_VCO.t6 514.134
R3479 F_VCO.n2 F_VCO.t4 289.2
R3480 F_VCO.n0 F_VCO.t7 273.134
R3481 F_VCO.n4 F_VCO.t1 233
R3482 F_VCO F_VCO.n0 216.9
R3483 F_VCO.n3 F_VCO.n2 208.868
R3484 F_VCO F_VCO.n1 194.333
R3485 F_VCO.n2 F_VCO.t5 176.733
R3486 F_VCO.n5 F_VCO.n4 40.3205
R3487 F_VCO F_VCO.n5 38.4005
R3488 F_VCO.n1 F_VCO 24.1005
R3489 F_VCO.n1 F_VCO 24.1005
R3490 VCO_FD_magic_0.div120_2_0.div5_2_0.I VCO_FD_magic_0.div120_2_0.div5_2_0.I.n0 279.933
R3491 VCO_FD_magic_0.div120_2_0.div5_2_0.I VCO_FD_magic_0.div120_2_0.div5_2_0.I.t2 251.133
R3492 VCO_FD_magic_0.div120_2_0.div5_2_0.I.n0 VCO_FD_magic_0.div120_2_0.div5_2_0.I.t1 48.0005
R3493 VCO_FD_magic_0.div120_2_0.div5_2_0.I.n0 VCO_FD_magic_0.div120_2_0.div5_2_0.I.t0 48.0005
R3494 VCO_FD_magic_0.div120_2_0.div5_2_0.H.t0 VCO_FD_magic_0.div120_2_0.div5_2_0.H.t1 96.0005
R3495 V_OSC.t2 V_OSC.t5 401.668
R3496 V_OSC.n1 V_OSC.t0 372.118
R3497 V_OSC.n3 V_OSC.t3 353.467
R3498 V_OSC V_OSC.n3 313.3
R3499 V_OSC.n3 V_OSC.t2 257.067
R3500 V_OSC.n1 V_OSC.t1 247.934
R3501 V_OSC.n2 V_OSC.n1 236.756
R3502 V_OSC.n0 V_OSC.t6 224.934
R3503 V_OSC.n2 V_OSC.n0 224.934
R3504 V_OSC.n0 V_OSC.t4 144.601
R3505 V_OSC V_OSC.n2 120.501
R3506 VCO_FD_magic_0.div120_2_0.div5_2_0.A.n2 VCO_FD_magic_0.div120_2_0.div5_2_0.A.t1 755.534
R3507 VCO_FD_magic_0.div120_2_0.div5_2_0.A.t2 VCO_FD_magic_0.div120_2_0.div5_2_0.A.n2 685.134
R3508 VCO_FD_magic_0.div120_2_0.div5_2_0.A.n1 VCO_FD_magic_0.div120_2_0.div5_2_0.A.n0 389.733
R3509 VCO_FD_magic_0.div120_2_0.div5_2_0.A.n1 VCO_FD_magic_0.div120_2_0.div5_2_0.A.t0 340.2
R3510 VCO_FD_magic_0.div120_2_0.div5_2_0.A.n0 VCO_FD_magic_0.div120_2_0.div5_2_0.A.t3 321.334
R3511 VCO_FD_magic_0.div120_2_0.div5_2_0.A.n0 VCO_FD_magic_0.div120_2_0.div5_2_0.A.t4 144.601
R3512 VCO_FD_magic_0.div120_2_0.div5_2_0.A.n2 VCO_FD_magic_0.div120_2_0.div5_2_0.A.n1 19.2005
R3513 VCO_FD_magic_0.div120_2_0.div5_2_0.C.t0 VCO_FD_magic_0.div120_2_0.div5_2_0.C.t1 96.0005
R3514 pfd_8_0.E.n4 pfd_8_0.E.n0 1319.38
R3515 pfd_8_0.E.n0 pfd_8_0.E.t3 562.333
R3516 pfd_8_0.E.n2 pfd_8_0.E.t5 388.813
R3517 pfd_8_0.E.n2 pfd_8_0.E.t4 356.68
R3518 pfd_8_0.E.n3 pfd_8_0.E.n2 232
R3519 pfd_8_0.E.n0 pfd_8_0.E.t6 224.934
R3520 pfd_8_0.E.t1 pfd_8_0.E.n4 221.411
R3521 pfd_8_0.E.n3 pfd_8_0.E.n1 157.278
R3522 pfd_8_0.E.n4 pfd_8_0.E.n3 90.64
R3523 pfd_8_0.E.n1 pfd_8_0.E.t0 24.0005
R3524 pfd_8_0.E.n1 pfd_8_0.E.t2 24.0005
R3525 pfd_8_0.E_b.n0 pfd_8_0.E_b.t4 517.347
R3526 pfd_8_0.E_b.n2 pfd_8_0.E_b.n0 417.574
R3527 pfd_8_0.E_b.n2 pfd_8_0.E_b.n1 244.716
R3528 pfd_8_0.E_b.n0 pfd_8_0.E_b.t3 228.148
R3529 pfd_8_0.E_b.t2 pfd_8_0.E_b.n2 221.411
R3530 pfd_8_0.E_b.n1 pfd_8_0.E_b.t0 24.0005
R3531 pfd_8_0.E_b.n1 pfd_8_0.E_b.t1 24.0005
R3532 a_1390_1400.t0 a_1390_1400.t1 39.4005
R3533 pfd_8_0.QB_b.t6 pfd_8_0.QB_b.t4 1188.93
R3534 pfd_8_0.QB_b pfd_8_0.QB_b.n2 899.734
R3535 pfd_8_0.QB_b.t4 pfd_8_0.QB_b.t3 835.467
R3536 pfd_8_0.QB_b.n2 pfd_8_0.QB_b.t5 562.333
R3537 pfd_8_0.QB_b pfd_8_0.QB_b.n1 419.647
R3538 pfd_8_0.QB_b.n1 pfd_8_0.QB_b.n0 247.917
R3539 pfd_8_0.QB_b.n2 pfd_8_0.QB_b.t6 224.934
R3540 pfd_8_0.QB_b.n1 pfd_8_0.QB_b.t1 221.411
R3541 pfd_8_0.QB_b.n0 pfd_8_0.QB_b.t0 24.0005
R3542 pfd_8_0.QB_b.n0 pfd_8_0.QB_b.t2 24.0005
R3543 a_870_640.t0 a_870_640.t1 39.4005
R3544 VCO_FD_magic_0.div120_2_0.div5_2_0.F.t0 VCO_FD_magic_0.div120_2_0.div5_2_0.F.t1 157.601
R3545 a_2530_190.t1 a_2530_190.n2 500.086
R3546 a_2530_190.n0 a_2530_190.t2 465.933
R3547 a_2530_190.t1 a_2530_190.n2 461.389
R3548 a_2530_190.n1 a_2530_190.n0 392.623
R3549 a_2530_190.n0 a_2530_190.t3 321.334
R3550 a_2530_190.n1 a_2530_190.t0 177.577
R3551 a_2530_190.n2 a_2530_190.n1 48.3899
R3552 a_2200_190.t1 a_2200_190.n2 500.086
R3553 a_2200_190.n1 a_2200_190.n0 473.334
R3554 a_2200_190.n0 a_2200_190.t2 465.933
R3555 a_2200_190.t1 a_2200_190.n2 461.389
R3556 a_2200_190.n0 a_2200_190.t3 321.334
R3557 a_2200_190.n1 a_2200_190.t0 177.577
R3558 a_2200_190.n2 a_2200_190.n1 48.3898
R3559 a_9360_3514.t1 a_9360_3514.t0 323.964
R3560 VCO_FD_magic_0.div120_2_0.div5_2_0.B.n0 VCO_FD_magic_0.div120_2_0.div5_2_0.B.t1 663.801
R3561 VCO_FD_magic_0.div120_2_0.div5_2_0.B.t0 VCO_FD_magic_0.div120_2_0.div5_2_0.B.n0 397.053
R3562 VCO_FD_magic_0.div120_2_0.div5_2_0.B.n0 VCO_FD_magic_0.div120_2_0.div5_2_0.B.t2 348.851
R3563 VCO_FD_magic_0.vco2_3_0.V9.n1 VCO_FD_magic_0.vco2_3_0.V9.n0 437.733
R3564 VCO_FD_magic_0.vco2_3_0.V9.t0 VCO_FD_magic_0.vco2_3_0.V9.n1 372.118
R3565 VCO_FD_magic_0.vco2_3_0.V9.n1 VCO_FD_magic_0.vco2_3_0.V9.t1 247.934
R3566 VCO_FD_magic_0.vco2_3_0.V9.n0 VCO_FD_magic_0.vco2_3_0.V9.t2 224.934
R3567 VCO_FD_magic_0.vco2_3_0.V9.n0 VCO_FD_magic_0.vco2_3_0.V9.t3 144.601
R3568 VCO_FD_magic_0.vco2_3_0.V8.n1 VCO_FD_magic_0.vco2_3_0.V8.n0 437.733
R3569 VCO_FD_magic_0.vco2_3_0.V8.t1 VCO_FD_magic_0.vco2_3_0.V8.n1 372.118
R3570 VCO_FD_magic_0.vco2_3_0.V8.n1 VCO_FD_magic_0.vco2_3_0.V8.t0 247.934
R3571 VCO_FD_magic_0.vco2_3_0.V8.n0 VCO_FD_magic_0.vco2_3_0.V8.t3 224.934
R3572 VCO_FD_magic_0.vco2_3_0.V8.n0 VCO_FD_magic_0.vco2_3_0.V8.t2 144.601
R3573 VCO_FD_magic_0.vco2_3_0.V3.n0 VCO_FD_magic_0.vco2_3_0.V3.t0 284.2
R3574 VCO_FD_magic_0.vco2_3_0.V3.n0 VCO_FD_magic_0.vco2_3_0.V3.t2 233
R3575 VCO_FD_magic_0.vco2_3_0.V3 VCO_FD_magic_0.vco2_3_0.V3.t1 162.857
R3576 VCO_FD_magic_0.vco2_3_0.V3 VCO_FD_magic_0.vco2_3_0.V3.n0 21.3338
R3577 pfd_8_0.F.n4 pfd_8_0.F.n0 1319.38
R3578 pfd_8_0.F.n0 pfd_8_0.F.t3 562.333
R3579 pfd_8_0.F.n2 pfd_8_0.F.t5 388.813
R3580 pfd_8_0.F.n2 pfd_8_0.F.t6 356.68
R3581 pfd_8_0.F.n3 pfd_8_0.F.n2 232
R3582 pfd_8_0.F.n0 pfd_8_0.F.t4 224.934
R3583 pfd_8_0.F.t0 pfd_8_0.F.n4 221.411
R3584 pfd_8_0.F.n3 pfd_8_0.F.n1 157.278
R3585 pfd_8_0.F.n4 pfd_8_0.F.n3 90.64
R3586 pfd_8_0.F.n1 pfd_8_0.F.t2 24.0005
R3587 pfd_8_0.F.n1 pfd_8_0.F.t1 24.0005
R3588 VCO_FD_magic_0.div120_2_0.div5_2_0.D VCO_FD_magic_0.div120_2_0.div5_2_0.D.t3 742.201
R3589 VCO_FD_magic_0.div120_2_0.div5_2_0.D.n1 VCO_FD_magic_0.div120_2_0.div5_2_0.D.t4 350.349
R3590 VCO_FD_magic_0.div120_2_0.div5_2_0.D.n2 VCO_FD_magic_0.div120_2_0.div5_2_0.D.t0 254.333
R3591 VCO_FD_magic_0.div120_2_0.div5_2_0.D.n1 VCO_FD_magic_0.div120_2_0.div5_2_0.D.n0 206.333
R3592 VCO_FD_magic_0.div120_2_0.div5_2_0.D.n2 VCO_FD_magic_0.div120_2_0.div5_2_0.D.n1 70.4005
R3593 VCO_FD_magic_0.div120_2_0.div5_2_0.D.n0 VCO_FD_magic_0.div120_2_0.div5_2_0.D.t2 48.0005
R3594 VCO_FD_magic_0.div120_2_0.div5_2_0.D.n0 VCO_FD_magic_0.div120_2_0.div5_2_0.D.t1 48.0005
R3595 VCO_FD_magic_0.div120_2_0.div5_2_0.D VCO_FD_magic_0.div120_2_0.div5_2_0.D.n2 19.2005
R3596 VCO_FD_magic_0.div120_2_0.div2_4_1.A.n0 VCO_FD_magic_0.div120_2_0.div2_4_1.A.t1 713.933
R3597 VCO_FD_magic_0.div120_2_0.div2_4_1.A VCO_FD_magic_0.div120_2_0.div2_4_1.A.t0 327.401
R3598 VCO_FD_magic_0.div120_2_0.div2_4_1.A.n0 VCO_FD_magic_0.div120_2_0.div2_4_1.A.t2 314.233
R3599 VCO_FD_magic_0.div120_2_0.div2_4_1.A VCO_FD_magic_0.div120_2_0.div2_4_1.A.n0 9.6005
R3600 VCO_FD_magic_0.div120_2_0.div2_4_1.B.t0 VCO_FD_magic_0.div120_2_0.div2_4_1.B.t1 96.0005
R3601 VCO_FD_magic_0.div120_2_0.div3_3_0.G.t0 VCO_FD_magic_0.div120_2_0.div3_3_0.G.t1 96.0005
R3602 VCO_FD_magic_0.div120_2_0.div5_2_0.M VCO_FD_magic_0.div120_2_0.div5_2_0.M.t3 739
R3603 VCO_FD_magic_0.div120_2_0.div5_2_0.M.n1 VCO_FD_magic_0.div120_2_0.div5_2_0.M.t4 349.433
R3604 VCO_FD_magic_0.div120_2_0.div5_2_0.M.n2 VCO_FD_magic_0.div120_2_0.div5_2_0.M.t1 254.333
R3605 VCO_FD_magic_0.div120_2_0.div5_2_0.M.n1 VCO_FD_magic_0.div120_2_0.div5_2_0.M.n0 206.333
R3606 VCO_FD_magic_0.div120_2_0.div5_2_0.M.n2 VCO_FD_magic_0.div120_2_0.div5_2_0.M.n1 70.4005
R3607 VCO_FD_magic_0.div120_2_0.div5_2_0.M.n0 VCO_FD_magic_0.div120_2_0.div5_2_0.M.t2 48.0005
R3608 VCO_FD_magic_0.div120_2_0.div5_2_0.M.n0 VCO_FD_magic_0.div120_2_0.div5_2_0.M.t0 48.0005
R3609 VCO_FD_magic_0.div120_2_0.div5_2_0.M VCO_FD_magic_0.div120_2_0.div5_2_0.M.n2 22.4005
R3610 a_9360_6440.t1 a_9360_6440.t0 245.883
R3611 VCO_FD_magic_0.div120_2_0.div2_4_0.A.n0 VCO_FD_magic_0.div120_2_0.div2_4_0.A.t1 713.933
R3612 VCO_FD_magic_0.div120_2_0.div2_4_0.A VCO_FD_magic_0.div120_2_0.div2_4_0.A.t0 327.401
R3613 VCO_FD_magic_0.div120_2_0.div2_4_0.A.n0 VCO_FD_magic_0.div120_2_0.div2_4_0.A.t2 314.233
R3614 VCO_FD_magic_0.div120_2_0.div2_4_0.A VCO_FD_magic_0.div120_2_0.div2_4_0.A.n0 9.6005
R3615 pfd_8_0.F_b.n0 pfd_8_0.F_b.t3 517.347
R3616 pfd_8_0.F_b.n2 pfd_8_0.F_b.n0 417.574
R3617 pfd_8_0.F_b.n2 pfd_8_0.F_b.n1 244.716
R3618 pfd_8_0.F_b.n0 pfd_8_0.F_b.t4 228.148
R3619 pfd_8_0.F_b.t1 pfd_8_0.F_b.n2 221.411
R3620 pfd_8_0.F_b.n1 pfd_8_0.F_b.t0 24.0005
R3621 pfd_8_0.F_b.n1 pfd_8_0.F_b.t2 24.0005
R3622 a_1390_640.t0 a_1390_640.t1 39.4005
R3623 VCO_FD_magic_0.div120_2_0.div5_2_0.L.t0 VCO_FD_magic_0.div120_2_0.div5_2_0.L.t1 96.0005
R3624 VCO_FD_magic_0.div120_2_0.div3_3_0.E.n0 VCO_FD_magic_0.div120_2_0.div3_3_0.E.t0 685.134
R3625 VCO_FD_magic_0.div120_2_0.div3_3_0.E.n1 VCO_FD_magic_0.div120_2_0.div3_3_0.E.t2 663.801
R3626 VCO_FD_magic_0.div120_2_0.div3_3_0.E.n0 VCO_FD_magic_0.div120_2_0.div3_3_0.E.t3 534.268
R3627 VCO_FD_magic_0.div120_2_0.div3_3_0.E.t1 VCO_FD_magic_0.div120_2_0.div3_3_0.E.n1 362.921
R3628 VCO_FD_magic_0.div120_2_0.div3_3_0.E.n1 VCO_FD_magic_0.div120_2_0.div3_3_0.E.n0 91.7338
R3629 VCO_FD_magic_0.div120_2_0.div5_2_0.K.n0 VCO_FD_magic_0.div120_2_0.div5_2_0.K.t1 663.801
R3630 VCO_FD_magic_0.div120_2_0.div5_2_0.K.n0 VCO_FD_magic_0.div120_2_0.div5_2_0.K.t2 355.378
R3631 VCO_FD_magic_0.div120_2_0.div5_2_0.K VCO_FD_magic_0.div120_2_0.div5_2_0.K.t0 276.521
R3632 VCO_FD_magic_0.div120_2_0.div5_2_0.K VCO_FD_magic_0.div120_2_0.div5_2_0.K.n0 120.534
R3633 a_490_640.t0 a_490_640.t1 39.4005
R3634 VCO_FD_magic_0.div120_2_0.div2_4_0.B.t0 VCO_FD_magic_0.div120_2_0.div2_4_0.B.t1 96.0005
R3635 VCO_FD_magic_0.vco2_3_0.V7.n0 VCO_FD_magic_0.vco2_3_0.V7.t0 284.2
R3636 VCO_FD_magic_0.vco2_3_0.V7.n0 VCO_FD_magic_0.vco2_3_0.V7.t2 233
R3637 VCO_FD_magic_0.vco2_3_0.V7 VCO_FD_magic_0.vco2_3_0.V7.t1 162.857
R3638 VCO_FD_magic_0.vco2_3_0.V7 VCO_FD_magic_0.vco2_3_0.V7.n0 21.3338
R3639 VCO_FD_magic_0.vco2_3_0.V5.n0 VCO_FD_magic_0.vco2_3_0.V5.t0 284.2
R3640 VCO_FD_magic_0.vco2_3_0.V5.n0 VCO_FD_magic_0.vco2_3_0.V5.t2 233
R3641 VCO_FD_magic_0.vco2_3_0.V5 VCO_FD_magic_0.vco2_3_0.V5.t1 162.857
R3642 VCO_FD_magic_0.vco2_3_0.V5 VCO_FD_magic_0.vco2_3_0.V5.n0 21.3338
R3643 VCO_FD_magic_0.vco2_3_0.V2.n0 VCO_FD_magic_0.vco2_3_0.V2.t1 421.027
R3644 VCO_FD_magic_0.vco2_3_0.V2.n0 VCO_FD_magic_0.vco2_3_0.V2.t2 348.81
R3645 VCO_FD_magic_0.vco2_3_0.V2 VCO_FD_magic_0.vco2_3_0.V2.t0 284.317
R3646 VCO_FD_magic_0.vco2_3_0.V2 VCO_FD_magic_0.vco2_3_0.V2.n0 31.8427
R3647 VCO_FD_magic_0.div120_2_0.div5_2_0.E.n0 VCO_FD_magic_0.div120_2_0.div5_2_0.E.t0 723
R3648 VCO_FD_magic_0.div120_2_0.div5_2_0.E.t3 VCO_FD_magic_0.div120_2_0.div5_2_0.E.t2 514.134
R3649 VCO_FD_magic_0.div120_2_0.div5_2_0.E.n1 VCO_FD_magic_0.div120_2_0.div5_2_0.E.t3 332.783
R3650 VCO_FD_magic_0.div120_2_0.div5_2_0.E.n0 VCO_FD_magic_0.div120_2_0.div5_2_0.E.t1 314.921
R3651 VCO_FD_magic_0.div120_2_0.div5_2_0.E VCO_FD_magic_0.div120_2_0.div5_2_0.E.n1 6.4005
R3652 VCO_FD_magic_0.div120_2_0.div5_2_0.E.n1 VCO_FD_magic_0.div120_2_0.div5_2_0.E.n0 3.2005
R3653 a_490_1400.t0 a_490_1400.t1 39.4005
R3654 pfd_8_0.Reset.n1 pfd_8_0.Reset.t3 562.333
R3655 pfd_8_0.Reset.n2 pfd_8_0.Reset.n1 480.45
R3656 pfd_8_0.Reset.n0 pfd_8_0.Reset.t4 417.733
R3657 pfd_8_0.Reset.n0 pfd_8_0.Reset.t5 369.534
R3658 pfd_8_0.Reset.n3 pfd_8_0.Reset.n2 328.733
R3659 pfd_8_0.Reset.t1 pfd_8_0.Reset.n3 288.37
R3660 pfd_8_0.Reset.n1 pfd_8_0.Reset.t2 224.934
R3661 pfd_8_0.Reset.n3 pfd_8_0.Reset.t0 177.577
R3662 pfd_8_0.Reset.n2 pfd_8_0.Reset.n0 176.733
R3663 VCO_FD_magic_0.div120_2_0.div3_3_0.B.t0 VCO_FD_magic_0.div120_2_0.div3_3_0.B.t1 96.0005
R3664 a_1870_190.t1 a_1870_190.n2 500.086
R3665 a_1870_190.n1 a_1870_190.n0 473.334
R3666 a_1870_190.n0 a_1870_190.t2 465.933
R3667 a_1870_190.t1 a_1870_190.n2 461.389
R3668 a_1870_190.n0 a_1870_190.t3 321.334
R3669 a_1870_190.n1 a_1870_190.t0 177.577
R3670 a_1870_190.n2 a_1870_190.n1 48.3898
R3671 VCO_FD_magic_0.div120_2_0.div3_3_0.A.n0 VCO_FD_magic_0.div120_2_0.div3_3_0.A.t0 713.933
R3672 VCO_FD_magic_0.div120_2_0.div3_3_0.A.n0 VCO_FD_magic_0.div120_2_0.div3_3_0.A.t2 314.233
R3673 VCO_FD_magic_0.div120_2_0.div3_3_0.A.t1 VCO_FD_magic_0.div120_2_0.div3_3_0.A.n0 308.2
R3674 VCO_FD_magic_0.vco2_3_0.V6.n0 VCO_FD_magic_0.vco2_3_0.V6.t0 421.027
R3675 VCO_FD_magic_0.vco2_3_0.V6.n0 VCO_FD_magic_0.vco2_3_0.V6.t2 348.81
R3676 VCO_FD_magic_0.vco2_3_0.V6 VCO_FD_magic_0.vco2_3_0.V6.t1 280.05
R3677 VCO_FD_magic_0.vco2_3_0.V6 VCO_FD_magic_0.vco2_3_0.V6.n0 36.1094
R3678 VCO_FD_magic_0.div120_2_0.div3_3_0.F.t0 VCO_FD_magic_0.div120_2_0.div3_3_0.F.t1 96.0005
R3679 a_n30_640.t0 a_n30_640.t1 39.4005
C0 VCO_FD_magic_0.div120_2_0.div5_2_0.I F_VCO 0.021863f
C1 VCO_FD_magic_0.div120_2_0.div5_2_0.I VCO_FD_magic_0.div120_2_0.div24 0.076865f
C2 VCO_FD_magic_0.div120_2_0.div3_3_0.C VCO_FD_magic_0.div120_2_0.div24 0.03648f
C3 VCO_FD_magic_0.div120_2_0.div3_3_0.D VCO_FD_magic_0.div120_2_0.div24 0.024014f
C4 VCO_FD_magic_0.div120_2_0.div5_2_0.E VCO_FD_magic_0.div120_2_0.div5_2_0.I 0.021344f
C5 VCO_FD_magic_0.div120_2_0.div5_2_0.G VCO_FD_magic_0.div120_2_0.div5_2_0.I 0.069172f
C6 VDDA VCO_FD_magic_0.div120_2_0.div2_4_2.C 0.111144f
C7 VCO_FD_magic_0.div120_2_0.div2_4_1.A VDDA 0.126015f
C8 VCO_FD_magic_0.div120_2_0.div5_2_0.M VDDA 0.157966f
C9 VCO_FD_magic_0.div120_2_0.div5_2_0.J VDDA 0.104998f
C10 pfd_8_0.QA F_REF 0.056f
C11 VCO_FD_magic_0.div120_2_0.div2_4_0.A VCO_FD_magic_0.div120_2_0.div2_4_0.C 0.122602f
C12 V_OSC VCO_FD_magic_0.vco2_3_0.V5 0.017652f
C13 pfd_8_0.QB F_VCO 0.060952f
C14 pfd_8_0.QA_b pfd_8_0.QA 0.422694f
C15 VCO_FD_magic_0.div120_2_0.div5_2_0.K VDDA 0.482256f
C16 VCO_FD_magic_0.div120_2_0.div3_3_0.H VDDA 0.106696f
C17 VCO_FD_magic_0.div120_2_0.div24 F_VCO 0.067501f
C18 VCO_FD_magic_0.div120_2_0.div5_2_0.D VCO_FD_magic_0.div120_2_0.div24 0.163145f
C19 VCO_FD_magic_0.div120_2_0.div5_2_0.E F_VCO 0.139506f
C20 VCO_FD_magic_0.div120_2_0.div5_2_0.G F_VCO 0.081976f
C21 VCO_FD_magic_0.div120_2_0.div5_2_0.E VCO_FD_magic_0.div120_2_0.div24 0.108607f
C22 pfd_8_0.DOWN_input I_IN 0.928029f
C23 VCO_FD_magic_0.div120_2_0.div5_2_0.G VCO_FD_magic_0.div120_2_0.div24 0.240642f
C24 VDDA F_REF 0.098433f
C25 VCO_FD_magic_0.div120_2_0.div5_2_0.K VCO_FD_magic_0.div120_2_0.div5_2_0.M 0.169071f
C26 V_OSC VDDA 0.627267f
C27 pfd_8_0.DOWN_input opamp_cell_4_0.VIN+ 0.080549f
C28 pfd_8_0.QA_b VDDA 0.52066f
C29 VCO_FD_magic_0.div120_2_0.div5_2_0.E VCO_FD_magic_0.div120_2_0.div5_2_0.D 0.070599f
C30 pfd_8_0.QB pfd_8_0.QB_b 0.388258f
C31 VDDA VCO_FD_magic_0.vco2_3_0.V6 0.281338f
C32 F_VCO pfd_8_0.QB_b 0.044529f
C33 opamp_cell_4_0.p_bias VDDA 2.86573f
C34 VCO_FD_magic_0.div120_2_0.div5_2_0.E VCO_FD_magic_0.div120_2_0.div5_2_0.G 0.112235f
C35 VCO_FD_magic_0.vco2_3_0.V3 VDDA 0.040599f
C36 VDDA VCO_FD_magic_0.div120_2_0.div3_3_0.C 0.125686f
C37 VCO_FD_magic_0.vco2_3_0.V7 VDDA 0.033517f
C38 VDDA VCO_FD_magic_0.vco2_3_0.V2 0.410554f
C39 pfd_8_0.QA pfd_8_0.QB 0.074487f
C40 VDDA VCO_FD_magic_0.div120_2_0.div3_3_0.D 0.311052f
C41 I_IN VDDA 0.541032f
C42 opamp_cell_4_0.VIN+ VDDA 0.832915f
C43 VCO_FD_magic_0.div120_2_0.div5_2_0.J VCO_FD_magic_0.div120_2_0.div5_2_0.I 0.016448f
C44 VCO_FD_magic_0.div120_2_0.div2_4_2.A VDDA 0.125335f
C45 VCO_FD_magic_0.div120_2_0.div2_4_0.A VDDA 0.125335f
C46 VDDA VCO_FD_magic_0.div120_2_0.div2_4_0.C 0.111144f
C47 pfd_8_0.QB VDDA 2.75013f
C48 VDDA F_VCO 1.25401f
C49 VDDA VCO_FD_magic_0.div120_2_0.div24 0.654009f
C50 pfd_8_0.QA_b F_REF 0.027208f
C51 VCO_FD_magic_0.div120_2_0.div2_4_1.C VDDA 0.111409f
C52 VCO_FD_magic_0.div120_2_0.div2_4_2.A VCO_FD_magic_0.div120_2_0.div2_4_2.C 0.122602f
C53 VCO_FD_magic_0.div120_2_0.div5_2_0.D VDDA 0.144695f
C54 V_OSC VCO_FD_magic_0.vco2_3_0.V6 0.019495f
C55 VCO_FD_magic_0.div120_2_0.div5_2_0.E VDDA 0.53342f
C56 VCO_FD_magic_0.div120_2_0.div5_2_0.G VDDA 0.25905f
C57 V_OSC VCO_FD_magic_0.vco2_3_0.V3 0.046941f
C58 VCO_FD_magic_0.div120_2_0.div5_2_0.M F_VCO 0.119081f
C59 VCO_FD_magic_0.div120_2_0.div5_2_0.J F_VCO 0.036046f
C60 VCO_FD_magic_0.vco2_3_0.V7 V_OSC 0.108092f
C61 VCO_FD_magic_0.div120_2_0.div2_4_1.A VCO_FD_magic_0.div120_2_0.div2_4_1.C 0.122602f
C62 VCO_FD_magic_0.div120_2_0.div5_2_0.J VCO_FD_magic_0.div120_2_0.div24 0.176046f
C63 V_OSC VCO_FD_magic_0.vco2_3_0.V2 0.063469f
C64 VCO_FD_magic_0.vco2_3_0.V5 VCO_FD_magic_0.vco2_3_0.V4 0.010316f
C65 VCO_FD_magic_0.div120_2_0.div5_2_0.K F_VCO 0.174679f
C66 VCO_FD_magic_0.vco2_3_0.V7 VCO_FD_magic_0.vco2_3_0.V6 0.010316f
C67 VCO_FD_magic_0.div120_2_0.div3_3_0.H VCO_FD_magic_0.div120_2_0.div24 0.038583f
C68 VDDA pfd_8_0.QB_b 0.512673f
C69 VCO_FD_magic_0.vco2_3_0.V3 VCO_FD_magic_0.vco2_3_0.V2 0.010316f
C70 VCO_FD_magic_0.div120_2_0.div5_2_0.J VCO_FD_magic_0.div120_2_0.div5_2_0.G 0.061186f
C71 pfd_8_0.DOWN_input VDDA 0.221484f
C72 opamp_cell_4_0.VIN+ opamp_cell_4_0.p_bias 0.100967f
C73 VCO_FD_magic_0.div120_2_0.div3_3_0.D VCO_FD_magic_0.div120_2_0.div3_3_0.C 0.060684f
C74 VCO_FD_magic_0.vco2_3_0.V5 VDDA 0.040599f
C75 pfd_8_0.QA VDDA 0.550605f
C76 VDDA VCO_FD_magic_0.vco2_3_0.V4 0.413959f
C77 I_IN opamp_cell_4_0.VIN+ 0.166322f
C78 V_OSC GNDA 2.90637f
C79 I_IN GNDA 2.82399f
C80 F_REF GNDA 0.277742f
C81 VDDA GNDA 71.3612f
C82 VCO_FD_magic_0.vco2_3_0.V2 GNDA 0.045471f
C83 VCO_FD_magic_0.vco2_3_0.V4 GNDA 0.045471f
C84 VCO_FD_magic_0.vco2_3_0.V6 GNDA 0.157087f
C85 VCO_FD_magic_0.div120_2_0.div2_4_1.A GNDA 0.200071f
C86 VCO_FD_magic_0.div120_2_0.div2_4_2.A GNDA 0.200074f
C87 VCO_FD_magic_0.div120_2_0.div2_4_0.A GNDA 0.200071f
C88 VCO_FD_magic_0.div120_2_0.div5_2_0.G GNDA 0.195152f
C89 VCO_FD_magic_0.div120_2_0.div5_2_0.I GNDA 0.152847f
C90 VCO_FD_magic_0.div120_2_0.div3_3_0.C GNDA 0.36191f
C91 VCO_FD_magic_0.div120_2_0.div3_3_0.D GNDA 0.301961f
C92 VCO_FD_magic_0.div120_2_0.div3_3_0.H GNDA 0.423425f
C93 VCO_FD_magic_0.div120_2_0.div5_2_0.D GNDA 0.366928f
C94 VCO_FD_magic_0.div120_2_0.div5_2_0.E GNDA 0.297109f
C95 VCO_FD_magic_0.div120_2_0.div5_2_0.J GNDA 0.398061f
C96 VCO_FD_magic_0.div120_2_0.div5_2_0.K GNDA 0.180033f
C97 VCO_FD_magic_0.div120_2_0.div5_2_0.M GNDA 0.397035f
C98 VCO_FD_magic_0.div120_2_0.div2_4_1.C GNDA 0.45763f
C99 VCO_FD_magic_0.div120_2_0.div2_4_2.C GNDA 0.457627f
C100 VCO_FD_magic_0.div120_2_0.div2_4_0.C GNDA 0.46146f
C101 VCO_FD_magic_0.div120_2_0.div24 GNDA 3.78529f
C102 VCO_FD_magic_0.vco2_3_0.V3 GNDA 0.300759f
C103 VCO_FD_magic_0.vco2_3_0.V5 GNDA 0.302737f
C104 VCO_FD_magic_0.vco2_3_0.V7 GNDA 0.314921f
C105 pfd_8_0.DOWN_input GNDA 3.02729f
C106 pfd_8_0.QB_b GNDA 1.04775f
C107 F_VCO GNDA 3.25572f
C108 pfd_8_0.QB GNDA 1.307779f
C109 pfd_8_0.QA GNDA 3.10102f
C110 pfd_8_0.QA_b GNDA 1.05138f
C111 opamp_cell_4_0.VIN+ GNDA 2.37749f
C112 opamp_cell_4_0.p_bias GNDA 3.954681f
C113 pfd_8_0.QB.t7 GNDA 0.069179f
C114 pfd_8_0.QB.t8 GNDA 0.032493f
C115 pfd_8_0.QB.n0 GNDA 0.099932f
C116 pfd_8_0.QB.t3 GNDA 0.069179f
C117 pfd_8_0.QB.t4 GNDA 0.104293f
C118 pfd_8_0.QB.n1 GNDA 1.25065f
C119 pfd_8_0.QB.t5 GNDA 0.069862f
C120 pfd_8_0.QB.t6 GNDA 0.030633f
C121 pfd_8_0.QB.n2 GNDA 0.176466f
C122 pfd_8_0.QB.t0 GNDA 0.147114f
C123 pfd_8_0.QB.t1 GNDA 0.027951f
C124 pfd_8_0.QB.t2 GNDA 0.027951f
C125 pfd_8_0.QB.n3 GNDA 0.149246f
C126 pfd_8_0.QB.n4 GNDA 0.265156f
C127 pfd_8_0.QB.n5 GNDA 0.226459f
C128 loop_filter_3_0.R1_C1.t1 GNDA 2.79887f
C129 opamp_cell_4_0.p_bias.t0 GNDA 1.66267f
C130 opamp_cell_4_0.p_bias.t2 GNDA 0.019693f
C131 opamp_cell_4_0.p_bias.t6 GNDA 0.019693f
C132 opamp_cell_4_0.p_bias.n0 GNDA 0.054067f
C133 opamp_cell_4_0.p_bias.t8 GNDA 0.019693f
C134 opamp_cell_4_0.p_bias.t4 GNDA 0.019693f
C135 opamp_cell_4_0.p_bias.n1 GNDA 0.054067f
C136 opamp_cell_4_0.p_bias.n2 GNDA 0.068502f
C137 opamp_cell_4_0.p_bias.t1 GNDA 0.054353f
C138 opamp_cell_4_0.p_bias.t3 GNDA 0.054353f
C139 opamp_cell_4_0.p_bias.t7 GNDA 0.054353f
C140 opamp_cell_4_0.p_bias.t11 GNDA 0.054353f
C141 opamp_cell_4_0.p_bias.t9 GNDA 0.074733f
C142 opamp_cell_4_0.p_bias.n3 GNDA 0.04185f
C143 opamp_cell_4_0.p_bias.n4 GNDA 0.029697f
C144 opamp_cell_4_0.p_bias.n5 GNDA 0.012761f
C145 opamp_cell_4_0.p_bias.n6 GNDA 0.029697f
C146 opamp_cell_4_0.p_bias.n7 GNDA 0.029697f
C147 opamp_cell_4_0.p_bias.t5 GNDA 0.054353f
C148 opamp_cell_4_0.p_bias.t12 GNDA 0.054353f
C149 opamp_cell_4_0.p_bias.t10 GNDA 0.074733f
C150 opamp_cell_4_0.p_bias.n8 GNDA 0.04185f
C151 opamp_cell_4_0.p_bias.n9 GNDA 0.029697f
C152 opamp_cell_4_0.p_bias.n10 GNDA 0.012761f
C153 opamp_cell_4_0.p_bias.n11 GNDA 0.120625f
C154 pfd_8_0.opamp_out.t12 GNDA 0.957954f
C155 pfd_8_0.opamp_out.t11 GNDA 0.957546f
C156 pfd_8_0.opamp_out.n6 GNDA 0.012958f
C157 pfd_8_0.opamp_out.t14 GNDA 0.012873f
C158 pfd_8_0.opamp_out.t0 GNDA 0.012026f
C159 pfd_8_0.opamp_out.n13 GNDA 0.015342f
C160 pfd_8_0.opamp_out.n14 GNDA 0.081091f
C161 pfd_8_0.opamp_out.n15 GNDA 0.047633f
C162 VCO_FD_magic_0.vco2_3_0.V1.t1 GNDA 0.104706f
C163 VCO_FD_magic_0.vco2_3_0.V1.n0 GNDA 0.184398f
C164 VCO_FD_magic_0.vco2_3_0.V1.t4 GNDA 0.298444f
C165 VCO_FD_magic_0.vco2_3_0.V1.t3 GNDA 0.298444f
C166 VCO_FD_magic_0.vco2_3_0.V1.t5 GNDA 0.497217f
C167 VCO_FD_magic_0.vco2_3_0.V1.n1 GNDA 0.243367f
C168 VCO_FD_magic_0.vco2_3_0.V1.n2 GNDA 0.217957f
C169 VCO_FD_magic_0.vco2_3_0.V1.t0 GNDA 0.298444f
C170 VCO_FD_magic_0.vco2_3_0.V1.n3 GNDA 0.169192f
C171 VCO_FD_magic_0.vco2_3_0.V1.n4 GNDA 0.045341f
C172 VCO_FD_magic_0.vco2_3_0.V1.n5 GNDA 0.177452f
C173 VCO_FD_magic_0.vco2_3_0.V1.t2 GNDA 0.165036f
C174 VDDA.n71 GNDA 0.051784f
C175 VDDA.t29 GNDA 0.173447f
C176 VDDA.n74 GNDA 0.115632f
C177 VDDA.n80 GNDA 0.01246f
C178 VDDA.n86 GNDA 0.014434f
C179 VDDA.n87 GNDA 0.03888f
C180 VDDA.t184 GNDA 0.089652f
C181 VDDA.t2 GNDA 0.070664f
C182 VDDA.t73 GNDA 0.033245f
C183 VDDA.n90 GNDA 0.014698f
C184 VDDA.t59 GNDA 0.015182f
C185 VDDA.t210 GNDA 0.025751f
C186 VDDA.t0 GNDA 0.025751f
C187 VDDA.t66 GNDA 0.016911f
C188 VDDA.t195 GNDA 0.016911f
C189 VDDA.t69 GNDA 0.028057f
C190 VDDA.t99 GNDA 0.029018f
C191 VDDA.n91 GNDA 0.014698f
C192 VDDA.t120 GNDA 0.015182f
C193 VDDA.t188 GNDA 0.017295f
C194 VDDA.t36 GNDA 0.017295f
C195 VDDA.t34 GNDA 0.013836f
C196 VDDA.t91 GNDA 0.013836f
C197 VDDA.t214 GNDA 0.022292f
C198 VDDA.t200 GNDA 0.022292f
C199 VDDA.t26 GNDA 0.016911f
C200 VDDA.t15 GNDA 0.016911f
C201 VDDA.t40 GNDA 0.023829f
C202 VDDA.t208 GNDA 0.02479f
C203 VDDA.n92 GNDA 0.011623f
C204 VDDA.t128 GNDA 0.012107f
C205 VDDA.t122 GNDA 0.013836f
C206 VDDA.t132 GNDA 0.013836f
C207 VDDA.t216 GNDA 0.02306f
C208 VDDA.t22 GNDA 0.024021f
C209 VDDA.n94 GNDA 0.011623f
C210 VDDA.t202 GNDA 0.012107f
C211 VDDA.t93 GNDA 0.013836f
C212 VDDA.t84 GNDA 0.013836f
C213 VDDA.t186 GNDA 0.02306f
C214 VDDA.t86 GNDA 0.024021f
C215 VDDA.n95 GNDA 0.011623f
C216 VDDA.t5 GNDA 0.012107f
C217 VDDA.t54 GNDA 0.013836f
C218 VDDA.t212 GNDA 0.013836f
C219 VDDA.t193 GNDA 0.02306f
C220 VDDA.t56 GNDA 0.024021f
C221 VDDA.n97 GNDA 0.011623f
C222 VDDA.t97 GNDA 0.012107f
C223 VDDA.t204 GNDA 0.013836f
C224 VDDA.t106 GNDA 0.013836f
C225 VDDA.t7 GNDA 0.0214f
C226 VDDA.t119 GNDA 0.100683f
C227 VDDA.t43 GNDA 0.089652f
C228 VDDA.n99 GNDA 0.038136f
C229 VDDA.n108 GNDA 0.099572f
C230 VDDA.t42 GNDA 0.070664f
C231 VDDA.t47 GNDA 0.089652f
C232 VDDA.n110 GNDA 0.038136f
C233 VDDA.n116 GNDA 0.099572f
C234 VDDA.n128 GNDA 0.05312f
C235 VDDA.n129 GNDA 0.039691f
C236 VDDA.n300 GNDA 0.093595f
C237 VDDA.t24 GNDA 0.030637f
C238 VDDA.t199 GNDA 0.011111f
C239 VDDA.n324 GNDA 0.012169f
C240 VDDA.t219 GNDA 0.030637f
C241 VDDA.n341 GNDA 0.028191f
C242 VDDA.n344 GNDA 0.010981f
C243 VDDA.t11 GNDA 0.10326f
C244 VDDA.n350 GNDA 0.010981f
C245 VDDA.n351 GNDA 0.010981f
C246 VDDA.n379 GNDA 0.010229f
C247 VDDA.n387 GNDA 0.050308f
C248 VDDA.t168 GNDA 0.123217f
C249 VDDA.t101 GNDA 0.062336f
C250 VDDA.t117 GNDA 0.062336f
C251 VDDA.t138 GNDA 0.062336f
C252 VDDA.t31 GNDA 0.062336f
C253 VDDA.t174 GNDA 0.070728f
C254 VDDA.n392 GNDA 0.013768f
C255 VDDA.t156 GNDA 0.018131f
C256 VDDA.n397 GNDA 0.013726f
C257 VDDA.n407 GNDA 0.099498f
C258 VDDA.t147 GNDA 0.047951f
C259 VDDA.t157 GNDA 0.031168f
C260 VDDA.t145 GNDA 0.037162f
C261 VDDA.t146 GNDA 0.041957f
C262 VDDA.t124 GNDA 0.031168f
C263 VDDA.t192 GNDA 0.047951f
C264 VDDA.t112 GNDA 0.031168f
C265 VDDA.t90 GNDA 0.034764f
C266 VDDA.t148 GNDA 0.044355f
C267 VDDA.t3 GNDA 0.061138f
C268 VDDA.t80 GNDA 0.064734f
C269 VDDA.n408 GNDA 0.051668f
C270 VDDA.t190 GNDA 0.03956f
C271 VDDA.t153 GNDA 0.03956f
C272 VDDA.t110 GNDA 0.03956f
C273 VDDA.t38 GNDA 0.031168f
C274 VDDA.t75 GNDA 0.047951f
C275 VDDA.t140 GNDA 0.031168f
C276 VDDA.t45 GNDA 0.037162f
C277 VDDA.t108 GNDA 0.041957f
C278 VDDA.t103 GNDA 0.031168f
C279 VDDA.t150 GNDA 0.047951f
C280 VDDA.t161 GNDA 0.03956f
C281 VDDA.n412 GNDA 0.016359f
C282 VDDA.n413 GNDA 0.046733f
C283 VDDA.t160 GNDA 0.018502f
C284 VDDA.n416 GNDA 0.013726f
C285 VDDA.n423 GNDA 0.012928f
C286 VDDA.n425 GNDA 0.037812f
C287 VDDA.n426 GNDA 0.045674f
C288 VDDA.n427 GNDA 0.013768f
C289 VDDA.n430 GNDA 0.011329f
C290 VDDA.n431 GNDA 0.032916f
C291 VDDA.n432 GNDA 0.033073f
C292 VDDA.n440 GNDA 0.032073f
C293 VDDA.n447 GNDA 0.032073f
C294 VDDA.n454 GNDA 0.032073f
C295 VDDA.n461 GNDA 0.032073f
C296 VDDA.n471 GNDA 0.021537f
C297 VDDA.n475 GNDA 0.010981f
C298 VDDA.t164 GNDA 0.045645f
C299 VDDA.n482 GNDA 0.010249f
C300 VDDA.n485 GNDA 0.010249f
C301 VDDA.n488 GNDA 0.010584f
C302 VDDA.n489 GNDA 0.014893f
C303 VDDA.n491 GNDA 0.010584f
C304 VDDA.n492 GNDA 0.014893f
C305 VDDA.n511 GNDA 0.010584f
C306 VDDA.n514 GNDA 0.010584f
C307 VDDA.t170 GNDA 0.018245f
C308 VDDA.t134 GNDA 0.046707f
C309 VDDA.t13 GNDA 0.046707f
C310 VDDA.t130 GNDA 0.046707f
C311 VDDA.t64 GNDA 0.046707f
C312 VDDA.t171 GNDA 0.045645f
C313 VDDA.n525 GNDA 0.041399f
C314 VDDA.n530 GNDA 0.010981f
C315 VDDA.n531 GNDA 0.010584f
C316 VDDA.n532 GNDA 0.015082f
C317 VDDA.n539 GNDA 0.014161f
C318 VDDA.n546 GNDA 0.014893f
C319 VDDA.n554 GNDA 0.014893f
C320 VDDA.n555 GNDA 0.010584f
C321 VDDA.n556 GNDA 0.010981f
C322 VDDA.t163 GNDA 0.017216f
C323 VDDA.t177 GNDA 0.017216f
C324 VDDA.n559 GNDA 0.013217f
C325 VDDA.n560 GNDA 0.010981f
C326 VDDA.n561 GNDA 0.012452f
C327 VDDA.n563 GNDA 0.044583f
C328 VDDA.t178 GNDA 0.045645f
C329 VDDA.t88 GNDA 0.046707f
C330 VDDA.t52 GNDA 0.046707f
C331 VDDA.t136 GNDA 0.046707f
C332 VDDA.t71 GNDA 0.046707f
C333 VDDA.t181 GNDA 0.045645f
C334 VDDA.n569 GNDA 0.041399f
C335 VDDA.t180 GNDA 0.018245f
C336 VDDA.n579 GNDA 0.014987f
C337 VDDA.n580 GNDA 0.156827f
C338 VDDA.n581 GNDA 0.028105f
C339 VDDA.n583 GNDA 0.010981f
C340 VDDA.t95 GNDA 0.107798f
C341 VDDA.t68 GNDA 0.116876f
C342 VDDA.n590 GNDA 0.088508f
C343 VDDA.n614 GNDA 0.088508f
C344 VDDA.t126 GNDA 0.088508f
C345 VDDA.t206 GNDA 0.030637f
C346 VDDA.n627 GNDA 0.044254f
C347 VDDA.n635 GNDA 0.044254f
C348 VDDA.t115 GNDA 0.030637f
C349 VDDA.t196 GNDA 0.030637f
C350 VDDA.n643 GNDA 0.06241f
C351 VDDA.n646 GNDA 0.010981f
C352 VDDA.n655 GNDA 0.010981f
C353 VDDA.n663 GNDA 0.096451f
C354 VDDA.t77 GNDA 0.088508f
C355 VDDA.n669 GNDA 0.088508f
C356 VDDA.n705 GNDA 0.044254f
C357 VDDA.t17 GNDA 0.027233f
C358 VDDA.t198 GNDA 0.028368f
C359 VDDA.n711 GNDA 0.044254f
C360 VDDA.n727 GNDA 0.06014f
C361 VDDA.n746 GNDA 0.066949f
C362 VDDA.t82 GNDA 0.055601f
C363 VDDA.t28 GNDA 0.118011f
C364 VDDA.t114 GNDA 0.118011f
C365 VDDA.t49 GNDA 0.055601f
C366 VDDA.n770 GNDA 0.061275f
C367 VDDA.t9 GNDA 0.055601f
C368 VDDA.t33 GNDA 0.118011f
C369 VDDA.t58 GNDA 0.118011f
C370 VDDA.t61 GNDA 0.055601f
C371 VDDA.n783 GNDA 0.06241f
C372 VDDA.n818 GNDA 0.082395f
C373 a_5970_4630.t10 GNDA 0.030769f
C374 a_5970_4630.n0 GNDA 0.124795f
C375 a_5970_4630.t0 GNDA 0.020325f
C376 a_5970_4630.t12 GNDA 0.020325f
C377 a_5970_4630.t6 GNDA 0.020325f
C378 a_5970_4630.n1 GNDA 0.044943f
C379 a_5970_4630.t5 GNDA 0.020325f
C380 a_5970_4630.t8 GNDA 0.020325f
C381 a_5970_4630.n2 GNDA 0.044943f
C382 a_5970_4630.t9 GNDA 0.077457f
C383 a_5970_4630.t7 GNDA 0.030769f
C384 a_5970_4630.n3 GNDA 0.097952f
C385 a_5970_4630.n4 GNDA 0.087903f
C386 a_5970_4630.n5 GNDA 0.089425f
C387 a_5970_4630.t1 GNDA 0.050813f
C388 a_5970_4630.t4 GNDA 0.050813f
C389 a_5970_4630.n6 GNDA 0.295522f
C390 a_5970_4630.t2 GNDA 0.050813f
C391 a_5970_4630.t3 GNDA 0.050813f
C392 a_5970_4630.n7 GNDA 0.144587f
C393 a_5970_4630.n8 GNDA 0.360746f
C394 a_5970_4630.n9 GNDA 0.13437f
C395 a_5970_4630.n10 GNDA 0.085474f
C396 a_5970_4630.n11 GNDA 0.045257f
C397 a_5970_4630.t11 GNDA 0.100208f
C398 V_CONT.n2 GNDA 0.012539f
C399 V_CONT.n5 GNDA 0.010782f
C400 V_CONT.n8 GNDA 0.073739f
C401 V_CONT.t6 GNDA 4.75017f
C402 V_CONT.n9 GNDA 0.038434f
C403 V_CONT.n15 GNDA 0.035035f
C404 opamp_cell_4_0.VIN- GNDA 0.018669f
.ends

