* NGSPICE file created from opamp_6_2.ext - technology: sky130A

**.subckt opamp_6_2
X0 a_2700_n50# VIN+ a_2130_1020# VDDA sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X1 GNDA a_2460_n1410# a_3060_n450# GNDA sky130_fd_pr__nfet_01v8 ad=5 pd=21 as=5 ps=21 w=10 l=0.5
X2 VDDA a_2930_n450# a_2930_n450# VDDA sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X3 a_2700_n50# a_2270_n450# GNDA GNDA sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X4 VOUT a_4140_1090# sky130_fd_pr__cap_mim_m3_1 l=8 w=8
X5 a_3390_n450# VIN- a_3060_n450# GNDA sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X6 a_2700_n50# a_4140_n1660# GNDA sky130_fd_pr__res_xhigh_po_0p35 l=1.01
X7 a_1920_n1410# a_2460_n1410# GNDA sky130_fd_pr__res_xhigh_po_2p85 l=0.66
X8 a_2130_1020# VIN- a_2270_n450# VDDA sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X9 a_3390_n450# a_2930_n450# VDDA VDDA sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X10 VOUT a_4140_n1660# sky130_fd_pr__cap_mim_m3_1 l=8 w=8
X11 a_4140_1090# a_3390_n450# GNDA sky130_fd_pr__res_xhigh_po_0p35 l=1.31
X12 VOUT a_2700_n50# GNDA GNDA sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X13 a_2460_n1410# a_2460_n1410# GNDA GNDA sky130_fd_pr__nfet_01v8 ad=5 pd=21 as=5 ps=21 w=10 l=0.5
X14 VOUT a_3390_n450# VDDA VDDA sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X15 a_3060_n450# VIN+ a_2930_n450# GNDA sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X16 VDDA a_1920_n1410# a_2130_1020# VDDA sky130_fd_pr__pfet_01v8 ad=10 pd=41 as=10 ps=41 w=20 l=0.5
X17 a_1920_n1410# a_1920_n1410# VDDA VDDA sky130_fd_pr__pfet_01v8 ad=10 pd=41 as=10 ps=41 w=20 l=0.5
X18 GNDA a_2270_n450# a_2270_n450# GNDA sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
.ends

