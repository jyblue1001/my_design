magic
tech sky130A
timestamp 1722703054
<< nwell >>
rect -75 335 465 695
<< nmos >>
rect 0 150 15 250
rect 40 150 55 250
rect 105 150 120 250
rect 250 150 265 250
rect 315 150 330 250
rect 380 150 395 250
rect 0 -65 15 35
rect 40 -65 55 35
rect 105 -65 120 35
rect 250 -65 265 35
rect 315 -65 330 35
rect 380 -65 395 35
<< pmos >>
rect 0 575 15 675
rect 65 575 80 675
rect 130 575 145 675
rect 275 575 290 675
rect 315 575 330 675
rect 380 575 395 675
rect 0 360 15 460
rect 65 360 80 460
rect 130 360 145 460
rect 275 360 290 460
rect 315 360 330 460
rect 380 360 395 460
<< ndiff >>
rect -50 235 0 250
rect -50 165 -35 235
rect -15 165 0 235
rect -50 150 0 165
rect 15 150 40 250
rect 55 235 105 250
rect 55 165 70 235
rect 90 165 105 235
rect 55 150 105 165
rect 120 235 170 250
rect 120 165 135 235
rect 155 165 170 235
rect 120 150 170 165
rect 200 235 250 250
rect 200 165 215 235
rect 235 165 250 235
rect 200 150 250 165
rect 265 235 315 250
rect 265 165 280 235
rect 300 165 315 235
rect 265 150 315 165
rect 330 235 380 250
rect 330 165 345 235
rect 365 165 380 235
rect 330 150 380 165
rect 395 235 445 250
rect 395 165 410 235
rect 430 165 445 235
rect 395 150 445 165
rect -50 20 0 35
rect -50 -50 -35 20
rect -15 -50 0 20
rect -50 -65 0 -50
rect 15 -65 40 35
rect 55 20 105 35
rect 55 -50 70 20
rect 90 -50 105 20
rect 55 -65 105 -50
rect 120 20 170 35
rect 120 -50 135 20
rect 155 -50 170 20
rect 120 -65 170 -50
rect 200 20 250 35
rect 200 -50 215 20
rect 235 -50 250 20
rect 200 -65 250 -50
rect 265 20 315 35
rect 265 -50 280 20
rect 300 -50 315 20
rect 265 -65 315 -50
rect 330 20 380 35
rect 330 -50 345 20
rect 365 -50 380 20
rect 330 -65 380 -50
rect 395 20 445 35
rect 395 -50 410 20
rect 430 -50 445 20
rect 395 -65 445 -50
<< pdiff >>
rect -50 660 0 675
rect -50 590 -35 660
rect -15 590 0 660
rect -50 575 0 590
rect 15 660 65 675
rect 15 590 30 660
rect 50 590 65 660
rect 15 575 65 590
rect 80 660 130 675
rect 80 590 95 660
rect 115 590 130 660
rect 80 575 130 590
rect 145 660 195 675
rect 145 590 160 660
rect 180 590 195 660
rect 145 575 195 590
rect 225 660 275 675
rect 225 590 240 660
rect 260 590 275 660
rect 225 575 275 590
rect 290 575 315 675
rect 330 660 380 675
rect 330 590 345 660
rect 365 590 380 660
rect 330 575 380 590
rect 395 660 445 675
rect 395 590 410 660
rect 430 590 445 660
rect 395 575 445 590
rect -50 445 0 460
rect -50 375 -35 445
rect -15 375 0 445
rect -50 360 0 375
rect 15 445 65 460
rect 15 375 30 445
rect 50 375 65 445
rect 15 360 65 375
rect 80 445 130 460
rect 80 375 95 445
rect 115 375 130 445
rect 80 360 130 375
rect 145 445 195 460
rect 145 375 160 445
rect 180 375 195 445
rect 145 360 195 375
rect 225 445 275 460
rect 225 375 240 445
rect 260 375 275 445
rect 225 360 275 375
rect 290 360 315 460
rect 330 445 380 460
rect 330 375 345 445
rect 365 375 380 445
rect 330 360 380 375
rect 395 445 445 460
rect 395 375 410 445
rect 430 375 445 445
rect 395 360 445 375
<< ndiffc >>
rect -35 165 -15 235
rect 70 165 90 235
rect 135 165 155 235
rect 215 165 235 235
rect 280 165 300 235
rect 345 165 365 235
rect 410 165 430 235
rect -35 -50 -15 20
rect 70 -50 90 20
rect 135 -50 155 20
rect 215 -50 235 20
rect 280 -50 300 20
rect 345 -50 365 20
rect 410 -50 430 20
<< pdiffc >>
rect -35 590 -15 660
rect 30 590 50 660
rect 95 590 115 660
rect 160 590 180 660
rect 240 590 260 660
rect 345 590 365 660
rect 410 590 430 660
rect -35 375 -15 445
rect 30 375 50 445
rect 95 375 115 445
rect 160 375 180 445
rect 240 375 260 445
rect 345 375 365 445
rect 410 375 430 445
<< psubdiff >>
rect 200 105 300 120
rect 200 85 215 105
rect 285 85 300 105
rect 200 70 300 85
<< nsubdiff >>
rect -50 525 50 540
rect -50 505 -35 525
rect 35 505 50 525
rect -50 490 50 505
<< psubdiffcont >>
rect 215 85 285 105
<< nsubdiffcont >>
rect -35 505 35 525
<< poly >>
rect 355 720 395 730
rect 355 700 365 720
rect 385 700 395 720
rect 355 690 395 700
rect 0 675 15 690
rect 65 675 80 690
rect 130 675 145 690
rect 275 675 290 690
rect 315 675 330 690
rect 380 675 395 690
rect 0 565 15 575
rect -60 550 15 565
rect 0 460 15 475
rect 65 460 80 575
rect 130 560 145 575
rect 275 560 290 575
rect 105 550 145 560
rect 105 530 115 550
rect 135 530 145 550
rect 105 520 145 530
rect 170 550 290 560
rect 170 530 180 550
rect 200 545 290 550
rect 200 530 210 545
rect 170 520 210 530
rect 170 490 185 520
rect 130 475 185 490
rect 130 460 145 475
rect 275 460 290 475
rect 315 460 330 575
rect 380 560 395 575
rect 420 550 465 565
rect 355 515 395 520
rect 420 515 435 550
rect 355 510 435 515
rect 355 490 365 510
rect 385 500 435 510
rect 385 490 395 500
rect 355 480 395 490
rect 380 460 395 480
rect 0 305 15 360
rect 65 350 80 360
rect 130 350 145 360
rect -25 295 15 305
rect -25 275 -15 295
rect 5 275 15 295
rect -25 265 15 275
rect 0 250 15 265
rect 40 335 80 350
rect 105 335 145 350
rect 275 345 290 360
rect 250 335 290 345
rect 40 250 55 335
rect 105 250 120 335
rect 250 315 260 335
rect 280 315 290 335
rect 250 305 290 315
rect 250 250 265 305
rect 315 250 330 360
rect 380 250 395 360
rect 0 135 15 150
rect -60 45 15 60
rect 0 35 15 45
rect 40 35 55 150
rect 105 135 120 150
rect 250 135 265 150
rect 80 125 120 135
rect 80 105 90 125
rect 110 110 120 125
rect 110 105 160 110
rect 80 95 160 105
rect 145 60 160 95
rect 105 35 120 50
rect 145 45 265 60
rect 250 35 265 45
rect 315 35 330 150
rect 380 140 395 150
rect 380 125 435 140
rect 355 80 395 90
rect 355 60 365 80
rect 385 60 395 80
rect 355 50 395 60
rect 380 35 395 50
rect 420 85 435 125
rect 420 75 460 85
rect 420 55 430 75
rect 450 60 460 75
rect 450 55 465 60
rect 420 45 465 55
rect 0 -80 15 -65
rect 40 -120 55 -65
rect 105 -80 120 -65
rect 250 -80 265 -65
rect 80 -90 120 -80
rect 80 -110 90 -90
rect 110 -110 120 -90
rect 80 -120 120 -110
rect 315 -120 330 -65
rect 380 -80 395 -65
rect 15 -130 55 -120
rect 15 -150 25 -130
rect 45 -150 55 -130
rect 15 -160 55 -150
rect 290 -130 330 -120
rect 290 -150 300 -130
rect 320 -150 330 -130
rect 290 -160 330 -150
<< polycont >>
rect 365 700 385 720
rect 115 530 135 550
rect 180 530 200 550
rect 365 490 385 510
rect -15 275 5 295
rect 260 315 280 335
rect 90 105 110 125
rect 365 60 385 80
rect 430 55 450 75
rect 90 -110 110 -90
rect 25 -150 45 -130
rect 300 -150 320 -130
<< locali >>
rect 355 720 395 730
rect 355 710 365 720
rect -25 690 105 710
rect -25 670 -5 690
rect 85 670 105 690
rect 295 700 365 710
rect 385 700 395 720
rect 295 690 395 700
rect -45 660 -5 670
rect -45 590 -35 660
rect -15 590 -5 660
rect -45 580 -5 590
rect 20 660 60 670
rect 20 590 30 660
rect 50 590 60 660
rect 20 580 60 590
rect 85 660 125 670
rect 85 590 95 660
rect 115 590 125 660
rect 85 580 125 590
rect 150 660 190 670
rect 150 590 160 660
rect 180 590 190 660
rect 150 580 190 590
rect 20 535 40 580
rect 170 560 190 580
rect 230 660 270 670
rect 230 590 240 660
rect 260 590 270 660
rect 230 580 270 590
rect 105 550 145 560
rect -45 525 45 535
rect -45 505 -35 525
rect 35 505 45 525
rect 105 530 115 550
rect 135 530 145 550
rect 105 520 145 530
rect 170 550 210 560
rect 170 530 180 550
rect 200 530 210 550
rect 170 520 210 530
rect -45 495 45 505
rect 125 500 145 520
rect 20 455 40 495
rect 125 480 170 500
rect 150 455 170 480
rect 230 455 250 580
rect 295 455 315 690
rect 335 660 375 670
rect 335 590 345 660
rect 365 590 375 660
rect 335 580 375 590
rect 400 660 440 670
rect 400 590 410 660
rect 430 590 440 660
rect 400 580 440 590
rect 355 520 375 580
rect 355 510 395 520
rect 355 490 365 510
rect 385 490 395 510
rect 355 480 395 490
rect 420 455 440 580
rect -45 445 -5 455
rect -45 375 -35 445
rect -15 375 -5 445
rect -45 365 -5 375
rect 20 445 60 455
rect 20 375 30 445
rect 50 375 60 445
rect 20 365 60 375
rect 85 445 125 455
rect 85 375 95 445
rect 115 375 125 445
rect 85 365 125 375
rect 150 445 190 455
rect 150 375 160 445
rect 180 375 190 445
rect 150 365 190 375
rect 230 445 270 455
rect 230 375 240 445
rect 260 375 270 445
rect 295 445 375 455
rect 295 435 345 445
rect 230 365 270 375
rect 335 375 345 435
rect 365 375 375 445
rect 335 365 375 375
rect 400 445 440 455
rect 400 375 410 445
rect 430 375 440 445
rect 400 365 440 375
rect -25 345 -5 365
rect 85 345 105 365
rect -25 325 105 345
rect 150 345 170 365
rect 355 345 375 365
rect 150 335 290 345
rect 150 325 260 335
rect -25 295 15 305
rect -25 285 -15 295
rect -50 275 -15 285
rect 5 275 15 295
rect 150 285 170 325
rect 250 315 260 325
rect 280 315 290 335
rect 355 325 440 345
rect 250 305 290 315
rect 420 285 440 325
rect -50 265 15 275
rect 80 265 170 285
rect 225 265 355 285
rect 80 245 100 265
rect 225 245 245 265
rect 335 245 355 265
rect 420 265 465 285
rect 420 245 440 265
rect -45 235 -5 245
rect -45 165 -35 235
rect -15 165 -5 235
rect 60 235 100 245
rect 60 175 70 235
rect -45 155 -5 165
rect 20 165 70 175
rect 90 165 100 235
rect 20 155 100 165
rect 125 235 165 245
rect 125 165 135 235
rect 155 165 165 235
rect 125 155 165 165
rect 205 235 245 245
rect 205 165 215 235
rect 235 165 245 235
rect 205 155 245 165
rect 270 235 310 245
rect 270 165 280 235
rect 300 165 310 235
rect 270 155 310 165
rect 335 235 375 245
rect 335 165 345 235
rect 365 165 375 235
rect 335 155 375 165
rect 400 235 440 245
rect 400 165 410 235
rect 430 165 440 235
rect 400 155 440 165
rect -45 30 -25 155
rect -45 20 -5 30
rect -45 -50 -35 20
rect -15 -50 -5 20
rect -45 -60 -5 -50
rect 20 -80 40 155
rect 80 125 120 135
rect 80 105 90 125
rect 110 105 120 125
rect 80 95 120 105
rect 80 30 100 95
rect 145 30 165 155
rect 270 115 290 155
rect 400 135 420 155
rect 375 115 420 135
rect 205 105 295 115
rect 205 85 215 105
rect 285 85 295 105
rect 375 90 395 115
rect 205 75 295 85
rect 355 80 395 90
rect 270 30 290 75
rect 355 60 365 80
rect 385 60 395 80
rect 355 50 395 60
rect 420 75 460 85
rect 420 55 430 75
rect 450 55 460 75
rect 420 45 460 55
rect 420 30 440 45
rect 60 20 100 30
rect 60 -50 70 20
rect 90 -50 100 20
rect 60 -60 100 -50
rect 125 20 165 30
rect 125 -50 135 20
rect 155 -50 165 20
rect 125 -60 165 -50
rect 205 20 245 30
rect 205 -50 215 20
rect 235 -50 245 20
rect 205 -60 245 -50
rect 270 20 310 30
rect 270 -50 280 20
rect 300 -50 310 20
rect 270 -60 310 -50
rect 335 20 375 30
rect 335 -50 345 20
rect 365 -50 375 20
rect 335 -60 375 -50
rect 400 20 440 30
rect 400 -50 410 20
rect 430 -50 440 20
rect 400 -60 440 -50
rect 225 -80 245 -60
rect 335 -80 355 -60
rect 20 -90 120 -80
rect 20 -100 90 -90
rect 80 -110 90 -100
rect 110 -110 120 -90
rect 225 -100 355 -80
rect 80 -120 120 -110
rect 15 -130 55 -120
rect 15 -150 25 -130
rect 45 -150 55 -130
rect 15 -160 55 -150
rect 290 -130 330 -120
rect 290 -150 300 -130
rect 320 -150 330 -130
rect 290 -160 330 -150
<< viali >>
rect 30 590 50 660
rect 240 590 260 660
rect -35 505 35 525
rect 410 590 430 660
rect 30 375 50 445
rect 240 375 260 445
rect 410 375 430 445
rect -35 165 -15 235
rect 135 165 155 235
rect 280 165 300 235
rect -35 -50 -15 20
rect 215 85 285 105
rect 135 -50 155 20
rect 280 -50 300 20
rect 25 -150 45 -130
rect 300 -150 320 -130
<< metal1 >>
rect -60 660 465 675
rect -60 590 30 660
rect 50 590 240 660
rect 260 590 410 660
rect 430 590 465 660
rect -60 525 465 590
rect -60 505 -35 525
rect 35 505 465 525
rect -60 445 465 505
rect -60 375 30 445
rect 50 375 240 445
rect 260 375 410 445
rect 430 375 465 445
rect -60 360 465 375
rect -60 235 465 250
rect -60 165 -35 235
rect -15 165 135 235
rect 155 165 280 235
rect 300 165 465 235
rect -60 105 465 165
rect -60 85 215 105
rect 285 85 465 105
rect -60 20 465 85
rect -60 -50 -35 20
rect -15 -50 135 20
rect 155 -50 280 20
rect 300 -50 465 20
rect -60 -65 465 -50
rect -60 -130 465 -120
rect -60 -150 25 -130
rect 45 -150 300 -130
rect 320 -150 465 -130
rect -60 -160 465 -150
<< labels >>
flabel poly -60 50 -60 50 7 FreeSans 80 0 -40 0 Dn2
flabel metal1 -60 95 -60 95 7 FreeSans 80 0 -80 0 VN
flabel metal1 -60 -140 -60 -140 7 FreeSans 80 0 -80 0 CLK
flabel poly -60 555 -60 555 7 FreeSans 80 0 -40 0 Dn1
flabel locali -50 275 -50 275 7 FreeSans 80 0 -40 0 D
flabel metal1 -60 515 -60 515 7 FreeSans 80 0 -40 0 VP
flabel locali 465 275 465 275 3 FreeSans 80 0 40 0 Q
flabel poly 465 555 465 555 3 FreeSans 80 0 40 0 Qb1
<< end >>
