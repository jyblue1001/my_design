magic
tech sky130A
timestamp 1753628751
<< metal1 >>
rect 2320 15410 2380 15425
rect 2320 15380 2335 15410
rect 2365 15380 2380 15410
rect 2320 15345 2380 15380
rect 2320 15315 2335 15345
rect 2365 15315 2380 15345
rect 2320 15275 2380 15315
rect 2320 15245 2335 15275
rect 2365 15245 2380 15275
rect 2320 15205 2380 15245
rect 2320 15175 2335 15205
rect 2365 15175 2380 15205
rect 2320 15135 2380 15175
rect 2320 15105 2335 15135
rect 2365 15105 2380 15135
rect 2320 15070 2380 15105
rect 2320 15040 2335 15070
rect 2365 15040 2380 15070
rect 2320 15025 2380 15040
rect 6690 15410 6750 15425
rect 6690 15380 6705 15410
rect 6735 15380 6750 15410
rect 6690 15345 6750 15380
rect 6690 15315 6705 15345
rect 6735 15315 6750 15345
rect 6690 15275 6750 15315
rect 6690 15245 6705 15275
rect 6735 15245 6750 15275
rect 6690 15205 6750 15245
rect 6690 15175 6705 15205
rect 6735 15175 6750 15205
rect 6690 15135 6750 15175
rect 6690 15105 6705 15135
rect 6735 15105 6750 15135
rect 6690 15070 6750 15105
rect 6690 15040 6705 15070
rect 6735 15040 6750 15070
rect 6690 15025 6750 15040
rect 2330 13080 2370 15025
rect 2330 13050 2335 13080
rect 2365 13050 2370 13080
rect 2330 9895 2370 13050
rect 2330 9865 2335 9895
rect 2365 9865 2370 9895
rect 2330 9660 2370 9865
rect 2330 9630 2335 9660
rect 2365 9630 2370 9660
rect 2330 9625 2370 9630
rect 2385 13225 2425 13230
rect 2385 13195 2390 13225
rect 2420 13195 2425 13225
rect 2385 6950 2425 13195
rect 6700 13005 6740 15025
rect 6700 12975 6705 13005
rect 6735 12975 6740 13005
rect 6700 10085 6740 12975
rect 6700 10055 6705 10085
rect 6735 10055 6740 10085
rect 6700 10050 6740 10055
rect 6590 9345 6630 9350
rect 6590 9315 6595 9345
rect 6625 9315 6630 9345
rect 6300 8630 6340 8635
rect 6300 8600 6305 8630
rect 6335 8600 6340 8630
rect 2375 6935 2435 6950
rect 2375 6905 2390 6935
rect 2420 6905 2435 6935
rect 2375 6870 2435 6905
rect 2375 6840 2390 6870
rect 2420 6840 2435 6870
rect 2375 6800 2435 6840
rect 2375 6770 2390 6800
rect 2420 6770 2435 6800
rect 2375 6730 2435 6770
rect 2375 6700 2390 6730
rect 2420 6700 2435 6730
rect 2375 6660 2435 6700
rect 2375 6630 2390 6660
rect 2420 6630 2435 6660
rect 2375 6595 2435 6630
rect 2375 6565 2390 6595
rect 2420 6565 2435 6595
rect 2375 6550 2435 6565
rect 2485 6390 2505 7190
rect 2395 6385 2435 6390
rect 2395 6355 2400 6385
rect 2430 6355 2435 6385
rect 2395 6350 2435 6355
rect 2475 6385 2515 6390
rect 2475 6355 2480 6385
rect 2510 6355 2515 6385
rect 2475 6350 2515 6355
rect 2350 6280 2390 6285
rect 2350 6250 2355 6280
rect 2385 6250 2390 6280
rect 2350 6245 2390 6250
rect 2360 2410 2380 6245
rect 2350 2405 2390 2410
rect 2350 2375 2355 2405
rect 2385 2375 2390 2405
rect 2350 2370 2390 2375
rect 2405 2205 2425 6350
rect 2725 6225 2745 7185
rect 2855 6350 2875 7185
rect 2845 6345 2885 6350
rect 2845 6315 2850 6345
rect 2880 6315 2885 6345
rect 2845 6310 2885 6315
rect 2715 6220 2755 6225
rect 2715 6190 2720 6220
rect 2750 6190 2755 6220
rect 2715 6185 2755 6190
rect 3000 6180 3020 7190
rect 3240 6950 3280 7970
rect 3230 6935 3290 6950
rect 3230 6905 3245 6935
rect 3275 6905 3290 6935
rect 3230 6870 3290 6905
rect 3230 6840 3245 6870
rect 3275 6840 3290 6870
rect 3230 6800 3290 6840
rect 3230 6770 3245 6800
rect 3275 6770 3290 6800
rect 3230 6730 3290 6770
rect 3230 6700 3245 6730
rect 3275 6700 3290 6730
rect 3230 6660 3290 6700
rect 3230 6630 3245 6660
rect 3275 6630 3290 6660
rect 3230 6595 3290 6630
rect 3230 6565 3245 6595
rect 3275 6565 3290 6595
rect 3230 6550 3290 6565
rect 3400 6345 3440 6350
rect 3400 6315 3405 6345
rect 3435 6315 3440 6345
rect 3400 6310 3440 6315
rect 2990 6175 3030 6180
rect 2990 6145 2995 6175
rect 3025 6145 3030 6175
rect 2990 6140 3030 6145
rect 3410 3060 3430 6310
rect 3785 6285 3805 7190
rect 4470 6950 4510 7505
rect 4465 6935 4515 6950
rect 4465 6905 4475 6935
rect 4505 6905 4515 6935
rect 4465 6870 4515 6905
rect 4465 6840 4475 6870
rect 4505 6840 4515 6870
rect 4465 6800 4515 6840
rect 4465 6770 4475 6800
rect 4505 6770 4515 6800
rect 4465 6730 4515 6770
rect 4465 6700 4475 6730
rect 4505 6700 4515 6730
rect 4465 6660 4515 6700
rect 4465 6630 4475 6660
rect 4505 6630 4515 6660
rect 4465 6595 4515 6630
rect 4465 6565 4475 6595
rect 4505 6565 4515 6595
rect 4465 6550 4515 6565
rect 4480 6355 4500 6550
rect 3775 6280 3815 6285
rect 3775 6250 3780 6280
rect 3810 6250 3815 6280
rect 3775 6245 3815 6250
rect 3450 6175 3490 6180
rect 3450 6145 3455 6175
rect 3485 6145 3490 6175
rect 3450 6140 3490 6145
rect 3400 3055 3440 3060
rect 3400 3025 3405 3055
rect 3435 3025 3440 3055
rect 3400 3020 3440 3025
rect 3460 2530 3480 6140
rect 4530 5165 4550 7190
rect 5175 6285 5195 7190
rect 6155 6390 6175 7190
rect 5490 6385 5530 6390
rect 5490 6355 5495 6385
rect 5525 6355 5530 6385
rect 5490 6350 5530 6355
rect 6145 6385 6185 6390
rect 6145 6355 6150 6385
rect 6180 6355 6185 6385
rect 6145 6350 6185 6355
rect 5165 6280 5205 6285
rect 5165 6250 5170 6280
rect 5200 6250 5205 6280
rect 5165 6245 5205 6250
rect 4820 6220 4860 6225
rect 4820 6190 4825 6220
rect 4855 6190 4860 6220
rect 4820 6185 4860 6190
rect 4520 5160 4560 5165
rect 4520 5130 4525 5160
rect 4555 5130 4560 5160
rect 4520 5125 4560 5130
rect 4830 5120 4850 6185
rect 4820 5115 4860 5120
rect 4820 5085 4825 5115
rect 4855 5085 4860 5115
rect 4820 5080 4860 5085
rect 4940 5115 4980 5120
rect 4940 5085 4945 5115
rect 4975 5085 4980 5115
rect 4940 5080 4980 5085
rect 4950 4505 4970 5080
rect 5166 4555 5196 4560
rect 5166 4520 5196 4525
rect 4940 4500 4980 4505
rect 4940 4470 4945 4500
rect 4975 4470 4980 4500
rect 4940 4465 4980 4470
rect 5500 3340 5520 6350
rect 5545 5160 5585 5165
rect 5545 5130 5550 5160
rect 5580 5130 5585 5160
rect 6230 5140 6250 7190
rect 6300 6950 6340 8600
rect 6290 6935 6350 6950
rect 6290 6905 6305 6935
rect 6335 6905 6350 6935
rect 6290 6870 6350 6905
rect 6290 6840 6305 6870
rect 6335 6840 6350 6870
rect 6290 6800 6350 6840
rect 6290 6770 6305 6800
rect 6335 6770 6350 6800
rect 6290 6730 6350 6770
rect 6290 6700 6305 6730
rect 6335 6700 6350 6730
rect 6290 6660 6350 6700
rect 6290 6630 6305 6660
rect 6335 6630 6350 6660
rect 6290 6595 6350 6630
rect 6290 6565 6305 6595
rect 6335 6565 6350 6595
rect 6290 6550 6350 6565
rect 6475 6390 6495 7190
rect 6590 6950 6630 9315
rect 6580 6935 6640 6950
rect 6580 6905 6595 6935
rect 6625 6905 6640 6935
rect 6580 6870 6640 6905
rect 6580 6840 6595 6870
rect 6625 6840 6640 6870
rect 6580 6800 6640 6840
rect 6580 6770 6595 6800
rect 6625 6770 6640 6800
rect 6580 6730 6640 6770
rect 6580 6700 6595 6730
rect 6625 6700 6640 6730
rect 6580 6660 6640 6700
rect 6580 6630 6595 6660
rect 6625 6630 6640 6660
rect 6580 6595 6640 6630
rect 6580 6565 6595 6595
rect 6625 6565 6640 6595
rect 6580 6550 6640 6565
rect 6465 6385 6505 6390
rect 6465 6355 6470 6385
rect 6500 6355 6505 6385
rect 6465 6350 6505 6355
rect 6545 6385 6585 6390
rect 6545 6355 6550 6385
rect 6580 6355 6585 6385
rect 6545 6350 6585 6355
rect 5545 5125 5585 5130
rect 5870 5135 5910 5140
rect 5490 3335 5530 3340
rect 4415 3330 4455 3335
rect 4415 3300 4420 3330
rect 4450 3300 4455 3330
rect 5490 3305 5495 3335
rect 5525 3305 5530 3335
rect 5490 3300 5530 3305
rect 4415 3295 4455 3300
rect 5555 2605 5575 5125
rect 5870 5105 5875 5135
rect 5905 5105 5910 5135
rect 5870 5100 5910 5105
rect 6220 5135 6260 5140
rect 6220 5105 6225 5135
rect 6255 5105 6260 5135
rect 6220 5100 6260 5105
rect 5880 4570 5900 5100
rect 5870 4565 5910 4570
rect 5870 4535 5875 4565
rect 5905 4535 5910 4565
rect 5870 4530 5910 4535
rect 4530 2600 4570 2605
rect 4530 2570 4535 2600
rect 4565 2570 4570 2600
rect 4530 2565 4570 2570
rect 5545 2600 5585 2605
rect 5545 2570 5550 2600
rect 5580 2570 5585 2600
rect 5545 2565 5585 2570
rect 3420 2525 3480 2530
rect 3420 2495 3425 2525
rect 3455 2495 3480 2525
rect 3420 2490 3480 2495
rect 2395 2200 2435 2205
rect 2395 2170 2400 2200
rect 2430 2170 2435 2200
rect 2395 2165 2435 2170
rect 4540 2110 4560 2565
rect 6555 2205 6575 6350
rect 6590 6280 6630 6285
rect 6590 6250 6595 6280
rect 6625 6250 6630 6280
rect 6590 6245 6630 6250
rect 6600 2410 6620 6245
rect 6590 2405 6630 2410
rect 6590 2375 6595 2405
rect 6625 2375 6630 2405
rect 6590 2370 6630 2375
rect 6545 2200 6585 2205
rect 6545 2170 6550 2200
rect 6580 2170 6585 2200
rect 6545 2165 6585 2170
rect 4460 -215 4520 -200
rect 4460 -245 4475 -215
rect 4505 -245 4520 -215
rect 4460 -280 4520 -245
rect 4460 -310 4475 -280
rect 4505 -310 4520 -280
rect 4460 -350 4520 -310
rect 4460 -380 4475 -350
rect 4505 -380 4520 -350
rect 4460 -420 4520 -380
rect 4460 -450 4475 -420
rect 4505 -450 4520 -420
rect 4460 -490 4520 -450
rect 4460 -520 4475 -490
rect 4505 -520 4520 -490
rect 4460 -555 4520 -520
rect 4460 -585 4475 -555
rect 4505 -585 4520 -555
rect 4460 -600 4520 -585
<< via1 >>
rect 2335 15380 2365 15410
rect 2335 15315 2365 15345
rect 2335 15245 2365 15275
rect 2335 15175 2365 15205
rect 2335 15105 2365 15135
rect 2335 15040 2365 15070
rect 6705 15380 6735 15410
rect 6705 15315 6735 15345
rect 6705 15245 6735 15275
rect 6705 15175 6735 15205
rect 6705 15105 6735 15135
rect 6705 15040 6735 15070
rect 2335 13050 2365 13080
rect 2335 9865 2365 9895
rect 2335 9630 2365 9660
rect 2390 13195 2420 13225
rect 6705 12975 6735 13005
rect 6705 10055 6735 10085
rect 6595 9315 6625 9345
rect 6305 8600 6335 8630
rect 2390 6905 2420 6935
rect 2390 6840 2420 6870
rect 2390 6770 2420 6800
rect 2390 6700 2420 6730
rect 2390 6630 2420 6660
rect 2390 6565 2420 6595
rect 2400 6355 2430 6385
rect 2480 6355 2510 6385
rect 2355 6250 2385 6280
rect 2355 2375 2385 2405
rect 2850 6315 2880 6345
rect 2720 6190 2750 6220
rect 3245 6905 3275 6935
rect 3245 6840 3275 6870
rect 3245 6770 3275 6800
rect 3245 6700 3275 6730
rect 3245 6630 3275 6660
rect 3245 6565 3275 6595
rect 3405 6315 3435 6345
rect 2995 6145 3025 6175
rect 4475 6905 4505 6935
rect 4475 6840 4505 6870
rect 4475 6770 4505 6800
rect 4475 6700 4505 6730
rect 4475 6630 4505 6660
rect 4475 6565 4505 6595
rect 3780 6250 3810 6280
rect 3455 6145 3485 6175
rect 3405 3025 3435 3055
rect 5495 6355 5525 6385
rect 6150 6355 6180 6385
rect 5170 6250 5200 6280
rect 4825 6190 4855 6220
rect 4525 5130 4555 5160
rect 4825 5085 4855 5115
rect 4945 5085 4975 5115
rect 5166 4525 5196 4555
rect 4945 4470 4975 4500
rect 5550 5130 5580 5160
rect 6305 6905 6335 6935
rect 6305 6840 6335 6870
rect 6305 6770 6335 6800
rect 6305 6700 6335 6730
rect 6305 6630 6335 6660
rect 6305 6565 6335 6595
rect 6595 6905 6625 6935
rect 6595 6840 6625 6870
rect 6595 6770 6625 6800
rect 6595 6700 6625 6730
rect 6595 6630 6625 6660
rect 6595 6565 6625 6595
rect 6470 6355 6500 6385
rect 6550 6355 6580 6385
rect 4420 3300 4450 3330
rect 5495 3305 5525 3335
rect 5875 5105 5905 5135
rect 6225 5105 6255 5135
rect 5875 4535 5905 4565
rect 4535 2570 4565 2600
rect 5550 2570 5580 2600
rect 3425 2495 3455 2525
rect 2400 2170 2430 2200
rect 6595 6250 6625 6280
rect 6595 2375 6625 2405
rect 6550 2170 6580 2200
rect 4475 -245 4505 -215
rect 4475 -310 4505 -280
rect 4475 -380 4505 -350
rect 4475 -450 4505 -420
rect 4475 -520 4505 -490
rect 4475 -585 4505 -555
<< metal2 >>
rect 2320 15410 2380 15425
rect 2320 15380 2335 15410
rect 2365 15380 2380 15410
rect 2320 15345 2380 15380
rect 2320 15315 2335 15345
rect 2365 15315 2380 15345
rect 2320 15275 2380 15315
rect 2320 15245 2335 15275
rect 2365 15245 2380 15275
rect 2320 15205 2380 15245
rect 2320 15175 2335 15205
rect 2365 15175 2380 15205
rect 2320 15135 2380 15175
rect 2320 15105 2335 15135
rect 2365 15105 2380 15135
rect 2320 15070 2380 15105
rect 2320 15040 2335 15070
rect 2365 15040 2380 15070
rect 2320 15025 2380 15040
rect 6690 15410 6750 15425
rect 6690 15380 6705 15410
rect 6735 15380 6750 15410
rect 6690 15345 6750 15380
rect 6690 15315 6705 15345
rect 6735 15315 6750 15345
rect 6690 15275 6750 15315
rect 6690 15245 6705 15275
rect 6735 15245 6750 15275
rect 6690 15205 6750 15245
rect 6690 15175 6705 15205
rect 6735 15175 6750 15205
rect 6690 15135 6750 15175
rect 6690 15105 6705 15135
rect 6735 15105 6750 15135
rect 6690 15070 6750 15105
rect 6690 15040 6705 15070
rect 6735 15040 6750 15070
rect 6690 15025 6750 15040
rect 2385 13225 2425 13230
rect 2385 13195 2390 13225
rect 2420 13195 2425 13225
rect 2385 13190 2425 13195
rect 2330 13080 2370 13085
rect 2330 13050 2335 13080
rect 2365 13075 2370 13080
rect 2365 13055 2970 13075
rect 2365 13050 2370 13055
rect 2330 13045 2370 13050
rect 6700 13005 6740 13010
rect 6700 13000 6705 13005
rect 6625 12980 6705 13000
rect 6700 12975 6705 12980
rect 6735 12975 6740 13005
rect 6700 12970 6740 12975
rect 6700 10085 6740 10090
rect 6700 10080 6705 10085
rect 5400 10060 6705 10080
rect 6700 10055 6705 10060
rect 6735 10055 6740 10085
rect 6700 10050 6740 10055
rect 2330 9895 2370 9900
rect 2330 9865 2335 9895
rect 2365 9890 2370 9895
rect 2365 9870 3355 9890
rect 2365 9865 2370 9870
rect 2330 9860 2370 9865
rect 2330 9660 2370 9665
rect 2330 9630 2335 9660
rect 2365 9655 2370 9660
rect 2365 9635 3800 9655
rect 2365 9630 2370 9635
rect 2330 9625 2370 9630
rect 6590 9345 6630 9350
rect 6590 9340 6595 9345
rect 5670 9320 6595 9340
rect 6590 9315 6595 9320
rect 6625 9315 6630 9345
rect 6590 9310 6630 9315
rect 6300 8630 6340 8635
rect 6300 8625 6305 8630
rect 5870 8605 6305 8625
rect 6300 8600 6305 8605
rect 6335 8600 6340 8630
rect 6300 8595 6340 8600
rect 2375 6935 2435 6950
rect 2375 6905 2390 6935
rect 2420 6905 2435 6935
rect 2375 6870 2435 6905
rect 2375 6840 2390 6870
rect 2420 6840 2435 6870
rect 2375 6800 2435 6840
rect 2375 6770 2390 6800
rect 2420 6770 2435 6800
rect 2375 6730 2435 6770
rect 2375 6700 2390 6730
rect 2420 6700 2435 6730
rect 2375 6660 2435 6700
rect 2375 6630 2390 6660
rect 2420 6630 2435 6660
rect 2375 6595 2435 6630
rect 2375 6565 2390 6595
rect 2420 6565 2435 6595
rect 2375 6550 2435 6565
rect 3230 6935 3290 6950
rect 3230 6905 3245 6935
rect 3275 6905 3290 6935
rect 3230 6870 3290 6905
rect 3230 6840 3245 6870
rect 3275 6840 3290 6870
rect 3230 6800 3290 6840
rect 3230 6770 3245 6800
rect 3275 6770 3290 6800
rect 3230 6730 3290 6770
rect 3230 6700 3245 6730
rect 3275 6700 3290 6730
rect 3230 6660 3290 6700
rect 3230 6630 3245 6660
rect 3275 6630 3290 6660
rect 3230 6595 3290 6630
rect 3230 6565 3245 6595
rect 3275 6565 3290 6595
rect 3230 6550 3290 6565
rect 4465 6935 4515 6950
rect 4465 6905 4475 6935
rect 4505 6905 4515 6935
rect 4465 6870 4515 6905
rect 4465 6840 4475 6870
rect 4505 6840 4515 6870
rect 4465 6800 4515 6840
rect 4465 6770 4475 6800
rect 4505 6770 4515 6800
rect 4465 6730 4515 6770
rect 4465 6700 4475 6730
rect 4505 6700 4515 6730
rect 4465 6660 4515 6700
rect 4465 6630 4475 6660
rect 4505 6630 4515 6660
rect 4465 6595 4515 6630
rect 4465 6565 4475 6595
rect 4505 6565 4515 6595
rect 4465 6550 4515 6565
rect 6290 6935 6350 6950
rect 6290 6905 6305 6935
rect 6335 6905 6350 6935
rect 6290 6870 6350 6905
rect 6290 6840 6305 6870
rect 6335 6840 6350 6870
rect 6290 6800 6350 6840
rect 6290 6770 6305 6800
rect 6335 6770 6350 6800
rect 6290 6730 6350 6770
rect 6290 6700 6305 6730
rect 6335 6700 6350 6730
rect 6290 6660 6350 6700
rect 6290 6630 6305 6660
rect 6335 6630 6350 6660
rect 6290 6595 6350 6630
rect 6290 6565 6305 6595
rect 6335 6565 6350 6595
rect 6290 6550 6350 6565
rect 6580 6935 6640 6950
rect 6580 6905 6595 6935
rect 6625 6905 6640 6935
rect 6580 6870 6640 6905
rect 6580 6840 6595 6870
rect 6625 6840 6640 6870
rect 6580 6800 6640 6840
rect 6580 6770 6595 6800
rect 6625 6770 6640 6800
rect 6580 6730 6640 6770
rect 6580 6700 6595 6730
rect 6625 6700 6640 6730
rect 6580 6660 6640 6700
rect 6580 6630 6595 6660
rect 6625 6630 6640 6660
rect 6580 6595 6640 6630
rect 6580 6565 6595 6595
rect 6625 6565 6640 6595
rect 6580 6550 6640 6565
rect 2395 6385 2435 6390
rect 2395 6355 2400 6385
rect 2430 6380 2435 6385
rect 2475 6385 2515 6390
rect 2475 6380 2480 6385
rect 2430 6360 2480 6380
rect 2430 6355 2435 6360
rect 2395 6350 2435 6355
rect 2475 6355 2480 6360
rect 2510 6355 2515 6385
rect 2475 6350 2515 6355
rect 5490 6385 5530 6390
rect 5490 6355 5495 6385
rect 5525 6380 5530 6385
rect 6145 6385 6185 6390
rect 6145 6380 6150 6385
rect 5525 6360 6150 6380
rect 5525 6355 5530 6360
rect 5490 6350 5530 6355
rect 6145 6355 6150 6360
rect 6180 6355 6185 6385
rect 6465 6385 6505 6390
rect 6465 6380 6470 6385
rect 6455 6360 6470 6380
rect 6145 6350 6185 6355
rect 6465 6355 6470 6360
rect 6500 6380 6505 6385
rect 6545 6385 6585 6390
rect 6545 6380 6550 6385
rect 6500 6360 6550 6380
rect 6500 6355 6505 6360
rect 6465 6350 6505 6355
rect 6545 6355 6550 6360
rect 6580 6355 6585 6385
rect 6545 6350 6585 6355
rect 2845 6345 2885 6350
rect 2845 6315 2850 6345
rect 2880 6340 2885 6345
rect 3400 6345 3440 6350
rect 3400 6340 3405 6345
rect 2880 6320 3405 6340
rect 2880 6315 2885 6320
rect 2845 6310 2885 6315
rect 3400 6315 3405 6320
rect 3435 6315 3440 6345
rect 3400 6310 3440 6315
rect 2350 6280 2390 6285
rect 2350 6250 2355 6280
rect 2385 6275 2390 6280
rect 3775 6280 3815 6285
rect 3775 6275 3780 6280
rect 2385 6255 3780 6275
rect 2385 6250 2390 6255
rect 2350 6245 2390 6250
rect 3775 6250 3780 6255
rect 3810 6250 3815 6280
rect 3775 6245 3815 6250
rect 5165 6280 5205 6285
rect 5165 6250 5170 6280
rect 5200 6275 5205 6280
rect 6590 6280 6630 6285
rect 6590 6275 6595 6280
rect 5200 6255 6595 6275
rect 5200 6250 5205 6255
rect 5165 6245 5205 6250
rect 6590 6250 6595 6255
rect 6625 6250 6630 6280
rect 6590 6245 6630 6250
rect 2715 6220 2755 6225
rect 2715 6190 2720 6220
rect 2750 6215 2755 6220
rect 4820 6220 4860 6225
rect 4820 6215 4825 6220
rect 2750 6195 4825 6215
rect 2750 6190 2755 6195
rect 2715 6185 2755 6190
rect 4820 6190 4825 6195
rect 4855 6190 4860 6220
rect 4820 6185 4860 6190
rect 2990 6175 3030 6180
rect 2990 6145 2995 6175
rect 3025 6170 3030 6175
rect 3450 6175 3490 6180
rect 3450 6170 3455 6175
rect 3025 6150 3455 6170
rect 3025 6145 3030 6150
rect 2990 6140 3030 6145
rect 3450 6145 3455 6150
rect 3485 6145 3490 6175
rect 3450 6140 3490 6145
rect 4520 5160 4560 5165
rect 4520 5130 4525 5160
rect 4555 5155 4560 5160
rect 5545 5160 5585 5165
rect 5545 5155 5550 5160
rect 4555 5135 5550 5155
rect 4555 5130 4560 5135
rect 4520 5125 4560 5130
rect 5545 5130 5550 5135
rect 5580 5130 5585 5160
rect 5545 5125 5585 5130
rect 5870 5135 5910 5140
rect 4820 5115 4860 5120
rect 4940 5115 4980 5120
rect 4820 5085 4825 5115
rect 4855 5090 4945 5115
rect 4855 5085 4860 5090
rect 4820 5080 4860 5085
rect 4940 5085 4945 5090
rect 4975 5085 4980 5115
rect 5870 5105 5875 5135
rect 5905 5130 5910 5135
rect 6220 5135 6260 5140
rect 6220 5130 6225 5135
rect 5905 5110 6225 5130
rect 5905 5105 5910 5110
rect 5870 5100 5910 5105
rect 6220 5105 6225 5110
rect 6255 5105 6260 5135
rect 6220 5100 6260 5105
rect 4940 5080 4980 5085
rect 5870 4565 5910 4570
rect 5870 4560 5875 4565
rect 4515 4555 5875 4560
rect 4515 4540 5166 4555
rect 5196 4540 5875 4555
rect 5870 4535 5875 4540
rect 5905 4535 5910 4565
rect 5870 4530 5910 4535
rect 5166 4520 5196 4525
rect 4940 4500 4980 4505
rect 4940 4470 4945 4500
rect 4975 4470 4980 4500
rect 4940 4465 4980 4470
rect 4515 4430 5595 4450
rect 5490 3335 5530 3340
rect 4415 3330 4455 3335
rect 4415 3300 4420 3330
rect 4450 3325 4455 3330
rect 5490 3325 5495 3335
rect 4450 3305 5495 3325
rect 5525 3305 5530 3335
rect 4450 3300 4455 3305
rect 5490 3300 5530 3305
rect 4415 3295 4455 3300
rect 3400 3055 3440 3060
rect 3400 3025 3405 3055
rect 3435 3040 3440 3055
rect 3435 3025 3545 3040
rect 3400 3020 3545 3025
rect 4530 2600 4570 2605
rect 4530 2570 4535 2600
rect 4565 2595 4570 2600
rect 5545 2600 5585 2605
rect 5545 2595 5550 2600
rect 4565 2575 5550 2595
rect 4565 2570 4570 2575
rect 4530 2565 4570 2570
rect 5545 2570 5550 2575
rect 5580 2570 5585 2600
rect 5545 2565 5585 2570
rect 3420 2525 3460 2530
rect 3420 2495 3425 2525
rect 3455 2520 3460 2525
rect 3455 2500 3510 2520
rect 3455 2495 3460 2500
rect 3420 2490 3460 2495
rect 2350 2405 2390 2410
rect 2350 2375 2355 2405
rect 2385 2400 2390 2405
rect 6590 2405 6630 2410
rect 2385 2380 2445 2400
rect 2385 2375 2390 2380
rect 2350 2370 2390 2375
rect 6590 2375 6595 2405
rect 6625 2375 6630 2405
rect 6590 2370 6630 2375
rect 2395 2200 2435 2205
rect 2395 2170 2400 2200
rect 2430 2195 2435 2200
rect 6545 2200 6585 2205
rect 2430 2175 2445 2195
rect 2430 2170 2435 2175
rect 2395 2165 2435 2170
rect 6545 2170 6550 2200
rect 6580 2170 6585 2200
rect 6545 2165 6585 2170
rect 3605 2015 3625 2035
rect 5355 2015 5375 2035
rect 2050 1485 2070 1505
rect 6865 1485 6885 1505
rect 4460 -215 4520 -200
rect 4460 -245 4475 -215
rect 4505 -245 4520 -215
rect 4460 -280 4520 -245
rect 4460 -310 4475 -280
rect 4505 -310 4520 -280
rect 4460 -350 4520 -310
rect 4460 -380 4475 -350
rect 4505 -380 4520 -350
rect 4460 -420 4520 -380
rect 4460 -450 4475 -420
rect 4505 -450 4520 -420
rect 4460 -490 4520 -450
rect 4460 -520 4475 -490
rect 4505 -520 4520 -490
rect 4460 -555 4520 -520
rect 4460 -585 4475 -555
rect 4505 -585 4520 -555
rect 4460 -600 4520 -585
<< via2 >>
rect 2335 15380 2365 15410
rect 2335 15315 2365 15345
rect 2335 15245 2365 15275
rect 2335 15175 2365 15205
rect 2335 15105 2365 15135
rect 2335 15040 2365 15070
rect 6705 15380 6735 15410
rect 6705 15315 6735 15345
rect 6705 15245 6735 15275
rect 6705 15175 6735 15205
rect 6705 15105 6735 15135
rect 6705 15040 6735 15070
rect 2390 6905 2420 6935
rect 2390 6840 2420 6870
rect 2390 6770 2420 6800
rect 2390 6700 2420 6730
rect 2390 6630 2420 6660
rect 2390 6565 2420 6595
rect 3245 6905 3275 6935
rect 3245 6840 3275 6870
rect 3245 6770 3275 6800
rect 3245 6700 3275 6730
rect 3245 6630 3275 6660
rect 3245 6565 3275 6595
rect 4475 6905 4505 6935
rect 4475 6840 4505 6870
rect 4475 6770 4505 6800
rect 4475 6700 4505 6730
rect 4475 6630 4505 6660
rect 4475 6565 4505 6595
rect 6305 6905 6335 6935
rect 6305 6840 6335 6870
rect 6305 6770 6335 6800
rect 6305 6700 6335 6730
rect 6305 6630 6335 6660
rect 6305 6565 6335 6595
rect 6595 6905 6625 6935
rect 6595 6840 6625 6870
rect 6595 6770 6625 6800
rect 6595 6700 6625 6730
rect 6595 6630 6625 6660
rect 6595 6565 6625 6595
rect 4475 -245 4505 -215
rect 4475 -310 4505 -280
rect 4475 -380 4505 -350
rect 4475 -450 4505 -420
rect 4475 -520 4505 -490
rect 4475 -585 4505 -555
<< metal3 >>
rect 2320 15415 2380 15425
rect 2320 15375 2330 15415
rect 2370 15375 2380 15415
rect 2320 15350 2380 15375
rect 2320 15310 2330 15350
rect 2370 15310 2380 15350
rect 2320 15280 2380 15310
rect 2320 15240 2330 15280
rect 2370 15240 2380 15280
rect 2320 15210 2380 15240
rect 2320 15170 2330 15210
rect 2370 15170 2380 15210
rect 2320 15140 2380 15170
rect 2320 15100 2330 15140
rect 2370 15100 2380 15140
rect 2320 15075 2380 15100
rect 2320 15035 2330 15075
rect 2370 15035 2380 15075
rect 2320 15025 2380 15035
rect 6690 15415 6750 15425
rect 6690 15375 6700 15415
rect 6740 15375 6750 15415
rect 6690 15350 6750 15375
rect 6690 15310 6700 15350
rect 6740 15310 6750 15350
rect 6690 15280 6750 15310
rect 6690 15240 6700 15280
rect 6740 15240 6750 15280
rect 6690 15210 6750 15240
rect 6690 15170 6700 15210
rect 6740 15170 6750 15210
rect 6690 15140 6750 15170
rect 6690 15100 6700 15140
rect 6740 15100 6750 15140
rect 6690 15075 6750 15100
rect 6690 15035 6700 15075
rect 6740 15035 6750 15075
rect 6690 15025 6750 15035
rect 10710 15390 11510 15425
rect 10710 15340 10745 15390
rect 10795 15340 10840 15390
rect 10890 15340 10935 15390
rect 10985 15340 11035 15390
rect 11085 15340 11135 15390
rect 11185 15340 11235 15390
rect 11285 15340 11330 15390
rect 11380 15340 11425 15390
rect 11475 15340 11510 15390
rect 10710 15300 11510 15340
rect 10710 15250 10745 15300
rect 10795 15250 10840 15300
rect 10890 15250 10935 15300
rect 10985 15250 11035 15300
rect 11085 15250 11135 15300
rect 11185 15250 11235 15300
rect 11285 15250 11330 15300
rect 11380 15250 11425 15300
rect 11475 15250 11510 15300
rect 10710 15200 11510 15250
rect 10710 15150 10745 15200
rect 10795 15150 10840 15200
rect 10890 15150 10935 15200
rect 10985 15150 11035 15200
rect 11085 15150 11135 15200
rect 11185 15150 11235 15200
rect 11285 15150 11330 15200
rect 11380 15150 11425 15200
rect 11475 15150 11510 15200
rect 10710 15110 11510 15150
rect 10710 15060 10745 15110
rect 10795 15060 10840 15110
rect 10890 15060 10935 15110
rect 10985 15060 11035 15110
rect 11085 15060 11135 15110
rect 11185 15060 11235 15110
rect 11285 15060 11330 15110
rect 11380 15060 11425 15110
rect 11475 15060 11510 15110
rect 6860 14850 7090 14935
rect 7210 14850 7440 14935
rect 7560 14850 7790 14935
rect 7910 14850 8140 14935
rect 8260 14850 8490 14935
rect 8610 14850 8840 14935
rect 8960 14850 9190 14935
rect 9310 14850 9540 14935
rect 9660 14850 9890 14935
rect 10010 14850 10240 14935
rect 10360 14850 10590 14935
rect 10710 14850 11510 15060
rect 6860 14800 11510 14850
rect 6860 14705 7090 14800
rect 7210 14705 7440 14800
rect 7560 14705 7790 14800
rect 7910 14705 8140 14800
rect 8260 14705 8490 14800
rect 8610 14705 8840 14800
rect 8960 14705 9190 14800
rect 9310 14705 9540 14800
rect 9660 14705 9890 14800
rect 10010 14705 10240 14800
rect 10360 14705 10590 14800
rect 8700 14585 8750 14705
rect 6860 14500 7090 14585
rect 7210 14500 7440 14585
rect 7560 14500 7790 14585
rect 7910 14500 8140 14585
rect 8260 14500 8490 14585
rect 8610 14500 8840 14585
rect 8960 14500 9190 14585
rect 9310 14500 9540 14585
rect 9660 14500 9890 14585
rect 10010 14500 10240 14585
rect 10360 14500 10590 14585
rect 6860 14450 10590 14500
rect 6860 14355 7090 14450
rect 7210 14355 7440 14450
rect 7560 14355 7790 14450
rect 7910 14355 8140 14450
rect 8260 14355 8490 14450
rect 8610 14355 8840 14450
rect 8960 14355 9190 14450
rect 9310 14355 9540 14450
rect 9660 14355 9890 14450
rect 10010 14355 10240 14450
rect 10360 14355 10590 14450
rect 8700 14235 8750 14355
rect 6860 14150 7090 14235
rect 7210 14150 7440 14235
rect 7560 14150 7790 14235
rect 7910 14150 8140 14235
rect 8260 14150 8490 14235
rect 8610 14150 8840 14235
rect 8960 14150 9190 14235
rect 9310 14150 9540 14235
rect 9660 14150 9890 14235
rect 10010 14150 10240 14235
rect 10360 14150 10590 14235
rect 6860 14100 10590 14150
rect 6860 14005 7090 14100
rect 7210 14005 7440 14100
rect 7560 14005 7790 14100
rect 7910 14005 8140 14100
rect 8260 14005 8490 14100
rect 8610 14005 8840 14100
rect 8960 14005 9190 14100
rect 9310 14005 9540 14100
rect 9660 14005 9890 14100
rect 10010 14005 10240 14100
rect 10360 14005 10590 14100
rect 8700 13885 8750 14005
rect 6860 13800 7090 13885
rect 7210 13800 7440 13885
rect 7560 13800 7790 13885
rect 7910 13800 8140 13885
rect 8260 13800 8490 13885
rect 8610 13800 8840 13885
rect 8960 13800 9190 13885
rect 9310 13800 9540 13885
rect 9660 13800 9890 13885
rect 10010 13800 10240 13885
rect 10360 13800 10590 13885
rect 6860 13750 10590 13800
rect 6860 13655 7090 13750
rect 7210 13655 7440 13750
rect 7560 13655 7790 13750
rect 7910 13655 8140 13750
rect 8260 13655 8490 13750
rect 8610 13655 8840 13750
rect 8960 13655 9190 13750
rect 9310 13655 9540 13750
rect 9660 13655 9890 13750
rect 10010 13655 10240 13750
rect 10360 13655 10590 13750
rect 8700 13535 8750 13655
rect 6860 13450 7090 13535
rect 7210 13450 7440 13535
rect 7560 13450 7790 13535
rect 7910 13450 8140 13535
rect 8260 13450 8490 13535
rect 8610 13450 8840 13535
rect 8960 13450 9190 13535
rect 9310 13450 9540 13535
rect 9660 13450 9890 13535
rect 10010 13450 10240 13535
rect 10360 13450 10590 13535
rect 6860 13400 10590 13450
rect 6860 13305 7090 13400
rect 7210 13305 7440 13400
rect 7560 13305 7790 13400
rect 7910 13305 8140 13400
rect 8260 13305 8490 13400
rect 8610 13305 8840 13400
rect 8960 13305 9190 13400
rect 9310 13305 9540 13400
rect 9660 13305 9890 13400
rect 10010 13305 10240 13400
rect 10360 13305 10590 13400
rect 8700 13185 8750 13305
rect 6860 13100 7090 13185
rect 7210 13100 7440 13185
rect 7560 13100 7790 13185
rect 7910 13100 8140 13185
rect 8260 13100 8490 13185
rect 8610 13100 8840 13185
rect 8960 13100 9190 13185
rect 9310 13100 9540 13185
rect 9660 13100 9890 13185
rect 10010 13100 10240 13185
rect 10360 13100 10590 13185
rect 6860 13050 10590 13100
rect 6860 12955 7090 13050
rect 7210 12955 7440 13050
rect 7560 12955 7790 13050
rect 7910 12955 8140 13050
rect 8260 12955 8490 13050
rect 8610 12955 8840 13050
rect 8960 12955 9190 13050
rect 9310 12955 9540 13050
rect 9660 12955 9890 13050
rect 10010 12955 10240 13050
rect 10360 12955 10590 13050
rect 8700 12835 8750 12955
rect 6860 12750 7090 12835
rect 7210 12750 7440 12835
rect 7560 12750 7790 12835
rect 7910 12750 8140 12835
rect 8260 12750 8490 12835
rect 8610 12750 8840 12835
rect 8960 12750 9190 12835
rect 9310 12750 9540 12835
rect 9660 12750 9890 12835
rect 10010 12750 10240 12835
rect 10360 12750 10590 12835
rect 6860 12700 10590 12750
rect 6860 12605 7090 12700
rect 7210 12605 7440 12700
rect 7560 12605 7790 12700
rect 7910 12605 8140 12700
rect 8260 12605 8490 12700
rect 8610 12605 8840 12700
rect 8960 12605 9190 12700
rect 9310 12605 9540 12700
rect 9660 12605 9890 12700
rect 10010 12605 10240 12700
rect 10360 12605 10590 12700
rect 8700 12485 8750 12605
rect 6860 12400 7090 12485
rect 7210 12400 7440 12485
rect 7560 12400 7790 12485
rect 7910 12400 8140 12485
rect 8260 12400 8490 12485
rect 8610 12400 8840 12485
rect 8960 12400 9190 12485
rect 9310 12400 9540 12485
rect 9660 12400 9890 12485
rect 10010 12400 10240 12485
rect 10360 12400 10590 12485
rect 6860 12350 10590 12400
rect 6860 12255 7090 12350
rect 7210 12255 7440 12350
rect 7560 12255 7790 12350
rect 7910 12255 8140 12350
rect 8260 12255 8490 12350
rect 8610 12255 8840 12350
rect 8960 12255 9190 12350
rect 9310 12255 9540 12350
rect 9660 12255 9890 12350
rect 10010 12255 10240 12350
rect 10360 12255 10590 12350
rect 8700 12135 8750 12255
rect 6860 12050 7090 12135
rect 7210 12050 7440 12135
rect 7560 12050 7790 12135
rect 7910 12050 8140 12135
rect 8260 12050 8490 12135
rect 8610 12050 8840 12135
rect 8960 12050 9190 12135
rect 9310 12050 9540 12135
rect 9660 12050 9890 12135
rect 10010 12050 10240 12135
rect 10360 12050 10590 12135
rect 6860 12000 10590 12050
rect 6860 11905 7090 12000
rect 7210 11905 7440 12000
rect 7560 11905 7790 12000
rect 7910 11905 8140 12000
rect 8260 11905 8490 12000
rect 8610 11905 8840 12000
rect 8960 11905 9190 12000
rect 9310 11905 9540 12000
rect 9660 11905 9890 12000
rect 10010 11905 10240 12000
rect 10360 11905 10590 12000
rect 8700 11785 8750 11905
rect 6860 11700 7090 11785
rect 7210 11700 7440 11785
rect 7560 11700 7790 11785
rect 7910 11700 8140 11785
rect 8260 11700 8490 11785
rect 8610 11700 8840 11785
rect 8960 11700 9190 11785
rect 9310 11700 9540 11785
rect 9660 11700 9890 11785
rect 10010 11700 10240 11785
rect 10360 11700 10590 11785
rect 6860 11650 10590 11700
rect 6860 11555 7090 11650
rect 7210 11555 7440 11650
rect 7560 11555 7790 11650
rect 7910 11555 8140 11650
rect 8260 11555 8490 11650
rect 8610 11555 8840 11650
rect 8960 11555 9190 11650
rect 9310 11555 9540 11650
rect 9660 11555 9890 11650
rect 10010 11555 10240 11650
rect 10360 11555 10590 11650
rect 8700 11435 8750 11555
rect 6860 11350 7090 11435
rect 7210 11350 7440 11435
rect 7560 11350 7790 11435
rect 7910 11350 8140 11435
rect 8260 11350 8490 11435
rect 8610 11350 8840 11435
rect 8960 11350 9190 11435
rect 9310 11350 9540 11435
rect 9660 11350 9890 11435
rect 10010 11350 10240 11435
rect 10360 11350 10590 11435
rect 6860 11300 10590 11350
rect 6860 11205 7090 11300
rect 7210 11205 7440 11300
rect 7560 11205 7790 11300
rect 7910 11205 8140 11300
rect 8260 11205 8490 11300
rect 8610 11205 8840 11300
rect 8960 11205 9190 11300
rect 9310 11205 9540 11300
rect 9660 11205 9890 11300
rect 10010 11205 10240 11300
rect 10360 11205 10590 11300
rect 8700 11085 8750 11205
rect 6860 11000 7090 11085
rect 7210 11000 7440 11085
rect 7560 11000 7790 11085
rect 7910 11000 8140 11085
rect 8260 11000 8490 11085
rect 8610 11000 8840 11085
rect 8960 11000 9190 11085
rect 9310 11000 9540 11085
rect 9660 11000 9890 11085
rect 10010 11000 10240 11085
rect 10360 11000 10590 11085
rect 6860 10950 10590 11000
rect 6860 10855 7090 10950
rect 7210 10855 7440 10950
rect 7560 10855 7790 10950
rect 7910 10855 8140 10950
rect 8260 10855 8490 10950
rect 8610 10855 8840 10950
rect 8960 10855 9190 10950
rect 9310 10855 9540 10950
rect 9660 10855 9890 10950
rect 10010 10855 10240 10950
rect 10360 10855 10590 10950
rect 8700 10735 8750 10855
rect 6860 10650 7090 10735
rect 7210 10650 7440 10735
rect 7560 10650 7790 10735
rect 7910 10650 8140 10735
rect 8260 10650 8490 10735
rect 8610 10650 8840 10735
rect 8960 10650 9190 10735
rect 9310 10650 9540 10735
rect 9660 10650 9890 10735
rect 10010 10650 10240 10735
rect 10360 10650 10590 10735
rect 6860 10600 10590 10650
rect 6860 10505 7090 10600
rect 7210 10505 7440 10600
rect 7560 10505 7790 10600
rect 7910 10505 8140 10600
rect 8260 10505 8490 10600
rect 8610 10505 8840 10600
rect 8960 10505 9190 10600
rect 9310 10505 9540 10600
rect 9660 10505 9890 10600
rect 10010 10505 10240 10600
rect 10360 10505 10590 10600
rect 8700 10385 8750 10505
rect 6860 10300 7090 10385
rect 7210 10300 7440 10385
rect 7560 10300 7790 10385
rect 7910 10300 8140 10385
rect 8260 10300 8490 10385
rect 8610 10300 8840 10385
rect 8960 10300 9190 10385
rect 9310 10300 9540 10385
rect 9660 10300 9890 10385
rect 10010 10300 10240 10385
rect 10360 10300 10590 10385
rect 6860 10250 10590 10300
rect 6860 10155 7090 10250
rect 7210 10155 7440 10250
rect 7560 10155 7790 10250
rect 7910 10155 8140 10250
rect 8260 10155 8490 10250
rect 8610 10155 8840 10250
rect 8960 10155 9190 10250
rect 9310 10155 9540 10250
rect 9660 10155 9890 10250
rect 10010 10155 10240 10250
rect 10360 10155 10590 10250
rect 8700 10035 8750 10155
rect 6860 9950 7090 10035
rect 7210 9950 7440 10035
rect 7560 9950 7790 10035
rect 7910 9950 8140 10035
rect 8260 9950 8490 10035
rect 8610 9950 8840 10035
rect 8960 9950 9190 10035
rect 9310 9950 9540 10035
rect 9660 9950 9890 10035
rect 10010 9950 10240 10035
rect 10360 9950 10590 10035
rect 6860 9900 10590 9950
rect 6860 9805 7090 9900
rect 7210 9805 7440 9900
rect 7560 9805 7790 9900
rect 7910 9805 8140 9900
rect 8260 9805 8490 9900
rect 8610 9805 8840 9900
rect 8960 9805 9190 9900
rect 9310 9805 9540 9900
rect 9660 9805 9890 9900
rect 10010 9805 10240 9900
rect 10360 9805 10590 9900
rect 8700 9685 8750 9805
rect 6860 9600 7090 9685
rect 7210 9600 7440 9685
rect 7560 9600 7790 9685
rect 7910 9600 8140 9685
rect 8260 9600 8490 9685
rect 8610 9600 8840 9685
rect 8960 9600 9190 9685
rect 9310 9600 9540 9685
rect 9660 9600 9890 9685
rect 10010 9600 10240 9685
rect 10360 9600 10590 9685
rect 6860 9550 10590 9600
rect 6860 9455 7090 9550
rect 7210 9455 7440 9550
rect 7560 9455 7790 9550
rect 7910 9455 8140 9550
rect 8260 9455 8490 9550
rect 8610 9455 8840 9550
rect 8960 9455 9190 9550
rect 9310 9455 9540 9550
rect 9660 9455 9890 9550
rect 10010 9455 10240 9550
rect 10360 9455 10590 9550
rect 8700 9335 8750 9455
rect 6860 9250 7090 9335
rect 7210 9250 7440 9335
rect 7560 9250 7790 9335
rect 7910 9250 8140 9335
rect 8260 9250 8490 9335
rect 8610 9250 8840 9335
rect 8960 9250 9190 9335
rect 9310 9250 9540 9335
rect 9660 9250 9890 9335
rect 10010 9250 10240 9335
rect 10360 9250 10590 9335
rect 6860 9200 10590 9250
rect 6860 9105 7090 9200
rect 7210 9105 7440 9200
rect 7560 9105 7790 9200
rect 7910 9105 8140 9200
rect 8260 9105 8490 9200
rect 8610 9105 8840 9200
rect 8960 9105 9190 9200
rect 9310 9105 9540 9200
rect 9660 9105 9890 9200
rect 10010 9105 10240 9200
rect 10360 9105 10590 9200
rect 8700 8985 8750 9105
rect 6860 8900 7090 8985
rect 7210 8900 7440 8985
rect 7560 8900 7790 8985
rect 7910 8900 8140 8985
rect 8260 8900 8490 8985
rect 8610 8900 8840 8985
rect 8960 8900 9190 8985
rect 9310 8900 9540 8985
rect 9660 8900 9890 8985
rect 10010 8900 10240 8985
rect 10360 8900 10590 8985
rect 6860 8850 10590 8900
rect 6860 8755 7090 8850
rect 7210 8755 7440 8850
rect 7560 8755 7790 8850
rect 7910 8755 8140 8850
rect 8260 8755 8490 8850
rect 8610 8755 8840 8850
rect 8960 8755 9190 8850
rect 9310 8755 9540 8850
rect 9660 8755 9890 8850
rect 10010 8755 10240 8850
rect 10360 8755 10590 8850
rect 8700 8635 8750 8755
rect 6860 8550 7090 8635
rect 7210 8550 7440 8635
rect 7560 8550 7790 8635
rect 7910 8550 8140 8635
rect 8260 8550 8490 8635
rect 8610 8550 8840 8635
rect 8960 8550 9190 8635
rect 9310 8550 9540 8635
rect 9660 8550 9890 8635
rect 10010 8550 10240 8635
rect 10360 8550 10590 8635
rect 6860 8500 10590 8550
rect 6860 8405 7090 8500
rect 7210 8405 7440 8500
rect 7560 8405 7790 8500
rect 7910 8405 8140 8500
rect 8260 8405 8490 8500
rect 8610 8405 8840 8500
rect 8960 8405 9190 8500
rect 9310 8405 9540 8500
rect 9660 8405 9890 8500
rect 10010 8405 10240 8500
rect 10360 8405 10590 8500
rect 8700 8285 8750 8405
rect -2440 6915 -1640 8255
rect 6860 8200 7090 8285
rect 7210 8200 7440 8285
rect 7560 8200 7790 8285
rect 7910 8200 8140 8285
rect 8260 8200 8490 8285
rect 8610 8200 8840 8285
rect 8960 8200 9190 8285
rect 9310 8200 9540 8285
rect 9660 8200 9890 8285
rect 10010 8200 10240 8285
rect 10360 8200 10590 8285
rect 6860 8150 10590 8200
rect 6860 8055 7090 8150
rect 7210 8055 7440 8150
rect 7560 8055 7790 8150
rect 7910 8055 8140 8150
rect 8260 8055 8490 8150
rect 8610 8055 8840 8150
rect 8960 8055 9190 8150
rect 9310 8055 9540 8150
rect 9660 8055 9890 8150
rect 10010 8055 10240 8150
rect 10360 8055 10590 8150
rect 8700 7935 8750 8055
rect 6860 7850 7090 7935
rect 7210 7850 7440 7935
rect 7560 7850 7790 7935
rect 7910 7850 8140 7935
rect 8260 7850 8490 7935
rect 8610 7850 8840 7935
rect 8960 7850 9190 7935
rect 9310 7850 9540 7935
rect 9660 7850 9890 7935
rect 10010 7850 10240 7935
rect 10360 7850 10590 7935
rect 6860 7800 10590 7850
rect 6860 7705 7090 7800
rect 7210 7705 7440 7800
rect 7560 7705 7790 7800
rect 7910 7705 8140 7800
rect 8260 7705 8490 7800
rect 8610 7705 8840 7800
rect 8960 7705 9190 7800
rect 9310 7705 9540 7800
rect 9660 7705 9890 7800
rect 10010 7705 10240 7800
rect 10360 7705 10590 7800
rect 8700 7585 8750 7705
rect 6860 7500 7090 7585
rect 7210 7500 7440 7585
rect 7560 7500 7790 7585
rect 7910 7500 8140 7585
rect 8260 7500 8490 7585
rect 8610 7500 8840 7585
rect 8960 7500 9190 7585
rect 9310 7500 9540 7585
rect 9660 7500 9890 7585
rect 10010 7500 10240 7585
rect 10360 7500 10590 7585
rect 6860 7450 10590 7500
rect 6860 7355 7090 7450
rect 7210 7355 7440 7450
rect 7560 7355 7790 7450
rect 7910 7355 8140 7450
rect 8260 7355 8490 7450
rect 8610 7355 8840 7450
rect 8960 7355 9190 7450
rect 9310 7355 9540 7450
rect 9660 7355 9890 7450
rect 10010 7355 10240 7450
rect 10360 7355 10590 7450
rect 8700 7235 8750 7355
rect 6860 7150 7090 7235
rect 7210 7150 7440 7235
rect 7560 7150 7790 7235
rect 7910 7150 8140 7235
rect 8260 7150 8490 7235
rect 8610 7150 8840 7235
rect 8960 7150 9190 7235
rect 9310 7150 9540 7235
rect 9660 7150 9890 7235
rect 10010 7150 10240 7235
rect 10360 7150 10590 7235
rect 6860 7100 10590 7150
rect 6860 7005 7090 7100
rect 7210 7005 7440 7100
rect 7560 7005 7790 7100
rect 7910 7005 8140 7100
rect 8260 7005 8490 7100
rect 8610 7005 8840 7100
rect 8960 7005 9190 7100
rect 9310 7005 9540 7100
rect 9660 7005 9890 7100
rect 10010 7005 10240 7100
rect 10360 7005 10590 7100
rect -2440 6865 -2405 6915
rect -2355 6865 -2310 6915
rect -2260 6865 -2215 6915
rect -2165 6865 -2115 6915
rect -2065 6865 -2015 6915
rect -1965 6865 -1915 6915
rect -1865 6865 -1820 6915
rect -1770 6865 -1725 6915
rect -1675 6865 -1640 6915
rect -2440 6825 -1640 6865
rect -2440 6775 -2405 6825
rect -2355 6775 -2310 6825
rect -2260 6775 -2215 6825
rect -2165 6775 -2115 6825
rect -2065 6775 -2015 6825
rect -1965 6775 -1915 6825
rect -1865 6775 -1820 6825
rect -1770 6775 -1725 6825
rect -1675 6775 -1640 6825
rect -2440 6725 -1640 6775
rect -2440 6675 -2405 6725
rect -2355 6675 -2310 6725
rect -2260 6675 -2215 6725
rect -2165 6675 -2115 6725
rect -2065 6675 -2015 6725
rect -1965 6675 -1915 6725
rect -1865 6675 -1820 6725
rect -1770 6675 -1725 6725
rect -1675 6675 -1640 6725
rect -2440 6635 -1640 6675
rect -2440 6585 -2405 6635
rect -2355 6585 -2310 6635
rect -2260 6585 -2215 6635
rect -2165 6585 -2115 6635
rect -2065 6585 -2015 6635
rect -1965 6585 -1915 6635
rect -1865 6585 -1820 6635
rect -1770 6585 -1725 6635
rect -1675 6585 -1640 6635
rect -2440 6550 -1640 6585
rect 2375 6940 2435 6950
rect 2375 6900 2385 6940
rect 2425 6900 2435 6940
rect 2375 6875 2435 6900
rect 2375 6835 2385 6875
rect 2425 6835 2435 6875
rect 2375 6805 2435 6835
rect 2375 6765 2385 6805
rect 2425 6765 2435 6805
rect 2375 6735 2435 6765
rect 2375 6695 2385 6735
rect 2425 6695 2435 6735
rect 2375 6665 2435 6695
rect 2375 6625 2385 6665
rect 2425 6625 2435 6665
rect 2375 6600 2435 6625
rect 2375 6560 2385 6600
rect 2425 6560 2435 6600
rect 2375 6550 2435 6560
rect 3230 6940 3290 6950
rect 3230 6900 3240 6940
rect 3280 6900 3290 6940
rect 3230 6875 3290 6900
rect 3230 6835 3240 6875
rect 3280 6835 3290 6875
rect 3230 6805 3290 6835
rect 3230 6765 3240 6805
rect 3280 6765 3290 6805
rect 3230 6735 3290 6765
rect 3230 6695 3240 6735
rect 3280 6695 3290 6735
rect 3230 6665 3290 6695
rect 3230 6625 3240 6665
rect 3280 6625 3290 6665
rect 3230 6600 3290 6625
rect 3230 6560 3240 6600
rect 3280 6560 3290 6600
rect 3230 6550 3290 6560
rect 4465 6940 4515 6950
rect 4465 6900 4470 6940
rect 4510 6900 4515 6940
rect 4465 6875 4515 6900
rect 4465 6835 4470 6875
rect 4510 6835 4515 6875
rect 4465 6805 4515 6835
rect 4465 6765 4470 6805
rect 4510 6765 4515 6805
rect 4465 6735 4515 6765
rect 4465 6695 4470 6735
rect 4510 6695 4515 6735
rect 4465 6665 4515 6695
rect 4465 6625 4470 6665
rect 4510 6625 4515 6665
rect 4465 6600 4515 6625
rect 4465 6560 4470 6600
rect 4510 6560 4515 6600
rect 4465 6550 4515 6560
rect 6290 6940 6350 6950
rect 6290 6900 6300 6940
rect 6340 6900 6350 6940
rect 6290 6875 6350 6900
rect 6290 6835 6300 6875
rect 6340 6835 6350 6875
rect 6290 6805 6350 6835
rect 6290 6765 6300 6805
rect 6340 6765 6350 6805
rect 6290 6735 6350 6765
rect 6290 6695 6300 6735
rect 6340 6695 6350 6735
rect 6290 6665 6350 6695
rect 6290 6625 6300 6665
rect 6340 6625 6350 6665
rect 6290 6600 6350 6625
rect 6290 6560 6300 6600
rect 6340 6560 6350 6600
rect 6290 6550 6350 6560
rect 6580 6940 6640 6950
rect 6580 6900 6590 6940
rect 6630 6900 6640 6940
rect 6580 6875 6640 6900
rect 8700 6885 8750 7005
rect 10710 6915 11510 14800
rect 6580 6835 6590 6875
rect 6630 6835 6640 6875
rect 6580 6805 6640 6835
rect 6580 6765 6590 6805
rect 6630 6765 6640 6805
rect 6580 6735 6640 6765
rect 6580 6695 6590 6735
rect 6630 6695 6640 6735
rect 6580 6665 6640 6695
rect 6580 6625 6590 6665
rect 6630 6625 6640 6665
rect 6860 6800 7090 6885
rect 7210 6800 7440 6885
rect 7560 6800 7790 6885
rect 7910 6800 8140 6885
rect 8260 6800 8490 6885
rect 8610 6800 8840 6885
rect 8960 6800 9190 6885
rect 9310 6800 9540 6885
rect 9660 6800 9890 6885
rect 10010 6800 10240 6885
rect 10360 6800 10590 6885
rect 6860 6750 10590 6800
rect 6860 6655 7090 6750
rect 7210 6655 7440 6750
rect 7560 6655 7790 6750
rect 7910 6655 8140 6750
rect 8260 6655 8490 6750
rect 8610 6655 8840 6750
rect 8960 6655 9190 6750
rect 9310 6655 9540 6750
rect 9660 6655 9890 6750
rect 10010 6655 10240 6750
rect 10360 6655 10590 6750
rect 10710 6865 10745 6915
rect 10795 6865 10840 6915
rect 10890 6865 10935 6915
rect 10985 6865 11035 6915
rect 11085 6865 11135 6915
rect 11185 6865 11235 6915
rect 11285 6865 11330 6915
rect 11380 6865 11425 6915
rect 11475 6865 11510 6915
rect 10710 6825 11510 6865
rect 10710 6775 10745 6825
rect 10795 6775 10840 6825
rect 10890 6775 10935 6825
rect 10985 6775 11035 6825
rect 11085 6775 11135 6825
rect 11185 6775 11235 6825
rect 11285 6775 11330 6825
rect 11380 6775 11425 6825
rect 11475 6775 11510 6825
rect 10710 6725 11510 6775
rect 10710 6675 10745 6725
rect 10795 6675 10840 6725
rect 10890 6675 10935 6725
rect 10985 6675 11035 6725
rect 11085 6675 11135 6725
rect 11185 6675 11235 6725
rect 11285 6675 11330 6725
rect 11380 6675 11425 6725
rect 11475 6675 11510 6725
rect 6580 6600 6640 6625
rect 6580 6560 6590 6600
rect 6630 6560 6640 6600
rect 6580 6550 6640 6560
rect 10710 6635 11510 6675
rect 10710 6585 10745 6635
rect 10795 6585 10840 6635
rect 10890 6585 10935 6635
rect 10985 6585 11035 6635
rect 11085 6585 11135 6635
rect 11185 6585 11235 6635
rect 11285 6585 11330 6635
rect 11380 6585 11425 6635
rect 11475 6585 11510 6635
rect 4460 -210 4520 -200
rect 4460 -250 4470 -210
rect 4510 -250 4520 -210
rect 4460 -275 4520 -250
rect 4460 -315 4470 -275
rect 4510 -315 4520 -275
rect 4460 -345 4520 -315
rect 4460 -385 4470 -345
rect 4510 -385 4520 -345
rect 4460 -415 4520 -385
rect 4460 -455 4470 -415
rect 4510 -455 4520 -415
rect 4460 -485 4520 -455
rect 4460 -525 4470 -485
rect 4510 -525 4520 -485
rect 4460 -550 4520 -525
rect 4460 -590 4470 -550
rect 4510 -590 4520 -550
rect 4460 -600 4520 -590
rect 10710 -235 11510 6585
rect 10710 -285 10745 -235
rect 10795 -285 10840 -235
rect 10890 -285 10935 -235
rect 10985 -285 11035 -235
rect 11085 -285 11135 -235
rect 11185 -285 11235 -235
rect 11285 -285 11330 -235
rect 11380 -285 11425 -235
rect 11475 -285 11510 -235
rect 10710 -325 11510 -285
rect 10710 -375 10745 -325
rect 10795 -375 10840 -325
rect 10890 -375 10935 -325
rect 10985 -375 11035 -325
rect 11085 -375 11135 -325
rect 11185 -375 11235 -325
rect 11285 -375 11330 -325
rect 11380 -375 11425 -325
rect 11475 -375 11510 -325
rect 10710 -425 11510 -375
rect 10710 -475 10745 -425
rect 10795 -475 10840 -425
rect 10890 -475 10935 -425
rect 10985 -475 11035 -425
rect 11085 -475 11135 -425
rect 11185 -475 11235 -425
rect 11285 -475 11330 -425
rect 11380 -475 11425 -425
rect 11475 -475 11510 -425
rect 10710 -515 11510 -475
rect 10710 -565 10745 -515
rect 10795 -565 10840 -515
rect 10890 -565 10935 -515
rect 10985 -565 11035 -515
rect 11085 -565 11135 -515
rect 11185 -565 11235 -515
rect 11285 -565 11330 -515
rect 11380 -565 11425 -515
rect 11475 -565 11510 -515
rect 10710 -600 11510 -565
<< via3 >>
rect 2330 15410 2370 15415
rect 2330 15380 2335 15410
rect 2335 15380 2365 15410
rect 2365 15380 2370 15410
rect 2330 15375 2370 15380
rect 2330 15345 2370 15350
rect 2330 15315 2335 15345
rect 2335 15315 2365 15345
rect 2365 15315 2370 15345
rect 2330 15310 2370 15315
rect 2330 15275 2370 15280
rect 2330 15245 2335 15275
rect 2335 15245 2365 15275
rect 2365 15245 2370 15275
rect 2330 15240 2370 15245
rect 2330 15205 2370 15210
rect 2330 15175 2335 15205
rect 2335 15175 2365 15205
rect 2365 15175 2370 15205
rect 2330 15170 2370 15175
rect 2330 15135 2370 15140
rect 2330 15105 2335 15135
rect 2335 15105 2365 15135
rect 2365 15105 2370 15135
rect 2330 15100 2370 15105
rect 2330 15070 2370 15075
rect 2330 15040 2335 15070
rect 2335 15040 2365 15070
rect 2365 15040 2370 15070
rect 2330 15035 2370 15040
rect 6700 15410 6740 15415
rect 6700 15380 6705 15410
rect 6705 15380 6735 15410
rect 6735 15380 6740 15410
rect 6700 15375 6740 15380
rect 6700 15345 6740 15350
rect 6700 15315 6705 15345
rect 6705 15315 6735 15345
rect 6735 15315 6740 15345
rect 6700 15310 6740 15315
rect 6700 15275 6740 15280
rect 6700 15245 6705 15275
rect 6705 15245 6735 15275
rect 6735 15245 6740 15275
rect 6700 15240 6740 15245
rect 6700 15205 6740 15210
rect 6700 15175 6705 15205
rect 6705 15175 6735 15205
rect 6735 15175 6740 15205
rect 6700 15170 6740 15175
rect 6700 15135 6740 15140
rect 6700 15105 6705 15135
rect 6705 15105 6735 15135
rect 6735 15105 6740 15135
rect 6700 15100 6740 15105
rect 6700 15070 6740 15075
rect 6700 15040 6705 15070
rect 6705 15040 6735 15070
rect 6735 15040 6740 15070
rect 6700 15035 6740 15040
rect 10745 15340 10795 15390
rect 10840 15340 10890 15390
rect 10935 15340 10985 15390
rect 11035 15340 11085 15390
rect 11135 15340 11185 15390
rect 11235 15340 11285 15390
rect 11330 15340 11380 15390
rect 11425 15340 11475 15390
rect 10745 15250 10795 15300
rect 10840 15250 10890 15300
rect 10935 15250 10985 15300
rect 11035 15250 11085 15300
rect 11135 15250 11185 15300
rect 11235 15250 11285 15300
rect 11330 15250 11380 15300
rect 11425 15250 11475 15300
rect 10745 15150 10795 15200
rect 10840 15150 10890 15200
rect 10935 15150 10985 15200
rect 11035 15150 11085 15200
rect 11135 15150 11185 15200
rect 11235 15150 11285 15200
rect 11330 15150 11380 15200
rect 11425 15150 11475 15200
rect 10745 15060 10795 15110
rect 10840 15060 10890 15110
rect 10935 15060 10985 15110
rect 11035 15060 11085 15110
rect 11135 15060 11185 15110
rect 11235 15060 11285 15110
rect 11330 15060 11380 15110
rect 11425 15060 11475 15110
rect -2405 6865 -2355 6915
rect -2310 6865 -2260 6915
rect -2215 6865 -2165 6915
rect -2115 6865 -2065 6915
rect -2015 6865 -1965 6915
rect -1915 6865 -1865 6915
rect -1820 6865 -1770 6915
rect -1725 6865 -1675 6915
rect -2405 6775 -2355 6825
rect -2310 6775 -2260 6825
rect -2215 6775 -2165 6825
rect -2115 6775 -2065 6825
rect -2015 6775 -1965 6825
rect -1915 6775 -1865 6825
rect -1820 6775 -1770 6825
rect -1725 6775 -1675 6825
rect -2405 6675 -2355 6725
rect -2310 6675 -2260 6725
rect -2215 6675 -2165 6725
rect -2115 6675 -2065 6725
rect -2015 6675 -1965 6725
rect -1915 6675 -1865 6725
rect -1820 6675 -1770 6725
rect -1725 6675 -1675 6725
rect -2405 6585 -2355 6635
rect -2310 6585 -2260 6635
rect -2215 6585 -2165 6635
rect -2115 6585 -2065 6635
rect -2015 6585 -1965 6635
rect -1915 6585 -1865 6635
rect -1820 6585 -1770 6635
rect -1725 6585 -1675 6635
rect 2385 6935 2425 6940
rect 2385 6905 2390 6935
rect 2390 6905 2420 6935
rect 2420 6905 2425 6935
rect 2385 6900 2425 6905
rect 2385 6870 2425 6875
rect 2385 6840 2390 6870
rect 2390 6840 2420 6870
rect 2420 6840 2425 6870
rect 2385 6835 2425 6840
rect 2385 6800 2425 6805
rect 2385 6770 2390 6800
rect 2390 6770 2420 6800
rect 2420 6770 2425 6800
rect 2385 6765 2425 6770
rect 2385 6730 2425 6735
rect 2385 6700 2390 6730
rect 2390 6700 2420 6730
rect 2420 6700 2425 6730
rect 2385 6695 2425 6700
rect 2385 6660 2425 6665
rect 2385 6630 2390 6660
rect 2390 6630 2420 6660
rect 2420 6630 2425 6660
rect 2385 6625 2425 6630
rect 2385 6595 2425 6600
rect 2385 6565 2390 6595
rect 2390 6565 2420 6595
rect 2420 6565 2425 6595
rect 2385 6560 2425 6565
rect 3240 6935 3280 6940
rect 3240 6905 3245 6935
rect 3245 6905 3275 6935
rect 3275 6905 3280 6935
rect 3240 6900 3280 6905
rect 3240 6870 3280 6875
rect 3240 6840 3245 6870
rect 3245 6840 3275 6870
rect 3275 6840 3280 6870
rect 3240 6835 3280 6840
rect 3240 6800 3280 6805
rect 3240 6770 3245 6800
rect 3245 6770 3275 6800
rect 3275 6770 3280 6800
rect 3240 6765 3280 6770
rect 3240 6730 3280 6735
rect 3240 6700 3245 6730
rect 3245 6700 3275 6730
rect 3275 6700 3280 6730
rect 3240 6695 3280 6700
rect 3240 6660 3280 6665
rect 3240 6630 3245 6660
rect 3245 6630 3275 6660
rect 3275 6630 3280 6660
rect 3240 6625 3280 6630
rect 3240 6595 3280 6600
rect 3240 6565 3245 6595
rect 3245 6565 3275 6595
rect 3275 6565 3280 6595
rect 3240 6560 3280 6565
rect 4470 6935 4510 6940
rect 4470 6905 4475 6935
rect 4475 6905 4505 6935
rect 4505 6905 4510 6935
rect 4470 6900 4510 6905
rect 4470 6870 4510 6875
rect 4470 6840 4475 6870
rect 4475 6840 4505 6870
rect 4505 6840 4510 6870
rect 4470 6835 4510 6840
rect 4470 6800 4510 6805
rect 4470 6770 4475 6800
rect 4475 6770 4505 6800
rect 4505 6770 4510 6800
rect 4470 6765 4510 6770
rect 4470 6730 4510 6735
rect 4470 6700 4475 6730
rect 4475 6700 4505 6730
rect 4505 6700 4510 6730
rect 4470 6695 4510 6700
rect 4470 6660 4510 6665
rect 4470 6630 4475 6660
rect 4475 6630 4505 6660
rect 4505 6630 4510 6660
rect 4470 6625 4510 6630
rect 4470 6595 4510 6600
rect 4470 6565 4475 6595
rect 4475 6565 4505 6595
rect 4505 6565 4510 6595
rect 4470 6560 4510 6565
rect 6300 6935 6340 6940
rect 6300 6905 6305 6935
rect 6305 6905 6335 6935
rect 6335 6905 6340 6935
rect 6300 6900 6340 6905
rect 6300 6870 6340 6875
rect 6300 6840 6305 6870
rect 6305 6840 6335 6870
rect 6335 6840 6340 6870
rect 6300 6835 6340 6840
rect 6300 6800 6340 6805
rect 6300 6770 6305 6800
rect 6305 6770 6335 6800
rect 6335 6770 6340 6800
rect 6300 6765 6340 6770
rect 6300 6730 6340 6735
rect 6300 6700 6305 6730
rect 6305 6700 6335 6730
rect 6335 6700 6340 6730
rect 6300 6695 6340 6700
rect 6300 6660 6340 6665
rect 6300 6630 6305 6660
rect 6305 6630 6335 6660
rect 6335 6630 6340 6660
rect 6300 6625 6340 6630
rect 6300 6595 6340 6600
rect 6300 6565 6305 6595
rect 6305 6565 6335 6595
rect 6335 6565 6340 6595
rect 6300 6560 6340 6565
rect 6590 6935 6630 6940
rect 6590 6905 6595 6935
rect 6595 6905 6625 6935
rect 6625 6905 6630 6935
rect 6590 6900 6630 6905
rect 6590 6870 6630 6875
rect 6590 6840 6595 6870
rect 6595 6840 6625 6870
rect 6625 6840 6630 6870
rect 6590 6835 6630 6840
rect 6590 6800 6630 6805
rect 6590 6770 6595 6800
rect 6595 6770 6625 6800
rect 6625 6770 6630 6800
rect 6590 6765 6630 6770
rect 6590 6730 6630 6735
rect 6590 6700 6595 6730
rect 6595 6700 6625 6730
rect 6625 6700 6630 6730
rect 6590 6695 6630 6700
rect 6590 6660 6630 6665
rect 6590 6630 6595 6660
rect 6595 6630 6625 6660
rect 6625 6630 6630 6660
rect 6590 6625 6630 6630
rect 10745 6865 10795 6915
rect 10840 6865 10890 6915
rect 10935 6865 10985 6915
rect 11035 6865 11085 6915
rect 11135 6865 11185 6915
rect 11235 6865 11285 6915
rect 11330 6865 11380 6915
rect 11425 6865 11475 6915
rect 10745 6775 10795 6825
rect 10840 6775 10890 6825
rect 10935 6775 10985 6825
rect 11035 6775 11085 6825
rect 11135 6775 11185 6825
rect 11235 6775 11285 6825
rect 11330 6775 11380 6825
rect 11425 6775 11475 6825
rect 10745 6675 10795 6725
rect 10840 6675 10890 6725
rect 10935 6675 10985 6725
rect 11035 6675 11085 6725
rect 11135 6675 11185 6725
rect 11235 6675 11285 6725
rect 11330 6675 11380 6725
rect 11425 6675 11475 6725
rect 6590 6595 6630 6600
rect 6590 6565 6595 6595
rect 6595 6565 6625 6595
rect 6625 6565 6630 6595
rect 6590 6560 6630 6565
rect 10745 6585 10795 6635
rect 10840 6585 10890 6635
rect 10935 6585 10985 6635
rect 11035 6585 11085 6635
rect 11135 6585 11185 6635
rect 11235 6585 11285 6635
rect 11330 6585 11380 6635
rect 11425 6585 11475 6635
rect 4470 -215 4510 -210
rect 4470 -245 4475 -215
rect 4475 -245 4505 -215
rect 4505 -245 4510 -215
rect 4470 -250 4510 -245
rect 4470 -280 4510 -275
rect 4470 -310 4475 -280
rect 4475 -310 4505 -280
rect 4505 -310 4510 -280
rect 4470 -315 4510 -310
rect 4470 -350 4510 -345
rect 4470 -380 4475 -350
rect 4475 -380 4505 -350
rect 4505 -380 4510 -350
rect 4470 -385 4510 -380
rect 4470 -420 4510 -415
rect 4470 -450 4475 -420
rect 4475 -450 4505 -420
rect 4505 -450 4510 -420
rect 4470 -455 4510 -450
rect 4470 -490 4510 -485
rect 4470 -520 4475 -490
rect 4475 -520 4505 -490
rect 4505 -520 4510 -490
rect 4470 -525 4510 -520
rect 4470 -555 4510 -550
rect 4470 -585 4475 -555
rect 4475 -585 4505 -555
rect 4505 -585 4510 -555
rect 4470 -590 4510 -585
rect 10745 -285 10795 -235
rect 10840 -285 10890 -235
rect 10935 -285 10985 -235
rect 11035 -285 11085 -235
rect 11135 -285 11185 -235
rect 11235 -285 11285 -235
rect 11330 -285 11380 -235
rect 11425 -285 11475 -235
rect 10745 -375 10795 -325
rect 10840 -375 10890 -325
rect 10935 -375 10985 -325
rect 11035 -375 11085 -325
rect 11135 -375 11185 -325
rect 11235 -375 11285 -325
rect 11330 -375 11380 -325
rect 11425 -375 11475 -325
rect 10745 -475 10795 -425
rect 10840 -475 10890 -425
rect 10935 -475 10985 -425
rect 11035 -475 11085 -425
rect 11135 -475 11185 -425
rect 11235 -475 11285 -425
rect 11330 -475 11380 -425
rect 11425 -475 11475 -425
rect 10745 -565 10795 -515
rect 10840 -565 10890 -515
rect 10935 -565 10985 -515
rect 11035 -565 11085 -515
rect 11135 -565 11185 -515
rect 11235 -565 11285 -515
rect 11330 -565 11380 -515
rect 11425 -565 11475 -515
<< mimcap >>
rect 6875 14845 7075 14920
rect 6875 14805 6955 14845
rect 6995 14805 7075 14845
rect 6875 14720 7075 14805
rect 7225 14845 7425 14920
rect 7225 14805 7305 14845
rect 7345 14805 7425 14845
rect 7225 14720 7425 14805
rect 7575 14845 7775 14920
rect 7575 14805 7655 14845
rect 7695 14805 7775 14845
rect 7575 14720 7775 14805
rect 7925 14845 8125 14920
rect 7925 14805 8005 14845
rect 8045 14805 8125 14845
rect 7925 14720 8125 14805
rect 8275 14845 8475 14920
rect 8275 14805 8355 14845
rect 8395 14805 8475 14845
rect 8275 14720 8475 14805
rect 8625 14845 8825 14920
rect 8625 14805 8705 14845
rect 8745 14805 8825 14845
rect 8625 14720 8825 14805
rect 8975 14845 9175 14920
rect 8975 14805 9055 14845
rect 9095 14805 9175 14845
rect 8975 14720 9175 14805
rect 9325 14845 9525 14920
rect 9325 14805 9405 14845
rect 9445 14805 9525 14845
rect 9325 14720 9525 14805
rect 9675 14845 9875 14920
rect 9675 14805 9755 14845
rect 9795 14805 9875 14845
rect 9675 14720 9875 14805
rect 10025 14845 10225 14920
rect 10025 14805 10105 14845
rect 10145 14805 10225 14845
rect 10025 14720 10225 14805
rect 10375 14845 10575 14920
rect 10375 14805 10455 14845
rect 10495 14805 10575 14845
rect 10375 14720 10575 14805
rect 6875 14495 7075 14570
rect 6875 14455 6955 14495
rect 6995 14455 7075 14495
rect 6875 14370 7075 14455
rect 7225 14495 7425 14570
rect 7225 14455 7305 14495
rect 7345 14455 7425 14495
rect 7225 14370 7425 14455
rect 7575 14495 7775 14570
rect 7575 14455 7655 14495
rect 7695 14455 7775 14495
rect 7575 14370 7775 14455
rect 7925 14495 8125 14570
rect 7925 14455 8005 14495
rect 8045 14455 8125 14495
rect 7925 14370 8125 14455
rect 8275 14495 8475 14570
rect 8275 14455 8355 14495
rect 8395 14455 8475 14495
rect 8275 14370 8475 14455
rect 8625 14495 8825 14570
rect 8625 14455 8705 14495
rect 8745 14455 8825 14495
rect 8625 14370 8825 14455
rect 8975 14495 9175 14570
rect 8975 14455 9055 14495
rect 9095 14455 9175 14495
rect 8975 14370 9175 14455
rect 9325 14495 9525 14570
rect 9325 14455 9405 14495
rect 9445 14455 9525 14495
rect 9325 14370 9525 14455
rect 9675 14495 9875 14570
rect 9675 14455 9755 14495
rect 9795 14455 9875 14495
rect 9675 14370 9875 14455
rect 10025 14495 10225 14570
rect 10025 14455 10105 14495
rect 10145 14455 10225 14495
rect 10025 14370 10225 14455
rect 10375 14495 10575 14570
rect 10375 14455 10455 14495
rect 10495 14455 10575 14495
rect 10375 14370 10575 14455
rect 6875 14145 7075 14220
rect 6875 14105 6955 14145
rect 6995 14105 7075 14145
rect 6875 14020 7075 14105
rect 7225 14145 7425 14220
rect 7225 14105 7305 14145
rect 7345 14105 7425 14145
rect 7225 14020 7425 14105
rect 7575 14145 7775 14220
rect 7575 14105 7655 14145
rect 7695 14105 7775 14145
rect 7575 14020 7775 14105
rect 7925 14145 8125 14220
rect 7925 14105 8005 14145
rect 8045 14105 8125 14145
rect 7925 14020 8125 14105
rect 8275 14145 8475 14220
rect 8275 14105 8355 14145
rect 8395 14105 8475 14145
rect 8275 14020 8475 14105
rect 8625 14145 8825 14220
rect 8625 14105 8705 14145
rect 8745 14105 8825 14145
rect 8625 14020 8825 14105
rect 8975 14145 9175 14220
rect 8975 14105 9055 14145
rect 9095 14105 9175 14145
rect 8975 14020 9175 14105
rect 9325 14145 9525 14220
rect 9325 14105 9405 14145
rect 9445 14105 9525 14145
rect 9325 14020 9525 14105
rect 9675 14145 9875 14220
rect 9675 14105 9755 14145
rect 9795 14105 9875 14145
rect 9675 14020 9875 14105
rect 10025 14145 10225 14220
rect 10025 14105 10105 14145
rect 10145 14105 10225 14145
rect 10025 14020 10225 14105
rect 10375 14145 10575 14220
rect 10375 14105 10455 14145
rect 10495 14105 10575 14145
rect 10375 14020 10575 14105
rect 6875 13795 7075 13870
rect 6875 13755 6955 13795
rect 6995 13755 7075 13795
rect 6875 13670 7075 13755
rect 7225 13795 7425 13870
rect 7225 13755 7305 13795
rect 7345 13755 7425 13795
rect 7225 13670 7425 13755
rect 7575 13795 7775 13870
rect 7575 13755 7655 13795
rect 7695 13755 7775 13795
rect 7575 13670 7775 13755
rect 7925 13795 8125 13870
rect 7925 13755 8005 13795
rect 8045 13755 8125 13795
rect 7925 13670 8125 13755
rect 8275 13795 8475 13870
rect 8275 13755 8355 13795
rect 8395 13755 8475 13795
rect 8275 13670 8475 13755
rect 8625 13795 8825 13870
rect 8625 13755 8705 13795
rect 8745 13755 8825 13795
rect 8625 13670 8825 13755
rect 8975 13795 9175 13870
rect 8975 13755 9055 13795
rect 9095 13755 9175 13795
rect 8975 13670 9175 13755
rect 9325 13795 9525 13870
rect 9325 13755 9405 13795
rect 9445 13755 9525 13795
rect 9325 13670 9525 13755
rect 9675 13795 9875 13870
rect 9675 13755 9755 13795
rect 9795 13755 9875 13795
rect 9675 13670 9875 13755
rect 10025 13795 10225 13870
rect 10025 13755 10105 13795
rect 10145 13755 10225 13795
rect 10025 13670 10225 13755
rect 10375 13795 10575 13870
rect 10375 13755 10455 13795
rect 10495 13755 10575 13795
rect 10375 13670 10575 13755
rect 6875 13445 7075 13520
rect 6875 13405 6955 13445
rect 6995 13405 7075 13445
rect 6875 13320 7075 13405
rect 7225 13445 7425 13520
rect 7225 13405 7305 13445
rect 7345 13405 7425 13445
rect 7225 13320 7425 13405
rect 7575 13445 7775 13520
rect 7575 13405 7655 13445
rect 7695 13405 7775 13445
rect 7575 13320 7775 13405
rect 7925 13445 8125 13520
rect 7925 13405 8005 13445
rect 8045 13405 8125 13445
rect 7925 13320 8125 13405
rect 8275 13445 8475 13520
rect 8275 13405 8355 13445
rect 8395 13405 8475 13445
rect 8275 13320 8475 13405
rect 8625 13445 8825 13520
rect 8625 13405 8705 13445
rect 8745 13405 8825 13445
rect 8625 13320 8825 13405
rect 8975 13445 9175 13520
rect 8975 13405 9055 13445
rect 9095 13405 9175 13445
rect 8975 13320 9175 13405
rect 9325 13445 9525 13520
rect 9325 13405 9405 13445
rect 9445 13405 9525 13445
rect 9325 13320 9525 13405
rect 9675 13445 9875 13520
rect 9675 13405 9755 13445
rect 9795 13405 9875 13445
rect 9675 13320 9875 13405
rect 10025 13445 10225 13520
rect 10025 13405 10105 13445
rect 10145 13405 10225 13445
rect 10025 13320 10225 13405
rect 10375 13445 10575 13520
rect 10375 13405 10455 13445
rect 10495 13405 10575 13445
rect 10375 13320 10575 13405
rect 6875 13095 7075 13170
rect 6875 13055 6955 13095
rect 6995 13055 7075 13095
rect 6875 12970 7075 13055
rect 7225 13095 7425 13170
rect 7225 13055 7305 13095
rect 7345 13055 7425 13095
rect 7225 12970 7425 13055
rect 7575 13095 7775 13170
rect 7575 13055 7655 13095
rect 7695 13055 7775 13095
rect 7575 12970 7775 13055
rect 7925 13095 8125 13170
rect 7925 13055 8005 13095
rect 8045 13055 8125 13095
rect 7925 12970 8125 13055
rect 8275 13095 8475 13170
rect 8275 13055 8355 13095
rect 8395 13055 8475 13095
rect 8275 12970 8475 13055
rect 8625 13095 8825 13170
rect 8625 13055 8705 13095
rect 8745 13055 8825 13095
rect 8625 12970 8825 13055
rect 8975 13095 9175 13170
rect 8975 13055 9055 13095
rect 9095 13055 9175 13095
rect 8975 12970 9175 13055
rect 9325 13095 9525 13170
rect 9325 13055 9405 13095
rect 9445 13055 9525 13095
rect 9325 12970 9525 13055
rect 9675 13095 9875 13170
rect 9675 13055 9755 13095
rect 9795 13055 9875 13095
rect 9675 12970 9875 13055
rect 10025 13095 10225 13170
rect 10025 13055 10105 13095
rect 10145 13055 10225 13095
rect 10025 12970 10225 13055
rect 10375 13095 10575 13170
rect 10375 13055 10455 13095
rect 10495 13055 10575 13095
rect 10375 12970 10575 13055
rect 6875 12745 7075 12820
rect 6875 12705 6955 12745
rect 6995 12705 7075 12745
rect 6875 12620 7075 12705
rect 7225 12745 7425 12820
rect 7225 12705 7305 12745
rect 7345 12705 7425 12745
rect 7225 12620 7425 12705
rect 7575 12745 7775 12820
rect 7575 12705 7655 12745
rect 7695 12705 7775 12745
rect 7575 12620 7775 12705
rect 7925 12745 8125 12820
rect 7925 12705 8005 12745
rect 8045 12705 8125 12745
rect 7925 12620 8125 12705
rect 8275 12745 8475 12820
rect 8275 12705 8355 12745
rect 8395 12705 8475 12745
rect 8275 12620 8475 12705
rect 8625 12745 8825 12820
rect 8625 12705 8705 12745
rect 8745 12705 8825 12745
rect 8625 12620 8825 12705
rect 8975 12745 9175 12820
rect 8975 12705 9055 12745
rect 9095 12705 9175 12745
rect 8975 12620 9175 12705
rect 9325 12745 9525 12820
rect 9325 12705 9405 12745
rect 9445 12705 9525 12745
rect 9325 12620 9525 12705
rect 9675 12745 9875 12820
rect 9675 12705 9755 12745
rect 9795 12705 9875 12745
rect 9675 12620 9875 12705
rect 10025 12745 10225 12820
rect 10025 12705 10105 12745
rect 10145 12705 10225 12745
rect 10025 12620 10225 12705
rect 10375 12745 10575 12820
rect 10375 12705 10455 12745
rect 10495 12705 10575 12745
rect 10375 12620 10575 12705
rect 6875 12395 7075 12470
rect 6875 12355 6955 12395
rect 6995 12355 7075 12395
rect 6875 12270 7075 12355
rect 7225 12395 7425 12470
rect 7225 12355 7305 12395
rect 7345 12355 7425 12395
rect 7225 12270 7425 12355
rect 7575 12395 7775 12470
rect 7575 12355 7655 12395
rect 7695 12355 7775 12395
rect 7575 12270 7775 12355
rect 7925 12395 8125 12470
rect 7925 12355 8005 12395
rect 8045 12355 8125 12395
rect 7925 12270 8125 12355
rect 8275 12395 8475 12470
rect 8275 12355 8355 12395
rect 8395 12355 8475 12395
rect 8275 12270 8475 12355
rect 8625 12395 8825 12470
rect 8625 12355 8705 12395
rect 8745 12355 8825 12395
rect 8625 12270 8825 12355
rect 8975 12395 9175 12470
rect 8975 12355 9055 12395
rect 9095 12355 9175 12395
rect 8975 12270 9175 12355
rect 9325 12395 9525 12470
rect 9325 12355 9405 12395
rect 9445 12355 9525 12395
rect 9325 12270 9525 12355
rect 9675 12395 9875 12470
rect 9675 12355 9755 12395
rect 9795 12355 9875 12395
rect 9675 12270 9875 12355
rect 10025 12395 10225 12470
rect 10025 12355 10105 12395
rect 10145 12355 10225 12395
rect 10025 12270 10225 12355
rect 10375 12395 10575 12470
rect 10375 12355 10455 12395
rect 10495 12355 10575 12395
rect 10375 12270 10575 12355
rect 6875 12045 7075 12120
rect 6875 12005 6955 12045
rect 6995 12005 7075 12045
rect 6875 11920 7075 12005
rect 7225 12045 7425 12120
rect 7225 12005 7305 12045
rect 7345 12005 7425 12045
rect 7225 11920 7425 12005
rect 7575 12045 7775 12120
rect 7575 12005 7655 12045
rect 7695 12005 7775 12045
rect 7575 11920 7775 12005
rect 7925 12045 8125 12120
rect 7925 12005 8005 12045
rect 8045 12005 8125 12045
rect 7925 11920 8125 12005
rect 8275 12045 8475 12120
rect 8275 12005 8355 12045
rect 8395 12005 8475 12045
rect 8275 11920 8475 12005
rect 8625 12045 8825 12120
rect 8625 12005 8705 12045
rect 8745 12005 8825 12045
rect 8625 11920 8825 12005
rect 8975 12045 9175 12120
rect 8975 12005 9055 12045
rect 9095 12005 9175 12045
rect 8975 11920 9175 12005
rect 9325 12045 9525 12120
rect 9325 12005 9405 12045
rect 9445 12005 9525 12045
rect 9325 11920 9525 12005
rect 9675 12045 9875 12120
rect 9675 12005 9755 12045
rect 9795 12005 9875 12045
rect 9675 11920 9875 12005
rect 10025 12045 10225 12120
rect 10025 12005 10105 12045
rect 10145 12005 10225 12045
rect 10025 11920 10225 12005
rect 10375 12045 10575 12120
rect 10375 12005 10455 12045
rect 10495 12005 10575 12045
rect 10375 11920 10575 12005
rect 6875 11695 7075 11770
rect 6875 11655 6955 11695
rect 6995 11655 7075 11695
rect 6875 11570 7075 11655
rect 7225 11695 7425 11770
rect 7225 11655 7305 11695
rect 7345 11655 7425 11695
rect 7225 11570 7425 11655
rect 7575 11695 7775 11770
rect 7575 11655 7655 11695
rect 7695 11655 7775 11695
rect 7575 11570 7775 11655
rect 7925 11695 8125 11770
rect 7925 11655 8005 11695
rect 8045 11655 8125 11695
rect 7925 11570 8125 11655
rect 8275 11695 8475 11770
rect 8275 11655 8355 11695
rect 8395 11655 8475 11695
rect 8275 11570 8475 11655
rect 8625 11695 8825 11770
rect 8625 11655 8705 11695
rect 8745 11655 8825 11695
rect 8625 11570 8825 11655
rect 8975 11695 9175 11770
rect 8975 11655 9055 11695
rect 9095 11655 9175 11695
rect 8975 11570 9175 11655
rect 9325 11695 9525 11770
rect 9325 11655 9405 11695
rect 9445 11655 9525 11695
rect 9325 11570 9525 11655
rect 9675 11695 9875 11770
rect 9675 11655 9755 11695
rect 9795 11655 9875 11695
rect 9675 11570 9875 11655
rect 10025 11695 10225 11770
rect 10025 11655 10105 11695
rect 10145 11655 10225 11695
rect 10025 11570 10225 11655
rect 10375 11695 10575 11770
rect 10375 11655 10455 11695
rect 10495 11655 10575 11695
rect 10375 11570 10575 11655
rect 6875 11345 7075 11420
rect 6875 11305 6955 11345
rect 6995 11305 7075 11345
rect 6875 11220 7075 11305
rect 7225 11345 7425 11420
rect 7225 11305 7305 11345
rect 7345 11305 7425 11345
rect 7225 11220 7425 11305
rect 7575 11345 7775 11420
rect 7575 11305 7655 11345
rect 7695 11305 7775 11345
rect 7575 11220 7775 11305
rect 7925 11345 8125 11420
rect 7925 11305 8005 11345
rect 8045 11305 8125 11345
rect 7925 11220 8125 11305
rect 8275 11345 8475 11420
rect 8275 11305 8355 11345
rect 8395 11305 8475 11345
rect 8275 11220 8475 11305
rect 8625 11345 8825 11420
rect 8625 11305 8705 11345
rect 8745 11305 8825 11345
rect 8625 11220 8825 11305
rect 8975 11345 9175 11420
rect 8975 11305 9055 11345
rect 9095 11305 9175 11345
rect 8975 11220 9175 11305
rect 9325 11345 9525 11420
rect 9325 11305 9405 11345
rect 9445 11305 9525 11345
rect 9325 11220 9525 11305
rect 9675 11345 9875 11420
rect 9675 11305 9755 11345
rect 9795 11305 9875 11345
rect 9675 11220 9875 11305
rect 10025 11345 10225 11420
rect 10025 11305 10105 11345
rect 10145 11305 10225 11345
rect 10025 11220 10225 11305
rect 10375 11345 10575 11420
rect 10375 11305 10455 11345
rect 10495 11305 10575 11345
rect 10375 11220 10575 11305
rect 6875 10995 7075 11070
rect 6875 10955 6955 10995
rect 6995 10955 7075 10995
rect 6875 10870 7075 10955
rect 7225 10995 7425 11070
rect 7225 10955 7305 10995
rect 7345 10955 7425 10995
rect 7225 10870 7425 10955
rect 7575 10995 7775 11070
rect 7575 10955 7655 10995
rect 7695 10955 7775 10995
rect 7575 10870 7775 10955
rect 7925 10995 8125 11070
rect 7925 10955 8005 10995
rect 8045 10955 8125 10995
rect 7925 10870 8125 10955
rect 8275 10995 8475 11070
rect 8275 10955 8355 10995
rect 8395 10955 8475 10995
rect 8275 10870 8475 10955
rect 8625 10995 8825 11070
rect 8625 10955 8705 10995
rect 8745 10955 8825 10995
rect 8625 10870 8825 10955
rect 8975 10995 9175 11070
rect 8975 10955 9055 10995
rect 9095 10955 9175 10995
rect 8975 10870 9175 10955
rect 9325 10995 9525 11070
rect 9325 10955 9405 10995
rect 9445 10955 9525 10995
rect 9325 10870 9525 10955
rect 9675 10995 9875 11070
rect 9675 10955 9755 10995
rect 9795 10955 9875 10995
rect 9675 10870 9875 10955
rect 10025 10995 10225 11070
rect 10025 10955 10105 10995
rect 10145 10955 10225 10995
rect 10025 10870 10225 10955
rect 10375 10995 10575 11070
rect 10375 10955 10455 10995
rect 10495 10955 10575 10995
rect 10375 10870 10575 10955
rect 6875 10645 7075 10720
rect 6875 10605 6955 10645
rect 6995 10605 7075 10645
rect 6875 10520 7075 10605
rect 7225 10645 7425 10720
rect 7225 10605 7305 10645
rect 7345 10605 7425 10645
rect 7225 10520 7425 10605
rect 7575 10645 7775 10720
rect 7575 10605 7655 10645
rect 7695 10605 7775 10645
rect 7575 10520 7775 10605
rect 7925 10645 8125 10720
rect 7925 10605 8005 10645
rect 8045 10605 8125 10645
rect 7925 10520 8125 10605
rect 8275 10645 8475 10720
rect 8275 10605 8355 10645
rect 8395 10605 8475 10645
rect 8275 10520 8475 10605
rect 8625 10645 8825 10720
rect 8625 10605 8705 10645
rect 8745 10605 8825 10645
rect 8625 10520 8825 10605
rect 8975 10645 9175 10720
rect 8975 10605 9055 10645
rect 9095 10605 9175 10645
rect 8975 10520 9175 10605
rect 9325 10645 9525 10720
rect 9325 10605 9405 10645
rect 9445 10605 9525 10645
rect 9325 10520 9525 10605
rect 9675 10645 9875 10720
rect 9675 10605 9755 10645
rect 9795 10605 9875 10645
rect 9675 10520 9875 10605
rect 10025 10645 10225 10720
rect 10025 10605 10105 10645
rect 10145 10605 10225 10645
rect 10025 10520 10225 10605
rect 10375 10645 10575 10720
rect 10375 10605 10455 10645
rect 10495 10605 10575 10645
rect 10375 10520 10575 10605
rect 6875 10295 7075 10370
rect 6875 10255 6955 10295
rect 6995 10255 7075 10295
rect 6875 10170 7075 10255
rect 7225 10295 7425 10370
rect 7225 10255 7305 10295
rect 7345 10255 7425 10295
rect 7225 10170 7425 10255
rect 7575 10295 7775 10370
rect 7575 10255 7655 10295
rect 7695 10255 7775 10295
rect 7575 10170 7775 10255
rect 7925 10295 8125 10370
rect 7925 10255 8005 10295
rect 8045 10255 8125 10295
rect 7925 10170 8125 10255
rect 8275 10295 8475 10370
rect 8275 10255 8355 10295
rect 8395 10255 8475 10295
rect 8275 10170 8475 10255
rect 8625 10295 8825 10370
rect 8625 10255 8705 10295
rect 8745 10255 8825 10295
rect 8625 10170 8825 10255
rect 8975 10295 9175 10370
rect 8975 10255 9055 10295
rect 9095 10255 9175 10295
rect 8975 10170 9175 10255
rect 9325 10295 9525 10370
rect 9325 10255 9405 10295
rect 9445 10255 9525 10295
rect 9325 10170 9525 10255
rect 9675 10295 9875 10370
rect 9675 10255 9755 10295
rect 9795 10255 9875 10295
rect 9675 10170 9875 10255
rect 10025 10295 10225 10370
rect 10025 10255 10105 10295
rect 10145 10255 10225 10295
rect 10025 10170 10225 10255
rect 10375 10295 10575 10370
rect 10375 10255 10455 10295
rect 10495 10255 10575 10295
rect 10375 10170 10575 10255
rect 6875 9945 7075 10020
rect 6875 9905 6955 9945
rect 6995 9905 7075 9945
rect 6875 9820 7075 9905
rect 7225 9945 7425 10020
rect 7225 9905 7305 9945
rect 7345 9905 7425 9945
rect 7225 9820 7425 9905
rect 7575 9945 7775 10020
rect 7575 9905 7655 9945
rect 7695 9905 7775 9945
rect 7575 9820 7775 9905
rect 7925 9945 8125 10020
rect 7925 9905 8005 9945
rect 8045 9905 8125 9945
rect 7925 9820 8125 9905
rect 8275 9945 8475 10020
rect 8275 9905 8355 9945
rect 8395 9905 8475 9945
rect 8275 9820 8475 9905
rect 8625 9945 8825 10020
rect 8625 9905 8705 9945
rect 8745 9905 8825 9945
rect 8625 9820 8825 9905
rect 8975 9945 9175 10020
rect 8975 9905 9055 9945
rect 9095 9905 9175 9945
rect 8975 9820 9175 9905
rect 9325 9945 9525 10020
rect 9325 9905 9405 9945
rect 9445 9905 9525 9945
rect 9325 9820 9525 9905
rect 9675 9945 9875 10020
rect 9675 9905 9755 9945
rect 9795 9905 9875 9945
rect 9675 9820 9875 9905
rect 10025 9945 10225 10020
rect 10025 9905 10105 9945
rect 10145 9905 10225 9945
rect 10025 9820 10225 9905
rect 10375 9945 10575 10020
rect 10375 9905 10455 9945
rect 10495 9905 10575 9945
rect 10375 9820 10575 9905
rect 6875 9595 7075 9670
rect 6875 9555 6955 9595
rect 6995 9555 7075 9595
rect 6875 9470 7075 9555
rect 7225 9595 7425 9670
rect 7225 9555 7305 9595
rect 7345 9555 7425 9595
rect 7225 9470 7425 9555
rect 7575 9595 7775 9670
rect 7575 9555 7655 9595
rect 7695 9555 7775 9595
rect 7575 9470 7775 9555
rect 7925 9595 8125 9670
rect 7925 9555 8005 9595
rect 8045 9555 8125 9595
rect 7925 9470 8125 9555
rect 8275 9595 8475 9670
rect 8275 9555 8355 9595
rect 8395 9555 8475 9595
rect 8275 9470 8475 9555
rect 8625 9595 8825 9670
rect 8625 9555 8705 9595
rect 8745 9555 8825 9595
rect 8625 9470 8825 9555
rect 8975 9595 9175 9670
rect 8975 9555 9055 9595
rect 9095 9555 9175 9595
rect 8975 9470 9175 9555
rect 9325 9595 9525 9670
rect 9325 9555 9405 9595
rect 9445 9555 9525 9595
rect 9325 9470 9525 9555
rect 9675 9595 9875 9670
rect 9675 9555 9755 9595
rect 9795 9555 9875 9595
rect 9675 9470 9875 9555
rect 10025 9595 10225 9670
rect 10025 9555 10105 9595
rect 10145 9555 10225 9595
rect 10025 9470 10225 9555
rect 10375 9595 10575 9670
rect 10375 9555 10455 9595
rect 10495 9555 10575 9595
rect 10375 9470 10575 9555
rect 6875 9245 7075 9320
rect 6875 9205 6955 9245
rect 6995 9205 7075 9245
rect 6875 9120 7075 9205
rect 7225 9245 7425 9320
rect 7225 9205 7305 9245
rect 7345 9205 7425 9245
rect 7225 9120 7425 9205
rect 7575 9245 7775 9320
rect 7575 9205 7655 9245
rect 7695 9205 7775 9245
rect 7575 9120 7775 9205
rect 7925 9245 8125 9320
rect 7925 9205 8005 9245
rect 8045 9205 8125 9245
rect 7925 9120 8125 9205
rect 8275 9245 8475 9320
rect 8275 9205 8355 9245
rect 8395 9205 8475 9245
rect 8275 9120 8475 9205
rect 8625 9245 8825 9320
rect 8625 9205 8705 9245
rect 8745 9205 8825 9245
rect 8625 9120 8825 9205
rect 8975 9245 9175 9320
rect 8975 9205 9055 9245
rect 9095 9205 9175 9245
rect 8975 9120 9175 9205
rect 9325 9245 9525 9320
rect 9325 9205 9405 9245
rect 9445 9205 9525 9245
rect 9325 9120 9525 9205
rect 9675 9245 9875 9320
rect 9675 9205 9755 9245
rect 9795 9205 9875 9245
rect 9675 9120 9875 9205
rect 10025 9245 10225 9320
rect 10025 9205 10105 9245
rect 10145 9205 10225 9245
rect 10025 9120 10225 9205
rect 10375 9245 10575 9320
rect 10375 9205 10455 9245
rect 10495 9205 10575 9245
rect 10375 9120 10575 9205
rect 6875 8895 7075 8970
rect 6875 8855 6955 8895
rect 6995 8855 7075 8895
rect 6875 8770 7075 8855
rect 7225 8895 7425 8970
rect 7225 8855 7305 8895
rect 7345 8855 7425 8895
rect 7225 8770 7425 8855
rect 7575 8895 7775 8970
rect 7575 8855 7655 8895
rect 7695 8855 7775 8895
rect 7575 8770 7775 8855
rect 7925 8895 8125 8970
rect 7925 8855 8005 8895
rect 8045 8855 8125 8895
rect 7925 8770 8125 8855
rect 8275 8895 8475 8970
rect 8275 8855 8355 8895
rect 8395 8855 8475 8895
rect 8275 8770 8475 8855
rect 8625 8895 8825 8970
rect 8625 8855 8705 8895
rect 8745 8855 8825 8895
rect 8625 8770 8825 8855
rect 8975 8895 9175 8970
rect 8975 8855 9055 8895
rect 9095 8855 9175 8895
rect 8975 8770 9175 8855
rect 9325 8895 9525 8970
rect 9325 8855 9405 8895
rect 9445 8855 9525 8895
rect 9325 8770 9525 8855
rect 9675 8895 9875 8970
rect 9675 8855 9755 8895
rect 9795 8855 9875 8895
rect 9675 8770 9875 8855
rect 10025 8895 10225 8970
rect 10025 8855 10105 8895
rect 10145 8855 10225 8895
rect 10025 8770 10225 8855
rect 10375 8895 10575 8970
rect 10375 8855 10455 8895
rect 10495 8855 10575 8895
rect 10375 8770 10575 8855
rect 6875 8545 7075 8620
rect 6875 8505 6955 8545
rect 6995 8505 7075 8545
rect 6875 8420 7075 8505
rect 7225 8545 7425 8620
rect 7225 8505 7305 8545
rect 7345 8505 7425 8545
rect 7225 8420 7425 8505
rect 7575 8545 7775 8620
rect 7575 8505 7655 8545
rect 7695 8505 7775 8545
rect 7575 8420 7775 8505
rect 7925 8545 8125 8620
rect 7925 8505 8005 8545
rect 8045 8505 8125 8545
rect 7925 8420 8125 8505
rect 8275 8545 8475 8620
rect 8275 8505 8355 8545
rect 8395 8505 8475 8545
rect 8275 8420 8475 8505
rect 8625 8545 8825 8620
rect 8625 8505 8705 8545
rect 8745 8505 8825 8545
rect 8625 8420 8825 8505
rect 8975 8545 9175 8620
rect 8975 8505 9055 8545
rect 9095 8505 9175 8545
rect 8975 8420 9175 8505
rect 9325 8545 9525 8620
rect 9325 8505 9405 8545
rect 9445 8505 9525 8545
rect 9325 8420 9525 8505
rect 9675 8545 9875 8620
rect 9675 8505 9755 8545
rect 9795 8505 9875 8545
rect 9675 8420 9875 8505
rect 10025 8545 10225 8620
rect 10025 8505 10105 8545
rect 10145 8505 10225 8545
rect 10025 8420 10225 8505
rect 10375 8545 10575 8620
rect 10375 8505 10455 8545
rect 10495 8505 10575 8545
rect 10375 8420 10575 8505
rect 6875 8195 7075 8270
rect 6875 8155 6955 8195
rect 6995 8155 7075 8195
rect 6875 8070 7075 8155
rect 7225 8195 7425 8270
rect 7225 8155 7305 8195
rect 7345 8155 7425 8195
rect 7225 8070 7425 8155
rect 7575 8195 7775 8270
rect 7575 8155 7655 8195
rect 7695 8155 7775 8195
rect 7575 8070 7775 8155
rect 7925 8195 8125 8270
rect 7925 8155 8005 8195
rect 8045 8155 8125 8195
rect 7925 8070 8125 8155
rect 8275 8195 8475 8270
rect 8275 8155 8355 8195
rect 8395 8155 8475 8195
rect 8275 8070 8475 8155
rect 8625 8195 8825 8270
rect 8625 8155 8705 8195
rect 8745 8155 8825 8195
rect 8625 8070 8825 8155
rect 8975 8195 9175 8270
rect 8975 8155 9055 8195
rect 9095 8155 9175 8195
rect 8975 8070 9175 8155
rect 9325 8195 9525 8270
rect 9325 8155 9405 8195
rect 9445 8155 9525 8195
rect 9325 8070 9525 8155
rect 9675 8195 9875 8270
rect 9675 8155 9755 8195
rect 9795 8155 9875 8195
rect 9675 8070 9875 8155
rect 10025 8195 10225 8270
rect 10025 8155 10105 8195
rect 10145 8155 10225 8195
rect 10025 8070 10225 8155
rect 10375 8195 10575 8270
rect 10375 8155 10455 8195
rect 10495 8155 10575 8195
rect 10375 8070 10575 8155
rect 6875 7845 7075 7920
rect 6875 7805 6955 7845
rect 6995 7805 7075 7845
rect 6875 7720 7075 7805
rect 7225 7845 7425 7920
rect 7225 7805 7305 7845
rect 7345 7805 7425 7845
rect 7225 7720 7425 7805
rect 7575 7845 7775 7920
rect 7575 7805 7655 7845
rect 7695 7805 7775 7845
rect 7575 7720 7775 7805
rect 7925 7845 8125 7920
rect 7925 7805 8005 7845
rect 8045 7805 8125 7845
rect 7925 7720 8125 7805
rect 8275 7845 8475 7920
rect 8275 7805 8355 7845
rect 8395 7805 8475 7845
rect 8275 7720 8475 7805
rect 8625 7845 8825 7920
rect 8625 7805 8705 7845
rect 8745 7805 8825 7845
rect 8625 7720 8825 7805
rect 8975 7845 9175 7920
rect 8975 7805 9055 7845
rect 9095 7805 9175 7845
rect 8975 7720 9175 7805
rect 9325 7845 9525 7920
rect 9325 7805 9405 7845
rect 9445 7805 9525 7845
rect 9325 7720 9525 7805
rect 9675 7845 9875 7920
rect 9675 7805 9755 7845
rect 9795 7805 9875 7845
rect 9675 7720 9875 7805
rect 10025 7845 10225 7920
rect 10025 7805 10105 7845
rect 10145 7805 10225 7845
rect 10025 7720 10225 7805
rect 10375 7845 10575 7920
rect 10375 7805 10455 7845
rect 10495 7805 10575 7845
rect 10375 7720 10575 7805
rect 6875 7495 7075 7570
rect 6875 7455 6955 7495
rect 6995 7455 7075 7495
rect 6875 7370 7075 7455
rect 7225 7495 7425 7570
rect 7225 7455 7305 7495
rect 7345 7455 7425 7495
rect 7225 7370 7425 7455
rect 7575 7495 7775 7570
rect 7575 7455 7655 7495
rect 7695 7455 7775 7495
rect 7575 7370 7775 7455
rect 7925 7495 8125 7570
rect 7925 7455 8005 7495
rect 8045 7455 8125 7495
rect 7925 7370 8125 7455
rect 8275 7495 8475 7570
rect 8275 7455 8355 7495
rect 8395 7455 8475 7495
rect 8275 7370 8475 7455
rect 8625 7495 8825 7570
rect 8625 7455 8705 7495
rect 8745 7455 8825 7495
rect 8625 7370 8825 7455
rect 8975 7495 9175 7570
rect 8975 7455 9055 7495
rect 9095 7455 9175 7495
rect 8975 7370 9175 7455
rect 9325 7495 9525 7570
rect 9325 7455 9405 7495
rect 9445 7455 9525 7495
rect 9325 7370 9525 7455
rect 9675 7495 9875 7570
rect 9675 7455 9755 7495
rect 9795 7455 9875 7495
rect 9675 7370 9875 7455
rect 10025 7495 10225 7570
rect 10025 7455 10105 7495
rect 10145 7455 10225 7495
rect 10025 7370 10225 7455
rect 10375 7495 10575 7570
rect 10375 7455 10455 7495
rect 10495 7455 10575 7495
rect 10375 7370 10575 7455
rect 6875 7145 7075 7220
rect 6875 7105 6955 7145
rect 6995 7105 7075 7145
rect 6875 7020 7075 7105
rect 7225 7145 7425 7220
rect 7225 7105 7305 7145
rect 7345 7105 7425 7145
rect 7225 7020 7425 7105
rect 7575 7145 7775 7220
rect 7575 7105 7655 7145
rect 7695 7105 7775 7145
rect 7575 7020 7775 7105
rect 7925 7145 8125 7220
rect 7925 7105 8005 7145
rect 8045 7105 8125 7145
rect 7925 7020 8125 7105
rect 8275 7145 8475 7220
rect 8275 7105 8355 7145
rect 8395 7105 8475 7145
rect 8275 7020 8475 7105
rect 8625 7145 8825 7220
rect 8625 7105 8705 7145
rect 8745 7105 8825 7145
rect 8625 7020 8825 7105
rect 8975 7145 9175 7220
rect 8975 7105 9055 7145
rect 9095 7105 9175 7145
rect 8975 7020 9175 7105
rect 9325 7145 9525 7220
rect 9325 7105 9405 7145
rect 9445 7105 9525 7145
rect 9325 7020 9525 7105
rect 9675 7145 9875 7220
rect 9675 7105 9755 7145
rect 9795 7105 9875 7145
rect 9675 7020 9875 7105
rect 10025 7145 10225 7220
rect 10025 7105 10105 7145
rect 10145 7105 10225 7145
rect 10025 7020 10225 7105
rect 10375 7145 10575 7220
rect 10375 7105 10455 7145
rect 10495 7105 10575 7145
rect 10375 7020 10575 7105
rect 6875 6795 7075 6870
rect 6875 6755 6955 6795
rect 6995 6755 7075 6795
rect 6875 6670 7075 6755
rect 7225 6795 7425 6870
rect 7225 6755 7305 6795
rect 7345 6755 7425 6795
rect 7225 6670 7425 6755
rect 7575 6795 7775 6870
rect 7575 6755 7655 6795
rect 7695 6755 7775 6795
rect 7575 6670 7775 6755
rect 7925 6795 8125 6870
rect 7925 6755 8005 6795
rect 8045 6755 8125 6795
rect 7925 6670 8125 6755
rect 8275 6795 8475 6870
rect 8275 6755 8355 6795
rect 8395 6755 8475 6795
rect 8275 6670 8475 6755
rect 8625 6795 8825 6870
rect 8625 6755 8705 6795
rect 8745 6755 8825 6795
rect 8625 6670 8825 6755
rect 8975 6795 9175 6870
rect 8975 6755 9055 6795
rect 9095 6755 9175 6795
rect 8975 6670 9175 6755
rect 9325 6795 9525 6870
rect 9325 6755 9405 6795
rect 9445 6755 9525 6795
rect 9325 6670 9525 6755
rect 9675 6795 9875 6870
rect 9675 6755 9755 6795
rect 9795 6755 9875 6795
rect 9675 6670 9875 6755
rect 10025 6795 10225 6870
rect 10025 6755 10105 6795
rect 10145 6755 10225 6795
rect 10025 6670 10225 6755
rect 10375 6795 10575 6870
rect 10375 6755 10455 6795
rect 10495 6755 10575 6795
rect 10375 6670 10575 6755
<< mimcapcontact >>
rect 6955 14805 6995 14845
rect 7305 14805 7345 14845
rect 7655 14805 7695 14845
rect 8005 14805 8045 14845
rect 8355 14805 8395 14845
rect 8705 14805 8745 14845
rect 9055 14805 9095 14845
rect 9405 14805 9445 14845
rect 9755 14805 9795 14845
rect 10105 14805 10145 14845
rect 10455 14805 10495 14845
rect 6955 14455 6995 14495
rect 7305 14455 7345 14495
rect 7655 14455 7695 14495
rect 8005 14455 8045 14495
rect 8355 14455 8395 14495
rect 8705 14455 8745 14495
rect 9055 14455 9095 14495
rect 9405 14455 9445 14495
rect 9755 14455 9795 14495
rect 10105 14455 10145 14495
rect 10455 14455 10495 14495
rect 6955 14105 6995 14145
rect 7305 14105 7345 14145
rect 7655 14105 7695 14145
rect 8005 14105 8045 14145
rect 8355 14105 8395 14145
rect 8705 14105 8745 14145
rect 9055 14105 9095 14145
rect 9405 14105 9445 14145
rect 9755 14105 9795 14145
rect 10105 14105 10145 14145
rect 10455 14105 10495 14145
rect 6955 13755 6995 13795
rect 7305 13755 7345 13795
rect 7655 13755 7695 13795
rect 8005 13755 8045 13795
rect 8355 13755 8395 13795
rect 8705 13755 8745 13795
rect 9055 13755 9095 13795
rect 9405 13755 9445 13795
rect 9755 13755 9795 13795
rect 10105 13755 10145 13795
rect 10455 13755 10495 13795
rect 6955 13405 6995 13445
rect 7305 13405 7345 13445
rect 7655 13405 7695 13445
rect 8005 13405 8045 13445
rect 8355 13405 8395 13445
rect 8705 13405 8745 13445
rect 9055 13405 9095 13445
rect 9405 13405 9445 13445
rect 9755 13405 9795 13445
rect 10105 13405 10145 13445
rect 10455 13405 10495 13445
rect 6955 13055 6995 13095
rect 7305 13055 7345 13095
rect 7655 13055 7695 13095
rect 8005 13055 8045 13095
rect 8355 13055 8395 13095
rect 8705 13055 8745 13095
rect 9055 13055 9095 13095
rect 9405 13055 9445 13095
rect 9755 13055 9795 13095
rect 10105 13055 10145 13095
rect 10455 13055 10495 13095
rect 6955 12705 6995 12745
rect 7305 12705 7345 12745
rect 7655 12705 7695 12745
rect 8005 12705 8045 12745
rect 8355 12705 8395 12745
rect 8705 12705 8745 12745
rect 9055 12705 9095 12745
rect 9405 12705 9445 12745
rect 9755 12705 9795 12745
rect 10105 12705 10145 12745
rect 10455 12705 10495 12745
rect 6955 12355 6995 12395
rect 7305 12355 7345 12395
rect 7655 12355 7695 12395
rect 8005 12355 8045 12395
rect 8355 12355 8395 12395
rect 8705 12355 8745 12395
rect 9055 12355 9095 12395
rect 9405 12355 9445 12395
rect 9755 12355 9795 12395
rect 10105 12355 10145 12395
rect 10455 12355 10495 12395
rect 6955 12005 6995 12045
rect 7305 12005 7345 12045
rect 7655 12005 7695 12045
rect 8005 12005 8045 12045
rect 8355 12005 8395 12045
rect 8705 12005 8745 12045
rect 9055 12005 9095 12045
rect 9405 12005 9445 12045
rect 9755 12005 9795 12045
rect 10105 12005 10145 12045
rect 10455 12005 10495 12045
rect 6955 11655 6995 11695
rect 7305 11655 7345 11695
rect 7655 11655 7695 11695
rect 8005 11655 8045 11695
rect 8355 11655 8395 11695
rect 8705 11655 8745 11695
rect 9055 11655 9095 11695
rect 9405 11655 9445 11695
rect 9755 11655 9795 11695
rect 10105 11655 10145 11695
rect 10455 11655 10495 11695
rect 6955 11305 6995 11345
rect 7305 11305 7345 11345
rect 7655 11305 7695 11345
rect 8005 11305 8045 11345
rect 8355 11305 8395 11345
rect 8705 11305 8745 11345
rect 9055 11305 9095 11345
rect 9405 11305 9445 11345
rect 9755 11305 9795 11345
rect 10105 11305 10145 11345
rect 10455 11305 10495 11345
rect 6955 10955 6995 10995
rect 7305 10955 7345 10995
rect 7655 10955 7695 10995
rect 8005 10955 8045 10995
rect 8355 10955 8395 10995
rect 8705 10955 8745 10995
rect 9055 10955 9095 10995
rect 9405 10955 9445 10995
rect 9755 10955 9795 10995
rect 10105 10955 10145 10995
rect 10455 10955 10495 10995
rect 6955 10605 6995 10645
rect 7305 10605 7345 10645
rect 7655 10605 7695 10645
rect 8005 10605 8045 10645
rect 8355 10605 8395 10645
rect 8705 10605 8745 10645
rect 9055 10605 9095 10645
rect 9405 10605 9445 10645
rect 9755 10605 9795 10645
rect 10105 10605 10145 10645
rect 10455 10605 10495 10645
rect 6955 10255 6995 10295
rect 7305 10255 7345 10295
rect 7655 10255 7695 10295
rect 8005 10255 8045 10295
rect 8355 10255 8395 10295
rect 8705 10255 8745 10295
rect 9055 10255 9095 10295
rect 9405 10255 9445 10295
rect 9755 10255 9795 10295
rect 10105 10255 10145 10295
rect 10455 10255 10495 10295
rect 6955 9905 6995 9945
rect 7305 9905 7345 9945
rect 7655 9905 7695 9945
rect 8005 9905 8045 9945
rect 8355 9905 8395 9945
rect 8705 9905 8745 9945
rect 9055 9905 9095 9945
rect 9405 9905 9445 9945
rect 9755 9905 9795 9945
rect 10105 9905 10145 9945
rect 10455 9905 10495 9945
rect 6955 9555 6995 9595
rect 7305 9555 7345 9595
rect 7655 9555 7695 9595
rect 8005 9555 8045 9595
rect 8355 9555 8395 9595
rect 8705 9555 8745 9595
rect 9055 9555 9095 9595
rect 9405 9555 9445 9595
rect 9755 9555 9795 9595
rect 10105 9555 10145 9595
rect 10455 9555 10495 9595
rect 6955 9205 6995 9245
rect 7305 9205 7345 9245
rect 7655 9205 7695 9245
rect 8005 9205 8045 9245
rect 8355 9205 8395 9245
rect 8705 9205 8745 9245
rect 9055 9205 9095 9245
rect 9405 9205 9445 9245
rect 9755 9205 9795 9245
rect 10105 9205 10145 9245
rect 10455 9205 10495 9245
rect 6955 8855 6995 8895
rect 7305 8855 7345 8895
rect 7655 8855 7695 8895
rect 8005 8855 8045 8895
rect 8355 8855 8395 8895
rect 8705 8855 8745 8895
rect 9055 8855 9095 8895
rect 9405 8855 9445 8895
rect 9755 8855 9795 8895
rect 10105 8855 10145 8895
rect 10455 8855 10495 8895
rect 6955 8505 6995 8545
rect 7305 8505 7345 8545
rect 7655 8505 7695 8545
rect 8005 8505 8045 8545
rect 8355 8505 8395 8545
rect 8705 8505 8745 8545
rect 9055 8505 9095 8545
rect 9405 8505 9445 8545
rect 9755 8505 9795 8545
rect 10105 8505 10145 8545
rect 10455 8505 10495 8545
rect 6955 8155 6995 8195
rect 7305 8155 7345 8195
rect 7655 8155 7695 8195
rect 8005 8155 8045 8195
rect 8355 8155 8395 8195
rect 8705 8155 8745 8195
rect 9055 8155 9095 8195
rect 9405 8155 9445 8195
rect 9755 8155 9795 8195
rect 10105 8155 10145 8195
rect 10455 8155 10495 8195
rect 6955 7805 6995 7845
rect 7305 7805 7345 7845
rect 7655 7805 7695 7845
rect 8005 7805 8045 7845
rect 8355 7805 8395 7845
rect 8705 7805 8745 7845
rect 9055 7805 9095 7845
rect 9405 7805 9445 7845
rect 9755 7805 9795 7845
rect 10105 7805 10145 7845
rect 10455 7805 10495 7845
rect 6955 7455 6995 7495
rect 7305 7455 7345 7495
rect 7655 7455 7695 7495
rect 8005 7455 8045 7495
rect 8355 7455 8395 7495
rect 8705 7455 8745 7495
rect 9055 7455 9095 7495
rect 9405 7455 9445 7495
rect 9755 7455 9795 7495
rect 10105 7455 10145 7495
rect 10455 7455 10495 7495
rect 6955 7105 6995 7145
rect 7305 7105 7345 7145
rect 7655 7105 7695 7145
rect 8005 7105 8045 7145
rect 8355 7105 8395 7145
rect 8705 7105 8745 7145
rect 9055 7105 9095 7145
rect 9405 7105 9445 7145
rect 9755 7105 9795 7145
rect 10105 7105 10145 7145
rect 10455 7105 10495 7145
rect 6955 6755 6995 6795
rect 7305 6755 7345 6795
rect 7655 6755 7695 6795
rect 8005 6755 8045 6795
rect 8355 6755 8395 6795
rect 8705 6755 8745 6795
rect 9055 6755 9095 6795
rect 9405 6755 9445 6795
rect 9755 6755 9795 6795
rect 10105 6755 10145 6795
rect 10455 6755 10495 6795
<< metal4 >>
rect 2320 15415 11510 15425
rect 2320 15375 2330 15415
rect 2370 15375 6700 15415
rect 6740 15390 11510 15415
rect 6740 15375 10745 15390
rect 2320 15350 10745 15375
rect 2320 15310 2330 15350
rect 2370 15310 6700 15350
rect 6740 15340 10745 15350
rect 10795 15340 10840 15390
rect 10890 15340 10935 15390
rect 10985 15340 11035 15390
rect 11085 15340 11135 15390
rect 11185 15340 11235 15390
rect 11285 15340 11330 15390
rect 11380 15340 11425 15390
rect 11475 15340 11510 15390
rect 6740 15310 11510 15340
rect 2320 15300 11510 15310
rect 2320 15280 10745 15300
rect 2320 15240 2330 15280
rect 2370 15240 6700 15280
rect 6740 15250 10745 15280
rect 10795 15250 10840 15300
rect 10890 15250 10935 15300
rect 10985 15250 11035 15300
rect 11085 15250 11135 15300
rect 11185 15250 11235 15300
rect 11285 15250 11330 15300
rect 11380 15250 11425 15300
rect 11475 15250 11510 15300
rect 6740 15240 11510 15250
rect 2320 15210 11510 15240
rect 2320 15170 2330 15210
rect 2370 15170 6700 15210
rect 6740 15200 11510 15210
rect 6740 15170 10745 15200
rect 2320 15150 10745 15170
rect 10795 15150 10840 15200
rect 10890 15150 10935 15200
rect 10985 15150 11035 15200
rect 11085 15150 11135 15200
rect 11185 15150 11235 15200
rect 11285 15150 11330 15200
rect 11380 15150 11425 15200
rect 11475 15150 11510 15200
rect 2320 15140 11510 15150
rect 2320 15100 2330 15140
rect 2370 15100 6700 15140
rect 6740 15110 11510 15140
rect 6740 15100 10745 15110
rect 2320 15075 10745 15100
rect 2320 15035 2330 15075
rect 2370 15035 6700 15075
rect 6740 15060 10745 15075
rect 10795 15060 10840 15110
rect 10890 15060 10935 15110
rect 10985 15060 11035 15110
rect 11085 15060 11135 15110
rect 11185 15060 11235 15110
rect 11285 15060 11330 15110
rect 11380 15060 11425 15110
rect 11475 15060 11510 15110
rect 6740 15035 11510 15060
rect 2320 15025 11510 15035
rect 6950 14845 10500 14850
rect 6950 14805 6955 14845
rect 6995 14805 7305 14845
rect 7345 14805 7655 14845
rect 7695 14805 8005 14845
rect 8045 14805 8355 14845
rect 8395 14805 8705 14845
rect 8745 14805 9055 14845
rect 9095 14805 9405 14845
rect 9445 14805 9755 14845
rect 9795 14805 10105 14845
rect 10145 14805 10455 14845
rect 10495 14805 10500 14845
rect 6950 14800 10500 14805
rect 8700 14500 8750 14800
rect 6950 14495 10500 14500
rect 6950 14455 6955 14495
rect 6995 14455 7305 14495
rect 7345 14455 7655 14495
rect 7695 14455 8005 14495
rect 8045 14455 8355 14495
rect 8395 14455 8705 14495
rect 8745 14455 9055 14495
rect 9095 14455 9405 14495
rect 9445 14455 9755 14495
rect 9795 14455 10105 14495
rect 10145 14455 10455 14495
rect 10495 14455 10500 14495
rect 6950 14450 10500 14455
rect 8700 14150 8750 14450
rect 6950 14145 10500 14150
rect 6950 14105 6955 14145
rect 6995 14105 7305 14145
rect 7345 14105 7655 14145
rect 7695 14105 8005 14145
rect 8045 14105 8355 14145
rect 8395 14105 8705 14145
rect 8745 14105 9055 14145
rect 9095 14105 9405 14145
rect 9445 14105 9755 14145
rect 9795 14105 10105 14145
rect 10145 14105 10455 14145
rect 10495 14105 10500 14145
rect 6950 14100 10500 14105
rect 8700 13800 8750 14100
rect 6950 13795 10500 13800
rect 6950 13755 6955 13795
rect 6995 13755 7305 13795
rect 7345 13755 7655 13795
rect 7695 13755 8005 13795
rect 8045 13755 8355 13795
rect 8395 13755 8705 13795
rect 8745 13755 9055 13795
rect 9095 13755 9405 13795
rect 9445 13755 9755 13795
rect 9795 13755 10105 13795
rect 10145 13755 10455 13795
rect 10495 13755 10500 13795
rect 6950 13750 10500 13755
rect 8700 13450 8750 13750
rect 6950 13445 10500 13450
rect 6950 13405 6955 13445
rect 6995 13405 7305 13445
rect 7345 13405 7655 13445
rect 7695 13405 8005 13445
rect 8045 13405 8355 13445
rect 8395 13405 8705 13445
rect 8745 13405 9055 13445
rect 9095 13405 9405 13445
rect 9445 13405 9755 13445
rect 9795 13405 10105 13445
rect 10145 13405 10455 13445
rect 10495 13405 10500 13445
rect 6950 13400 10500 13405
rect 8700 13100 8750 13400
rect 6950 13095 10500 13100
rect 6950 13055 6955 13095
rect 6995 13055 7305 13095
rect 7345 13055 7655 13095
rect 7695 13055 8005 13095
rect 8045 13055 8355 13095
rect 8395 13055 8705 13095
rect 8745 13055 9055 13095
rect 9095 13055 9405 13095
rect 9445 13055 9755 13095
rect 9795 13055 10105 13095
rect 10145 13055 10455 13095
rect 10495 13055 10500 13095
rect 6950 13050 10500 13055
rect 8700 12750 8750 13050
rect 6950 12745 10500 12750
rect 6950 12705 6955 12745
rect 6995 12705 7305 12745
rect 7345 12705 7655 12745
rect 7695 12705 8005 12745
rect 8045 12705 8355 12745
rect 8395 12705 8705 12745
rect 8745 12705 9055 12745
rect 9095 12705 9405 12745
rect 9445 12705 9755 12745
rect 9795 12705 10105 12745
rect 10145 12705 10455 12745
rect 10495 12705 10500 12745
rect 6950 12700 10500 12705
rect 8700 12400 8750 12700
rect 6950 12395 10500 12400
rect 6950 12355 6955 12395
rect 6995 12355 7305 12395
rect 7345 12355 7655 12395
rect 7695 12355 8005 12395
rect 8045 12355 8355 12395
rect 8395 12355 8705 12395
rect 8745 12355 9055 12395
rect 9095 12355 9405 12395
rect 9445 12355 9755 12395
rect 9795 12355 10105 12395
rect 10145 12355 10455 12395
rect 10495 12355 10500 12395
rect 6950 12350 10500 12355
rect 8700 12050 8750 12350
rect 6950 12045 10500 12050
rect 6950 12005 6955 12045
rect 6995 12005 7305 12045
rect 7345 12005 7655 12045
rect 7695 12005 8005 12045
rect 8045 12005 8355 12045
rect 8395 12005 8705 12045
rect 8745 12005 9055 12045
rect 9095 12005 9405 12045
rect 9445 12005 9755 12045
rect 9795 12005 10105 12045
rect 10145 12005 10455 12045
rect 10495 12005 10500 12045
rect 6950 12000 10500 12005
rect 8700 11700 8750 12000
rect 6950 11695 10500 11700
rect 6950 11655 6955 11695
rect 6995 11655 7305 11695
rect 7345 11655 7655 11695
rect 7695 11655 8005 11695
rect 8045 11655 8355 11695
rect 8395 11655 8705 11695
rect 8745 11655 9055 11695
rect 9095 11655 9405 11695
rect 9445 11655 9755 11695
rect 9795 11655 10105 11695
rect 10145 11655 10455 11695
rect 10495 11655 10500 11695
rect 6950 11650 10500 11655
rect 8700 11350 8750 11650
rect 6950 11345 10500 11350
rect 6950 11305 6955 11345
rect 6995 11305 7305 11345
rect 7345 11305 7655 11345
rect 7695 11305 8005 11345
rect 8045 11305 8355 11345
rect 8395 11305 8705 11345
rect 8745 11305 9055 11345
rect 9095 11305 9405 11345
rect 9445 11305 9755 11345
rect 9795 11305 10105 11345
rect 10145 11305 10455 11345
rect 10495 11305 10500 11345
rect 6950 11300 10500 11305
rect 8700 11000 8750 11300
rect 6950 10995 10500 11000
rect 6950 10955 6955 10995
rect 6995 10955 7305 10995
rect 7345 10955 7655 10995
rect 7695 10955 8005 10995
rect 8045 10955 8355 10995
rect 8395 10955 8705 10995
rect 8745 10955 9055 10995
rect 9095 10955 9405 10995
rect 9445 10955 9755 10995
rect 9795 10955 10105 10995
rect 10145 10955 10455 10995
rect 10495 10955 10500 10995
rect 6950 10950 10500 10955
rect 8700 10650 8750 10950
rect 6950 10645 10500 10650
rect 6950 10605 6955 10645
rect 6995 10605 7305 10645
rect 7345 10605 7655 10645
rect 7695 10605 8005 10645
rect 8045 10605 8355 10645
rect 8395 10605 8705 10645
rect 8745 10605 9055 10645
rect 9095 10605 9405 10645
rect 9445 10605 9755 10645
rect 9795 10605 10105 10645
rect 10145 10605 10455 10645
rect 10495 10605 10500 10645
rect 6950 10600 10500 10605
rect 8700 10300 8750 10600
rect 6950 10295 10500 10300
rect 6950 10255 6955 10295
rect 6995 10255 7305 10295
rect 7345 10255 7655 10295
rect 7695 10255 8005 10295
rect 8045 10255 8355 10295
rect 8395 10255 8705 10295
rect 8745 10255 9055 10295
rect 9095 10255 9405 10295
rect 9445 10255 9755 10295
rect 9795 10255 10105 10295
rect 10145 10255 10455 10295
rect 10495 10255 10500 10295
rect 6950 10250 10500 10255
rect 8700 9950 8750 10250
rect 6950 9945 10500 9950
rect 6950 9905 6955 9945
rect 6995 9905 7305 9945
rect 7345 9905 7655 9945
rect 7695 9905 8005 9945
rect 8045 9905 8355 9945
rect 8395 9905 8705 9945
rect 8745 9905 9055 9945
rect 9095 9905 9405 9945
rect 9445 9905 9755 9945
rect 9795 9905 10105 9945
rect 10145 9905 10455 9945
rect 10495 9905 10500 9945
rect 6950 9900 10500 9905
rect 8700 9600 8750 9900
rect 6950 9595 10500 9600
rect 6950 9555 6955 9595
rect 6995 9555 7305 9595
rect 7345 9555 7655 9595
rect 7695 9555 8005 9595
rect 8045 9555 8355 9595
rect 8395 9555 8705 9595
rect 8745 9555 9055 9595
rect 9095 9555 9405 9595
rect 9445 9555 9755 9595
rect 9795 9555 10105 9595
rect 10145 9555 10455 9595
rect 10495 9555 10500 9595
rect 6950 9550 10500 9555
rect 8700 9250 8750 9550
rect 6950 9245 10500 9250
rect 6950 9205 6955 9245
rect 6995 9205 7305 9245
rect 7345 9205 7655 9245
rect 7695 9205 8005 9245
rect 8045 9205 8355 9245
rect 8395 9205 8705 9245
rect 8745 9205 9055 9245
rect 9095 9205 9405 9245
rect 9445 9205 9755 9245
rect 9795 9205 10105 9245
rect 10145 9205 10455 9245
rect 10495 9205 10500 9245
rect 6950 9200 10500 9205
rect 8700 8900 8750 9200
rect 6950 8895 10500 8900
rect 6950 8855 6955 8895
rect 6995 8855 7305 8895
rect 7345 8855 7655 8895
rect 7695 8855 8005 8895
rect 8045 8855 8355 8895
rect 8395 8855 8705 8895
rect 8745 8855 9055 8895
rect 9095 8855 9405 8895
rect 9445 8855 9755 8895
rect 9795 8855 10105 8895
rect 10145 8855 10455 8895
rect 10495 8855 10500 8895
rect 6950 8850 10500 8855
rect 8700 8550 8750 8850
rect 6950 8545 10500 8550
rect 6950 8505 6955 8545
rect 6995 8505 7305 8545
rect 7345 8505 7655 8545
rect 7695 8505 8005 8545
rect 8045 8505 8355 8545
rect 8395 8505 8705 8545
rect 8745 8505 9055 8545
rect 9095 8505 9405 8545
rect 9445 8505 9755 8545
rect 9795 8505 10105 8545
rect 10145 8505 10455 8545
rect 10495 8505 10500 8545
rect 6950 8500 10500 8505
rect 8700 8200 8750 8500
rect 6950 8195 10500 8200
rect 6950 8155 6955 8195
rect 6995 8155 7305 8195
rect 7345 8155 7655 8195
rect 7695 8155 8005 8195
rect 8045 8155 8355 8195
rect 8395 8155 8705 8195
rect 8745 8155 9055 8195
rect 9095 8155 9405 8195
rect 9445 8155 9755 8195
rect 9795 8155 10105 8195
rect 10145 8155 10455 8195
rect 10495 8155 10500 8195
rect 6950 8150 10500 8155
rect 8700 7850 8750 8150
rect 6950 7845 10500 7850
rect 6950 7805 6955 7845
rect 6995 7805 7305 7845
rect 7345 7805 7655 7845
rect 7695 7805 8005 7845
rect 8045 7805 8355 7845
rect 8395 7805 8705 7845
rect 8745 7805 9055 7845
rect 9095 7805 9405 7845
rect 9445 7805 9755 7845
rect 9795 7805 10105 7845
rect 10145 7805 10455 7845
rect 10495 7805 10500 7845
rect 6950 7800 10500 7805
rect 8700 7500 8750 7800
rect 6950 7495 10500 7500
rect 6950 7455 6955 7495
rect 6995 7455 7305 7495
rect 7345 7455 7655 7495
rect 7695 7455 8005 7495
rect 8045 7455 8355 7495
rect 8395 7455 8705 7495
rect 8745 7455 9055 7495
rect 9095 7455 9405 7495
rect 9445 7455 9755 7495
rect 9795 7455 10105 7495
rect 10145 7455 10455 7495
rect 10495 7455 10500 7495
rect 6950 7450 10500 7455
rect 8700 7150 8750 7450
rect 6950 7145 10500 7150
rect 6950 7105 6955 7145
rect 6995 7105 7305 7145
rect 7345 7105 7655 7145
rect 7695 7105 8005 7145
rect 8045 7105 8355 7145
rect 8395 7105 8705 7145
rect 8745 7105 9055 7145
rect 9095 7105 9405 7145
rect 9445 7105 9755 7145
rect 9795 7105 10105 7145
rect 10145 7105 10455 7145
rect 10495 7105 10500 7145
rect 6950 7100 10500 7105
rect -2440 6940 6640 6950
rect -2440 6915 2385 6940
rect -2440 6865 -2405 6915
rect -2355 6865 -2310 6915
rect -2260 6865 -2215 6915
rect -2165 6865 -2115 6915
rect -2065 6865 -2015 6915
rect -1965 6865 -1915 6915
rect -1865 6865 -1820 6915
rect -1770 6865 -1725 6915
rect -1675 6900 2385 6915
rect 2425 6900 3240 6940
rect 3280 6900 4470 6940
rect 4510 6900 6300 6940
rect 6340 6900 6590 6940
rect 6630 6900 6640 6940
rect -1675 6875 6640 6900
rect -1675 6865 2385 6875
rect -2440 6835 2385 6865
rect 2425 6835 3240 6875
rect 3280 6835 4470 6875
rect 4510 6835 6300 6875
rect 6340 6835 6590 6875
rect 6630 6835 6640 6875
rect -2440 6825 6640 6835
rect -2440 6775 -2405 6825
rect -2355 6775 -2310 6825
rect -2260 6775 -2215 6825
rect -2165 6775 -2115 6825
rect -2065 6775 -2015 6825
rect -1965 6775 -1915 6825
rect -1865 6775 -1820 6825
rect -1770 6775 -1725 6825
rect -1675 6805 6640 6825
rect -1675 6775 2385 6805
rect -2440 6765 2385 6775
rect 2425 6765 3240 6805
rect 3280 6765 4470 6805
rect 4510 6765 6300 6805
rect 6340 6765 6590 6805
rect 6630 6800 6640 6805
rect 8700 6800 8750 7100
rect 10710 6915 15040 6950
rect 10710 6865 10745 6915
rect 10795 6865 10840 6915
rect 10890 6865 10935 6915
rect 10985 6865 11035 6915
rect 11085 6865 11135 6915
rect 11185 6865 11235 6915
rect 11285 6865 11330 6915
rect 11380 6865 11425 6915
rect 11475 6865 15040 6915
rect 10710 6825 15040 6865
rect 6630 6795 10500 6800
rect 6630 6765 6955 6795
rect -2440 6755 6955 6765
rect 6995 6755 7305 6795
rect 7345 6755 7655 6795
rect 7695 6755 8005 6795
rect 8045 6755 8355 6795
rect 8395 6755 8705 6795
rect 8745 6755 9055 6795
rect 9095 6755 9405 6795
rect 9445 6755 9755 6795
rect 9795 6755 10105 6795
rect 10145 6755 10455 6795
rect 10495 6755 10500 6795
rect -2440 6750 10500 6755
rect 10710 6775 10745 6825
rect 10795 6775 10840 6825
rect 10890 6775 10935 6825
rect 10985 6775 11035 6825
rect 11085 6775 11135 6825
rect 11185 6775 11235 6825
rect 11285 6775 11330 6825
rect 11380 6775 11425 6825
rect 11475 6775 15040 6825
rect -2440 6735 6640 6750
rect -2440 6725 2385 6735
rect -2440 6675 -2405 6725
rect -2355 6675 -2310 6725
rect -2260 6675 -2215 6725
rect -2165 6675 -2115 6725
rect -2065 6675 -2015 6725
rect -1965 6675 -1915 6725
rect -1865 6675 -1820 6725
rect -1770 6675 -1725 6725
rect -1675 6695 2385 6725
rect 2425 6695 3240 6735
rect 3280 6695 4470 6735
rect 4510 6695 6300 6735
rect 6340 6695 6590 6735
rect 6630 6695 6640 6735
rect -1675 6675 6640 6695
rect -2440 6665 6640 6675
rect -2440 6635 2385 6665
rect -2440 6585 -2405 6635
rect -2355 6585 -2310 6635
rect -2260 6585 -2215 6635
rect -2165 6585 -2115 6635
rect -2065 6585 -2015 6635
rect -1965 6585 -1915 6635
rect -1865 6585 -1820 6635
rect -1770 6585 -1725 6635
rect -1675 6625 2385 6635
rect 2425 6625 3240 6665
rect 3280 6625 4470 6665
rect 4510 6625 6300 6665
rect 6340 6625 6590 6665
rect 6630 6625 6640 6665
rect -1675 6600 6640 6625
rect -1675 6585 2385 6600
rect -2440 6560 2385 6585
rect 2425 6560 3240 6600
rect 3280 6560 4470 6600
rect 4510 6560 6300 6600
rect 6340 6560 6590 6600
rect 6630 6560 6640 6600
rect -2440 6550 6640 6560
rect 10710 6725 15040 6775
rect 10710 6675 10745 6725
rect 10795 6675 10840 6725
rect 10890 6675 10935 6725
rect 10985 6675 11035 6725
rect 11085 6675 11135 6725
rect 11185 6675 11235 6725
rect 11285 6675 11330 6725
rect 11380 6675 11425 6725
rect 11475 6675 15040 6725
rect 10710 6635 15040 6675
rect 10710 6585 10745 6635
rect 10795 6585 10840 6635
rect 10890 6585 10935 6635
rect 10985 6585 11035 6635
rect 11085 6585 11135 6635
rect 11185 6585 11235 6635
rect 11285 6585 11330 6635
rect 11380 6585 11425 6635
rect 11475 6585 15040 6635
rect 10710 6550 15040 6585
rect 4460 -210 11510 -200
rect 4460 -250 4470 -210
rect 4510 -235 11510 -210
rect 4510 -250 10745 -235
rect 4460 -275 10745 -250
rect 4460 -315 4470 -275
rect 4510 -285 10745 -275
rect 10795 -285 10840 -235
rect 10890 -285 10935 -235
rect 10985 -285 11035 -235
rect 11085 -285 11135 -235
rect 11185 -285 11235 -235
rect 11285 -285 11330 -235
rect 11380 -285 11425 -235
rect 11475 -285 11510 -235
rect 4510 -315 11510 -285
rect 4460 -325 11510 -315
rect 4460 -345 10745 -325
rect 4460 -385 4470 -345
rect 4510 -375 10745 -345
rect 10795 -375 10840 -325
rect 10890 -375 10935 -325
rect 10985 -375 11035 -325
rect 11085 -375 11135 -325
rect 11185 -375 11235 -325
rect 11285 -375 11330 -325
rect 11380 -375 11425 -325
rect 11475 -375 11510 -325
rect 4510 -385 11510 -375
rect 4460 -415 11510 -385
rect 4460 -455 4470 -415
rect 4510 -425 11510 -415
rect 4510 -455 10745 -425
rect 4460 -475 10745 -455
rect 10795 -475 10840 -425
rect 10890 -475 10935 -425
rect 10985 -475 11035 -425
rect 11085 -475 11135 -425
rect 11185 -475 11235 -425
rect 11285 -475 11330 -425
rect 11380 -475 11425 -425
rect 11475 -475 11510 -425
rect 4460 -485 11510 -475
rect 4460 -525 4470 -485
rect 4510 -515 11510 -485
rect 4510 -525 10745 -515
rect 4460 -550 10745 -525
rect 4460 -590 4470 -550
rect 4510 -565 10745 -550
rect 10795 -565 10840 -515
rect 10890 -565 10935 -515
rect 10985 -565 11035 -515
rect 11085 -565 11135 -515
rect 11185 -565 11235 -515
rect 11285 -565 11330 -515
rect 11380 -565 11425 -515
rect 11475 -565 11510 -515
rect 4510 -590 11510 -565
rect 4460 -600 11510 -590
use bgr_11  bgr_11_0
timestamp 1753627268
transform -1 0 22290 0 -1 8785
box 15665 -6150 19905 1600
use two_stage_opamp_dummy_magic_23  two_stage_opamp_dummy_magic_23_0
timestamp 1753589008
transform 1 0 -52410 0 1 255
box 52410 -455 61390 6101
<< labels >>
flabel metal3 -2040 8255 -2040 8255 1 FreeSans 800 0 0 320 VDDA
port 1 n
flabel metal2 5375 2025 5375 2025 3 FreeSans 400 0 160 0 VIN-
port 6 e
flabel metal2 3605 2025 3605 2025 7 FreeSans 400 0 -160 0 VIN+
port 5 w
flabel metal2 2060 1485 2060 1485 5 FreeSans 400 0 0 -160 VOUT+
port 3 s
flabel metal2 6875 1485 6875 1485 5 FreeSans 400 0 0 -160 VOUT-
port 4 s
flabel metal4 15040 6750 15040 6750 3 FreeSans 800 0 320 0 GNDA
port 2 e
<< end >>
