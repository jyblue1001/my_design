magic
tech sky130A
timestamp 1739811012
<< nwell >>
rect 3005 1875 4725 2070
rect 3005 900 4645 1875
rect 2340 610 3055 900
rect 3265 640 3325 655
<< poly >>
rect 2645 2790 3005 2800
rect 2645 2770 2655 2790
rect 2675 2785 3005 2790
rect 2675 2770 2685 2785
rect 2645 2760 2685 2770
rect -130 960 -90 975
rect 2180 945 2220 955
rect 2180 930 2190 945
rect 2090 925 2190 930
rect 2210 925 2220 945
rect 2090 915 2220 925
rect 3030 650 3070 660
rect 3030 630 3040 650
rect 3060 640 3070 650
rect 3265 640 3325 655
rect 3060 630 3325 640
rect 3030 620 3325 630
rect 4025 640 4065 650
rect 4025 620 4035 640
rect 4055 620 4065 640
rect 4025 610 4065 620
rect 4245 455 4285 465
rect 4245 435 4255 455
rect 4275 435 4285 455
rect 4245 425 4285 435
rect -130 245 -90 260
rect 2075 85 2115 95
rect 2075 65 2085 85
rect 2105 65 2115 85
rect 2075 55 2115 65
<< polycont >>
rect 2655 2770 2675 2790
rect 2190 925 2210 945
rect 3040 630 3060 650
rect 4035 620 4055 640
rect 4255 435 4275 455
rect 2085 65 2105 85
<< locali >>
rect 2865 3045 2915 3060
rect 2865 3025 2880 3045
rect 2900 3025 2915 3045
rect 2865 3010 2915 3025
rect 2705 2810 2745 2820
rect 2645 2790 2685 2800
rect 2645 2770 2655 2790
rect 2675 2770 2685 2790
rect 2645 1575 2685 2770
rect 2645 1555 2655 1575
rect 2675 1555 2685 1575
rect 2645 1545 2685 1555
rect 2705 2790 2715 2810
rect 2735 2790 2745 2810
rect 2380 1210 2430 1220
rect 2355 1190 2390 1210
rect 2380 1180 2390 1190
rect 2420 1180 2430 1210
rect 2380 1170 2430 1180
rect 2040 1130 2680 1150
rect 2040 1105 2060 1130
rect 2180 945 2220 955
rect 2180 925 2190 945
rect 2210 925 2220 945
rect 2180 915 2220 925
rect 2300 945 2340 955
rect 2300 925 2310 945
rect 2330 925 2340 945
rect 2300 915 2340 925
rect 2660 660 2680 1130
rect 2640 650 2680 660
rect 2500 625 2550 640
rect 2500 620 2515 625
rect 2355 600 2385 620
rect 2405 600 2440 620
rect 2460 605 2515 620
rect 2535 605 2550 625
rect 2640 630 2650 650
rect 2670 630 2680 650
rect 2640 620 2680 630
rect 2460 600 2550 605
rect 2500 590 2550 600
rect 2705 585 2745 2790
rect 4910 2755 5950 2775
rect 2865 2450 2915 2465
rect 2865 2430 2880 2450
rect 2900 2430 2915 2450
rect 2865 2415 2915 2430
rect 5930 1625 5950 2755
rect 2785 1605 5950 1625
rect 2785 660 2805 1605
rect 2910 975 2960 990
rect 2910 955 2925 975
rect 2945 955 2960 975
rect 2910 940 2960 955
rect 2765 650 2805 660
rect 2765 630 2775 650
rect 2795 640 2805 650
rect 3030 650 3070 660
rect 3030 640 3040 650
rect 2795 630 3040 640
rect 3060 630 3070 650
rect 2765 620 3070 630
rect 4025 640 4065 650
rect 3330 585 3370 625
rect 4025 620 4035 640
rect 4055 620 4065 640
rect 4025 610 4065 620
rect 2040 540 2200 560
rect 2705 545 3370 585
rect 4625 555 4665 565
rect 2040 505 2060 540
rect 2180 520 2200 540
rect 4625 535 4635 555
rect 4655 535 4665 555
rect 4625 525 4665 535
rect 2180 500 2900 520
rect 2650 455 2690 465
rect 2650 435 2660 455
rect 2680 435 2690 455
rect 2650 425 2690 435
rect 4245 455 4285 465
rect 4245 435 4255 455
rect 4275 435 4285 455
rect 4245 425 4285 435
rect 2650 265 2670 425
rect 2320 245 2670 265
rect 2910 135 2960 150
rect 2910 115 2925 135
rect 2945 115 2960 135
rect 2910 100 2960 115
rect 2075 85 2115 95
rect 2075 65 2085 85
rect 2105 65 2115 85
rect 2075 55 2115 65
rect 2380 40 2430 50
rect 2380 30 2390 40
rect 2355 10 2390 30
rect 2420 10 2430 40
rect 2380 0 2430 10
<< viali >>
rect 2880 3025 2900 3045
rect 2655 1555 2675 1575
rect 2715 2790 2735 2810
rect 2390 1180 2420 1210
rect 2190 925 2210 945
rect 2310 925 2330 945
rect 2385 600 2405 620
rect 2440 600 2460 620
rect 2515 605 2535 625
rect 2650 630 2670 650
rect 2880 2430 2900 2450
rect 2925 955 2945 975
rect 2775 630 2795 650
rect 4035 620 4055 640
rect 4635 535 4655 555
rect 2660 435 2680 455
rect 4255 435 4275 455
rect 2925 115 2945 135
rect 2085 65 2105 85
rect 2390 10 2420 40
<< metal1 >>
rect 2865 3050 2915 3060
rect 2865 3020 2875 3050
rect 2905 3020 2915 3050
rect 2865 3010 2915 3020
rect 2705 2810 3005 2820
rect 2705 2790 2715 2810
rect 2735 2805 3005 2810
rect 2735 2790 2745 2805
rect 2705 2780 2745 2790
rect 2865 2455 2915 2465
rect 2865 2425 2875 2455
rect 2905 2425 2915 2455
rect 2865 2415 2915 2425
rect 2645 1575 5650 1585
rect 2645 1555 2655 1575
rect 2675 1555 5650 1575
rect 2645 1545 5650 1555
rect 2520 1445 2910 1500
rect 2355 1210 2430 1220
rect 2355 1180 2390 1210
rect 2420 1180 2430 1210
rect 2380 1170 2430 1180
rect 2520 1020 2565 1445
rect 2180 980 2565 1020
rect 2910 980 2960 990
rect 2180 945 2220 980
rect 2180 925 2190 945
rect 2210 925 2220 945
rect 2180 915 2220 925
rect 2300 945 2340 955
rect 2300 925 2310 945
rect 2330 935 2340 945
rect 2910 950 2920 980
rect 2950 950 2960 980
rect 2910 940 2960 950
rect 2330 925 2595 935
rect 2300 915 2595 925
rect 2500 630 2550 640
rect -140 590 -115 630
rect 2355 620 2510 630
rect 2355 600 2385 620
rect 2405 600 2440 620
rect 2460 600 2510 620
rect 2540 600 2550 630
rect 2355 590 2550 600
rect 2575 605 2595 915
rect 2640 650 2680 660
rect 2640 630 2650 650
rect 2670 640 2680 650
rect 2765 650 2805 660
rect 2765 640 2775 650
rect 2670 630 2775 640
rect 2795 630 2805 650
rect 2640 620 2805 630
rect 4025 640 4065 650
rect 4025 620 4035 640
rect 4055 620 4065 640
rect 4025 605 4065 620
rect 2575 585 4065 605
rect 5610 565 5650 1545
rect 4625 555 5650 565
rect 4625 535 4635 555
rect 4655 535 5650 555
rect 4625 525 5650 535
rect 2650 455 4285 465
rect 2650 435 2660 455
rect 2680 445 4255 455
rect 2680 435 2690 445
rect 2650 425 2690 435
rect 4245 435 4255 445
rect 4275 435 4285 455
rect 4245 425 4285 435
rect 2910 140 2960 150
rect 2910 110 2920 140
rect 2950 110 2960 140
rect 2910 100 2960 110
rect 2075 85 2775 95
rect 2075 65 2085 85
rect 2105 75 2775 85
rect 2105 65 2115 75
rect 2075 55 2115 65
rect 2380 40 2430 50
rect 2355 10 2390 40
rect 2420 10 2430 40
rect 2355 0 2430 10
rect 2735 5 2775 75
rect 2735 -50 2910 5
<< via1 >>
rect 2875 3045 2905 3050
rect 2875 3025 2880 3045
rect 2880 3025 2900 3045
rect 2900 3025 2905 3045
rect 2875 3020 2905 3025
rect 2875 2450 2905 2455
rect 2875 2430 2880 2450
rect 2880 2430 2900 2450
rect 2900 2430 2905 2450
rect 2875 2425 2905 2430
rect 2390 1180 2420 1210
rect 2920 975 2950 980
rect 2920 955 2925 975
rect 2925 955 2945 975
rect 2945 955 2950 975
rect 2920 950 2950 955
rect 2510 625 2540 630
rect 2510 605 2515 625
rect 2515 605 2535 625
rect 2535 605 2540 625
rect 2510 600 2540 605
rect 2920 135 2950 140
rect 2920 115 2925 135
rect 2925 115 2945 135
rect 2945 115 2950 135
rect 2920 110 2950 115
rect 2390 10 2420 40
<< metal2 >>
rect 2865 3050 2915 3060
rect 2865 3020 2875 3050
rect 2905 3020 2915 3050
rect 2865 3010 2915 3020
rect 2865 2455 2915 2465
rect 2865 2425 2875 2455
rect 2905 2425 2915 2455
rect 2865 2415 2915 2425
rect 2380 1210 2430 1220
rect 2380 1180 2390 1210
rect 2420 1180 2430 1210
rect 2380 1170 2430 1180
rect 2910 980 2960 990
rect 2910 950 2920 980
rect 2950 950 2960 980
rect 2910 940 2960 950
rect 2500 630 2550 640
rect 2500 600 2510 630
rect 2540 600 2550 630
rect 2500 590 2550 600
rect 2910 140 2960 150
rect 2910 110 2920 140
rect 2950 110 2960 140
rect 2910 100 2960 110
rect 2380 40 2430 50
rect 2380 10 2390 40
rect 2420 10 2430 40
rect 2380 0 2430 10
<< via2 >>
rect 2875 3020 2905 3050
rect 2875 2425 2905 2455
rect 2390 1180 2420 1210
rect 2920 950 2950 980
rect 2510 600 2540 630
rect 2920 110 2950 140
rect 2390 10 2420 40
<< metal3 >>
rect 2380 3055 2915 3060
rect 2380 3015 2385 3055
rect 2425 3050 2915 3055
rect 2425 3020 2875 3050
rect 2905 3020 2915 3050
rect 2425 3015 2915 3020
rect 2380 3010 2915 3015
rect 2500 2460 2915 2465
rect 2500 2420 2505 2460
rect 2545 2455 2915 2460
rect 2545 2425 2875 2455
rect 2905 2425 2915 2455
rect 2545 2420 2915 2425
rect 2500 2415 2915 2420
rect 2380 1215 2430 1220
rect 2380 1175 2385 1215
rect 2425 1175 2430 1215
rect 2380 1170 2430 1175
rect 2500 985 2960 990
rect 2500 945 2505 985
rect 2545 980 2960 985
rect 2545 950 2920 980
rect 2950 950 2960 980
rect 2545 945 2960 950
rect 2500 940 2960 945
rect 2500 635 2550 640
rect 2500 595 2505 635
rect 2545 595 2550 635
rect 2500 590 2550 595
rect 2380 145 2960 150
rect 2380 105 2385 145
rect 2425 140 2960 145
rect 2425 110 2920 140
rect 2950 110 2960 140
rect 2425 105 2960 110
rect 2380 100 2960 105
rect 2380 45 2430 50
rect 2380 5 2385 45
rect 2425 5 2430 45
rect 2380 0 2430 5
<< via3 >>
rect 2385 3015 2425 3055
rect 2505 2420 2545 2460
rect 2385 1210 2425 1215
rect 2385 1180 2390 1210
rect 2390 1180 2420 1210
rect 2420 1180 2425 1210
rect 2385 1175 2425 1180
rect 2505 945 2545 985
rect 2505 630 2545 635
rect 2505 600 2510 630
rect 2510 600 2540 630
rect 2540 600 2545 630
rect 2505 595 2545 600
rect 2385 105 2425 145
rect 2385 40 2425 45
rect 2385 10 2390 40
rect 2390 10 2420 40
rect 2420 10 2425 40
rect 2385 5 2425 10
<< metal4 >>
rect 2380 3055 2430 3060
rect 2380 3015 2385 3055
rect 2425 3015 2430 3055
rect 2380 1215 2430 3015
rect 2380 1175 2385 1215
rect 2425 1175 2430 1215
rect -280 105 -230 155
rect 2380 145 2430 1175
rect 2500 2460 2550 2465
rect 2500 2420 2505 2460
rect 2545 2420 2550 2460
rect 2500 985 2550 2420
rect 2500 945 2505 985
rect 2545 945 2550 985
rect 2500 635 2550 945
rect 2500 595 2505 635
rect 2545 595 2550 635
rect 2500 590 2550 595
rect 2380 105 2385 145
rect 2425 105 2430 145
rect 2380 45 2430 105
rect 2380 5 2385 45
rect 2425 5 2430 45
rect 2380 0 2430 5
use charge_pump_cell_6  charge_pump_cell_6_0
timestamp 1739810861
transform 1 0 -6195 0 1 -1605
box 9095 1555 11740 3105
use opamp_cell_4  opamp_cell_4_0
timestamp 1739772381
transform 1 0 -335 0 -1 4855
box 3110 897 6365 3205
use pfd_8  pfd_8_0
timestamp 1739770731
transform 1 0 -930 0 1 4655
box 650 -4655 3290 -3435
<< labels >>
flabel locali 2880 510 2880 510 5 FreeSans 400 0 0 -200 I_IN
port 6 s
flabel metal1 -140 610 -140 610 7 FreeSans 400 0 -200 0 VDDA
port 2 w
flabel metal4 -280 130 -280 130 7 FreeSans 400 0 -200 0 GNDA
port 3 w
flabel poly -130 250 -130 250 7 FreeSans 400 0 -200 0 F_VCO
port 5 w
flabel poly -130 965 -130 965 7 FreeSans 400 0 -200 0 F_REF
port 4 w
flabel metal1 5650 545 5650 545 3 FreeSans 400 0 200 0 V_OUT
port 1 e
<< end >>
