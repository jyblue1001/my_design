* NGSPICE file created from passgate_4.ext - technology: sky130A

.subckt passgate_4
X0 B GNDA A VDDA sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X1 B VDDA A GNDA sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
.ends

