magic
tech sky130A
magscale 1 2
timestamp 1746510996
<< nwell >>
rect 4300 3700 9310 5500
<< pwell >>
rect 5620 3120 7300 3320
rect 1500 1320 2550 1340
rect 2630 1320 2670 1340
rect 1370 1187 2670 1320
rect 1370 153 1503 1187
rect 2537 153 2670 1187
rect 40 50 80 90
rect 1370 20 2670 153
rect 2710 1320 2770 1340
rect 2850 1320 4050 1340
rect 2710 1187 4050 1320
rect 2710 153 2863 1187
rect 3897 153 4050 1187
rect 2710 20 4050 153
rect 4070 1187 5390 1340
rect 4070 153 4223 1187
rect 5257 153 5390 1187
rect 4070 20 5390 153
rect 5430 1187 6750 1340
rect 5430 153 5583 1187
rect 6617 153 6750 1187
rect 5430 20 6750 153
rect 6790 1187 8110 1340
rect 6790 153 6943 1187
rect 7977 153 8110 1187
rect 6790 20 8110 153
rect 8150 1187 9470 1340
rect 8150 153 8303 1187
rect 9337 153 9470 1187
rect 8150 20 9470 153
<< nbase >>
rect 1503 153 2537 1187
rect 2863 153 3897 1187
rect 4223 153 5257 1187
rect 5583 153 6617 1187
rect 6943 153 7977 1187
rect 8303 153 9337 1187
<< nmos >>
rect 5700 3120 5820 3320
rect 5900 3120 6020 3320
rect 6100 3120 6220 3320
rect 6300 3120 6420 3320
rect 6500 3120 6620 3320
rect 6700 3120 6820 3320
rect 6900 3120 7020 3320
rect 7100 3120 7220 3320
rect 5540 1970 6340 2770
rect 6580 1970 7380 2770
rect 5440 1510 7440 1710
<< pmos >>
rect 4700 4660 4820 5460
rect 4900 4660 5020 5460
rect 5100 4660 5220 5460
rect 5300 4660 5420 5460
rect 5500 4660 5620 5460
rect 5700 4660 5820 5460
rect 5900 4660 6020 5460
rect 6100 4660 6220 5460
rect 6300 4660 6420 5460
rect 6500 4660 6620 5460
rect 6700 4660 6820 5460
rect 6900 4660 7020 5460
rect 7100 4660 7220 5460
rect 7300 4660 7420 5460
rect 7500 4660 7620 5460
rect 7700 4660 7820 5460
rect 7900 4660 8020 5460
rect 8100 4660 8220 5460
rect 5300 3820 5420 4220
rect 5500 3820 5620 4220
rect 5700 3820 5820 4220
rect 5900 3820 6020 4220
rect 6100 3820 6220 4220
rect 6300 3820 6420 4220
rect 6500 3820 6620 4220
rect 6700 3820 6820 4220
rect 6900 3820 7020 4220
rect 7100 3820 7220 4220
rect 7300 3820 7420 4220
rect 7500 3820 7620 4220
rect 8830 3820 8860 4220
rect 9080 3820 9110 4220
<< ndiff >>
rect 5620 3290 5700 3320
rect 5620 3250 5640 3290
rect 5680 3250 5700 3290
rect 5620 3190 5700 3250
rect 5620 3150 5640 3190
rect 5680 3150 5700 3190
rect 5620 3120 5700 3150
rect 5820 3290 5900 3320
rect 5820 3250 5840 3290
rect 5880 3250 5900 3290
rect 5820 3190 5900 3250
rect 5820 3150 5840 3190
rect 5880 3150 5900 3190
rect 5820 3120 5900 3150
rect 6020 3290 6100 3320
rect 6020 3250 6040 3290
rect 6080 3250 6100 3290
rect 6020 3190 6100 3250
rect 6020 3150 6040 3190
rect 6080 3150 6100 3190
rect 6020 3120 6100 3150
rect 6220 3290 6300 3320
rect 6220 3250 6240 3290
rect 6280 3250 6300 3290
rect 6220 3190 6300 3250
rect 6220 3150 6240 3190
rect 6280 3150 6300 3190
rect 6220 3120 6300 3150
rect 6420 3290 6500 3320
rect 6420 3250 6440 3290
rect 6480 3250 6500 3290
rect 6420 3190 6500 3250
rect 6420 3150 6440 3190
rect 6480 3150 6500 3190
rect 6420 3120 6500 3150
rect 6620 3290 6700 3320
rect 6620 3250 6640 3290
rect 6680 3250 6700 3290
rect 6620 3190 6700 3250
rect 6620 3150 6640 3190
rect 6680 3150 6700 3190
rect 6620 3120 6700 3150
rect 6820 3290 6900 3320
rect 6820 3250 6840 3290
rect 6880 3250 6900 3290
rect 6820 3190 6900 3250
rect 6820 3150 6840 3190
rect 6880 3150 6900 3190
rect 6820 3120 6900 3150
rect 7020 3290 7100 3320
rect 7020 3250 7040 3290
rect 7080 3250 7100 3290
rect 7020 3190 7100 3250
rect 7020 3150 7040 3190
rect 7080 3150 7100 3190
rect 7020 3120 7100 3150
rect 7220 3290 7300 3320
rect 7220 3250 7240 3290
rect 7280 3250 7300 3290
rect 7220 3190 7300 3250
rect 7220 3150 7240 3190
rect 7280 3150 7300 3190
rect 7220 3120 7300 3150
rect 5460 2740 5540 2770
rect 5460 2700 5480 2740
rect 5520 2700 5540 2740
rect 5460 2640 5540 2700
rect 5460 2600 5480 2640
rect 5520 2600 5540 2640
rect 5460 2540 5540 2600
rect 5460 2500 5480 2540
rect 5520 2500 5540 2540
rect 5460 2440 5540 2500
rect 5460 2400 5480 2440
rect 5520 2400 5540 2440
rect 5460 2340 5540 2400
rect 5460 2300 5480 2340
rect 5520 2300 5540 2340
rect 5460 2240 5540 2300
rect 5460 2200 5480 2240
rect 5520 2200 5540 2240
rect 5460 2140 5540 2200
rect 5460 2100 5480 2140
rect 5520 2100 5540 2140
rect 5460 2040 5540 2100
rect 5460 2000 5480 2040
rect 5520 2000 5540 2040
rect 5460 1970 5540 2000
rect 6340 2740 6420 2770
rect 6500 2740 6580 2770
rect 6340 2700 6360 2740
rect 6400 2700 6420 2740
rect 6500 2700 6520 2740
rect 6560 2700 6580 2740
rect 6340 2640 6420 2700
rect 6500 2640 6580 2700
rect 6340 2600 6360 2640
rect 6400 2600 6420 2640
rect 6500 2600 6520 2640
rect 6560 2600 6580 2640
rect 6340 2540 6420 2600
rect 6500 2540 6580 2600
rect 6340 2500 6360 2540
rect 6400 2500 6420 2540
rect 6500 2500 6520 2540
rect 6560 2500 6580 2540
rect 6340 2440 6420 2500
rect 6500 2440 6580 2500
rect 6340 2400 6360 2440
rect 6400 2400 6420 2440
rect 6500 2400 6520 2440
rect 6560 2400 6580 2440
rect 6340 2340 6420 2400
rect 6500 2340 6580 2400
rect 6340 2300 6360 2340
rect 6400 2300 6420 2340
rect 6500 2300 6520 2340
rect 6560 2300 6580 2340
rect 6340 2240 6420 2300
rect 6500 2240 6580 2300
rect 6340 2200 6360 2240
rect 6400 2200 6420 2240
rect 6500 2200 6520 2240
rect 6560 2200 6580 2240
rect 6340 2140 6420 2200
rect 6500 2140 6580 2200
rect 6340 2100 6360 2140
rect 6400 2100 6420 2140
rect 6500 2100 6520 2140
rect 6560 2100 6580 2140
rect 6340 2040 6420 2100
rect 6500 2040 6580 2100
rect 6340 2000 6360 2040
rect 6400 2000 6420 2040
rect 6500 2000 6520 2040
rect 6560 2000 6580 2040
rect 6340 1970 6420 2000
rect 6500 1970 6580 2000
rect 7380 2740 7460 2770
rect 7380 2700 7400 2740
rect 7440 2700 7460 2740
rect 7380 2640 7460 2700
rect 7380 2600 7400 2640
rect 7440 2600 7460 2640
rect 7380 2540 7460 2600
rect 7380 2500 7400 2540
rect 7440 2500 7460 2540
rect 7380 2440 7460 2500
rect 7380 2400 7400 2440
rect 7440 2400 7460 2440
rect 7380 2340 7460 2400
rect 7380 2300 7400 2340
rect 7440 2300 7460 2340
rect 7380 2240 7460 2300
rect 7380 2200 7400 2240
rect 7440 2200 7460 2240
rect 7380 2140 7460 2200
rect 7380 2100 7400 2140
rect 7440 2100 7460 2140
rect 7380 2040 7460 2100
rect 7380 2000 7400 2040
rect 7440 2000 7460 2040
rect 7380 1970 7460 2000
rect 5360 1680 5440 1710
rect 5360 1640 5380 1680
rect 5420 1640 5440 1680
rect 5360 1580 5440 1640
rect 5360 1540 5380 1580
rect 5420 1540 5440 1580
rect 5360 1510 5440 1540
rect 7440 1680 7520 1710
rect 7440 1640 7460 1680
rect 7500 1640 7520 1680
rect 7440 1580 7520 1640
rect 7440 1540 7460 1580
rect 7500 1540 7520 1580
rect 7440 1510 7520 1540
<< pdiff >>
rect 4620 5430 4700 5460
rect 4620 5390 4640 5430
rect 4680 5390 4700 5430
rect 4620 5330 4700 5390
rect 4620 5290 4640 5330
rect 4680 5290 4700 5330
rect 4620 5230 4700 5290
rect 4620 5190 4640 5230
rect 4680 5190 4700 5230
rect 4620 5130 4700 5190
rect 4620 5090 4640 5130
rect 4680 5090 4700 5130
rect 4620 5030 4700 5090
rect 4620 4990 4640 5030
rect 4680 4990 4700 5030
rect 4620 4930 4700 4990
rect 4620 4890 4640 4930
rect 4680 4890 4700 4930
rect 4620 4830 4700 4890
rect 4620 4790 4640 4830
rect 4680 4790 4700 4830
rect 4620 4730 4700 4790
rect 4620 4690 4640 4730
rect 4680 4690 4700 4730
rect 4620 4660 4700 4690
rect 4820 5430 4900 5460
rect 4820 5390 4840 5430
rect 4880 5390 4900 5430
rect 4820 5330 4900 5390
rect 4820 5290 4840 5330
rect 4880 5290 4900 5330
rect 4820 5230 4900 5290
rect 4820 5190 4840 5230
rect 4880 5190 4900 5230
rect 4820 5130 4900 5190
rect 4820 5090 4840 5130
rect 4880 5090 4900 5130
rect 4820 5030 4900 5090
rect 4820 4990 4840 5030
rect 4880 4990 4900 5030
rect 4820 4930 4900 4990
rect 4820 4890 4840 4930
rect 4880 4890 4900 4930
rect 4820 4830 4900 4890
rect 4820 4790 4840 4830
rect 4880 4790 4900 4830
rect 4820 4730 4900 4790
rect 4820 4690 4840 4730
rect 4880 4690 4900 4730
rect 4820 4660 4900 4690
rect 5020 5430 5100 5460
rect 5020 5390 5040 5430
rect 5080 5390 5100 5430
rect 5020 5330 5100 5390
rect 5020 5290 5040 5330
rect 5080 5290 5100 5330
rect 5020 5230 5100 5290
rect 5020 5190 5040 5230
rect 5080 5190 5100 5230
rect 5020 5130 5100 5190
rect 5020 5090 5040 5130
rect 5080 5090 5100 5130
rect 5020 5030 5100 5090
rect 5020 4990 5040 5030
rect 5080 4990 5100 5030
rect 5020 4930 5100 4990
rect 5020 4890 5040 4930
rect 5080 4890 5100 4930
rect 5020 4830 5100 4890
rect 5020 4790 5040 4830
rect 5080 4790 5100 4830
rect 5020 4730 5100 4790
rect 5020 4690 5040 4730
rect 5080 4690 5100 4730
rect 5020 4660 5100 4690
rect 5220 5430 5300 5460
rect 5220 5390 5240 5430
rect 5280 5390 5300 5430
rect 5220 5330 5300 5390
rect 5220 5290 5240 5330
rect 5280 5290 5300 5330
rect 5220 5230 5300 5290
rect 5220 5190 5240 5230
rect 5280 5190 5300 5230
rect 5220 5130 5300 5190
rect 5220 5090 5240 5130
rect 5280 5090 5300 5130
rect 5220 5030 5300 5090
rect 5220 4990 5240 5030
rect 5280 4990 5300 5030
rect 5220 4930 5300 4990
rect 5220 4890 5240 4930
rect 5280 4890 5300 4930
rect 5220 4830 5300 4890
rect 5220 4790 5240 4830
rect 5280 4790 5300 4830
rect 5220 4730 5300 4790
rect 5220 4690 5240 4730
rect 5280 4690 5300 4730
rect 5220 4660 5300 4690
rect 5420 5430 5500 5460
rect 5420 5390 5440 5430
rect 5480 5390 5500 5430
rect 5420 5330 5500 5390
rect 5420 5290 5440 5330
rect 5480 5290 5500 5330
rect 5420 5230 5500 5290
rect 5420 5190 5440 5230
rect 5480 5190 5500 5230
rect 5420 5130 5500 5190
rect 5420 5090 5440 5130
rect 5480 5090 5500 5130
rect 5420 5030 5500 5090
rect 5420 4990 5440 5030
rect 5480 4990 5500 5030
rect 5420 4930 5500 4990
rect 5420 4890 5440 4930
rect 5480 4890 5500 4930
rect 5420 4830 5500 4890
rect 5420 4790 5440 4830
rect 5480 4790 5500 4830
rect 5420 4730 5500 4790
rect 5420 4690 5440 4730
rect 5480 4690 5500 4730
rect 5420 4660 5500 4690
rect 5620 5430 5700 5460
rect 5620 5390 5640 5430
rect 5680 5390 5700 5430
rect 5620 5330 5700 5390
rect 5620 5290 5640 5330
rect 5680 5290 5700 5330
rect 5620 5230 5700 5290
rect 5620 5190 5640 5230
rect 5680 5190 5700 5230
rect 5620 5130 5700 5190
rect 5620 5090 5640 5130
rect 5680 5090 5700 5130
rect 5620 5030 5700 5090
rect 5620 4990 5640 5030
rect 5680 4990 5700 5030
rect 5620 4930 5700 4990
rect 5620 4890 5640 4930
rect 5680 4890 5700 4930
rect 5620 4830 5700 4890
rect 5620 4790 5640 4830
rect 5680 4790 5700 4830
rect 5620 4730 5700 4790
rect 5620 4690 5640 4730
rect 5680 4690 5700 4730
rect 5620 4660 5700 4690
rect 5820 5430 5900 5460
rect 5820 5390 5840 5430
rect 5880 5390 5900 5430
rect 5820 5330 5900 5390
rect 5820 5290 5840 5330
rect 5880 5290 5900 5330
rect 5820 5230 5900 5290
rect 5820 5190 5840 5230
rect 5880 5190 5900 5230
rect 5820 5130 5900 5190
rect 5820 5090 5840 5130
rect 5880 5090 5900 5130
rect 5820 5030 5900 5090
rect 5820 4990 5840 5030
rect 5880 4990 5900 5030
rect 5820 4930 5900 4990
rect 5820 4890 5840 4930
rect 5880 4890 5900 4930
rect 5820 4830 5900 4890
rect 5820 4790 5840 4830
rect 5880 4790 5900 4830
rect 5820 4730 5900 4790
rect 5820 4690 5840 4730
rect 5880 4690 5900 4730
rect 5820 4660 5900 4690
rect 6020 5430 6100 5460
rect 6020 5390 6040 5430
rect 6080 5390 6100 5430
rect 6020 5330 6100 5390
rect 6020 5290 6040 5330
rect 6080 5290 6100 5330
rect 6020 5230 6100 5290
rect 6020 5190 6040 5230
rect 6080 5190 6100 5230
rect 6020 5130 6100 5190
rect 6020 5090 6040 5130
rect 6080 5090 6100 5130
rect 6020 5030 6100 5090
rect 6020 4990 6040 5030
rect 6080 4990 6100 5030
rect 6020 4930 6100 4990
rect 6020 4890 6040 4930
rect 6080 4890 6100 4930
rect 6020 4830 6100 4890
rect 6020 4790 6040 4830
rect 6080 4790 6100 4830
rect 6020 4730 6100 4790
rect 6020 4690 6040 4730
rect 6080 4690 6100 4730
rect 6020 4660 6100 4690
rect 6220 5430 6300 5460
rect 6220 5390 6240 5430
rect 6280 5390 6300 5430
rect 6220 5330 6300 5390
rect 6220 5290 6240 5330
rect 6280 5290 6300 5330
rect 6220 5230 6300 5290
rect 6220 5190 6240 5230
rect 6280 5190 6300 5230
rect 6220 5130 6300 5190
rect 6220 5090 6240 5130
rect 6280 5090 6300 5130
rect 6220 5030 6300 5090
rect 6220 4990 6240 5030
rect 6280 4990 6300 5030
rect 6220 4930 6300 4990
rect 6220 4890 6240 4930
rect 6280 4890 6300 4930
rect 6220 4830 6300 4890
rect 6220 4790 6240 4830
rect 6280 4790 6300 4830
rect 6220 4730 6300 4790
rect 6220 4690 6240 4730
rect 6280 4690 6300 4730
rect 6220 4660 6300 4690
rect 6420 5430 6500 5460
rect 6420 5390 6440 5430
rect 6480 5390 6500 5430
rect 6420 5330 6500 5390
rect 6420 5290 6440 5330
rect 6480 5290 6500 5330
rect 6420 5230 6500 5290
rect 6420 5190 6440 5230
rect 6480 5190 6500 5230
rect 6420 5130 6500 5190
rect 6420 5090 6440 5130
rect 6480 5090 6500 5130
rect 6420 5030 6500 5090
rect 6420 4990 6440 5030
rect 6480 4990 6500 5030
rect 6420 4930 6500 4990
rect 6420 4890 6440 4930
rect 6480 4890 6500 4930
rect 6420 4830 6500 4890
rect 6420 4790 6440 4830
rect 6480 4790 6500 4830
rect 6420 4730 6500 4790
rect 6420 4690 6440 4730
rect 6480 4690 6500 4730
rect 6420 4660 6500 4690
rect 6620 5430 6700 5460
rect 6620 5390 6640 5430
rect 6680 5390 6700 5430
rect 6620 5330 6700 5390
rect 6620 5290 6640 5330
rect 6680 5290 6700 5330
rect 6620 5230 6700 5290
rect 6620 5190 6640 5230
rect 6680 5190 6700 5230
rect 6620 5130 6700 5190
rect 6620 5090 6640 5130
rect 6680 5090 6700 5130
rect 6620 5030 6700 5090
rect 6620 4990 6640 5030
rect 6680 4990 6700 5030
rect 6620 4930 6700 4990
rect 6620 4890 6640 4930
rect 6680 4890 6700 4930
rect 6620 4830 6700 4890
rect 6620 4790 6640 4830
rect 6680 4790 6700 4830
rect 6620 4730 6700 4790
rect 6620 4690 6640 4730
rect 6680 4690 6700 4730
rect 6620 4660 6700 4690
rect 6820 5430 6900 5460
rect 6820 5390 6840 5430
rect 6880 5390 6900 5430
rect 6820 5330 6900 5390
rect 6820 5290 6840 5330
rect 6880 5290 6900 5330
rect 6820 5230 6900 5290
rect 6820 5190 6840 5230
rect 6880 5190 6900 5230
rect 6820 5130 6900 5190
rect 6820 5090 6840 5130
rect 6880 5090 6900 5130
rect 6820 5030 6900 5090
rect 6820 4990 6840 5030
rect 6880 4990 6900 5030
rect 6820 4930 6900 4990
rect 6820 4890 6840 4930
rect 6880 4890 6900 4930
rect 6820 4830 6900 4890
rect 6820 4790 6840 4830
rect 6880 4790 6900 4830
rect 6820 4730 6900 4790
rect 6820 4690 6840 4730
rect 6880 4690 6900 4730
rect 6820 4660 6900 4690
rect 7020 5430 7100 5460
rect 7020 5390 7040 5430
rect 7080 5390 7100 5430
rect 7020 5330 7100 5390
rect 7020 5290 7040 5330
rect 7080 5290 7100 5330
rect 7020 5230 7100 5290
rect 7020 5190 7040 5230
rect 7080 5190 7100 5230
rect 7020 5130 7100 5190
rect 7020 5090 7040 5130
rect 7080 5090 7100 5130
rect 7020 5030 7100 5090
rect 7020 4990 7040 5030
rect 7080 4990 7100 5030
rect 7020 4930 7100 4990
rect 7020 4890 7040 4930
rect 7080 4890 7100 4930
rect 7020 4830 7100 4890
rect 7020 4790 7040 4830
rect 7080 4790 7100 4830
rect 7020 4730 7100 4790
rect 7020 4690 7040 4730
rect 7080 4690 7100 4730
rect 7020 4660 7100 4690
rect 7220 5430 7300 5460
rect 7220 5390 7240 5430
rect 7280 5390 7300 5430
rect 7220 5330 7300 5390
rect 7220 5290 7240 5330
rect 7280 5290 7300 5330
rect 7220 5230 7300 5290
rect 7220 5190 7240 5230
rect 7280 5190 7300 5230
rect 7220 5130 7300 5190
rect 7220 5090 7240 5130
rect 7280 5090 7300 5130
rect 7220 5030 7300 5090
rect 7220 4990 7240 5030
rect 7280 4990 7300 5030
rect 7220 4930 7300 4990
rect 7220 4890 7240 4930
rect 7280 4890 7300 4930
rect 7220 4830 7300 4890
rect 7220 4790 7240 4830
rect 7280 4790 7300 4830
rect 7220 4730 7300 4790
rect 7220 4690 7240 4730
rect 7280 4690 7300 4730
rect 7220 4660 7300 4690
rect 7420 5430 7500 5460
rect 7420 5390 7440 5430
rect 7480 5390 7500 5430
rect 7420 5330 7500 5390
rect 7420 5290 7440 5330
rect 7480 5290 7500 5330
rect 7420 5230 7500 5290
rect 7420 5190 7440 5230
rect 7480 5190 7500 5230
rect 7420 5130 7500 5190
rect 7420 5090 7440 5130
rect 7480 5090 7500 5130
rect 7420 5030 7500 5090
rect 7420 4990 7440 5030
rect 7480 4990 7500 5030
rect 7420 4930 7500 4990
rect 7420 4890 7440 4930
rect 7480 4890 7500 4930
rect 7420 4830 7500 4890
rect 7420 4790 7440 4830
rect 7480 4790 7500 4830
rect 7420 4730 7500 4790
rect 7420 4690 7440 4730
rect 7480 4690 7500 4730
rect 7420 4660 7500 4690
rect 7620 5430 7700 5460
rect 7620 5390 7640 5430
rect 7680 5390 7700 5430
rect 7620 5330 7700 5390
rect 7620 5290 7640 5330
rect 7680 5290 7700 5330
rect 7620 5230 7700 5290
rect 7620 5190 7640 5230
rect 7680 5190 7700 5230
rect 7620 5130 7700 5190
rect 7620 5090 7640 5130
rect 7680 5090 7700 5130
rect 7620 5030 7700 5090
rect 7620 4990 7640 5030
rect 7680 4990 7700 5030
rect 7620 4930 7700 4990
rect 7620 4890 7640 4930
rect 7680 4890 7700 4930
rect 7620 4830 7700 4890
rect 7620 4790 7640 4830
rect 7680 4790 7700 4830
rect 7620 4730 7700 4790
rect 7620 4690 7640 4730
rect 7680 4690 7700 4730
rect 7620 4660 7700 4690
rect 7820 5430 7900 5460
rect 7820 5390 7840 5430
rect 7880 5390 7900 5430
rect 7820 5330 7900 5390
rect 7820 5290 7840 5330
rect 7880 5290 7900 5330
rect 7820 5230 7900 5290
rect 7820 5190 7840 5230
rect 7880 5190 7900 5230
rect 7820 5130 7900 5190
rect 7820 5090 7840 5130
rect 7880 5090 7900 5130
rect 7820 5030 7900 5090
rect 7820 4990 7840 5030
rect 7880 4990 7900 5030
rect 7820 4930 7900 4990
rect 7820 4890 7840 4930
rect 7880 4890 7900 4930
rect 7820 4830 7900 4890
rect 7820 4790 7840 4830
rect 7880 4790 7900 4830
rect 7820 4730 7900 4790
rect 7820 4690 7840 4730
rect 7880 4690 7900 4730
rect 7820 4660 7900 4690
rect 8020 5430 8100 5460
rect 8020 5390 8040 5430
rect 8080 5390 8100 5430
rect 8020 5330 8100 5390
rect 8020 5290 8040 5330
rect 8080 5290 8100 5330
rect 8020 5230 8100 5290
rect 8020 5190 8040 5230
rect 8080 5190 8100 5230
rect 8020 5130 8100 5190
rect 8020 5090 8040 5130
rect 8080 5090 8100 5130
rect 8020 5030 8100 5090
rect 8020 4990 8040 5030
rect 8080 4990 8100 5030
rect 8020 4930 8100 4990
rect 8020 4890 8040 4930
rect 8080 4890 8100 4930
rect 8020 4830 8100 4890
rect 8020 4790 8040 4830
rect 8080 4790 8100 4830
rect 8020 4730 8100 4790
rect 8020 4690 8040 4730
rect 8080 4690 8100 4730
rect 8020 4660 8100 4690
rect 8220 5430 8300 5460
rect 8220 5390 8240 5430
rect 8280 5390 8300 5430
rect 8220 5330 8300 5390
rect 8220 5290 8240 5330
rect 8280 5290 8300 5330
rect 8220 5230 8300 5290
rect 8220 5190 8240 5230
rect 8280 5190 8300 5230
rect 8220 5130 8300 5190
rect 8220 5090 8240 5130
rect 8280 5090 8300 5130
rect 8220 5030 8300 5090
rect 8220 4990 8240 5030
rect 8280 4990 8300 5030
rect 8220 4930 8300 4990
rect 8220 4890 8240 4930
rect 8280 4890 8300 4930
rect 8220 4830 8300 4890
rect 8220 4790 8240 4830
rect 8280 4790 8300 4830
rect 8220 4730 8300 4790
rect 8220 4690 8240 4730
rect 8280 4690 8300 4730
rect 8220 4660 8300 4690
rect 5220 4190 5300 4220
rect 5220 4150 5240 4190
rect 5280 4150 5300 4190
rect 5220 4090 5300 4150
rect 5220 4050 5240 4090
rect 5280 4050 5300 4090
rect 5220 3990 5300 4050
rect 5220 3950 5240 3990
rect 5280 3950 5300 3990
rect 5220 3890 5300 3950
rect 5220 3850 5240 3890
rect 5280 3850 5300 3890
rect 5220 3820 5300 3850
rect 5420 4190 5500 4220
rect 5420 4150 5440 4190
rect 5480 4150 5500 4190
rect 5420 4090 5500 4150
rect 5420 4050 5440 4090
rect 5480 4050 5500 4090
rect 5420 3990 5500 4050
rect 5420 3950 5440 3990
rect 5480 3950 5500 3990
rect 5420 3890 5500 3950
rect 5420 3850 5440 3890
rect 5480 3850 5500 3890
rect 5420 3820 5500 3850
rect 5620 4190 5700 4220
rect 5620 4150 5640 4190
rect 5680 4150 5700 4190
rect 5620 4090 5700 4150
rect 5620 4050 5640 4090
rect 5680 4050 5700 4090
rect 5620 3990 5700 4050
rect 5620 3950 5640 3990
rect 5680 3950 5700 3990
rect 5620 3890 5700 3950
rect 5620 3850 5640 3890
rect 5680 3850 5700 3890
rect 5620 3820 5700 3850
rect 5820 4190 5900 4220
rect 5820 4150 5840 4190
rect 5880 4150 5900 4190
rect 5820 4090 5900 4150
rect 5820 4050 5840 4090
rect 5880 4050 5900 4090
rect 5820 3990 5900 4050
rect 5820 3950 5840 3990
rect 5880 3950 5900 3990
rect 5820 3890 5900 3950
rect 5820 3850 5840 3890
rect 5880 3850 5900 3890
rect 5820 3820 5900 3850
rect 6020 4190 6100 4220
rect 6020 4150 6040 4190
rect 6080 4150 6100 4190
rect 6020 4090 6100 4150
rect 6020 4050 6040 4090
rect 6080 4050 6100 4090
rect 6020 3990 6100 4050
rect 6020 3950 6040 3990
rect 6080 3950 6100 3990
rect 6020 3890 6100 3950
rect 6020 3850 6040 3890
rect 6080 3850 6100 3890
rect 6020 3820 6100 3850
rect 6220 4190 6300 4220
rect 6220 4150 6240 4190
rect 6280 4150 6300 4190
rect 6220 4090 6300 4150
rect 6220 4050 6240 4090
rect 6280 4050 6300 4090
rect 6220 3990 6300 4050
rect 6220 3950 6240 3990
rect 6280 3950 6300 3990
rect 6220 3890 6300 3950
rect 6220 3850 6240 3890
rect 6280 3850 6300 3890
rect 6220 3820 6300 3850
rect 6420 4190 6500 4220
rect 6420 4150 6440 4190
rect 6480 4150 6500 4190
rect 6420 4090 6500 4150
rect 6420 4050 6440 4090
rect 6480 4050 6500 4090
rect 6420 3990 6500 4050
rect 6420 3950 6440 3990
rect 6480 3950 6500 3990
rect 6420 3890 6500 3950
rect 6420 3850 6440 3890
rect 6480 3850 6500 3890
rect 6420 3820 6500 3850
rect 6620 4190 6700 4220
rect 6620 4150 6640 4190
rect 6680 4150 6700 4190
rect 6620 4090 6700 4150
rect 6620 4050 6640 4090
rect 6680 4050 6700 4090
rect 6620 3990 6700 4050
rect 6620 3950 6640 3990
rect 6680 3950 6700 3990
rect 6620 3890 6700 3950
rect 6620 3850 6640 3890
rect 6680 3850 6700 3890
rect 6620 3820 6700 3850
rect 6820 4190 6900 4220
rect 6820 4150 6840 4190
rect 6880 4150 6900 4190
rect 6820 4090 6900 4150
rect 6820 4050 6840 4090
rect 6880 4050 6900 4090
rect 6820 3990 6900 4050
rect 6820 3950 6840 3990
rect 6880 3950 6900 3990
rect 6820 3890 6900 3950
rect 6820 3850 6840 3890
rect 6880 3850 6900 3890
rect 6820 3820 6900 3850
rect 7020 4190 7100 4220
rect 7020 4150 7040 4190
rect 7080 4150 7100 4190
rect 7020 4090 7100 4150
rect 7020 4050 7040 4090
rect 7080 4050 7100 4090
rect 7020 3990 7100 4050
rect 7020 3950 7040 3990
rect 7080 3950 7100 3990
rect 7020 3890 7100 3950
rect 7020 3850 7040 3890
rect 7080 3850 7100 3890
rect 7020 3820 7100 3850
rect 7220 4190 7300 4220
rect 7220 4150 7240 4190
rect 7280 4150 7300 4190
rect 7220 4090 7300 4150
rect 7220 4050 7240 4090
rect 7280 4050 7300 4090
rect 7220 3990 7300 4050
rect 7220 3950 7240 3990
rect 7280 3950 7300 3990
rect 7220 3890 7300 3950
rect 7220 3850 7240 3890
rect 7280 3850 7300 3890
rect 7220 3820 7300 3850
rect 7420 4190 7500 4220
rect 7420 4150 7440 4190
rect 7480 4150 7500 4190
rect 7420 4090 7500 4150
rect 7420 4050 7440 4090
rect 7480 4050 7500 4090
rect 7420 3990 7500 4050
rect 7420 3950 7440 3990
rect 7480 3950 7500 3990
rect 7420 3890 7500 3950
rect 7420 3850 7440 3890
rect 7480 3850 7500 3890
rect 7420 3820 7500 3850
rect 7620 4190 7700 4220
rect 7620 4150 7640 4190
rect 7680 4150 7700 4190
rect 7620 4090 7700 4150
rect 7620 4050 7640 4090
rect 7680 4050 7700 4090
rect 7620 3990 7700 4050
rect 7620 3950 7640 3990
rect 7680 3950 7700 3990
rect 7620 3890 7700 3950
rect 7620 3850 7640 3890
rect 7680 3850 7700 3890
rect 7620 3820 7700 3850
rect 8750 4190 8830 4220
rect 8750 4150 8770 4190
rect 8810 4150 8830 4190
rect 8750 4090 8830 4150
rect 8750 4050 8770 4090
rect 8810 4050 8830 4090
rect 8750 3990 8830 4050
rect 8750 3950 8770 3990
rect 8810 3950 8830 3990
rect 8750 3890 8830 3950
rect 8750 3850 8770 3890
rect 8810 3850 8830 3890
rect 8750 3820 8830 3850
rect 8860 4190 8940 4220
rect 8860 4150 8880 4190
rect 8920 4150 8940 4190
rect 8860 4090 8940 4150
rect 8860 4050 8880 4090
rect 8920 4050 8940 4090
rect 8860 3990 8940 4050
rect 8860 3950 8880 3990
rect 8920 3950 8940 3990
rect 8860 3890 8940 3950
rect 8860 3850 8880 3890
rect 8920 3850 8940 3890
rect 8860 3820 8940 3850
rect 9000 4190 9080 4220
rect 9000 4150 9020 4190
rect 9060 4150 9080 4190
rect 9000 4090 9080 4150
rect 9000 4050 9020 4090
rect 9060 4050 9080 4090
rect 9000 3990 9080 4050
rect 9000 3950 9020 3990
rect 9060 3950 9080 3990
rect 9000 3890 9080 3950
rect 9000 3850 9020 3890
rect 9060 3850 9080 3890
rect 9000 3820 9080 3850
rect 9110 4190 9190 4220
rect 9110 4150 9130 4190
rect 9170 4150 9190 4190
rect 9110 4090 9190 4150
rect 9110 4050 9130 4090
rect 9170 4050 9190 4090
rect 9110 3990 9190 4050
rect 9110 3950 9130 3990
rect 9170 3950 9190 3990
rect 9110 3890 9190 3950
rect 9110 3850 9130 3890
rect 9170 3850 9190 3890
rect 9110 3820 9190 3850
rect 1680 958 2360 1010
rect 1680 924 1734 958
rect 1768 924 1824 958
rect 1858 924 1914 958
rect 1948 924 2004 958
rect 2038 924 2094 958
rect 2128 924 2184 958
rect 2218 924 2274 958
rect 2308 924 2360 958
rect 1680 868 2360 924
rect 1680 834 1734 868
rect 1768 834 1824 868
rect 1858 834 1914 868
rect 1948 834 2004 868
rect 2038 834 2094 868
rect 2128 834 2184 868
rect 2218 834 2274 868
rect 2308 834 2360 868
rect 1680 778 2360 834
rect 1680 744 1734 778
rect 1768 744 1824 778
rect 1858 744 1914 778
rect 1948 744 2004 778
rect 2038 744 2094 778
rect 2128 744 2184 778
rect 2218 744 2274 778
rect 2308 744 2360 778
rect 1680 688 2360 744
rect 1680 654 1734 688
rect 1768 654 1824 688
rect 1858 654 1914 688
rect 1948 654 2004 688
rect 2038 654 2094 688
rect 2128 654 2184 688
rect 2218 654 2274 688
rect 2308 654 2360 688
rect 1680 598 2360 654
rect 1680 564 1734 598
rect 1768 564 1824 598
rect 1858 564 1914 598
rect 1948 564 2004 598
rect 2038 564 2094 598
rect 2128 564 2184 598
rect 2218 564 2274 598
rect 2308 564 2360 598
rect 1680 508 2360 564
rect 1680 474 1734 508
rect 1768 474 1824 508
rect 1858 474 1914 508
rect 1948 474 2004 508
rect 2038 474 2094 508
rect 2128 474 2184 508
rect 2218 474 2274 508
rect 2308 474 2360 508
rect 1680 418 2360 474
rect 1680 384 1734 418
rect 1768 384 1824 418
rect 1858 384 1914 418
rect 1948 384 2004 418
rect 2038 384 2094 418
rect 2128 384 2184 418
rect 2218 384 2274 418
rect 2308 384 2360 418
rect 1680 330 2360 384
rect 3040 958 3720 1010
rect 3040 924 3094 958
rect 3128 924 3184 958
rect 3218 924 3274 958
rect 3308 924 3364 958
rect 3398 924 3454 958
rect 3488 924 3544 958
rect 3578 924 3634 958
rect 3668 924 3720 958
rect 3040 868 3720 924
rect 3040 834 3094 868
rect 3128 834 3184 868
rect 3218 834 3274 868
rect 3308 834 3364 868
rect 3398 834 3454 868
rect 3488 834 3544 868
rect 3578 834 3634 868
rect 3668 834 3720 868
rect 3040 778 3720 834
rect 3040 744 3094 778
rect 3128 744 3184 778
rect 3218 744 3274 778
rect 3308 744 3364 778
rect 3398 744 3454 778
rect 3488 744 3544 778
rect 3578 744 3634 778
rect 3668 744 3720 778
rect 3040 688 3720 744
rect 3040 654 3094 688
rect 3128 654 3184 688
rect 3218 654 3274 688
rect 3308 654 3364 688
rect 3398 654 3454 688
rect 3488 654 3544 688
rect 3578 654 3634 688
rect 3668 654 3720 688
rect 3040 598 3720 654
rect 3040 564 3094 598
rect 3128 564 3184 598
rect 3218 564 3274 598
rect 3308 564 3364 598
rect 3398 564 3454 598
rect 3488 564 3544 598
rect 3578 564 3634 598
rect 3668 564 3720 598
rect 3040 508 3720 564
rect 3040 474 3094 508
rect 3128 474 3184 508
rect 3218 474 3274 508
rect 3308 474 3364 508
rect 3398 474 3454 508
rect 3488 474 3544 508
rect 3578 474 3634 508
rect 3668 474 3720 508
rect 3040 418 3720 474
rect 3040 384 3094 418
rect 3128 384 3184 418
rect 3218 384 3274 418
rect 3308 384 3364 418
rect 3398 384 3454 418
rect 3488 384 3544 418
rect 3578 384 3634 418
rect 3668 384 3720 418
rect 3040 330 3720 384
rect 4400 958 5080 1010
rect 4400 924 4454 958
rect 4488 924 4544 958
rect 4578 924 4634 958
rect 4668 924 4724 958
rect 4758 924 4814 958
rect 4848 924 4904 958
rect 4938 924 4994 958
rect 5028 924 5080 958
rect 4400 868 5080 924
rect 4400 834 4454 868
rect 4488 834 4544 868
rect 4578 834 4634 868
rect 4668 834 4724 868
rect 4758 834 4814 868
rect 4848 834 4904 868
rect 4938 834 4994 868
rect 5028 834 5080 868
rect 4400 778 5080 834
rect 4400 744 4454 778
rect 4488 744 4544 778
rect 4578 744 4634 778
rect 4668 744 4724 778
rect 4758 744 4814 778
rect 4848 744 4904 778
rect 4938 744 4994 778
rect 5028 744 5080 778
rect 4400 688 5080 744
rect 4400 654 4454 688
rect 4488 654 4544 688
rect 4578 654 4634 688
rect 4668 654 4724 688
rect 4758 654 4814 688
rect 4848 654 4904 688
rect 4938 654 4994 688
rect 5028 654 5080 688
rect 4400 598 5080 654
rect 4400 564 4454 598
rect 4488 564 4544 598
rect 4578 564 4634 598
rect 4668 564 4724 598
rect 4758 564 4814 598
rect 4848 564 4904 598
rect 4938 564 4994 598
rect 5028 564 5080 598
rect 4400 508 5080 564
rect 4400 474 4454 508
rect 4488 474 4544 508
rect 4578 474 4634 508
rect 4668 474 4724 508
rect 4758 474 4814 508
rect 4848 474 4904 508
rect 4938 474 4994 508
rect 5028 474 5080 508
rect 4400 418 5080 474
rect 4400 384 4454 418
rect 4488 384 4544 418
rect 4578 384 4634 418
rect 4668 384 4724 418
rect 4758 384 4814 418
rect 4848 384 4904 418
rect 4938 384 4994 418
rect 5028 384 5080 418
rect 4400 330 5080 384
rect 5760 958 6440 1010
rect 5760 924 5814 958
rect 5848 924 5904 958
rect 5938 924 5994 958
rect 6028 924 6084 958
rect 6118 924 6174 958
rect 6208 924 6264 958
rect 6298 924 6354 958
rect 6388 924 6440 958
rect 5760 868 6440 924
rect 5760 834 5814 868
rect 5848 834 5904 868
rect 5938 834 5994 868
rect 6028 834 6084 868
rect 6118 834 6174 868
rect 6208 834 6264 868
rect 6298 834 6354 868
rect 6388 834 6440 868
rect 5760 778 6440 834
rect 5760 744 5814 778
rect 5848 744 5904 778
rect 5938 744 5994 778
rect 6028 744 6084 778
rect 6118 744 6174 778
rect 6208 744 6264 778
rect 6298 744 6354 778
rect 6388 744 6440 778
rect 5760 688 6440 744
rect 5760 654 5814 688
rect 5848 654 5904 688
rect 5938 654 5994 688
rect 6028 654 6084 688
rect 6118 654 6174 688
rect 6208 654 6264 688
rect 6298 654 6354 688
rect 6388 654 6440 688
rect 5760 598 6440 654
rect 5760 564 5814 598
rect 5848 564 5904 598
rect 5938 564 5994 598
rect 6028 564 6084 598
rect 6118 564 6174 598
rect 6208 564 6264 598
rect 6298 564 6354 598
rect 6388 564 6440 598
rect 5760 508 6440 564
rect 5760 474 5814 508
rect 5848 474 5904 508
rect 5938 474 5994 508
rect 6028 474 6084 508
rect 6118 474 6174 508
rect 6208 474 6264 508
rect 6298 474 6354 508
rect 6388 474 6440 508
rect 5760 418 6440 474
rect 5760 384 5814 418
rect 5848 384 5904 418
rect 5938 384 5994 418
rect 6028 384 6084 418
rect 6118 384 6174 418
rect 6208 384 6264 418
rect 6298 384 6354 418
rect 6388 384 6440 418
rect 5760 330 6440 384
rect 7120 958 7800 1010
rect 7120 924 7174 958
rect 7208 924 7264 958
rect 7298 924 7354 958
rect 7388 924 7444 958
rect 7478 924 7534 958
rect 7568 924 7624 958
rect 7658 924 7714 958
rect 7748 924 7800 958
rect 7120 868 7800 924
rect 7120 834 7174 868
rect 7208 834 7264 868
rect 7298 834 7354 868
rect 7388 834 7444 868
rect 7478 834 7534 868
rect 7568 834 7624 868
rect 7658 834 7714 868
rect 7748 834 7800 868
rect 7120 778 7800 834
rect 7120 744 7174 778
rect 7208 744 7264 778
rect 7298 744 7354 778
rect 7388 744 7444 778
rect 7478 744 7534 778
rect 7568 744 7624 778
rect 7658 744 7714 778
rect 7748 744 7800 778
rect 7120 688 7800 744
rect 7120 654 7174 688
rect 7208 654 7264 688
rect 7298 654 7354 688
rect 7388 654 7444 688
rect 7478 654 7534 688
rect 7568 654 7624 688
rect 7658 654 7714 688
rect 7748 654 7800 688
rect 7120 598 7800 654
rect 7120 564 7174 598
rect 7208 564 7264 598
rect 7298 564 7354 598
rect 7388 564 7444 598
rect 7478 564 7534 598
rect 7568 564 7624 598
rect 7658 564 7714 598
rect 7748 564 7800 598
rect 7120 508 7800 564
rect 7120 474 7174 508
rect 7208 474 7264 508
rect 7298 474 7354 508
rect 7388 474 7444 508
rect 7478 474 7534 508
rect 7568 474 7624 508
rect 7658 474 7714 508
rect 7748 474 7800 508
rect 7120 418 7800 474
rect 7120 384 7174 418
rect 7208 384 7264 418
rect 7298 384 7354 418
rect 7388 384 7444 418
rect 7478 384 7534 418
rect 7568 384 7624 418
rect 7658 384 7714 418
rect 7748 384 7800 418
rect 7120 330 7800 384
rect 8480 958 9160 1010
rect 8480 924 8534 958
rect 8568 924 8624 958
rect 8658 924 8714 958
rect 8748 924 8804 958
rect 8838 924 8894 958
rect 8928 924 8984 958
rect 9018 924 9074 958
rect 9108 924 9160 958
rect 8480 868 9160 924
rect 8480 834 8534 868
rect 8568 834 8624 868
rect 8658 834 8714 868
rect 8748 834 8804 868
rect 8838 834 8894 868
rect 8928 834 8984 868
rect 9018 834 9074 868
rect 9108 834 9160 868
rect 8480 778 9160 834
rect 8480 744 8534 778
rect 8568 744 8624 778
rect 8658 744 8714 778
rect 8748 744 8804 778
rect 8838 744 8894 778
rect 8928 744 8984 778
rect 9018 744 9074 778
rect 9108 744 9160 778
rect 8480 688 9160 744
rect 8480 654 8534 688
rect 8568 654 8624 688
rect 8658 654 8714 688
rect 8748 654 8804 688
rect 8838 654 8894 688
rect 8928 654 8984 688
rect 9018 654 9074 688
rect 9108 654 9160 688
rect 8480 598 9160 654
rect 8480 564 8534 598
rect 8568 564 8624 598
rect 8658 564 8714 598
rect 8748 564 8804 598
rect 8838 564 8894 598
rect 8928 564 8984 598
rect 9018 564 9074 598
rect 9108 564 9160 598
rect 8480 508 9160 564
rect 8480 474 8534 508
rect 8568 474 8624 508
rect 8658 474 8714 508
rect 8748 474 8804 508
rect 8838 474 8894 508
rect 8928 474 8984 508
rect 9018 474 9074 508
rect 9108 474 9160 508
rect 8480 418 9160 474
rect 8480 384 8534 418
rect 8568 384 8624 418
rect 8658 384 8714 418
rect 8748 384 8804 418
rect 8838 384 8894 418
rect 8928 384 8984 418
rect 9018 384 9074 418
rect 9108 384 9160 418
rect 8480 330 9160 384
<< ndiffc >>
rect 5640 3250 5680 3290
rect 5640 3150 5680 3190
rect 5840 3250 5880 3290
rect 5840 3150 5880 3190
rect 6040 3250 6080 3290
rect 6040 3150 6080 3190
rect 6240 3250 6280 3290
rect 6240 3150 6280 3190
rect 6440 3250 6480 3290
rect 6440 3150 6480 3190
rect 6640 3250 6680 3290
rect 6640 3150 6680 3190
rect 6840 3250 6880 3290
rect 6840 3150 6880 3190
rect 7040 3250 7080 3290
rect 7040 3150 7080 3190
rect 7240 3250 7280 3290
rect 7240 3150 7280 3190
rect 5480 2700 5520 2740
rect 5480 2600 5520 2640
rect 5480 2500 5520 2540
rect 5480 2400 5520 2440
rect 5480 2300 5520 2340
rect 5480 2200 5520 2240
rect 5480 2100 5520 2140
rect 5480 2000 5520 2040
rect 6360 2700 6400 2740
rect 6520 2700 6560 2740
rect 6360 2600 6400 2640
rect 6520 2600 6560 2640
rect 6360 2500 6400 2540
rect 6520 2500 6560 2540
rect 6360 2400 6400 2440
rect 6520 2400 6560 2440
rect 6360 2300 6400 2340
rect 6520 2300 6560 2340
rect 6360 2200 6400 2240
rect 6520 2200 6560 2240
rect 6360 2100 6400 2140
rect 6520 2100 6560 2140
rect 6360 2000 6400 2040
rect 6520 2000 6560 2040
rect 7400 2700 7440 2740
rect 7400 2600 7440 2640
rect 7400 2500 7440 2540
rect 7400 2400 7440 2440
rect 7400 2300 7440 2340
rect 7400 2200 7440 2240
rect 7400 2100 7440 2140
rect 7400 2000 7440 2040
rect 5380 1640 5420 1680
rect 5380 1540 5420 1580
rect 7460 1640 7500 1680
rect 7460 1540 7500 1580
<< pdiffc >>
rect 4640 5390 4680 5430
rect 4640 5290 4680 5330
rect 4640 5190 4680 5230
rect 4640 5090 4680 5130
rect 4640 4990 4680 5030
rect 4640 4890 4680 4930
rect 4640 4790 4680 4830
rect 4640 4690 4680 4730
rect 4840 5390 4880 5430
rect 4840 5290 4880 5330
rect 4840 5190 4880 5230
rect 4840 5090 4880 5130
rect 4840 4990 4880 5030
rect 4840 4890 4880 4930
rect 4840 4790 4880 4830
rect 4840 4690 4880 4730
rect 5040 5390 5080 5430
rect 5040 5290 5080 5330
rect 5040 5190 5080 5230
rect 5040 5090 5080 5130
rect 5040 4990 5080 5030
rect 5040 4890 5080 4930
rect 5040 4790 5080 4830
rect 5040 4690 5080 4730
rect 5240 5390 5280 5430
rect 5240 5290 5280 5330
rect 5240 5190 5280 5230
rect 5240 5090 5280 5130
rect 5240 4990 5280 5030
rect 5240 4890 5280 4930
rect 5240 4790 5280 4830
rect 5240 4690 5280 4730
rect 5440 5390 5480 5430
rect 5440 5290 5480 5330
rect 5440 5190 5480 5230
rect 5440 5090 5480 5130
rect 5440 4990 5480 5030
rect 5440 4890 5480 4930
rect 5440 4790 5480 4830
rect 5440 4690 5480 4730
rect 5640 5390 5680 5430
rect 5640 5290 5680 5330
rect 5640 5190 5680 5230
rect 5640 5090 5680 5130
rect 5640 4990 5680 5030
rect 5640 4890 5680 4930
rect 5640 4790 5680 4830
rect 5640 4690 5680 4730
rect 5840 5390 5880 5430
rect 5840 5290 5880 5330
rect 5840 5190 5880 5230
rect 5840 5090 5880 5130
rect 5840 4990 5880 5030
rect 5840 4890 5880 4930
rect 5840 4790 5880 4830
rect 5840 4690 5880 4730
rect 6040 5390 6080 5430
rect 6040 5290 6080 5330
rect 6040 5190 6080 5230
rect 6040 5090 6080 5130
rect 6040 4990 6080 5030
rect 6040 4890 6080 4930
rect 6040 4790 6080 4830
rect 6040 4690 6080 4730
rect 6240 5390 6280 5430
rect 6240 5290 6280 5330
rect 6240 5190 6280 5230
rect 6240 5090 6280 5130
rect 6240 4990 6280 5030
rect 6240 4890 6280 4930
rect 6240 4790 6280 4830
rect 6240 4690 6280 4730
rect 6440 5390 6480 5430
rect 6440 5290 6480 5330
rect 6440 5190 6480 5230
rect 6440 5090 6480 5130
rect 6440 4990 6480 5030
rect 6440 4890 6480 4930
rect 6440 4790 6480 4830
rect 6440 4690 6480 4730
rect 6640 5390 6680 5430
rect 6640 5290 6680 5330
rect 6640 5190 6680 5230
rect 6640 5090 6680 5130
rect 6640 4990 6680 5030
rect 6640 4890 6680 4930
rect 6640 4790 6680 4830
rect 6640 4690 6680 4730
rect 6840 5390 6880 5430
rect 6840 5290 6880 5330
rect 6840 5190 6880 5230
rect 6840 5090 6880 5130
rect 6840 4990 6880 5030
rect 6840 4890 6880 4930
rect 6840 4790 6880 4830
rect 6840 4690 6880 4730
rect 7040 5390 7080 5430
rect 7040 5290 7080 5330
rect 7040 5190 7080 5230
rect 7040 5090 7080 5130
rect 7040 4990 7080 5030
rect 7040 4890 7080 4930
rect 7040 4790 7080 4830
rect 7040 4690 7080 4730
rect 7240 5390 7280 5430
rect 7240 5290 7280 5330
rect 7240 5190 7280 5230
rect 7240 5090 7280 5130
rect 7240 4990 7280 5030
rect 7240 4890 7280 4930
rect 7240 4790 7280 4830
rect 7240 4690 7280 4730
rect 7440 5390 7480 5430
rect 7440 5290 7480 5330
rect 7440 5190 7480 5230
rect 7440 5090 7480 5130
rect 7440 4990 7480 5030
rect 7440 4890 7480 4930
rect 7440 4790 7480 4830
rect 7440 4690 7480 4730
rect 7640 5390 7680 5430
rect 7640 5290 7680 5330
rect 7640 5190 7680 5230
rect 7640 5090 7680 5130
rect 7640 4990 7680 5030
rect 7640 4890 7680 4930
rect 7640 4790 7680 4830
rect 7640 4690 7680 4730
rect 7840 5390 7880 5430
rect 7840 5290 7880 5330
rect 7840 5190 7880 5230
rect 7840 5090 7880 5130
rect 7840 4990 7880 5030
rect 7840 4890 7880 4930
rect 7840 4790 7880 4830
rect 7840 4690 7880 4730
rect 8040 5390 8080 5430
rect 8040 5290 8080 5330
rect 8040 5190 8080 5230
rect 8040 5090 8080 5130
rect 8040 4990 8080 5030
rect 8040 4890 8080 4930
rect 8040 4790 8080 4830
rect 8040 4690 8080 4730
rect 8240 5390 8280 5430
rect 8240 5290 8280 5330
rect 8240 5190 8280 5230
rect 8240 5090 8280 5130
rect 8240 4990 8280 5030
rect 8240 4890 8280 4930
rect 8240 4790 8280 4830
rect 8240 4690 8280 4730
rect 5240 4150 5280 4190
rect 5240 4050 5280 4090
rect 5240 3950 5280 3990
rect 5240 3850 5280 3890
rect 5440 4150 5480 4190
rect 5440 4050 5480 4090
rect 5440 3950 5480 3990
rect 5440 3850 5480 3890
rect 5640 4150 5680 4190
rect 5640 4050 5680 4090
rect 5640 3950 5680 3990
rect 5640 3850 5680 3890
rect 5840 4150 5880 4190
rect 5840 4050 5880 4090
rect 5840 3950 5880 3990
rect 5840 3850 5880 3890
rect 6040 4150 6080 4190
rect 6040 4050 6080 4090
rect 6040 3950 6080 3990
rect 6040 3850 6080 3890
rect 6240 4150 6280 4190
rect 6240 4050 6280 4090
rect 6240 3950 6280 3990
rect 6240 3850 6280 3890
rect 6440 4150 6480 4190
rect 6440 4050 6480 4090
rect 6440 3950 6480 3990
rect 6440 3850 6480 3890
rect 6640 4150 6680 4190
rect 6640 4050 6680 4090
rect 6640 3950 6680 3990
rect 6640 3850 6680 3890
rect 6840 4150 6880 4190
rect 6840 4050 6880 4090
rect 6840 3950 6880 3990
rect 6840 3850 6880 3890
rect 7040 4150 7080 4190
rect 7040 4050 7080 4090
rect 7040 3950 7080 3990
rect 7040 3850 7080 3890
rect 7240 4150 7280 4190
rect 7240 4050 7280 4090
rect 7240 3950 7280 3990
rect 7240 3850 7280 3890
rect 7440 4150 7480 4190
rect 7440 4050 7480 4090
rect 7440 3950 7480 3990
rect 7440 3850 7480 3890
rect 7640 4150 7680 4190
rect 7640 4050 7680 4090
rect 7640 3950 7680 3990
rect 7640 3850 7680 3890
rect 8770 4150 8810 4190
rect 8770 4050 8810 4090
rect 8770 3950 8810 3990
rect 8770 3850 8810 3890
rect 8880 4150 8920 4190
rect 8880 4050 8920 4090
rect 8880 3950 8920 3990
rect 8880 3850 8920 3890
rect 9020 4150 9060 4190
rect 9020 4050 9060 4090
rect 9020 3950 9060 3990
rect 9020 3850 9060 3890
rect 9130 4150 9170 4190
rect 9130 4050 9170 4090
rect 9130 3950 9170 3990
rect 9130 3850 9170 3890
rect 1734 924 1768 958
rect 1824 924 1858 958
rect 1914 924 1948 958
rect 2004 924 2038 958
rect 2094 924 2128 958
rect 2184 924 2218 958
rect 2274 924 2308 958
rect 1734 834 1768 868
rect 1824 834 1858 868
rect 1914 834 1948 868
rect 2004 834 2038 868
rect 2094 834 2128 868
rect 2184 834 2218 868
rect 2274 834 2308 868
rect 1734 744 1768 778
rect 1824 744 1858 778
rect 1914 744 1948 778
rect 2004 744 2038 778
rect 2094 744 2128 778
rect 2184 744 2218 778
rect 2274 744 2308 778
rect 1734 654 1768 688
rect 1824 654 1858 688
rect 1914 654 1948 688
rect 2004 654 2038 688
rect 2094 654 2128 688
rect 2184 654 2218 688
rect 2274 654 2308 688
rect 1734 564 1768 598
rect 1824 564 1858 598
rect 1914 564 1948 598
rect 2004 564 2038 598
rect 2094 564 2128 598
rect 2184 564 2218 598
rect 2274 564 2308 598
rect 1734 474 1768 508
rect 1824 474 1858 508
rect 1914 474 1948 508
rect 2004 474 2038 508
rect 2094 474 2128 508
rect 2184 474 2218 508
rect 2274 474 2308 508
rect 1734 384 1768 418
rect 1824 384 1858 418
rect 1914 384 1948 418
rect 2004 384 2038 418
rect 2094 384 2128 418
rect 2184 384 2218 418
rect 2274 384 2308 418
rect 3094 924 3128 958
rect 3184 924 3218 958
rect 3274 924 3308 958
rect 3364 924 3398 958
rect 3454 924 3488 958
rect 3544 924 3578 958
rect 3634 924 3668 958
rect 3094 834 3128 868
rect 3184 834 3218 868
rect 3274 834 3308 868
rect 3364 834 3398 868
rect 3454 834 3488 868
rect 3544 834 3578 868
rect 3634 834 3668 868
rect 3094 744 3128 778
rect 3184 744 3218 778
rect 3274 744 3308 778
rect 3364 744 3398 778
rect 3454 744 3488 778
rect 3544 744 3578 778
rect 3634 744 3668 778
rect 3094 654 3128 688
rect 3184 654 3218 688
rect 3274 654 3308 688
rect 3364 654 3398 688
rect 3454 654 3488 688
rect 3544 654 3578 688
rect 3634 654 3668 688
rect 3094 564 3128 598
rect 3184 564 3218 598
rect 3274 564 3308 598
rect 3364 564 3398 598
rect 3454 564 3488 598
rect 3544 564 3578 598
rect 3634 564 3668 598
rect 3094 474 3128 508
rect 3184 474 3218 508
rect 3274 474 3308 508
rect 3364 474 3398 508
rect 3454 474 3488 508
rect 3544 474 3578 508
rect 3634 474 3668 508
rect 3094 384 3128 418
rect 3184 384 3218 418
rect 3274 384 3308 418
rect 3364 384 3398 418
rect 3454 384 3488 418
rect 3544 384 3578 418
rect 3634 384 3668 418
rect 4454 924 4488 958
rect 4544 924 4578 958
rect 4634 924 4668 958
rect 4724 924 4758 958
rect 4814 924 4848 958
rect 4904 924 4938 958
rect 4994 924 5028 958
rect 4454 834 4488 868
rect 4544 834 4578 868
rect 4634 834 4668 868
rect 4724 834 4758 868
rect 4814 834 4848 868
rect 4904 834 4938 868
rect 4994 834 5028 868
rect 4454 744 4488 778
rect 4544 744 4578 778
rect 4634 744 4668 778
rect 4724 744 4758 778
rect 4814 744 4848 778
rect 4904 744 4938 778
rect 4994 744 5028 778
rect 4454 654 4488 688
rect 4544 654 4578 688
rect 4634 654 4668 688
rect 4724 654 4758 688
rect 4814 654 4848 688
rect 4904 654 4938 688
rect 4994 654 5028 688
rect 4454 564 4488 598
rect 4544 564 4578 598
rect 4634 564 4668 598
rect 4724 564 4758 598
rect 4814 564 4848 598
rect 4904 564 4938 598
rect 4994 564 5028 598
rect 4454 474 4488 508
rect 4544 474 4578 508
rect 4634 474 4668 508
rect 4724 474 4758 508
rect 4814 474 4848 508
rect 4904 474 4938 508
rect 4994 474 5028 508
rect 4454 384 4488 418
rect 4544 384 4578 418
rect 4634 384 4668 418
rect 4724 384 4758 418
rect 4814 384 4848 418
rect 4904 384 4938 418
rect 4994 384 5028 418
rect 5814 924 5848 958
rect 5904 924 5938 958
rect 5994 924 6028 958
rect 6084 924 6118 958
rect 6174 924 6208 958
rect 6264 924 6298 958
rect 6354 924 6388 958
rect 5814 834 5848 868
rect 5904 834 5938 868
rect 5994 834 6028 868
rect 6084 834 6118 868
rect 6174 834 6208 868
rect 6264 834 6298 868
rect 6354 834 6388 868
rect 5814 744 5848 778
rect 5904 744 5938 778
rect 5994 744 6028 778
rect 6084 744 6118 778
rect 6174 744 6208 778
rect 6264 744 6298 778
rect 6354 744 6388 778
rect 5814 654 5848 688
rect 5904 654 5938 688
rect 5994 654 6028 688
rect 6084 654 6118 688
rect 6174 654 6208 688
rect 6264 654 6298 688
rect 6354 654 6388 688
rect 5814 564 5848 598
rect 5904 564 5938 598
rect 5994 564 6028 598
rect 6084 564 6118 598
rect 6174 564 6208 598
rect 6264 564 6298 598
rect 6354 564 6388 598
rect 5814 474 5848 508
rect 5904 474 5938 508
rect 5994 474 6028 508
rect 6084 474 6118 508
rect 6174 474 6208 508
rect 6264 474 6298 508
rect 6354 474 6388 508
rect 5814 384 5848 418
rect 5904 384 5938 418
rect 5994 384 6028 418
rect 6084 384 6118 418
rect 6174 384 6208 418
rect 6264 384 6298 418
rect 6354 384 6388 418
rect 7174 924 7208 958
rect 7264 924 7298 958
rect 7354 924 7388 958
rect 7444 924 7478 958
rect 7534 924 7568 958
rect 7624 924 7658 958
rect 7714 924 7748 958
rect 7174 834 7208 868
rect 7264 834 7298 868
rect 7354 834 7388 868
rect 7444 834 7478 868
rect 7534 834 7568 868
rect 7624 834 7658 868
rect 7714 834 7748 868
rect 7174 744 7208 778
rect 7264 744 7298 778
rect 7354 744 7388 778
rect 7444 744 7478 778
rect 7534 744 7568 778
rect 7624 744 7658 778
rect 7714 744 7748 778
rect 7174 654 7208 688
rect 7264 654 7298 688
rect 7354 654 7388 688
rect 7444 654 7478 688
rect 7534 654 7568 688
rect 7624 654 7658 688
rect 7714 654 7748 688
rect 7174 564 7208 598
rect 7264 564 7298 598
rect 7354 564 7388 598
rect 7444 564 7478 598
rect 7534 564 7568 598
rect 7624 564 7658 598
rect 7714 564 7748 598
rect 7174 474 7208 508
rect 7264 474 7298 508
rect 7354 474 7388 508
rect 7444 474 7478 508
rect 7534 474 7568 508
rect 7624 474 7658 508
rect 7714 474 7748 508
rect 7174 384 7208 418
rect 7264 384 7298 418
rect 7354 384 7388 418
rect 7444 384 7478 418
rect 7534 384 7568 418
rect 7624 384 7658 418
rect 7714 384 7748 418
rect 8534 924 8568 958
rect 8624 924 8658 958
rect 8714 924 8748 958
rect 8804 924 8838 958
rect 8894 924 8928 958
rect 8984 924 9018 958
rect 9074 924 9108 958
rect 8534 834 8568 868
rect 8624 834 8658 868
rect 8714 834 8748 868
rect 8804 834 8838 868
rect 8894 834 8928 868
rect 8984 834 9018 868
rect 9074 834 9108 868
rect 8534 744 8568 778
rect 8624 744 8658 778
rect 8714 744 8748 778
rect 8804 744 8838 778
rect 8894 744 8928 778
rect 8984 744 9018 778
rect 9074 744 9108 778
rect 8534 654 8568 688
rect 8624 654 8658 688
rect 8714 654 8748 688
rect 8804 654 8838 688
rect 8894 654 8928 688
rect 8984 654 9018 688
rect 9074 654 9108 688
rect 8534 564 8568 598
rect 8624 564 8658 598
rect 8714 564 8748 598
rect 8804 564 8838 598
rect 8894 564 8928 598
rect 8984 564 9018 598
rect 9074 564 9108 598
rect 8534 474 8568 508
rect 8624 474 8658 508
rect 8714 474 8748 508
rect 8804 474 8838 508
rect 8894 474 8928 508
rect 8984 474 9018 508
rect 9074 474 9108 508
rect 8534 384 8568 418
rect 8624 384 8658 418
rect 8714 384 8748 418
rect 8804 384 8838 418
rect 8894 384 8928 418
rect 8984 384 9018 418
rect 9074 384 9108 418
<< psubdiff >>
rect 6420 2740 6500 2770
rect 6420 2700 6440 2740
rect 6480 2700 6500 2740
rect 6420 2640 6500 2700
rect 6420 2600 6440 2640
rect 6480 2600 6500 2640
rect 6420 2540 6500 2600
rect 6420 2500 6440 2540
rect 6480 2500 6500 2540
rect 6420 2440 6500 2500
rect 6420 2400 6440 2440
rect 6480 2400 6500 2440
rect 6420 2340 6500 2400
rect 6420 2300 6440 2340
rect 6480 2300 6500 2340
rect 6420 2240 6500 2300
rect 6420 2200 6440 2240
rect 6480 2200 6500 2240
rect 6420 2140 6500 2200
rect 6420 2100 6440 2140
rect 6480 2100 6500 2140
rect 6420 2040 6500 2100
rect 6420 2000 6440 2040
rect 6480 2000 6500 2040
rect 6420 1970 6500 2000
rect 1290 1640 1390 1670
rect 1290 1600 1320 1640
rect 1360 1600 1390 1640
rect 1290 1540 1390 1600
rect 1290 1500 1320 1540
rect 1360 1500 1390 1540
rect 7520 1680 7600 1710
rect 7520 1640 7540 1680
rect 7580 1640 7600 1680
rect 7520 1580 7600 1640
rect 7520 1540 7540 1580
rect 7580 1540 7600 1580
rect 7520 1510 7600 1540
rect 1290 1440 1390 1500
rect 1290 1400 1320 1440
rect 1360 1400 1390 1440
rect 1290 1370 1390 1400
rect 1376 1279 2664 1314
rect 1376 1256 1506 1279
rect 1376 1222 1410 1256
rect 1444 1245 1506 1256
rect 1540 1245 1596 1279
rect 1630 1245 1686 1279
rect 1720 1245 1776 1279
rect 1810 1245 1866 1279
rect 1900 1245 1956 1279
rect 1990 1245 2046 1279
rect 2080 1245 2136 1279
rect 2170 1245 2226 1279
rect 2260 1245 2316 1279
rect 2350 1245 2406 1279
rect 2440 1245 2496 1279
rect 2530 1256 2664 1279
rect 2530 1245 2597 1256
rect 1444 1222 2597 1245
rect 2631 1222 2664 1256
rect 1376 1213 2664 1222
rect 1376 1166 1477 1213
rect 1376 1132 1410 1166
rect 1444 1132 1477 1166
rect 2563 1166 2664 1213
rect 1376 1076 1477 1132
rect 1376 1042 1410 1076
rect 1444 1042 1477 1076
rect 1376 986 1477 1042
rect 1376 952 1410 986
rect 1444 952 1477 986
rect 1376 896 1477 952
rect 1376 862 1410 896
rect 1444 862 1477 896
rect 1376 806 1477 862
rect 1376 772 1410 806
rect 1444 772 1477 806
rect 1376 716 1477 772
rect 1376 682 1410 716
rect 1444 682 1477 716
rect 1376 626 1477 682
rect 1376 592 1410 626
rect 1444 592 1477 626
rect 1376 536 1477 592
rect 1376 502 1410 536
rect 1444 502 1477 536
rect 1376 446 1477 502
rect 1376 412 1410 446
rect 1444 412 1477 446
rect 1376 356 1477 412
rect 1376 322 1410 356
rect 1444 322 1477 356
rect 1376 266 1477 322
rect 1376 232 1410 266
rect 1444 232 1477 266
rect 1376 176 1477 232
rect 2563 1132 2597 1166
rect 2631 1132 2664 1166
rect 2563 1076 2664 1132
rect 2563 1042 2597 1076
rect 2631 1042 2664 1076
rect 2563 986 2664 1042
rect 2563 952 2597 986
rect 2631 952 2664 986
rect 2563 896 2664 952
rect 2563 862 2597 896
rect 2631 862 2664 896
rect 2563 806 2664 862
rect 2563 772 2597 806
rect 2631 772 2664 806
rect 2563 716 2664 772
rect 2563 682 2597 716
rect 2631 682 2664 716
rect 2563 626 2664 682
rect 2563 592 2597 626
rect 2631 592 2664 626
rect 2563 536 2664 592
rect 2563 502 2597 536
rect 2631 502 2664 536
rect 2563 446 2664 502
rect 2563 412 2597 446
rect 2631 412 2664 446
rect 2563 356 2664 412
rect 2563 322 2597 356
rect 2631 322 2664 356
rect 2563 266 2664 322
rect 2563 232 2597 266
rect 2631 232 2664 266
rect 1376 142 1410 176
rect 1444 142 1477 176
rect 1376 127 1477 142
rect 2563 176 2664 232
rect 2563 142 2597 176
rect 2631 142 2664 176
rect 2563 127 2664 142
rect 1376 92 2664 127
rect 40 50 80 90
rect 1376 58 1506 92
rect 1540 58 1596 92
rect 1630 58 1686 92
rect 1720 58 1776 92
rect 1810 58 1866 92
rect 1900 58 1956 92
rect 1990 58 2046 92
rect 2080 58 2136 92
rect 2170 58 2226 92
rect 2260 58 2316 92
rect 2350 58 2406 92
rect 2440 58 2496 92
rect 2530 58 2664 92
rect 1376 26 2664 58
rect 2736 1279 4024 1314
rect 2736 1256 2866 1279
rect 2736 1222 2770 1256
rect 2804 1245 2866 1256
rect 2900 1245 2956 1279
rect 2990 1245 3046 1279
rect 3080 1245 3136 1279
rect 3170 1245 3226 1279
rect 3260 1245 3316 1279
rect 3350 1245 3406 1279
rect 3440 1245 3496 1279
rect 3530 1245 3586 1279
rect 3620 1245 3676 1279
rect 3710 1245 3766 1279
rect 3800 1245 3856 1279
rect 3890 1256 4024 1279
rect 3890 1245 3957 1256
rect 2804 1222 3957 1245
rect 3991 1222 4024 1256
rect 2736 1213 4024 1222
rect 2736 1166 2837 1213
rect 2736 1132 2770 1166
rect 2804 1132 2837 1166
rect 3923 1166 4024 1213
rect 2736 1076 2837 1132
rect 2736 1042 2770 1076
rect 2804 1042 2837 1076
rect 2736 986 2837 1042
rect 2736 952 2770 986
rect 2804 952 2837 986
rect 2736 896 2837 952
rect 2736 862 2770 896
rect 2804 862 2837 896
rect 2736 806 2837 862
rect 2736 772 2770 806
rect 2804 772 2837 806
rect 2736 716 2837 772
rect 2736 682 2770 716
rect 2804 682 2837 716
rect 2736 626 2837 682
rect 2736 592 2770 626
rect 2804 592 2837 626
rect 2736 536 2837 592
rect 2736 502 2770 536
rect 2804 502 2837 536
rect 2736 446 2837 502
rect 2736 412 2770 446
rect 2804 412 2837 446
rect 2736 356 2837 412
rect 2736 322 2770 356
rect 2804 322 2837 356
rect 2736 266 2837 322
rect 2736 232 2770 266
rect 2804 232 2837 266
rect 2736 176 2837 232
rect 3923 1132 3957 1166
rect 3991 1132 4024 1166
rect 3923 1076 4024 1132
rect 3923 1042 3957 1076
rect 3991 1042 4024 1076
rect 3923 986 4024 1042
rect 3923 952 3957 986
rect 3991 952 4024 986
rect 3923 896 4024 952
rect 3923 862 3957 896
rect 3991 862 4024 896
rect 3923 806 4024 862
rect 3923 772 3957 806
rect 3991 772 4024 806
rect 3923 716 4024 772
rect 3923 682 3957 716
rect 3991 682 4024 716
rect 3923 626 4024 682
rect 3923 592 3957 626
rect 3991 592 4024 626
rect 3923 536 4024 592
rect 3923 502 3957 536
rect 3991 502 4024 536
rect 3923 446 4024 502
rect 3923 412 3957 446
rect 3991 412 4024 446
rect 3923 356 4024 412
rect 3923 322 3957 356
rect 3991 322 4024 356
rect 3923 266 4024 322
rect 3923 232 3957 266
rect 3991 232 4024 266
rect 2736 142 2770 176
rect 2804 142 2837 176
rect 2736 127 2837 142
rect 3923 176 4024 232
rect 3923 142 3957 176
rect 3991 142 4024 176
rect 3923 127 4024 142
rect 2736 92 4024 127
rect 2736 58 2866 92
rect 2900 58 2956 92
rect 2990 58 3046 92
rect 3080 58 3136 92
rect 3170 58 3226 92
rect 3260 58 3316 92
rect 3350 58 3406 92
rect 3440 58 3496 92
rect 3530 58 3586 92
rect 3620 58 3676 92
rect 3710 58 3766 92
rect 3800 58 3856 92
rect 3890 58 4024 92
rect 2736 26 4024 58
rect 4096 1279 5384 1314
rect 4096 1256 4226 1279
rect 4096 1222 4130 1256
rect 4164 1245 4226 1256
rect 4260 1245 4316 1279
rect 4350 1245 4406 1279
rect 4440 1245 4496 1279
rect 4530 1245 4586 1279
rect 4620 1245 4676 1279
rect 4710 1245 4766 1279
rect 4800 1245 4856 1279
rect 4890 1245 4946 1279
rect 4980 1245 5036 1279
rect 5070 1245 5126 1279
rect 5160 1245 5216 1279
rect 5250 1256 5384 1279
rect 5250 1245 5317 1256
rect 4164 1222 5317 1245
rect 5351 1222 5384 1256
rect 4096 1213 5384 1222
rect 4096 1166 4197 1213
rect 4096 1132 4130 1166
rect 4164 1132 4197 1166
rect 5283 1166 5384 1213
rect 4096 1076 4197 1132
rect 4096 1042 4130 1076
rect 4164 1042 4197 1076
rect 4096 986 4197 1042
rect 4096 952 4130 986
rect 4164 952 4197 986
rect 4096 896 4197 952
rect 4096 862 4130 896
rect 4164 862 4197 896
rect 4096 806 4197 862
rect 4096 772 4130 806
rect 4164 772 4197 806
rect 4096 716 4197 772
rect 4096 682 4130 716
rect 4164 682 4197 716
rect 4096 626 4197 682
rect 4096 592 4130 626
rect 4164 592 4197 626
rect 4096 536 4197 592
rect 4096 502 4130 536
rect 4164 502 4197 536
rect 4096 446 4197 502
rect 4096 412 4130 446
rect 4164 412 4197 446
rect 4096 356 4197 412
rect 4096 322 4130 356
rect 4164 322 4197 356
rect 4096 266 4197 322
rect 4096 232 4130 266
rect 4164 232 4197 266
rect 4096 176 4197 232
rect 5283 1132 5317 1166
rect 5351 1132 5384 1166
rect 5283 1076 5384 1132
rect 5283 1042 5317 1076
rect 5351 1042 5384 1076
rect 5283 986 5384 1042
rect 5283 952 5317 986
rect 5351 952 5384 986
rect 5283 896 5384 952
rect 5283 862 5317 896
rect 5351 862 5384 896
rect 5283 806 5384 862
rect 5283 772 5317 806
rect 5351 772 5384 806
rect 5283 716 5384 772
rect 5283 682 5317 716
rect 5351 682 5384 716
rect 5283 626 5384 682
rect 5283 592 5317 626
rect 5351 592 5384 626
rect 5283 536 5384 592
rect 5283 502 5317 536
rect 5351 502 5384 536
rect 5283 446 5384 502
rect 5283 412 5317 446
rect 5351 412 5384 446
rect 5283 356 5384 412
rect 5283 322 5317 356
rect 5351 322 5384 356
rect 5283 266 5384 322
rect 5283 232 5317 266
rect 5351 232 5384 266
rect 4096 142 4130 176
rect 4164 142 4197 176
rect 4096 127 4197 142
rect 5283 176 5384 232
rect 5283 142 5317 176
rect 5351 142 5384 176
rect 5283 127 5384 142
rect 4096 92 5384 127
rect 4096 58 4226 92
rect 4260 58 4316 92
rect 4350 58 4406 92
rect 4440 58 4496 92
rect 4530 58 4586 92
rect 4620 58 4676 92
rect 4710 58 4766 92
rect 4800 58 4856 92
rect 4890 58 4946 92
rect 4980 58 5036 92
rect 5070 58 5126 92
rect 5160 58 5216 92
rect 5250 58 5384 92
rect 4096 26 5384 58
rect 5456 1279 6744 1314
rect 5456 1256 5586 1279
rect 5456 1222 5490 1256
rect 5524 1245 5586 1256
rect 5620 1245 5676 1279
rect 5710 1245 5766 1279
rect 5800 1245 5856 1279
rect 5890 1245 5946 1279
rect 5980 1245 6036 1279
rect 6070 1245 6126 1279
rect 6160 1245 6216 1279
rect 6250 1245 6306 1279
rect 6340 1245 6396 1279
rect 6430 1245 6486 1279
rect 6520 1245 6576 1279
rect 6610 1256 6744 1279
rect 6610 1245 6677 1256
rect 5524 1222 6677 1245
rect 6711 1222 6744 1256
rect 5456 1213 6744 1222
rect 5456 1166 5557 1213
rect 5456 1132 5490 1166
rect 5524 1132 5557 1166
rect 6643 1166 6744 1213
rect 5456 1076 5557 1132
rect 5456 1042 5490 1076
rect 5524 1042 5557 1076
rect 5456 986 5557 1042
rect 5456 952 5490 986
rect 5524 952 5557 986
rect 5456 896 5557 952
rect 5456 862 5490 896
rect 5524 862 5557 896
rect 5456 806 5557 862
rect 5456 772 5490 806
rect 5524 772 5557 806
rect 5456 716 5557 772
rect 5456 682 5490 716
rect 5524 682 5557 716
rect 5456 626 5557 682
rect 5456 592 5490 626
rect 5524 592 5557 626
rect 5456 536 5557 592
rect 5456 502 5490 536
rect 5524 502 5557 536
rect 5456 446 5557 502
rect 5456 412 5490 446
rect 5524 412 5557 446
rect 5456 356 5557 412
rect 5456 322 5490 356
rect 5524 322 5557 356
rect 5456 266 5557 322
rect 5456 232 5490 266
rect 5524 232 5557 266
rect 5456 176 5557 232
rect 6643 1132 6677 1166
rect 6711 1132 6744 1166
rect 6643 1076 6744 1132
rect 6643 1042 6677 1076
rect 6711 1042 6744 1076
rect 6643 986 6744 1042
rect 6643 952 6677 986
rect 6711 952 6744 986
rect 6643 896 6744 952
rect 6643 862 6677 896
rect 6711 862 6744 896
rect 6643 806 6744 862
rect 6643 772 6677 806
rect 6711 772 6744 806
rect 6643 716 6744 772
rect 6643 682 6677 716
rect 6711 682 6744 716
rect 6643 626 6744 682
rect 6643 592 6677 626
rect 6711 592 6744 626
rect 6643 536 6744 592
rect 6643 502 6677 536
rect 6711 502 6744 536
rect 6643 446 6744 502
rect 6643 412 6677 446
rect 6711 412 6744 446
rect 6643 356 6744 412
rect 6643 322 6677 356
rect 6711 322 6744 356
rect 6643 266 6744 322
rect 6643 232 6677 266
rect 6711 232 6744 266
rect 5456 142 5490 176
rect 5524 142 5557 176
rect 5456 127 5557 142
rect 6643 176 6744 232
rect 6643 142 6677 176
rect 6711 142 6744 176
rect 6643 127 6744 142
rect 5456 92 6744 127
rect 5456 58 5586 92
rect 5620 58 5676 92
rect 5710 58 5766 92
rect 5800 58 5856 92
rect 5890 58 5946 92
rect 5980 58 6036 92
rect 6070 58 6126 92
rect 6160 58 6216 92
rect 6250 58 6306 92
rect 6340 58 6396 92
rect 6430 58 6486 92
rect 6520 58 6576 92
rect 6610 58 6744 92
rect 5456 26 6744 58
rect 6816 1279 8104 1314
rect 6816 1256 6946 1279
rect 6816 1222 6850 1256
rect 6884 1245 6946 1256
rect 6980 1245 7036 1279
rect 7070 1245 7126 1279
rect 7160 1245 7216 1279
rect 7250 1245 7306 1279
rect 7340 1245 7396 1279
rect 7430 1245 7486 1279
rect 7520 1245 7576 1279
rect 7610 1245 7666 1279
rect 7700 1245 7756 1279
rect 7790 1245 7846 1279
rect 7880 1245 7936 1279
rect 7970 1256 8104 1279
rect 7970 1245 8037 1256
rect 6884 1222 8037 1245
rect 8071 1222 8104 1256
rect 6816 1213 8104 1222
rect 6816 1166 6917 1213
rect 6816 1132 6850 1166
rect 6884 1132 6917 1166
rect 8003 1166 8104 1213
rect 6816 1076 6917 1132
rect 6816 1042 6850 1076
rect 6884 1042 6917 1076
rect 6816 986 6917 1042
rect 6816 952 6850 986
rect 6884 952 6917 986
rect 6816 896 6917 952
rect 6816 862 6850 896
rect 6884 862 6917 896
rect 6816 806 6917 862
rect 6816 772 6850 806
rect 6884 772 6917 806
rect 6816 716 6917 772
rect 6816 682 6850 716
rect 6884 682 6917 716
rect 6816 626 6917 682
rect 6816 592 6850 626
rect 6884 592 6917 626
rect 6816 536 6917 592
rect 6816 502 6850 536
rect 6884 502 6917 536
rect 6816 446 6917 502
rect 6816 412 6850 446
rect 6884 412 6917 446
rect 6816 356 6917 412
rect 6816 322 6850 356
rect 6884 322 6917 356
rect 6816 266 6917 322
rect 6816 232 6850 266
rect 6884 232 6917 266
rect 6816 176 6917 232
rect 8003 1132 8037 1166
rect 8071 1132 8104 1166
rect 8003 1076 8104 1132
rect 8003 1042 8037 1076
rect 8071 1042 8104 1076
rect 8003 986 8104 1042
rect 8003 952 8037 986
rect 8071 952 8104 986
rect 8003 896 8104 952
rect 8003 862 8037 896
rect 8071 862 8104 896
rect 8003 806 8104 862
rect 8003 772 8037 806
rect 8071 772 8104 806
rect 8003 716 8104 772
rect 8003 682 8037 716
rect 8071 682 8104 716
rect 8003 626 8104 682
rect 8003 592 8037 626
rect 8071 592 8104 626
rect 8003 536 8104 592
rect 8003 502 8037 536
rect 8071 502 8104 536
rect 8003 446 8104 502
rect 8003 412 8037 446
rect 8071 412 8104 446
rect 8003 356 8104 412
rect 8003 322 8037 356
rect 8071 322 8104 356
rect 8003 266 8104 322
rect 8003 232 8037 266
rect 8071 232 8104 266
rect 6816 142 6850 176
rect 6884 142 6917 176
rect 6816 127 6917 142
rect 8003 176 8104 232
rect 8003 142 8037 176
rect 8071 142 8104 176
rect 8003 127 8104 142
rect 6816 92 8104 127
rect 6816 58 6946 92
rect 6980 58 7036 92
rect 7070 58 7126 92
rect 7160 58 7216 92
rect 7250 58 7306 92
rect 7340 58 7396 92
rect 7430 58 7486 92
rect 7520 58 7576 92
rect 7610 58 7666 92
rect 7700 58 7756 92
rect 7790 58 7846 92
rect 7880 58 7936 92
rect 7970 58 8104 92
rect 6816 26 8104 58
rect 8176 1279 9464 1314
rect 8176 1256 8306 1279
rect 8176 1222 8210 1256
rect 8244 1245 8306 1256
rect 8340 1245 8396 1279
rect 8430 1245 8486 1279
rect 8520 1245 8576 1279
rect 8610 1245 8666 1279
rect 8700 1245 8756 1279
rect 8790 1245 8846 1279
rect 8880 1245 8936 1279
rect 8970 1245 9026 1279
rect 9060 1245 9116 1279
rect 9150 1245 9206 1279
rect 9240 1245 9296 1279
rect 9330 1256 9464 1279
rect 9330 1245 9397 1256
rect 8244 1222 9397 1245
rect 9431 1222 9464 1256
rect 8176 1213 9464 1222
rect 8176 1166 8277 1213
rect 8176 1132 8210 1166
rect 8244 1132 8277 1166
rect 9363 1166 9464 1213
rect 8176 1076 8277 1132
rect 8176 1042 8210 1076
rect 8244 1042 8277 1076
rect 8176 986 8277 1042
rect 8176 952 8210 986
rect 8244 952 8277 986
rect 8176 896 8277 952
rect 8176 862 8210 896
rect 8244 862 8277 896
rect 8176 806 8277 862
rect 8176 772 8210 806
rect 8244 772 8277 806
rect 8176 716 8277 772
rect 8176 682 8210 716
rect 8244 682 8277 716
rect 8176 626 8277 682
rect 8176 592 8210 626
rect 8244 592 8277 626
rect 8176 536 8277 592
rect 8176 502 8210 536
rect 8244 502 8277 536
rect 8176 446 8277 502
rect 8176 412 8210 446
rect 8244 412 8277 446
rect 8176 356 8277 412
rect 8176 322 8210 356
rect 8244 322 8277 356
rect 8176 266 8277 322
rect 8176 232 8210 266
rect 8244 232 8277 266
rect 8176 176 8277 232
rect 9363 1132 9397 1166
rect 9431 1132 9464 1166
rect 9363 1076 9464 1132
rect 9363 1042 9397 1076
rect 9431 1042 9464 1076
rect 9363 986 9464 1042
rect 9363 952 9397 986
rect 9431 952 9464 986
rect 9363 896 9464 952
rect 9363 862 9397 896
rect 9431 862 9464 896
rect 9363 806 9464 862
rect 9363 772 9397 806
rect 9431 772 9464 806
rect 9363 716 9464 772
rect 9363 682 9397 716
rect 9431 682 9464 716
rect 9363 626 9464 682
rect 9363 592 9397 626
rect 9431 592 9464 626
rect 9363 536 9464 592
rect 9363 502 9397 536
rect 9431 502 9464 536
rect 9363 446 9464 502
rect 9363 412 9397 446
rect 9431 412 9464 446
rect 9363 356 9464 412
rect 9363 322 9397 356
rect 9431 322 9464 356
rect 9363 266 9464 322
rect 9363 232 9397 266
rect 9431 232 9464 266
rect 8176 142 8210 176
rect 8244 142 8277 176
rect 8176 127 8277 142
rect 9363 176 9464 232
rect 9363 142 9397 176
rect 9431 142 9464 176
rect 9363 127 9464 142
rect 8176 92 9464 127
rect 8176 58 8306 92
rect 8340 58 8396 92
rect 8430 58 8486 92
rect 8520 58 8576 92
rect 8610 58 8666 92
rect 8700 58 8756 92
rect 8790 58 8846 92
rect 8880 58 8936 92
rect 8970 58 9026 92
rect 9060 58 9116 92
rect 9150 58 9206 92
rect 9240 58 9296 92
rect 9330 58 9464 92
rect 8176 26 9464 58
<< nsubdiff >>
rect 4540 5430 4620 5460
rect 4540 5390 4560 5430
rect 4600 5390 4620 5430
rect 4540 5330 4620 5390
rect 4540 5290 4560 5330
rect 4600 5290 4620 5330
rect 4540 5230 4620 5290
rect 4540 5190 4560 5230
rect 4600 5190 4620 5230
rect 4540 5130 4620 5190
rect 4540 5090 4560 5130
rect 4600 5090 4620 5130
rect 4540 5030 4620 5090
rect 4540 4990 4560 5030
rect 4600 4990 4620 5030
rect 4540 4930 4620 4990
rect 4540 4890 4560 4930
rect 4600 4890 4620 4930
rect 4540 4830 4620 4890
rect 4540 4790 4560 4830
rect 4600 4790 4620 4830
rect 4540 4730 4620 4790
rect 4540 4690 4560 4730
rect 4600 4690 4620 4730
rect 4540 4660 4620 4690
rect 8300 5430 8380 5460
rect 8300 5390 8320 5430
rect 8360 5390 8380 5430
rect 8300 5330 8380 5390
rect 8300 5290 8320 5330
rect 8360 5290 8380 5330
rect 8300 5230 8380 5290
rect 8300 5190 8320 5230
rect 8360 5190 8380 5230
rect 8300 5130 8380 5190
rect 8300 5090 8320 5130
rect 8360 5090 8380 5130
rect 8300 5030 8380 5090
rect 8300 4990 8320 5030
rect 8360 4990 8380 5030
rect 8300 4930 8380 4990
rect 8300 4890 8320 4930
rect 8360 4890 8380 4930
rect 8300 4830 8380 4890
rect 8300 4790 8320 4830
rect 8360 4790 8380 4830
rect 8300 4730 8380 4790
rect 8300 4690 8320 4730
rect 8360 4690 8380 4730
rect 8300 4660 8380 4690
rect 5140 4190 5220 4220
rect 5140 4150 5160 4190
rect 5200 4150 5220 4190
rect 5140 4090 5220 4150
rect 5140 4050 5160 4090
rect 5200 4050 5220 4090
rect 5140 3990 5220 4050
rect 5140 3950 5160 3990
rect 5200 3950 5220 3990
rect 5140 3890 5220 3950
rect 5140 3850 5160 3890
rect 5200 3850 5220 3890
rect 5140 3820 5220 3850
rect 7700 4190 7780 4220
rect 7700 4150 7720 4190
rect 7760 4150 7780 4190
rect 7700 4090 7780 4150
rect 7700 4050 7720 4090
rect 7760 4050 7780 4090
rect 7700 3990 7780 4050
rect 7700 3950 7720 3990
rect 7760 3950 7780 3990
rect 7700 3890 7780 3950
rect 7700 3850 7720 3890
rect 7760 3850 7780 3890
rect 7700 3820 7780 3850
rect 1539 1132 2501 1151
rect 1539 1098 1670 1132
rect 1704 1098 1760 1132
rect 1794 1098 1850 1132
rect 1884 1098 1940 1132
rect 1974 1098 2030 1132
rect 2064 1098 2120 1132
rect 2154 1098 2210 1132
rect 2244 1098 2300 1132
rect 2334 1098 2390 1132
rect 2424 1098 2501 1132
rect 1539 1079 2501 1098
rect 1539 1075 1611 1079
rect 1539 1041 1558 1075
rect 1592 1041 1611 1075
rect 1539 985 1611 1041
rect 2429 1056 2501 1079
rect 2429 1022 2448 1056
rect 2482 1022 2501 1056
rect 1539 951 1558 985
rect 1592 951 1611 985
rect 1539 895 1611 951
rect 1539 861 1558 895
rect 1592 861 1611 895
rect 1539 805 1611 861
rect 1539 771 1558 805
rect 1592 771 1611 805
rect 1539 715 1611 771
rect 1539 681 1558 715
rect 1592 681 1611 715
rect 1539 625 1611 681
rect 1539 591 1558 625
rect 1592 591 1611 625
rect 1539 535 1611 591
rect 1539 501 1558 535
rect 1592 501 1611 535
rect 1539 445 1611 501
rect 1539 411 1558 445
rect 1592 411 1611 445
rect 1539 355 1611 411
rect 1539 321 1558 355
rect 1592 321 1611 355
rect 2429 966 2501 1022
rect 2429 932 2448 966
rect 2482 932 2501 966
rect 2429 876 2501 932
rect 2429 842 2448 876
rect 2482 842 2501 876
rect 2429 786 2501 842
rect 2429 752 2448 786
rect 2482 752 2501 786
rect 2429 696 2501 752
rect 2429 662 2448 696
rect 2482 662 2501 696
rect 2429 606 2501 662
rect 2429 572 2448 606
rect 2482 572 2501 606
rect 2429 516 2501 572
rect 2429 482 2448 516
rect 2482 482 2501 516
rect 2429 426 2501 482
rect 2429 392 2448 426
rect 2482 392 2501 426
rect 2429 336 2501 392
rect 1539 261 1611 321
rect 2429 302 2448 336
rect 2482 302 2501 336
rect 2429 261 2501 302
rect 1539 242 2501 261
rect 1539 208 1636 242
rect 1670 208 1726 242
rect 1760 208 1816 242
rect 1850 208 1906 242
rect 1940 208 1996 242
rect 2030 208 2086 242
rect 2120 208 2176 242
rect 2210 208 2266 242
rect 2300 208 2356 242
rect 2390 208 2501 242
rect 1539 189 2501 208
rect 2899 1132 3861 1151
rect 2899 1098 3030 1132
rect 3064 1098 3120 1132
rect 3154 1098 3210 1132
rect 3244 1098 3300 1132
rect 3334 1098 3390 1132
rect 3424 1098 3480 1132
rect 3514 1098 3570 1132
rect 3604 1098 3660 1132
rect 3694 1098 3750 1132
rect 3784 1098 3861 1132
rect 2899 1079 3861 1098
rect 2899 1075 2971 1079
rect 2899 1041 2918 1075
rect 2952 1041 2971 1075
rect 2899 985 2971 1041
rect 3789 1056 3861 1079
rect 3789 1022 3808 1056
rect 3842 1022 3861 1056
rect 2899 951 2918 985
rect 2952 951 2971 985
rect 2899 895 2971 951
rect 2899 861 2918 895
rect 2952 861 2971 895
rect 2899 805 2971 861
rect 2899 771 2918 805
rect 2952 771 2971 805
rect 2899 715 2971 771
rect 2899 681 2918 715
rect 2952 681 2971 715
rect 2899 625 2971 681
rect 2899 591 2918 625
rect 2952 591 2971 625
rect 2899 535 2971 591
rect 2899 501 2918 535
rect 2952 501 2971 535
rect 2899 445 2971 501
rect 2899 411 2918 445
rect 2952 411 2971 445
rect 2899 355 2971 411
rect 2899 321 2918 355
rect 2952 321 2971 355
rect 3789 966 3861 1022
rect 3789 932 3808 966
rect 3842 932 3861 966
rect 3789 876 3861 932
rect 3789 842 3808 876
rect 3842 842 3861 876
rect 3789 786 3861 842
rect 3789 752 3808 786
rect 3842 752 3861 786
rect 3789 696 3861 752
rect 3789 662 3808 696
rect 3842 662 3861 696
rect 3789 606 3861 662
rect 3789 572 3808 606
rect 3842 572 3861 606
rect 3789 516 3861 572
rect 3789 482 3808 516
rect 3842 482 3861 516
rect 3789 426 3861 482
rect 3789 392 3808 426
rect 3842 392 3861 426
rect 3789 336 3861 392
rect 2899 261 2971 321
rect 3789 302 3808 336
rect 3842 302 3861 336
rect 3789 261 3861 302
rect 2899 242 3861 261
rect 2899 208 2996 242
rect 3030 208 3086 242
rect 3120 208 3176 242
rect 3210 208 3266 242
rect 3300 208 3356 242
rect 3390 208 3446 242
rect 3480 208 3536 242
rect 3570 208 3626 242
rect 3660 208 3716 242
rect 3750 208 3861 242
rect 2899 189 3861 208
rect 4259 1132 5221 1151
rect 4259 1098 4390 1132
rect 4424 1098 4480 1132
rect 4514 1098 4570 1132
rect 4604 1098 4660 1132
rect 4694 1098 4750 1132
rect 4784 1098 4840 1132
rect 4874 1098 4930 1132
rect 4964 1098 5020 1132
rect 5054 1098 5110 1132
rect 5144 1098 5221 1132
rect 4259 1079 5221 1098
rect 4259 1075 4331 1079
rect 4259 1041 4278 1075
rect 4312 1041 4331 1075
rect 4259 985 4331 1041
rect 5149 1056 5221 1079
rect 5149 1022 5168 1056
rect 5202 1022 5221 1056
rect 4259 951 4278 985
rect 4312 951 4331 985
rect 4259 895 4331 951
rect 4259 861 4278 895
rect 4312 861 4331 895
rect 4259 805 4331 861
rect 4259 771 4278 805
rect 4312 771 4331 805
rect 4259 715 4331 771
rect 4259 681 4278 715
rect 4312 681 4331 715
rect 4259 625 4331 681
rect 4259 591 4278 625
rect 4312 591 4331 625
rect 4259 535 4331 591
rect 4259 501 4278 535
rect 4312 501 4331 535
rect 4259 445 4331 501
rect 4259 411 4278 445
rect 4312 411 4331 445
rect 4259 355 4331 411
rect 4259 321 4278 355
rect 4312 321 4331 355
rect 5149 966 5221 1022
rect 5149 932 5168 966
rect 5202 932 5221 966
rect 5149 876 5221 932
rect 5149 842 5168 876
rect 5202 842 5221 876
rect 5149 786 5221 842
rect 5149 752 5168 786
rect 5202 752 5221 786
rect 5149 696 5221 752
rect 5149 662 5168 696
rect 5202 662 5221 696
rect 5149 606 5221 662
rect 5149 572 5168 606
rect 5202 572 5221 606
rect 5149 516 5221 572
rect 5149 482 5168 516
rect 5202 482 5221 516
rect 5149 426 5221 482
rect 5149 392 5168 426
rect 5202 392 5221 426
rect 5149 336 5221 392
rect 4259 261 4331 321
rect 5149 302 5168 336
rect 5202 302 5221 336
rect 5149 261 5221 302
rect 4259 242 5221 261
rect 4259 208 4356 242
rect 4390 208 4446 242
rect 4480 208 4536 242
rect 4570 208 4626 242
rect 4660 208 4716 242
rect 4750 208 4806 242
rect 4840 208 4896 242
rect 4930 208 4986 242
rect 5020 208 5076 242
rect 5110 208 5221 242
rect 4259 189 5221 208
rect 5619 1132 6581 1151
rect 5619 1098 5750 1132
rect 5784 1098 5840 1132
rect 5874 1098 5930 1132
rect 5964 1098 6020 1132
rect 6054 1098 6110 1132
rect 6144 1098 6200 1132
rect 6234 1098 6290 1132
rect 6324 1098 6380 1132
rect 6414 1098 6470 1132
rect 6504 1098 6581 1132
rect 5619 1079 6581 1098
rect 5619 1075 5691 1079
rect 5619 1041 5638 1075
rect 5672 1041 5691 1075
rect 5619 985 5691 1041
rect 6509 1056 6581 1079
rect 6509 1022 6528 1056
rect 6562 1022 6581 1056
rect 5619 951 5638 985
rect 5672 951 5691 985
rect 5619 895 5691 951
rect 5619 861 5638 895
rect 5672 861 5691 895
rect 5619 805 5691 861
rect 5619 771 5638 805
rect 5672 771 5691 805
rect 5619 715 5691 771
rect 5619 681 5638 715
rect 5672 681 5691 715
rect 5619 625 5691 681
rect 5619 591 5638 625
rect 5672 591 5691 625
rect 5619 535 5691 591
rect 5619 501 5638 535
rect 5672 501 5691 535
rect 5619 445 5691 501
rect 5619 411 5638 445
rect 5672 411 5691 445
rect 5619 355 5691 411
rect 5619 321 5638 355
rect 5672 321 5691 355
rect 6509 966 6581 1022
rect 6509 932 6528 966
rect 6562 932 6581 966
rect 6509 876 6581 932
rect 6509 842 6528 876
rect 6562 842 6581 876
rect 6509 786 6581 842
rect 6509 752 6528 786
rect 6562 752 6581 786
rect 6509 696 6581 752
rect 6509 662 6528 696
rect 6562 662 6581 696
rect 6509 606 6581 662
rect 6509 572 6528 606
rect 6562 572 6581 606
rect 6509 516 6581 572
rect 6509 482 6528 516
rect 6562 482 6581 516
rect 6509 426 6581 482
rect 6509 392 6528 426
rect 6562 392 6581 426
rect 6509 336 6581 392
rect 5619 261 5691 321
rect 6509 302 6528 336
rect 6562 302 6581 336
rect 6509 261 6581 302
rect 5619 242 6581 261
rect 5619 208 5716 242
rect 5750 208 5806 242
rect 5840 208 5896 242
rect 5930 208 5986 242
rect 6020 208 6076 242
rect 6110 208 6166 242
rect 6200 208 6256 242
rect 6290 208 6346 242
rect 6380 208 6436 242
rect 6470 208 6581 242
rect 5619 189 6581 208
rect 6979 1132 7941 1151
rect 6979 1098 7110 1132
rect 7144 1098 7200 1132
rect 7234 1098 7290 1132
rect 7324 1098 7380 1132
rect 7414 1098 7470 1132
rect 7504 1098 7560 1132
rect 7594 1098 7650 1132
rect 7684 1098 7740 1132
rect 7774 1098 7830 1132
rect 7864 1098 7941 1132
rect 6979 1079 7941 1098
rect 6979 1075 7051 1079
rect 6979 1041 6998 1075
rect 7032 1041 7051 1075
rect 6979 985 7051 1041
rect 7869 1056 7941 1079
rect 7869 1022 7888 1056
rect 7922 1022 7941 1056
rect 6979 951 6998 985
rect 7032 951 7051 985
rect 6979 895 7051 951
rect 6979 861 6998 895
rect 7032 861 7051 895
rect 6979 805 7051 861
rect 6979 771 6998 805
rect 7032 771 7051 805
rect 6979 715 7051 771
rect 6979 681 6998 715
rect 7032 681 7051 715
rect 6979 625 7051 681
rect 6979 591 6998 625
rect 7032 591 7051 625
rect 6979 535 7051 591
rect 6979 501 6998 535
rect 7032 501 7051 535
rect 6979 445 7051 501
rect 6979 411 6998 445
rect 7032 411 7051 445
rect 6979 355 7051 411
rect 6979 321 6998 355
rect 7032 321 7051 355
rect 7869 966 7941 1022
rect 7869 932 7888 966
rect 7922 932 7941 966
rect 7869 876 7941 932
rect 7869 842 7888 876
rect 7922 842 7941 876
rect 7869 786 7941 842
rect 7869 752 7888 786
rect 7922 752 7941 786
rect 7869 696 7941 752
rect 7869 662 7888 696
rect 7922 662 7941 696
rect 7869 606 7941 662
rect 7869 572 7888 606
rect 7922 572 7941 606
rect 7869 516 7941 572
rect 7869 482 7888 516
rect 7922 482 7941 516
rect 7869 426 7941 482
rect 7869 392 7888 426
rect 7922 392 7941 426
rect 7869 336 7941 392
rect 6979 261 7051 321
rect 7869 302 7888 336
rect 7922 302 7941 336
rect 7869 261 7941 302
rect 6979 242 7941 261
rect 6979 208 7076 242
rect 7110 208 7166 242
rect 7200 208 7256 242
rect 7290 208 7346 242
rect 7380 208 7436 242
rect 7470 208 7526 242
rect 7560 208 7616 242
rect 7650 208 7706 242
rect 7740 208 7796 242
rect 7830 208 7941 242
rect 6979 189 7941 208
rect 8339 1132 9301 1151
rect 8339 1098 8470 1132
rect 8504 1098 8560 1132
rect 8594 1098 8650 1132
rect 8684 1098 8740 1132
rect 8774 1098 8830 1132
rect 8864 1098 8920 1132
rect 8954 1098 9010 1132
rect 9044 1098 9100 1132
rect 9134 1098 9190 1132
rect 9224 1098 9301 1132
rect 8339 1079 9301 1098
rect 8339 1075 8411 1079
rect 8339 1041 8358 1075
rect 8392 1041 8411 1075
rect 8339 985 8411 1041
rect 9229 1056 9301 1079
rect 9229 1022 9248 1056
rect 9282 1022 9301 1056
rect 8339 951 8358 985
rect 8392 951 8411 985
rect 8339 895 8411 951
rect 8339 861 8358 895
rect 8392 861 8411 895
rect 8339 805 8411 861
rect 8339 771 8358 805
rect 8392 771 8411 805
rect 8339 715 8411 771
rect 8339 681 8358 715
rect 8392 681 8411 715
rect 8339 625 8411 681
rect 8339 591 8358 625
rect 8392 591 8411 625
rect 8339 535 8411 591
rect 8339 501 8358 535
rect 8392 501 8411 535
rect 8339 445 8411 501
rect 8339 411 8358 445
rect 8392 411 8411 445
rect 8339 355 8411 411
rect 8339 321 8358 355
rect 8392 321 8411 355
rect 9229 966 9301 1022
rect 9229 932 9248 966
rect 9282 932 9301 966
rect 9229 876 9301 932
rect 9229 842 9248 876
rect 9282 842 9301 876
rect 9229 786 9301 842
rect 9229 752 9248 786
rect 9282 752 9301 786
rect 9229 696 9301 752
rect 9229 662 9248 696
rect 9282 662 9301 696
rect 9229 606 9301 662
rect 9229 572 9248 606
rect 9282 572 9301 606
rect 9229 516 9301 572
rect 9229 482 9248 516
rect 9282 482 9301 516
rect 9229 426 9301 482
rect 9229 392 9248 426
rect 9282 392 9301 426
rect 9229 336 9301 392
rect 8339 261 8411 321
rect 9229 302 9248 336
rect 9282 302 9301 336
rect 9229 261 9301 302
rect 8339 242 9301 261
rect 8339 208 8436 242
rect 8470 208 8526 242
rect 8560 208 8616 242
rect 8650 208 8706 242
rect 8740 208 8796 242
rect 8830 208 8886 242
rect 8920 208 8976 242
rect 9010 208 9066 242
rect 9100 208 9156 242
rect 9190 208 9301 242
rect 8339 189 9301 208
<< psubdiffcont >>
rect 6440 2700 6480 2740
rect 6440 2600 6480 2640
rect 6440 2500 6480 2540
rect 6440 2400 6480 2440
rect 6440 2300 6480 2340
rect 6440 2200 6480 2240
rect 6440 2100 6480 2140
rect 6440 2000 6480 2040
rect 1320 1600 1360 1640
rect 1320 1500 1360 1540
rect 7540 1640 7580 1680
rect 7540 1540 7580 1580
rect 1320 1400 1360 1440
rect 1410 1222 1444 1256
rect 1506 1245 1540 1279
rect 1596 1245 1630 1279
rect 1686 1245 1720 1279
rect 1776 1245 1810 1279
rect 1866 1245 1900 1279
rect 1956 1245 1990 1279
rect 2046 1245 2080 1279
rect 2136 1245 2170 1279
rect 2226 1245 2260 1279
rect 2316 1245 2350 1279
rect 2406 1245 2440 1279
rect 2496 1245 2530 1279
rect 2597 1222 2631 1256
rect 1410 1132 1444 1166
rect 1410 1042 1444 1076
rect 1410 952 1444 986
rect 1410 862 1444 896
rect 1410 772 1444 806
rect 1410 682 1444 716
rect 1410 592 1444 626
rect 1410 502 1444 536
rect 1410 412 1444 446
rect 1410 322 1444 356
rect 1410 232 1444 266
rect 2597 1132 2631 1166
rect 2597 1042 2631 1076
rect 2597 952 2631 986
rect 2597 862 2631 896
rect 2597 772 2631 806
rect 2597 682 2631 716
rect 2597 592 2631 626
rect 2597 502 2631 536
rect 2597 412 2631 446
rect 2597 322 2631 356
rect 2597 232 2631 266
rect 1410 142 1444 176
rect 2597 142 2631 176
rect 1506 58 1540 92
rect 1596 58 1630 92
rect 1686 58 1720 92
rect 1776 58 1810 92
rect 1866 58 1900 92
rect 1956 58 1990 92
rect 2046 58 2080 92
rect 2136 58 2170 92
rect 2226 58 2260 92
rect 2316 58 2350 92
rect 2406 58 2440 92
rect 2496 58 2530 92
rect 2770 1222 2804 1256
rect 2866 1245 2900 1279
rect 2956 1245 2990 1279
rect 3046 1245 3080 1279
rect 3136 1245 3170 1279
rect 3226 1245 3260 1279
rect 3316 1245 3350 1279
rect 3406 1245 3440 1279
rect 3496 1245 3530 1279
rect 3586 1245 3620 1279
rect 3676 1245 3710 1279
rect 3766 1245 3800 1279
rect 3856 1245 3890 1279
rect 3957 1222 3991 1256
rect 2770 1132 2804 1166
rect 2770 1042 2804 1076
rect 2770 952 2804 986
rect 2770 862 2804 896
rect 2770 772 2804 806
rect 2770 682 2804 716
rect 2770 592 2804 626
rect 2770 502 2804 536
rect 2770 412 2804 446
rect 2770 322 2804 356
rect 2770 232 2804 266
rect 3957 1132 3991 1166
rect 3957 1042 3991 1076
rect 3957 952 3991 986
rect 3957 862 3991 896
rect 3957 772 3991 806
rect 3957 682 3991 716
rect 3957 592 3991 626
rect 3957 502 3991 536
rect 3957 412 3991 446
rect 3957 322 3991 356
rect 3957 232 3991 266
rect 2770 142 2804 176
rect 3957 142 3991 176
rect 2866 58 2900 92
rect 2956 58 2990 92
rect 3046 58 3080 92
rect 3136 58 3170 92
rect 3226 58 3260 92
rect 3316 58 3350 92
rect 3406 58 3440 92
rect 3496 58 3530 92
rect 3586 58 3620 92
rect 3676 58 3710 92
rect 3766 58 3800 92
rect 3856 58 3890 92
rect 4130 1222 4164 1256
rect 4226 1245 4260 1279
rect 4316 1245 4350 1279
rect 4406 1245 4440 1279
rect 4496 1245 4530 1279
rect 4586 1245 4620 1279
rect 4676 1245 4710 1279
rect 4766 1245 4800 1279
rect 4856 1245 4890 1279
rect 4946 1245 4980 1279
rect 5036 1245 5070 1279
rect 5126 1245 5160 1279
rect 5216 1245 5250 1279
rect 5317 1222 5351 1256
rect 4130 1132 4164 1166
rect 4130 1042 4164 1076
rect 4130 952 4164 986
rect 4130 862 4164 896
rect 4130 772 4164 806
rect 4130 682 4164 716
rect 4130 592 4164 626
rect 4130 502 4164 536
rect 4130 412 4164 446
rect 4130 322 4164 356
rect 4130 232 4164 266
rect 5317 1132 5351 1166
rect 5317 1042 5351 1076
rect 5317 952 5351 986
rect 5317 862 5351 896
rect 5317 772 5351 806
rect 5317 682 5351 716
rect 5317 592 5351 626
rect 5317 502 5351 536
rect 5317 412 5351 446
rect 5317 322 5351 356
rect 5317 232 5351 266
rect 4130 142 4164 176
rect 5317 142 5351 176
rect 4226 58 4260 92
rect 4316 58 4350 92
rect 4406 58 4440 92
rect 4496 58 4530 92
rect 4586 58 4620 92
rect 4676 58 4710 92
rect 4766 58 4800 92
rect 4856 58 4890 92
rect 4946 58 4980 92
rect 5036 58 5070 92
rect 5126 58 5160 92
rect 5216 58 5250 92
rect 5490 1222 5524 1256
rect 5586 1245 5620 1279
rect 5676 1245 5710 1279
rect 5766 1245 5800 1279
rect 5856 1245 5890 1279
rect 5946 1245 5980 1279
rect 6036 1245 6070 1279
rect 6126 1245 6160 1279
rect 6216 1245 6250 1279
rect 6306 1245 6340 1279
rect 6396 1245 6430 1279
rect 6486 1245 6520 1279
rect 6576 1245 6610 1279
rect 6677 1222 6711 1256
rect 5490 1132 5524 1166
rect 5490 1042 5524 1076
rect 5490 952 5524 986
rect 5490 862 5524 896
rect 5490 772 5524 806
rect 5490 682 5524 716
rect 5490 592 5524 626
rect 5490 502 5524 536
rect 5490 412 5524 446
rect 5490 322 5524 356
rect 5490 232 5524 266
rect 6677 1132 6711 1166
rect 6677 1042 6711 1076
rect 6677 952 6711 986
rect 6677 862 6711 896
rect 6677 772 6711 806
rect 6677 682 6711 716
rect 6677 592 6711 626
rect 6677 502 6711 536
rect 6677 412 6711 446
rect 6677 322 6711 356
rect 6677 232 6711 266
rect 5490 142 5524 176
rect 6677 142 6711 176
rect 5586 58 5620 92
rect 5676 58 5710 92
rect 5766 58 5800 92
rect 5856 58 5890 92
rect 5946 58 5980 92
rect 6036 58 6070 92
rect 6126 58 6160 92
rect 6216 58 6250 92
rect 6306 58 6340 92
rect 6396 58 6430 92
rect 6486 58 6520 92
rect 6576 58 6610 92
rect 6850 1222 6884 1256
rect 6946 1245 6980 1279
rect 7036 1245 7070 1279
rect 7126 1245 7160 1279
rect 7216 1245 7250 1279
rect 7306 1245 7340 1279
rect 7396 1245 7430 1279
rect 7486 1245 7520 1279
rect 7576 1245 7610 1279
rect 7666 1245 7700 1279
rect 7756 1245 7790 1279
rect 7846 1245 7880 1279
rect 7936 1245 7970 1279
rect 8037 1222 8071 1256
rect 6850 1132 6884 1166
rect 6850 1042 6884 1076
rect 6850 952 6884 986
rect 6850 862 6884 896
rect 6850 772 6884 806
rect 6850 682 6884 716
rect 6850 592 6884 626
rect 6850 502 6884 536
rect 6850 412 6884 446
rect 6850 322 6884 356
rect 6850 232 6884 266
rect 8037 1132 8071 1166
rect 8037 1042 8071 1076
rect 8037 952 8071 986
rect 8037 862 8071 896
rect 8037 772 8071 806
rect 8037 682 8071 716
rect 8037 592 8071 626
rect 8037 502 8071 536
rect 8037 412 8071 446
rect 8037 322 8071 356
rect 8037 232 8071 266
rect 6850 142 6884 176
rect 8037 142 8071 176
rect 6946 58 6980 92
rect 7036 58 7070 92
rect 7126 58 7160 92
rect 7216 58 7250 92
rect 7306 58 7340 92
rect 7396 58 7430 92
rect 7486 58 7520 92
rect 7576 58 7610 92
rect 7666 58 7700 92
rect 7756 58 7790 92
rect 7846 58 7880 92
rect 7936 58 7970 92
rect 8210 1222 8244 1256
rect 8306 1245 8340 1279
rect 8396 1245 8430 1279
rect 8486 1245 8520 1279
rect 8576 1245 8610 1279
rect 8666 1245 8700 1279
rect 8756 1245 8790 1279
rect 8846 1245 8880 1279
rect 8936 1245 8970 1279
rect 9026 1245 9060 1279
rect 9116 1245 9150 1279
rect 9206 1245 9240 1279
rect 9296 1245 9330 1279
rect 9397 1222 9431 1256
rect 8210 1132 8244 1166
rect 8210 1042 8244 1076
rect 8210 952 8244 986
rect 8210 862 8244 896
rect 8210 772 8244 806
rect 8210 682 8244 716
rect 8210 592 8244 626
rect 8210 502 8244 536
rect 8210 412 8244 446
rect 8210 322 8244 356
rect 8210 232 8244 266
rect 9397 1132 9431 1166
rect 9397 1042 9431 1076
rect 9397 952 9431 986
rect 9397 862 9431 896
rect 9397 772 9431 806
rect 9397 682 9431 716
rect 9397 592 9431 626
rect 9397 502 9431 536
rect 9397 412 9431 446
rect 9397 322 9431 356
rect 9397 232 9431 266
rect 8210 142 8244 176
rect 9397 142 9431 176
rect 8306 58 8340 92
rect 8396 58 8430 92
rect 8486 58 8520 92
rect 8576 58 8610 92
rect 8666 58 8700 92
rect 8756 58 8790 92
rect 8846 58 8880 92
rect 8936 58 8970 92
rect 9026 58 9060 92
rect 9116 58 9150 92
rect 9206 58 9240 92
rect 9296 58 9330 92
<< nsubdiffcont >>
rect 4560 5390 4600 5430
rect 4560 5290 4600 5330
rect 4560 5190 4600 5230
rect 4560 5090 4600 5130
rect 4560 4990 4600 5030
rect 4560 4890 4600 4930
rect 4560 4790 4600 4830
rect 4560 4690 4600 4730
rect 8320 5390 8360 5430
rect 8320 5290 8360 5330
rect 8320 5190 8360 5230
rect 8320 5090 8360 5130
rect 8320 4990 8360 5030
rect 8320 4890 8360 4930
rect 8320 4790 8360 4830
rect 8320 4690 8360 4730
rect 5160 4150 5200 4190
rect 5160 4050 5200 4090
rect 5160 3950 5200 3990
rect 5160 3850 5200 3890
rect 7720 4150 7760 4190
rect 7720 4050 7760 4090
rect 7720 3950 7760 3990
rect 7720 3850 7760 3890
rect 1670 1098 1704 1132
rect 1760 1098 1794 1132
rect 1850 1098 1884 1132
rect 1940 1098 1974 1132
rect 2030 1098 2064 1132
rect 2120 1098 2154 1132
rect 2210 1098 2244 1132
rect 2300 1098 2334 1132
rect 2390 1098 2424 1132
rect 1558 1041 1592 1075
rect 2448 1022 2482 1056
rect 1558 951 1592 985
rect 1558 861 1592 895
rect 1558 771 1592 805
rect 1558 681 1592 715
rect 1558 591 1592 625
rect 1558 501 1592 535
rect 1558 411 1592 445
rect 1558 321 1592 355
rect 2448 932 2482 966
rect 2448 842 2482 876
rect 2448 752 2482 786
rect 2448 662 2482 696
rect 2448 572 2482 606
rect 2448 482 2482 516
rect 2448 392 2482 426
rect 2448 302 2482 336
rect 1636 208 1670 242
rect 1726 208 1760 242
rect 1816 208 1850 242
rect 1906 208 1940 242
rect 1996 208 2030 242
rect 2086 208 2120 242
rect 2176 208 2210 242
rect 2266 208 2300 242
rect 2356 208 2390 242
rect 3030 1098 3064 1132
rect 3120 1098 3154 1132
rect 3210 1098 3244 1132
rect 3300 1098 3334 1132
rect 3390 1098 3424 1132
rect 3480 1098 3514 1132
rect 3570 1098 3604 1132
rect 3660 1098 3694 1132
rect 3750 1098 3784 1132
rect 2918 1041 2952 1075
rect 3808 1022 3842 1056
rect 2918 951 2952 985
rect 2918 861 2952 895
rect 2918 771 2952 805
rect 2918 681 2952 715
rect 2918 591 2952 625
rect 2918 501 2952 535
rect 2918 411 2952 445
rect 2918 321 2952 355
rect 3808 932 3842 966
rect 3808 842 3842 876
rect 3808 752 3842 786
rect 3808 662 3842 696
rect 3808 572 3842 606
rect 3808 482 3842 516
rect 3808 392 3842 426
rect 3808 302 3842 336
rect 2996 208 3030 242
rect 3086 208 3120 242
rect 3176 208 3210 242
rect 3266 208 3300 242
rect 3356 208 3390 242
rect 3446 208 3480 242
rect 3536 208 3570 242
rect 3626 208 3660 242
rect 3716 208 3750 242
rect 4390 1098 4424 1132
rect 4480 1098 4514 1132
rect 4570 1098 4604 1132
rect 4660 1098 4694 1132
rect 4750 1098 4784 1132
rect 4840 1098 4874 1132
rect 4930 1098 4964 1132
rect 5020 1098 5054 1132
rect 5110 1098 5144 1132
rect 4278 1041 4312 1075
rect 5168 1022 5202 1056
rect 4278 951 4312 985
rect 4278 861 4312 895
rect 4278 771 4312 805
rect 4278 681 4312 715
rect 4278 591 4312 625
rect 4278 501 4312 535
rect 4278 411 4312 445
rect 4278 321 4312 355
rect 5168 932 5202 966
rect 5168 842 5202 876
rect 5168 752 5202 786
rect 5168 662 5202 696
rect 5168 572 5202 606
rect 5168 482 5202 516
rect 5168 392 5202 426
rect 5168 302 5202 336
rect 4356 208 4390 242
rect 4446 208 4480 242
rect 4536 208 4570 242
rect 4626 208 4660 242
rect 4716 208 4750 242
rect 4806 208 4840 242
rect 4896 208 4930 242
rect 4986 208 5020 242
rect 5076 208 5110 242
rect 5750 1098 5784 1132
rect 5840 1098 5874 1132
rect 5930 1098 5964 1132
rect 6020 1098 6054 1132
rect 6110 1098 6144 1132
rect 6200 1098 6234 1132
rect 6290 1098 6324 1132
rect 6380 1098 6414 1132
rect 6470 1098 6504 1132
rect 5638 1041 5672 1075
rect 6528 1022 6562 1056
rect 5638 951 5672 985
rect 5638 861 5672 895
rect 5638 771 5672 805
rect 5638 681 5672 715
rect 5638 591 5672 625
rect 5638 501 5672 535
rect 5638 411 5672 445
rect 5638 321 5672 355
rect 6528 932 6562 966
rect 6528 842 6562 876
rect 6528 752 6562 786
rect 6528 662 6562 696
rect 6528 572 6562 606
rect 6528 482 6562 516
rect 6528 392 6562 426
rect 6528 302 6562 336
rect 5716 208 5750 242
rect 5806 208 5840 242
rect 5896 208 5930 242
rect 5986 208 6020 242
rect 6076 208 6110 242
rect 6166 208 6200 242
rect 6256 208 6290 242
rect 6346 208 6380 242
rect 6436 208 6470 242
rect 7110 1098 7144 1132
rect 7200 1098 7234 1132
rect 7290 1098 7324 1132
rect 7380 1098 7414 1132
rect 7470 1098 7504 1132
rect 7560 1098 7594 1132
rect 7650 1098 7684 1132
rect 7740 1098 7774 1132
rect 7830 1098 7864 1132
rect 6998 1041 7032 1075
rect 7888 1022 7922 1056
rect 6998 951 7032 985
rect 6998 861 7032 895
rect 6998 771 7032 805
rect 6998 681 7032 715
rect 6998 591 7032 625
rect 6998 501 7032 535
rect 6998 411 7032 445
rect 6998 321 7032 355
rect 7888 932 7922 966
rect 7888 842 7922 876
rect 7888 752 7922 786
rect 7888 662 7922 696
rect 7888 572 7922 606
rect 7888 482 7922 516
rect 7888 392 7922 426
rect 7888 302 7922 336
rect 7076 208 7110 242
rect 7166 208 7200 242
rect 7256 208 7290 242
rect 7346 208 7380 242
rect 7436 208 7470 242
rect 7526 208 7560 242
rect 7616 208 7650 242
rect 7706 208 7740 242
rect 7796 208 7830 242
rect 8470 1098 8504 1132
rect 8560 1098 8594 1132
rect 8650 1098 8684 1132
rect 8740 1098 8774 1132
rect 8830 1098 8864 1132
rect 8920 1098 8954 1132
rect 9010 1098 9044 1132
rect 9100 1098 9134 1132
rect 9190 1098 9224 1132
rect 8358 1041 8392 1075
rect 9248 1022 9282 1056
rect 8358 951 8392 985
rect 8358 861 8392 895
rect 8358 771 8392 805
rect 8358 681 8392 715
rect 8358 591 8392 625
rect 8358 501 8392 535
rect 8358 411 8392 445
rect 8358 321 8392 355
rect 9248 932 9282 966
rect 9248 842 9282 876
rect 9248 752 9282 786
rect 9248 662 9282 696
rect 9248 572 9282 606
rect 9248 482 9282 516
rect 9248 392 9282 426
rect 9248 302 9282 336
rect 8436 208 8470 242
rect 8526 208 8560 242
rect 8616 208 8650 242
rect 8706 208 8740 242
rect 8796 208 8830 242
rect 8886 208 8920 242
rect 8976 208 9010 242
rect 9066 208 9100 242
rect 9156 208 9190 242
<< poly >>
rect 4700 5460 4820 5490
rect 4900 5460 5020 5490
rect 5100 5460 5220 5490
rect 5300 5460 5420 5490
rect 5500 5460 5620 5490
rect 5700 5460 5820 5490
rect 5900 5460 6020 5490
rect 6100 5460 6220 5490
rect 6300 5460 6420 5490
rect 6500 5460 6620 5490
rect 6700 5460 6820 5490
rect 6900 5460 7020 5490
rect 7100 5460 7220 5490
rect 7300 5460 7420 5490
rect 7500 5460 7620 5490
rect 7700 5460 7820 5490
rect 7900 5460 8020 5490
rect 8100 5460 8220 5490
rect 4700 4640 4820 4660
rect 4900 4640 5020 4660
rect 5100 4640 5220 4660
rect 5300 4640 5420 4660
rect 5500 4640 5620 4660
rect 5700 4640 5820 4660
rect 5900 4640 6020 4660
rect 6100 4640 6220 4660
rect 6300 4640 6420 4660
rect 6500 4640 6620 4660
rect 6700 4640 6820 4660
rect 6900 4640 7020 4660
rect 7100 4640 7220 4660
rect 7300 4640 7420 4660
rect 7500 4640 7620 4660
rect 7700 4640 7820 4660
rect 7900 4640 8020 4660
rect 8100 4640 8220 4660
rect 4700 4610 8220 4640
rect 6220 4570 6240 4610
rect 6280 4570 6300 4610
rect 6220 4550 6300 4570
rect 6620 4570 6640 4610
rect 6680 4570 6700 4610
rect 6620 4550 6700 4570
rect 8140 4570 8160 4610
rect 8200 4570 8220 4610
rect 8140 4550 8220 4570
rect 9030 4390 9110 4410
rect 9030 4350 9050 4390
rect 9090 4350 9110 4390
rect 9030 4330 9110 4350
rect 5300 4220 5420 4250
rect 5500 4220 5620 4250
rect 5700 4220 5820 4250
rect 5900 4220 6020 4250
rect 6100 4220 6220 4250
rect 6300 4220 6420 4250
rect 6500 4220 6620 4250
rect 6700 4220 6820 4250
rect 6900 4220 7020 4250
rect 7100 4220 7220 4250
rect 7300 4220 7420 4250
rect 7500 4220 7620 4250
rect 8830 4220 8860 4250
rect 9080 4220 9110 4330
rect 5300 3800 5420 3820
rect 5500 3800 5620 3820
rect 5700 3800 5820 3820
rect 5900 3800 6020 3820
rect 5300 3770 6020 3800
rect 6100 3800 6220 3820
rect 6300 3800 6420 3820
rect 6500 3800 6620 3820
rect 6700 3800 6820 3820
rect 6100 3770 6820 3800
rect 6900 3800 7020 3820
rect 7100 3800 7220 3820
rect 7300 3800 7420 3820
rect 7500 3800 7620 3820
rect 6900 3770 7620 3800
rect 5820 3730 5840 3770
rect 5880 3730 5900 3770
rect 5820 3710 5900 3730
rect 6350 3700 6390 3770
rect 7020 3730 7040 3770
rect 7080 3730 7100 3770
rect 7020 3710 7100 3730
rect 8830 3740 8860 3820
rect 9080 3790 9110 3820
rect 8970 3740 9050 3760
rect 8830 3700 8990 3740
rect 9030 3700 9050 3740
rect 6330 3680 6410 3700
rect 8970 3680 9050 3700
rect 6330 3640 6350 3680
rect 6390 3640 6410 3680
rect 6330 3620 6410 3640
rect 6100 3410 6180 3430
rect 6100 3370 6120 3410
rect 6160 3370 6180 3410
rect 6740 3410 6820 3430
rect 6740 3370 6760 3410
rect 6800 3370 6820 3410
rect 5700 3320 5820 3350
rect 5900 3320 6020 3350
rect 6100 3340 6820 3370
rect 6100 3320 6220 3340
rect 6300 3320 6420 3340
rect 6500 3320 6620 3340
rect 6700 3320 6820 3340
rect 6900 3320 7020 3350
rect 7100 3320 7220 3350
rect 5700 3100 5820 3120
rect 5900 3100 6020 3120
rect 5700 3070 6020 3100
rect 6100 3090 6220 3120
rect 6300 3090 6420 3120
rect 6500 3090 6620 3120
rect 6700 3090 6820 3120
rect 6900 3100 7020 3120
rect 7100 3100 7220 3120
rect 6900 3070 7220 3100
rect 5820 3030 5840 3070
rect 5880 3030 5900 3070
rect 5820 3010 5900 3030
rect 7020 3030 7040 3070
rect 7080 3030 7100 3070
rect 7020 3010 7100 3030
rect 5540 2860 6340 2880
rect 5540 2820 5560 2860
rect 5600 2820 5640 2860
rect 5680 2820 5720 2860
rect 5760 2820 5800 2860
rect 5840 2820 5880 2860
rect 5920 2820 5960 2860
rect 6000 2820 6040 2860
rect 6080 2820 6120 2860
rect 6160 2820 6200 2860
rect 6240 2820 6280 2860
rect 6320 2820 6340 2860
rect 5540 2770 6340 2820
rect 6580 2860 7380 2880
rect 6580 2820 6600 2860
rect 6640 2820 6680 2860
rect 6720 2820 6760 2860
rect 6800 2820 6840 2860
rect 6880 2820 6920 2860
rect 6960 2820 7000 2860
rect 7040 2820 7080 2860
rect 7120 2820 7160 2860
rect 7200 2820 7240 2860
rect 7280 2820 7320 2860
rect 7360 2820 7380 2860
rect 6580 2770 7380 2820
rect 5540 1940 6340 1970
rect 6580 1940 7380 1970
rect 5440 1800 5520 1820
rect 5440 1760 5460 1800
rect 5500 1760 5520 1800
rect 5440 1740 5520 1760
rect 5600 1800 5680 1820
rect 5600 1760 5620 1800
rect 5660 1760 5680 1800
rect 5600 1740 5680 1760
rect 5760 1800 5840 1820
rect 5760 1760 5780 1800
rect 5820 1760 5840 1800
rect 5760 1740 5840 1760
rect 5920 1800 6000 1820
rect 5920 1760 5940 1800
rect 5980 1760 6000 1800
rect 5920 1740 6000 1760
rect 6080 1800 6160 1820
rect 6080 1760 6100 1800
rect 6140 1760 6160 1800
rect 6080 1740 6160 1760
rect 6240 1800 6320 1820
rect 6240 1760 6260 1800
rect 6300 1760 6320 1800
rect 6240 1740 6320 1760
rect 6400 1800 6480 1820
rect 6400 1760 6420 1800
rect 6460 1760 6480 1800
rect 6400 1740 6480 1760
rect 6560 1800 6640 1820
rect 6560 1760 6580 1800
rect 6620 1760 6640 1800
rect 6560 1740 6640 1760
rect 6720 1800 6800 1820
rect 6720 1760 6740 1800
rect 6780 1760 6800 1800
rect 6720 1740 6800 1760
rect 6880 1800 6960 1820
rect 6880 1760 6900 1800
rect 6940 1760 6960 1800
rect 6880 1740 6960 1760
rect 7040 1800 7120 1820
rect 7040 1760 7060 1800
rect 7100 1760 7120 1800
rect 7040 1740 7120 1760
rect 7200 1800 7280 1820
rect 7200 1760 7220 1800
rect 7260 1760 7280 1800
rect 7200 1740 7280 1760
rect 7360 1800 7440 1820
rect 7360 1760 7380 1800
rect 7420 1760 7440 1800
rect 7360 1740 7440 1760
rect 5440 1710 7440 1740
rect 5440 1480 7440 1510
<< polycont >>
rect 6240 4570 6280 4610
rect 6640 4570 6680 4610
rect 8160 4570 8200 4610
rect 9050 4350 9090 4390
rect 5840 3730 5880 3770
rect 7040 3730 7080 3770
rect 8990 3700 9030 3740
rect 6350 3640 6390 3680
rect 6120 3370 6160 3410
rect 6760 3370 6800 3410
rect 5840 3030 5880 3070
rect 7040 3030 7080 3070
rect 5560 2820 5600 2860
rect 5640 2820 5680 2860
rect 5720 2820 5760 2860
rect 5800 2820 5840 2860
rect 5880 2820 5920 2860
rect 5960 2820 6000 2860
rect 6040 2820 6080 2860
rect 6120 2820 6160 2860
rect 6200 2820 6240 2860
rect 6280 2820 6320 2860
rect 6600 2820 6640 2860
rect 6680 2820 6720 2860
rect 6760 2820 6800 2860
rect 6840 2820 6880 2860
rect 6920 2820 6960 2860
rect 7000 2820 7040 2860
rect 7080 2820 7120 2860
rect 7160 2820 7200 2860
rect 7240 2820 7280 2860
rect 7320 2820 7360 2860
rect 5460 1760 5500 1800
rect 5620 1760 5660 1800
rect 5780 1760 5820 1800
rect 5940 1760 5980 1800
rect 6100 1760 6140 1800
rect 6260 1760 6300 1800
rect 6420 1760 6460 1800
rect 6580 1760 6620 1800
rect 6740 1760 6780 1800
rect 6900 1760 6940 1800
rect 7060 1760 7100 1800
rect 7220 1760 7260 1800
rect 7380 1760 7420 1800
<< xpolycontact >>
rect 2010 4980 2450 5050
rect 3790 4980 4230 5050
rect 2010 4860 2450 4930
rect 3790 4860 4230 4930
rect 2010 4740 2450 4810
rect 3790 4740 4230 4810
rect 2010 4620 2450 4690
rect 3790 4620 4230 4690
rect 2010 4500 2450 4570
rect 3790 4500 4230 4570
rect 2010 3960 2450 4030
rect 3790 3960 4230 4030
rect 2010 3840 2450 3910
rect 3790 3840 4230 3910
rect 2010 3720 2450 3790
rect 3790 3720 4230 3790
rect 2010 3600 2450 3670
rect 3790 3600 4230 3670
rect 2010 3480 2450 3550
rect 3790 3480 4230 3550
rect 2010 3010 2450 3080
rect 3150 3010 3590 3080
rect 2010 2890 2450 2960
rect 3790 2890 4230 2960
rect 2010 2770 2450 2840
rect 3790 2770 4230 2840
rect 2010 2650 2450 2720
rect 3790 2650 4230 2720
rect 2010 2530 2450 2600
rect 3790 2530 4230 2600
rect 2010 2410 2450 2480
rect 3790 2410 4230 2480
<< xpolyres >>
rect 2450 4980 3790 5050
rect 2450 4860 3790 4930
rect 2450 4740 3790 4810
rect 2450 4620 3790 4690
rect 2450 4500 3790 4570
rect 2450 3960 3790 4030
rect 2450 3840 3790 3910
rect 2450 3720 3790 3790
rect 2450 3600 3790 3670
rect 2450 3480 3790 3550
rect 2450 3010 3150 3080
rect 2450 2890 3790 2960
rect 2450 2770 3790 2840
rect 2450 2650 3790 2720
rect 2450 2530 3790 2600
rect 2450 2410 3790 2480
<< locali >>
rect 4620 5550 4700 5570
rect 4620 5510 4640 5550
rect 4680 5510 4700 5550
rect 4620 5490 4700 5510
rect 5020 5550 5100 5570
rect 5020 5510 5040 5550
rect 5080 5510 5100 5550
rect 5020 5490 5100 5510
rect 5420 5550 5500 5570
rect 5420 5510 5440 5550
rect 5480 5510 5500 5550
rect 5420 5490 5500 5510
rect 5820 5550 5900 5570
rect 5820 5510 5840 5550
rect 5880 5510 5900 5550
rect 5820 5490 5900 5510
rect 6220 5550 6300 5570
rect 6220 5510 6240 5550
rect 6280 5510 6300 5550
rect 6220 5490 6300 5510
rect 6420 5550 6500 5570
rect 6420 5510 6440 5550
rect 6480 5510 6500 5550
rect 6420 5490 6500 5510
rect 6620 5550 6700 5570
rect 6620 5510 6640 5550
rect 6680 5510 6700 5550
rect 6620 5490 6700 5510
rect 7020 5550 7100 5570
rect 7020 5510 7040 5550
rect 7080 5510 7100 5550
rect 7020 5490 7100 5510
rect 7420 5550 7500 5570
rect 7420 5510 7440 5550
rect 7480 5510 7500 5550
rect 7420 5490 7500 5510
rect 7820 5550 7900 5570
rect 7820 5510 7840 5550
rect 7880 5510 7900 5550
rect 7820 5490 7900 5510
rect 8220 5550 8300 5570
rect 8220 5510 8240 5550
rect 8280 5510 8300 5550
rect 8220 5490 8300 5510
rect 4640 5450 4680 5490
rect 5040 5450 5080 5490
rect 5440 5450 5480 5490
rect 5840 5450 5880 5490
rect 6240 5450 6280 5490
rect 4550 5430 4690 5450
rect 4550 5390 4560 5430
rect 4600 5390 4640 5430
rect 4680 5390 4690 5430
rect 4550 5330 4690 5390
rect 4550 5290 4560 5330
rect 4600 5290 4640 5330
rect 4680 5290 4690 5330
rect 4550 5230 4690 5290
rect 4550 5190 4560 5230
rect 4600 5190 4640 5230
rect 4680 5190 4690 5230
rect 4550 5130 4690 5190
rect 4550 5090 4560 5130
rect 4600 5090 4640 5130
rect 4680 5090 4690 5130
rect 1890 5030 2010 5050
rect 1890 4990 1910 5030
rect 1950 4990 2010 5030
rect 1890 4980 2010 4990
rect 1890 4970 1970 4980
rect 3790 4930 4230 4980
rect 4550 5030 4690 5090
rect 4550 4990 4560 5030
rect 4600 4990 4640 5030
rect 4680 4990 4690 5030
rect 4550 4930 4690 4990
rect 4550 4890 4560 4930
rect 4600 4890 4640 4930
rect 4680 4890 4690 4930
rect 2010 4810 2450 4860
rect 4550 4830 4690 4890
rect 3790 4690 4230 4740
rect 4550 4790 4560 4830
rect 4600 4790 4640 4830
rect 4680 4790 4690 4830
rect 4550 4730 4690 4790
rect 4550 4690 4560 4730
rect 4600 4690 4640 4730
rect 4680 4690 4690 4730
rect 4550 4670 4690 4690
rect 4830 5430 4890 5450
rect 4830 5390 4840 5430
rect 4880 5390 4890 5430
rect 4830 5330 4890 5390
rect 4830 5290 4840 5330
rect 4880 5290 4890 5330
rect 4830 5230 4890 5290
rect 4830 5190 4840 5230
rect 4880 5190 4890 5230
rect 4830 5130 4890 5190
rect 4830 5090 4840 5130
rect 4880 5090 4890 5130
rect 4830 5030 4890 5090
rect 4830 4990 4840 5030
rect 4880 4990 4890 5030
rect 4830 4930 4890 4990
rect 4830 4890 4840 4930
rect 4880 4890 4890 4930
rect 4830 4830 4890 4890
rect 4830 4790 4840 4830
rect 4880 4790 4890 4830
rect 4830 4730 4890 4790
rect 4830 4690 4840 4730
rect 4880 4690 4890 4730
rect 4830 4670 4890 4690
rect 5030 5430 5090 5450
rect 5030 5390 5040 5430
rect 5080 5390 5090 5430
rect 5030 5330 5090 5390
rect 5030 5290 5040 5330
rect 5080 5290 5090 5330
rect 5030 5230 5090 5290
rect 5030 5190 5040 5230
rect 5080 5190 5090 5230
rect 5030 5130 5090 5190
rect 5030 5090 5040 5130
rect 5080 5090 5090 5130
rect 5030 5030 5090 5090
rect 5030 4990 5040 5030
rect 5080 4990 5090 5030
rect 5030 4930 5090 4990
rect 5030 4890 5040 4930
rect 5080 4890 5090 4930
rect 5030 4830 5090 4890
rect 5030 4790 5040 4830
rect 5080 4790 5090 4830
rect 5030 4730 5090 4790
rect 5030 4690 5040 4730
rect 5080 4690 5090 4730
rect 5030 4670 5090 4690
rect 5230 5430 5290 5450
rect 5230 5390 5240 5430
rect 5280 5390 5290 5430
rect 5230 5330 5290 5390
rect 5230 5290 5240 5330
rect 5280 5290 5290 5330
rect 5230 5230 5290 5290
rect 5230 5190 5240 5230
rect 5280 5190 5290 5230
rect 5230 5130 5290 5190
rect 5230 5090 5240 5130
rect 5280 5090 5290 5130
rect 5230 5030 5290 5090
rect 5230 4990 5240 5030
rect 5280 4990 5290 5030
rect 5230 4930 5290 4990
rect 5230 4890 5240 4930
rect 5280 4890 5290 4930
rect 5230 4830 5290 4890
rect 5230 4790 5240 4830
rect 5280 4790 5290 4830
rect 5230 4730 5290 4790
rect 5230 4690 5240 4730
rect 5280 4690 5290 4730
rect 5230 4670 5290 4690
rect 5430 5430 5490 5450
rect 5430 5390 5440 5430
rect 5480 5390 5490 5430
rect 5430 5330 5490 5390
rect 5430 5290 5440 5330
rect 5480 5290 5490 5330
rect 5430 5230 5490 5290
rect 5430 5190 5440 5230
rect 5480 5190 5490 5230
rect 5430 5130 5490 5190
rect 5430 5090 5440 5130
rect 5480 5090 5490 5130
rect 5430 5030 5490 5090
rect 5430 4990 5440 5030
rect 5480 4990 5490 5030
rect 5430 4930 5490 4990
rect 5430 4890 5440 4930
rect 5480 4890 5490 4930
rect 5430 4830 5490 4890
rect 5430 4790 5440 4830
rect 5480 4790 5490 4830
rect 5430 4730 5490 4790
rect 5430 4690 5440 4730
rect 5480 4690 5490 4730
rect 5430 4670 5490 4690
rect 5630 5430 5690 5450
rect 5630 5390 5640 5430
rect 5680 5390 5690 5430
rect 5630 5330 5690 5390
rect 5630 5290 5640 5330
rect 5680 5290 5690 5330
rect 5630 5230 5690 5290
rect 5630 5190 5640 5230
rect 5680 5190 5690 5230
rect 5630 5130 5690 5190
rect 5630 5090 5640 5130
rect 5680 5090 5690 5130
rect 5630 5030 5690 5090
rect 5630 4990 5640 5030
rect 5680 4990 5690 5030
rect 5630 4930 5690 4990
rect 5630 4890 5640 4930
rect 5680 4890 5690 4930
rect 5630 4830 5690 4890
rect 5630 4790 5640 4830
rect 5680 4790 5690 4830
rect 5630 4730 5690 4790
rect 5630 4690 5640 4730
rect 5680 4690 5690 4730
rect 5630 4670 5690 4690
rect 5830 5430 5890 5450
rect 5830 5390 5840 5430
rect 5880 5390 5890 5430
rect 5830 5330 5890 5390
rect 5830 5290 5840 5330
rect 5880 5290 5890 5330
rect 5830 5230 5890 5290
rect 5830 5190 5840 5230
rect 5880 5190 5890 5230
rect 5830 5130 5890 5190
rect 5830 5090 5840 5130
rect 5880 5090 5890 5130
rect 5830 5030 5890 5090
rect 5830 4990 5840 5030
rect 5880 4990 5890 5030
rect 5830 4930 5890 4990
rect 5830 4890 5840 4930
rect 5880 4890 5890 4930
rect 5830 4830 5890 4890
rect 5830 4790 5840 4830
rect 5880 4790 5890 4830
rect 5830 4730 5890 4790
rect 5830 4690 5840 4730
rect 5880 4690 5890 4730
rect 5830 4670 5890 4690
rect 6030 5430 6090 5450
rect 6030 5390 6040 5430
rect 6080 5390 6090 5430
rect 6030 5330 6090 5390
rect 6030 5290 6040 5330
rect 6080 5290 6090 5330
rect 6030 5230 6090 5290
rect 6030 5190 6040 5230
rect 6080 5190 6090 5230
rect 6030 5130 6090 5190
rect 6030 5090 6040 5130
rect 6080 5090 6090 5130
rect 6030 5030 6090 5090
rect 6030 4990 6040 5030
rect 6080 4990 6090 5030
rect 6030 4930 6090 4990
rect 6030 4890 6040 4930
rect 6080 4890 6090 4930
rect 6030 4830 6090 4890
rect 6030 4790 6040 4830
rect 6080 4790 6090 4830
rect 6030 4730 6090 4790
rect 6030 4690 6040 4730
rect 6080 4690 6090 4730
rect 6030 4670 6090 4690
rect 6230 5430 6290 5450
rect 6230 5390 6240 5430
rect 6280 5390 6290 5430
rect 6230 5330 6290 5390
rect 6230 5290 6240 5330
rect 6280 5290 6290 5330
rect 6230 5230 6290 5290
rect 6230 5190 6240 5230
rect 6280 5190 6290 5230
rect 6230 5130 6290 5190
rect 6230 5090 6240 5130
rect 6280 5090 6290 5130
rect 6230 5030 6290 5090
rect 6230 4990 6240 5030
rect 6280 4990 6290 5030
rect 6230 4930 6290 4990
rect 6230 4890 6240 4930
rect 6280 4890 6290 4930
rect 6230 4830 6290 4890
rect 6230 4790 6240 4830
rect 6280 4790 6290 4830
rect 6230 4730 6290 4790
rect 6230 4690 6240 4730
rect 6280 4690 6290 4730
rect 6230 4670 6290 4690
rect 6430 5430 6490 5490
rect 6640 5450 6680 5490
rect 7040 5450 7080 5490
rect 7440 5450 7480 5490
rect 7840 5450 7880 5490
rect 8240 5450 8280 5490
rect 6430 5390 6440 5430
rect 6480 5390 6490 5430
rect 6430 5330 6490 5390
rect 6430 5290 6440 5330
rect 6480 5290 6490 5330
rect 6430 5230 6490 5290
rect 6430 5190 6440 5230
rect 6480 5190 6490 5230
rect 6430 5130 6490 5190
rect 6430 5090 6440 5130
rect 6480 5090 6490 5130
rect 6430 5030 6490 5090
rect 6430 4990 6440 5030
rect 6480 4990 6490 5030
rect 6430 4930 6490 4990
rect 6430 4890 6440 4930
rect 6480 4890 6490 4930
rect 6430 4830 6490 4890
rect 6430 4790 6440 4830
rect 6480 4790 6490 4830
rect 6430 4730 6490 4790
rect 6430 4690 6440 4730
rect 6480 4690 6490 4730
rect 6430 4670 6490 4690
rect 6630 5430 6690 5450
rect 6630 5390 6640 5430
rect 6680 5390 6690 5430
rect 6630 5330 6690 5390
rect 6630 5290 6640 5330
rect 6680 5290 6690 5330
rect 6630 5230 6690 5290
rect 6630 5190 6640 5230
rect 6680 5190 6690 5230
rect 6630 5130 6690 5190
rect 6630 5090 6640 5130
rect 6680 5090 6690 5130
rect 6630 5030 6690 5090
rect 6630 4990 6640 5030
rect 6680 4990 6690 5030
rect 6630 4930 6690 4990
rect 6630 4890 6640 4930
rect 6680 4890 6690 4930
rect 6630 4830 6690 4890
rect 6630 4790 6640 4830
rect 6680 4790 6690 4830
rect 6630 4730 6690 4790
rect 6630 4690 6640 4730
rect 6680 4690 6690 4730
rect 6630 4670 6690 4690
rect 6830 5430 6890 5450
rect 6830 5390 6840 5430
rect 6880 5390 6890 5430
rect 6830 5330 6890 5390
rect 6830 5290 6840 5330
rect 6880 5290 6890 5330
rect 6830 5230 6890 5290
rect 6830 5190 6840 5230
rect 6880 5190 6890 5230
rect 6830 5130 6890 5190
rect 6830 5090 6840 5130
rect 6880 5090 6890 5130
rect 6830 5030 6890 5090
rect 6830 4990 6840 5030
rect 6880 4990 6890 5030
rect 6830 4930 6890 4990
rect 6830 4890 6840 4930
rect 6880 4890 6890 4930
rect 6830 4830 6890 4890
rect 6830 4790 6840 4830
rect 6880 4790 6890 4830
rect 6830 4730 6890 4790
rect 6830 4690 6840 4730
rect 6880 4690 6890 4730
rect 6830 4670 6890 4690
rect 7030 5430 7090 5450
rect 7030 5390 7040 5430
rect 7080 5390 7090 5430
rect 7030 5330 7090 5390
rect 7030 5290 7040 5330
rect 7080 5290 7090 5330
rect 7030 5230 7090 5290
rect 7030 5190 7040 5230
rect 7080 5190 7090 5230
rect 7030 5130 7090 5190
rect 7030 5090 7040 5130
rect 7080 5090 7090 5130
rect 7030 5030 7090 5090
rect 7030 4990 7040 5030
rect 7080 4990 7090 5030
rect 7030 4930 7090 4990
rect 7030 4890 7040 4930
rect 7080 4890 7090 4930
rect 7030 4830 7090 4890
rect 7030 4790 7040 4830
rect 7080 4790 7090 4830
rect 7030 4730 7090 4790
rect 7030 4690 7040 4730
rect 7080 4690 7090 4730
rect 7030 4670 7090 4690
rect 7230 5430 7290 5450
rect 7230 5390 7240 5430
rect 7280 5390 7290 5430
rect 7230 5330 7290 5390
rect 7230 5290 7240 5330
rect 7280 5290 7290 5330
rect 7230 5230 7290 5290
rect 7230 5190 7240 5230
rect 7280 5190 7290 5230
rect 7230 5130 7290 5190
rect 7230 5090 7240 5130
rect 7280 5090 7290 5130
rect 7230 5030 7290 5090
rect 7230 4990 7240 5030
rect 7280 4990 7290 5030
rect 7230 4930 7290 4990
rect 7230 4890 7240 4930
rect 7280 4890 7290 4930
rect 7230 4830 7290 4890
rect 7230 4790 7240 4830
rect 7280 4790 7290 4830
rect 7230 4730 7290 4790
rect 7230 4690 7240 4730
rect 7280 4690 7290 4730
rect 7230 4670 7290 4690
rect 7430 5430 7490 5450
rect 7430 5390 7440 5430
rect 7480 5390 7490 5430
rect 7430 5330 7490 5390
rect 7430 5290 7440 5330
rect 7480 5290 7490 5330
rect 7430 5230 7490 5290
rect 7430 5190 7440 5230
rect 7480 5190 7490 5230
rect 7430 5130 7490 5190
rect 7430 5090 7440 5130
rect 7480 5090 7490 5130
rect 7430 5030 7490 5090
rect 7430 4990 7440 5030
rect 7480 4990 7490 5030
rect 7430 4930 7490 4990
rect 7430 4890 7440 4930
rect 7480 4890 7490 4930
rect 7430 4830 7490 4890
rect 7430 4790 7440 4830
rect 7480 4790 7490 4830
rect 7430 4730 7490 4790
rect 7430 4690 7440 4730
rect 7480 4690 7490 4730
rect 7430 4670 7490 4690
rect 7630 5430 7690 5450
rect 7630 5390 7640 5430
rect 7680 5390 7690 5430
rect 7630 5330 7690 5390
rect 7630 5290 7640 5330
rect 7680 5290 7690 5330
rect 7630 5230 7690 5290
rect 7630 5190 7640 5230
rect 7680 5190 7690 5230
rect 7630 5130 7690 5190
rect 7630 5090 7640 5130
rect 7680 5090 7690 5130
rect 7630 5030 7690 5090
rect 7630 4990 7640 5030
rect 7680 4990 7690 5030
rect 7630 4930 7690 4990
rect 7630 4890 7640 4930
rect 7680 4890 7690 4930
rect 7630 4830 7690 4890
rect 7630 4790 7640 4830
rect 7680 4790 7690 4830
rect 7630 4730 7690 4790
rect 7630 4690 7640 4730
rect 7680 4690 7690 4730
rect 7630 4670 7690 4690
rect 7830 5430 7890 5450
rect 7830 5390 7840 5430
rect 7880 5390 7890 5430
rect 7830 5330 7890 5390
rect 7830 5290 7840 5330
rect 7880 5290 7890 5330
rect 7830 5230 7890 5290
rect 7830 5190 7840 5230
rect 7880 5190 7890 5230
rect 7830 5130 7890 5190
rect 7830 5090 7840 5130
rect 7880 5090 7890 5130
rect 7830 5030 7890 5090
rect 7830 4990 7840 5030
rect 7880 4990 7890 5030
rect 7830 4930 7890 4990
rect 7830 4890 7840 4930
rect 7880 4890 7890 4930
rect 7830 4830 7890 4890
rect 7830 4790 7840 4830
rect 7880 4790 7890 4830
rect 7830 4730 7890 4790
rect 7830 4690 7840 4730
rect 7880 4690 7890 4730
rect 7830 4670 7890 4690
rect 8030 5430 8090 5450
rect 8030 5390 8040 5430
rect 8080 5390 8090 5430
rect 8030 5330 8090 5390
rect 8030 5290 8040 5330
rect 8080 5290 8090 5330
rect 8030 5230 8090 5290
rect 8030 5190 8040 5230
rect 8080 5190 8090 5230
rect 8030 5130 8090 5190
rect 8030 5090 8040 5130
rect 8080 5090 8090 5130
rect 8030 5030 8090 5090
rect 8030 4990 8040 5030
rect 8080 4990 8090 5030
rect 8030 4930 8090 4990
rect 8030 4890 8040 4930
rect 8080 4890 8090 4930
rect 8030 4830 8090 4890
rect 8030 4790 8040 4830
rect 8080 4790 8090 4830
rect 8030 4730 8090 4790
rect 8030 4690 8040 4730
rect 8080 4690 8090 4730
rect 8030 4670 8090 4690
rect 8230 5430 8370 5450
rect 8230 5390 8240 5430
rect 8280 5390 8320 5430
rect 8360 5390 8370 5430
rect 8230 5330 8370 5390
rect 8230 5290 8240 5330
rect 8280 5290 8320 5330
rect 8360 5290 8370 5330
rect 8230 5230 8370 5290
rect 8230 5190 8240 5230
rect 8280 5190 8320 5230
rect 8360 5190 8370 5230
rect 8230 5130 8370 5190
rect 8230 5090 8240 5130
rect 8280 5090 8320 5130
rect 8360 5090 8370 5130
rect 8230 5030 8370 5090
rect 8230 4990 8240 5030
rect 8280 4990 8320 5030
rect 8360 4990 8370 5030
rect 8230 4930 8370 4990
rect 8230 4890 8240 4930
rect 8280 4890 8320 4930
rect 8360 4890 8370 4930
rect 8230 4830 8370 4890
rect 8230 4790 8240 4830
rect 8280 4790 8320 4830
rect 8360 4790 8370 4830
rect 8230 4730 8370 4790
rect 8230 4690 8240 4730
rect 8280 4690 8320 4730
rect 8360 4690 8370 4730
rect 8230 4670 8370 4690
rect 4840 4630 4880 4670
rect 2010 4570 2450 4620
rect 4820 4610 4900 4630
rect 4820 4570 4840 4610
rect 4880 4570 4900 4610
rect 4820 4550 4900 4570
rect 5240 4540 5280 4670
rect 3790 4440 4230 4500
rect 5220 4520 5300 4540
rect 5220 4480 5240 4520
rect 5280 4480 5300 4520
rect 5220 4460 5300 4480
rect 5640 4450 5680 4670
rect 6040 4540 6080 4670
rect 6220 4610 6300 4630
rect 6220 4570 6240 4610
rect 6280 4570 6300 4610
rect 6220 4550 6300 4570
rect 6020 4520 6100 4540
rect 6020 4480 6040 4520
rect 6080 4480 6100 4520
rect 6020 4460 6100 4480
rect 6440 4450 6480 4670
rect 6840 4630 6880 4670
rect 6620 4610 6700 4630
rect 6620 4570 6640 4610
rect 6680 4570 6700 4610
rect 6620 4550 6700 4570
rect 6820 4610 6900 4630
rect 6820 4570 6840 4610
rect 6880 4570 6900 4610
rect 6820 4550 6900 4570
rect 7240 4450 7280 4670
rect 7640 4630 7680 4670
rect 7620 4610 7700 4630
rect 7620 4570 7640 4610
rect 7680 4570 7700 4610
rect 7620 4550 7700 4570
rect 8040 4540 8080 4670
rect 8140 4610 8220 4630
rect 8140 4570 8160 4610
rect 8200 4570 8220 4610
rect 8140 4550 8220 4570
rect 8020 4520 8100 4540
rect 8020 4480 8040 4520
rect 8080 4480 8100 4520
rect 8020 4460 8100 4480
rect 3790 4400 3810 4440
rect 3850 4400 3900 4440
rect 3940 4400 3990 4440
rect 4030 4400 4080 4440
rect 4120 4400 4170 4440
rect 4210 4400 4230 4440
rect 3790 4380 4230 4400
rect 5620 4430 5700 4450
rect 5620 4390 5640 4430
rect 5680 4390 5700 4430
rect 5620 4370 5700 4390
rect 6420 4430 6500 4450
rect 6420 4390 6440 4430
rect 6480 4390 6500 4430
rect 6420 4370 6500 4390
rect 7220 4430 7300 4450
rect 7220 4390 7240 4430
rect 7280 4390 7300 4430
rect 7220 4370 7300 4390
rect 8750 4410 8830 4420
rect 8750 4370 8770 4410
rect 8810 4390 9110 4410
rect 8810 4370 9050 4390
rect 8750 4350 8830 4370
rect 9030 4350 9050 4370
rect 9090 4350 9110 4390
rect 5220 4310 5300 4330
rect 5220 4270 5240 4310
rect 5280 4270 5300 4310
rect 5220 4250 5300 4270
rect 5620 4310 5700 4330
rect 5620 4270 5640 4310
rect 5680 4270 5700 4310
rect 5620 4250 5700 4270
rect 6020 4310 6100 4330
rect 6020 4270 6040 4310
rect 6080 4270 6100 4310
rect 6020 4250 6100 4270
rect 6220 4310 6300 4330
rect 6220 4270 6240 4310
rect 6280 4270 6300 4310
rect 6220 4250 6300 4270
rect 6420 4310 6500 4330
rect 6420 4270 6440 4310
rect 6480 4270 6500 4310
rect 6420 4250 6500 4270
rect 6620 4310 6700 4330
rect 6620 4270 6640 4310
rect 6680 4270 6700 4310
rect 6620 4250 6700 4270
rect 6820 4310 6900 4330
rect 6820 4270 6840 4310
rect 6880 4270 6900 4310
rect 6820 4250 6900 4270
rect 7220 4310 7300 4330
rect 7220 4270 7240 4310
rect 7280 4270 7300 4310
rect 7220 4250 7300 4270
rect 7620 4310 7700 4330
rect 7620 4270 7640 4310
rect 7680 4270 7700 4310
rect 7620 4250 7700 4270
rect 5240 4210 5280 4250
rect 5640 4210 5680 4250
rect 6040 4210 6080 4250
rect 6240 4210 6280 4250
rect 6440 4210 6480 4250
rect 6640 4210 6680 4250
rect 6840 4210 6880 4250
rect 7240 4210 7280 4250
rect 7640 4210 7680 4250
rect 8770 4210 8810 4350
rect 9030 4330 9110 4350
rect 9170 4310 9250 4330
rect 9170 4270 9190 4310
rect 9230 4270 9250 4310
rect 9170 4250 9250 4270
rect 9190 4210 9230 4250
rect 5150 4190 5290 4210
rect 5150 4150 5160 4190
rect 5200 4150 5240 4190
rect 5280 4150 5290 4190
rect 5150 4090 5290 4150
rect 5150 4050 5160 4090
rect 5200 4050 5240 4090
rect 5280 4050 5290 4090
rect 1890 4010 2010 4030
rect 1890 3970 1910 4010
rect 1950 3970 2010 4010
rect 1890 3960 2010 3970
rect 1890 3950 1970 3960
rect 3790 3910 4230 3960
rect 5150 3990 5290 4050
rect 5150 3950 5160 3990
rect 5200 3950 5240 3990
rect 5280 3950 5290 3990
rect 5150 3890 5290 3950
rect 5150 3850 5160 3890
rect 5200 3850 5240 3890
rect 5280 3850 5290 3890
rect 2010 3790 2450 3840
rect 5150 3830 5290 3850
rect 5430 4190 5490 4210
rect 5430 4150 5440 4190
rect 5480 4150 5490 4190
rect 5430 4090 5490 4150
rect 5430 4050 5440 4090
rect 5480 4050 5490 4090
rect 5430 3990 5490 4050
rect 5430 3950 5440 3990
rect 5480 3950 5490 3990
rect 5430 3890 5490 3950
rect 5430 3850 5440 3890
rect 5480 3850 5490 3890
rect 5430 3830 5490 3850
rect 5630 4190 5690 4210
rect 5630 4150 5640 4190
rect 5680 4150 5690 4190
rect 5630 4090 5690 4150
rect 5630 4050 5640 4090
rect 5680 4050 5690 4090
rect 5630 3990 5690 4050
rect 5630 3950 5640 3990
rect 5680 3950 5690 3990
rect 5630 3890 5690 3950
rect 5630 3850 5640 3890
rect 5680 3850 5690 3890
rect 5630 3830 5690 3850
rect 5830 4190 5890 4210
rect 5830 4150 5840 4190
rect 5880 4150 5890 4190
rect 5830 4090 5890 4150
rect 5830 4050 5840 4090
rect 5880 4050 5890 4090
rect 5830 3990 5890 4050
rect 5830 3950 5840 3990
rect 5880 3950 5890 3990
rect 5830 3890 5890 3950
rect 5830 3850 5840 3890
rect 5880 3850 5890 3890
rect 5830 3830 5890 3850
rect 6030 4190 6090 4210
rect 6030 4150 6040 4190
rect 6080 4150 6090 4190
rect 6030 4090 6090 4150
rect 6030 4050 6040 4090
rect 6080 4050 6090 4090
rect 6030 3990 6090 4050
rect 6030 3950 6040 3990
rect 6080 3950 6090 3990
rect 6030 3890 6090 3950
rect 6030 3850 6040 3890
rect 6080 3850 6090 3890
rect 6030 3830 6090 3850
rect 6230 4190 6290 4210
rect 6230 4150 6240 4190
rect 6280 4150 6290 4190
rect 6230 4090 6290 4150
rect 6230 4050 6240 4090
rect 6280 4050 6290 4090
rect 6230 3990 6290 4050
rect 6230 3950 6240 3990
rect 6280 3950 6290 3990
rect 6230 3890 6290 3950
rect 6230 3850 6240 3890
rect 6280 3850 6290 3890
rect 6230 3830 6290 3850
rect 6430 4190 6490 4210
rect 6430 4150 6440 4190
rect 6480 4150 6490 4190
rect 6430 4090 6490 4150
rect 6430 4050 6440 4090
rect 6480 4050 6490 4090
rect 6430 3990 6490 4050
rect 6430 3950 6440 3990
rect 6480 3950 6490 3990
rect 6430 3890 6490 3950
rect 6430 3850 6440 3890
rect 6480 3850 6490 3890
rect 6430 3830 6490 3850
rect 6630 4190 6690 4210
rect 6630 4150 6640 4190
rect 6680 4150 6690 4190
rect 6630 4090 6690 4150
rect 6630 4050 6640 4090
rect 6680 4050 6690 4090
rect 6630 3990 6690 4050
rect 6630 3950 6640 3990
rect 6680 3950 6690 3990
rect 6630 3890 6690 3950
rect 6630 3850 6640 3890
rect 6680 3850 6690 3890
rect 6630 3830 6690 3850
rect 6830 4190 6890 4210
rect 6830 4150 6840 4190
rect 6880 4150 6890 4190
rect 6830 4090 6890 4150
rect 6830 4050 6840 4090
rect 6880 4050 6890 4090
rect 6830 3990 6890 4050
rect 6830 3950 6840 3990
rect 6880 3950 6890 3990
rect 6830 3890 6890 3950
rect 6830 3850 6840 3890
rect 6880 3850 6890 3890
rect 6830 3830 6890 3850
rect 7030 4190 7090 4210
rect 7030 4150 7040 4190
rect 7080 4150 7090 4190
rect 7030 4090 7090 4150
rect 7030 4050 7040 4090
rect 7080 4050 7090 4090
rect 7030 3990 7090 4050
rect 7030 3950 7040 3990
rect 7080 3950 7090 3990
rect 7030 3890 7090 3950
rect 7030 3850 7040 3890
rect 7080 3850 7090 3890
rect 7030 3830 7090 3850
rect 7230 4190 7290 4210
rect 7230 4150 7240 4190
rect 7280 4150 7290 4190
rect 7230 4090 7290 4150
rect 7230 4050 7240 4090
rect 7280 4050 7290 4090
rect 7230 3990 7290 4050
rect 7230 3950 7240 3990
rect 7280 3950 7290 3990
rect 7230 3890 7290 3950
rect 7230 3850 7240 3890
rect 7280 3850 7290 3890
rect 7230 3830 7290 3850
rect 7430 4190 7490 4210
rect 7430 4150 7440 4190
rect 7480 4150 7490 4190
rect 7430 4090 7490 4150
rect 7430 4050 7440 4090
rect 7480 4050 7490 4090
rect 7430 3990 7490 4050
rect 7430 3950 7440 3990
rect 7480 3950 7490 3990
rect 7430 3890 7490 3950
rect 7430 3850 7440 3890
rect 7480 3850 7490 3890
rect 7430 3830 7490 3850
rect 7630 4190 7770 4210
rect 7630 4150 7640 4190
rect 7680 4150 7720 4190
rect 7760 4150 7770 4190
rect 7630 4090 7770 4150
rect 7630 4050 7640 4090
rect 7680 4050 7720 4090
rect 7760 4050 7770 4090
rect 7630 3990 7770 4050
rect 7630 3950 7640 3990
rect 7680 3950 7720 3990
rect 7760 3950 7770 3990
rect 7630 3890 7770 3950
rect 7630 3850 7640 3890
rect 7680 3850 7720 3890
rect 7760 3850 7770 3890
rect 7630 3830 7770 3850
rect 8760 4190 8820 4210
rect 8760 4150 8770 4190
rect 8810 4150 8820 4190
rect 8760 4090 8820 4150
rect 8760 4050 8770 4090
rect 8810 4050 8820 4090
rect 8760 3990 8820 4050
rect 8760 3950 8770 3990
rect 8810 3950 8820 3990
rect 8760 3890 8820 3950
rect 8760 3850 8770 3890
rect 8810 3850 8820 3890
rect 8760 3830 8820 3850
rect 8870 4190 8930 4210
rect 8870 4150 8880 4190
rect 8920 4150 8930 4190
rect 8870 4090 8930 4150
rect 8870 4050 8880 4090
rect 8920 4050 8930 4090
rect 8870 3990 8930 4050
rect 8870 3950 8880 3990
rect 8920 3950 8930 3990
rect 8870 3890 8930 3950
rect 8870 3850 8880 3890
rect 8920 3850 8930 3890
rect 8870 3830 8930 3850
rect 9010 4190 9070 4210
rect 9010 4150 9020 4190
rect 9060 4150 9070 4190
rect 9010 4090 9070 4150
rect 9010 4050 9020 4090
rect 9060 4050 9070 4090
rect 9010 3990 9070 4050
rect 9010 3950 9020 3990
rect 9060 3950 9070 3990
rect 9010 3890 9070 3950
rect 9010 3850 9020 3890
rect 9060 3850 9070 3890
rect 9010 3830 9070 3850
rect 9120 4190 9230 4210
rect 9120 4150 9130 4190
rect 9170 4150 9230 4190
rect 9120 4090 9190 4150
rect 9120 4050 9130 4090
rect 9170 4050 9190 4090
rect 9120 3990 9190 4050
rect 9120 3950 9130 3990
rect 9170 3950 9190 3990
rect 9120 3890 9190 3950
rect 9120 3850 9130 3890
rect 9170 3850 9190 3890
rect 9120 3830 9190 3850
rect 3790 3670 4230 3720
rect 5440 3700 5480 3830
rect 5840 3790 5880 3830
rect 6240 3790 6280 3830
rect 6640 3790 6680 3830
rect 7040 3790 7080 3830
rect 5820 3770 5900 3790
rect 5820 3730 5840 3770
rect 5880 3730 5900 3770
rect 6240 3770 6680 3790
rect 6240 3750 6480 3770
rect 5820 3710 5900 3730
rect 6460 3730 6480 3750
rect 6520 3750 6680 3770
rect 7020 3770 7100 3790
rect 6520 3730 6540 3750
rect 6460 3710 6540 3730
rect 7020 3730 7040 3770
rect 7080 3730 7100 3770
rect 7020 3710 7100 3730
rect 7440 3700 7480 3830
rect 5420 3680 5500 3700
rect 5420 3640 5440 3680
rect 5480 3640 5500 3680
rect 5420 3620 5500 3640
rect 6330 3680 6410 3700
rect 6330 3640 6350 3680
rect 6390 3640 6410 3680
rect 6330 3620 6410 3640
rect 7420 3680 7500 3700
rect 7420 3640 7440 3680
rect 7480 3640 7500 3680
rect 7420 3620 7500 3640
rect 2010 3550 2450 3600
rect 6460 3590 6540 3610
rect 6460 3550 6480 3590
rect 6520 3550 6540 3590
rect 6460 3530 6540 3550
rect 3790 3420 4230 3480
rect 5820 3500 5900 3520
rect 5820 3460 5840 3500
rect 5880 3460 5900 3500
rect 5820 3440 5900 3460
rect 7020 3500 7100 3520
rect 7020 3460 7040 3500
rect 7080 3460 7100 3500
rect 7020 3440 7100 3460
rect 3790 3380 3810 3420
rect 3850 3380 3900 3420
rect 3940 3380 3990 3420
rect 4030 3380 4080 3420
rect 4120 3380 4170 3420
rect 4210 3380 4230 3420
rect 3790 3360 4230 3380
rect 5840 3310 5880 3440
rect 6100 3410 6180 3430
rect 6100 3370 6120 3410
rect 6160 3370 6180 3410
rect 6100 3350 6180 3370
rect 6220 3410 6300 3430
rect 6220 3370 6240 3410
rect 6280 3370 6300 3410
rect 6220 3350 6300 3370
rect 6620 3410 6700 3430
rect 6620 3370 6640 3410
rect 6680 3370 6700 3410
rect 6620 3350 6700 3370
rect 6740 3410 6820 3430
rect 6740 3370 6760 3410
rect 6800 3370 6820 3410
rect 6740 3350 6820 3370
rect 6240 3310 6280 3350
rect 6640 3310 6680 3350
rect 7040 3310 7080 3440
rect 8880 3430 8920 3830
rect 9010 3760 9050 3830
rect 8970 3740 9050 3760
rect 8970 3700 8990 3740
rect 9030 3700 9050 3740
rect 8970 3680 9050 3700
rect 8860 3410 8940 3430
rect 8860 3370 8880 3410
rect 8920 3370 8940 3410
rect 8860 3350 8940 3370
rect 5620 3290 5690 3310
rect 5620 3250 5640 3290
rect 5680 3250 5690 3290
rect 5620 3190 5690 3250
rect 5620 3150 5640 3190
rect 5680 3150 5690 3190
rect 5620 3130 5690 3150
rect 5830 3290 5890 3310
rect 5830 3250 5840 3290
rect 5880 3250 5890 3290
rect 5830 3190 5890 3250
rect 5830 3150 5840 3190
rect 5880 3150 5890 3190
rect 5830 3130 5890 3150
rect 6030 3290 6090 3310
rect 6030 3250 6040 3290
rect 6080 3250 6090 3290
rect 6030 3190 6090 3250
rect 6030 3150 6040 3190
rect 6080 3150 6090 3190
rect 6030 3130 6090 3150
rect 6230 3290 6290 3310
rect 6230 3250 6240 3290
rect 6280 3250 6290 3290
rect 6230 3190 6290 3250
rect 6230 3150 6240 3190
rect 6280 3150 6290 3190
rect 6230 3130 6290 3150
rect 6430 3290 6490 3310
rect 6430 3250 6440 3290
rect 6480 3250 6490 3290
rect 6430 3190 6490 3250
rect 6430 3150 6440 3190
rect 6480 3150 6490 3190
rect 6430 3130 6490 3150
rect 6630 3290 6690 3310
rect 6630 3250 6640 3290
rect 6680 3250 6690 3290
rect 6630 3190 6690 3250
rect 6630 3150 6640 3190
rect 6680 3150 6690 3190
rect 6630 3130 6690 3150
rect 6830 3290 6890 3310
rect 6830 3250 6840 3290
rect 6880 3250 6890 3290
rect 6830 3190 6890 3250
rect 6830 3150 6840 3190
rect 6880 3150 6890 3190
rect 6830 3130 6890 3150
rect 7030 3290 7090 3310
rect 7030 3250 7040 3290
rect 7080 3250 7090 3290
rect 7030 3190 7090 3250
rect 7030 3150 7040 3190
rect 7080 3150 7090 3190
rect 7030 3130 7090 3150
rect 7230 3290 7300 3310
rect 7230 3250 7240 3290
rect 7280 3250 7300 3290
rect 7230 3190 7300 3250
rect 7230 3150 7240 3190
rect 7280 3150 7300 3190
rect 7230 3130 7300 3150
rect 1890 3060 2010 3080
rect 1890 3020 1910 3060
rect 1950 3020 2010 3060
rect 1890 3010 2010 3020
rect 3590 3060 4230 3080
rect 3590 3020 3810 3060
rect 3850 3020 3900 3060
rect 3940 3020 3990 3060
rect 4030 3020 4080 3060
rect 4120 3020 4170 3060
rect 4210 3020 4230 3060
rect 3590 3010 4230 3020
rect 1890 3000 1970 3010
rect 3790 2960 4230 3010
rect 5640 3000 5680 3130
rect 5820 3070 5900 3090
rect 5820 3030 5840 3070
rect 5880 3030 5900 3070
rect 5820 3010 5900 3030
rect 6040 3000 6080 3130
rect 6440 3000 6480 3130
rect 6840 3000 6880 3130
rect 7020 3070 7100 3090
rect 7020 3030 7040 3070
rect 7080 3030 7100 3070
rect 7020 3010 7100 3030
rect 7240 3000 7280 3130
rect 5620 2980 5700 3000
rect 5620 2940 5640 2980
rect 5680 2940 5700 2980
rect 5620 2920 5700 2940
rect 6020 2980 6100 3000
rect 6020 2940 6040 2980
rect 6080 2940 6100 2980
rect 6020 2920 6100 2940
rect 6420 2980 6500 3000
rect 6420 2940 6440 2980
rect 6480 2940 6500 2980
rect 6420 2920 6500 2940
rect 6820 2980 6900 3000
rect 6820 2940 6840 2980
rect 6880 2940 6900 2980
rect 6820 2920 6900 2940
rect 7220 2980 7300 3000
rect 7220 2940 7240 2980
rect 7280 2940 7300 2980
rect 7220 2920 7300 2940
rect 2010 2840 2450 2890
rect 5640 2880 5680 2920
rect 6040 2880 6080 2920
rect 5470 2860 6340 2880
rect 3790 2720 4230 2770
rect 5470 2820 5560 2860
rect 5600 2820 5640 2860
rect 5680 2820 5720 2860
rect 5760 2820 5800 2860
rect 5840 2820 5880 2860
rect 5920 2820 5960 2860
rect 6000 2820 6040 2860
rect 6080 2820 6120 2860
rect 6160 2820 6200 2860
rect 6240 2820 6280 2860
rect 6320 2820 6340 2860
rect 5470 2800 6340 2820
rect 6580 2860 7460 2880
rect 6580 2820 6600 2860
rect 6640 2820 6680 2860
rect 6720 2820 6760 2860
rect 6800 2820 6840 2860
rect 6880 2820 6920 2860
rect 6960 2820 7000 2860
rect 7040 2820 7080 2860
rect 7120 2820 7160 2860
rect 7200 2820 7240 2860
rect 7280 2820 7320 2860
rect 7360 2820 7400 2860
rect 7440 2820 7460 2860
rect 6580 2800 7460 2820
rect 5470 2740 5530 2800
rect 5470 2700 5480 2740
rect 5520 2700 5530 2740
rect 2010 2600 2450 2650
rect 5470 2640 5530 2700
rect 5470 2600 5480 2640
rect 5520 2600 5530 2640
rect 1890 2480 1970 2490
rect 3790 2480 4230 2530
rect 1890 2470 2010 2480
rect 1890 2430 1910 2470
rect 1950 2430 2010 2470
rect 1890 2410 2010 2430
rect 5470 2540 5530 2600
rect 5470 2500 5480 2540
rect 5520 2500 5530 2540
rect 5470 2440 5530 2500
rect 5470 2400 5480 2440
rect 5520 2400 5530 2440
rect 5470 2340 5530 2400
rect 5470 2300 5480 2340
rect 5520 2300 5530 2340
rect 5470 2240 5530 2300
rect 5470 2200 5480 2240
rect 5520 2200 5530 2240
rect 5470 2140 5530 2200
rect 5470 2100 5480 2140
rect 5520 2100 5530 2140
rect 5470 2040 5530 2100
rect 5470 2000 5480 2040
rect 5520 2000 5530 2040
rect 5470 1980 5530 2000
rect 6350 2740 6570 2760
rect 6350 2700 6360 2740
rect 6400 2700 6440 2740
rect 6480 2700 6520 2740
rect 6560 2700 6570 2740
rect 6350 2640 6570 2700
rect 6350 2600 6360 2640
rect 6400 2600 6440 2640
rect 6480 2600 6520 2640
rect 6560 2600 6570 2640
rect 6350 2540 6570 2600
rect 6350 2500 6360 2540
rect 6400 2500 6440 2540
rect 6480 2500 6520 2540
rect 6560 2500 6570 2540
rect 6350 2440 6570 2500
rect 6350 2400 6360 2440
rect 6400 2400 6440 2440
rect 6480 2400 6520 2440
rect 6560 2400 6570 2440
rect 6350 2340 6570 2400
rect 6350 2300 6360 2340
rect 6400 2300 6440 2340
rect 6480 2300 6520 2340
rect 6560 2300 6570 2340
rect 6350 2240 6570 2300
rect 6350 2200 6360 2240
rect 6400 2200 6440 2240
rect 6480 2200 6520 2240
rect 6560 2200 6570 2240
rect 6350 2140 6570 2200
rect 6350 2100 6360 2140
rect 6400 2100 6440 2140
rect 6480 2100 6520 2140
rect 6560 2100 6570 2140
rect 6350 2040 6570 2100
rect 6350 2000 6360 2040
rect 6400 2000 6440 2040
rect 6480 2000 6520 2040
rect 6560 2000 6570 2040
rect 6350 1980 6570 2000
rect 7390 2740 7450 2800
rect 7390 2700 7400 2740
rect 7440 2700 7450 2740
rect 7390 2640 7450 2700
rect 7390 2600 7400 2640
rect 7440 2600 7450 2640
rect 7390 2540 7450 2600
rect 7390 2500 7400 2540
rect 7440 2500 7450 2540
rect 7390 2440 7450 2500
rect 7390 2400 7400 2440
rect 7440 2400 7450 2440
rect 7390 2340 7450 2400
rect 7390 2300 7400 2340
rect 7440 2300 7450 2340
rect 7390 2240 7450 2300
rect 7390 2200 7400 2240
rect 7440 2200 7450 2240
rect 7390 2140 7450 2200
rect 7390 2100 7400 2140
rect 7440 2100 7450 2140
rect 7390 2040 7450 2100
rect 7390 2000 7400 2040
rect 7440 2000 7450 2040
rect 7390 1980 7450 2000
rect 6360 1940 6400 1980
rect 6440 1940 6480 1980
rect 6520 1940 6560 1980
rect 6340 1920 6580 1940
rect 6340 1880 6360 1920
rect 6400 1880 6440 1920
rect 6480 1880 6520 1920
rect 6560 1880 6580 1920
rect 6340 1860 6580 1880
rect 5380 1800 7520 1820
rect 5380 1760 5460 1800
rect 5500 1760 5620 1800
rect 5660 1760 5780 1800
rect 5820 1760 5940 1800
rect 5980 1760 6100 1800
rect 6140 1760 6260 1800
rect 6300 1760 6420 1800
rect 6460 1760 6580 1800
rect 6620 1760 6740 1800
rect 6780 1760 6900 1800
rect 6940 1760 7060 1800
rect 7100 1760 7220 1800
rect 7260 1760 7380 1800
rect 7420 1760 7460 1800
rect 7500 1760 7520 1800
rect 5380 1740 7520 1760
rect 5380 1700 5420 1740
rect 5370 1680 5430 1700
rect 1300 1640 1380 1660
rect 1300 1600 1320 1640
rect 1360 1600 1380 1640
rect 1300 1540 1380 1600
rect 1300 1500 1320 1540
rect 1360 1500 1380 1540
rect 5370 1640 5380 1680
rect 5420 1640 5430 1680
rect 5370 1580 5430 1640
rect 5370 1540 5380 1580
rect 5420 1540 5430 1580
rect 5370 1520 5430 1540
rect 7450 1680 7590 1700
rect 7450 1640 7460 1680
rect 7500 1640 7540 1680
rect 7580 1650 7590 1680
rect 7580 1640 7670 1650
rect 7450 1630 7670 1640
rect 7450 1590 7610 1630
rect 7650 1590 7670 1630
rect 7450 1580 7670 1590
rect 7450 1540 7460 1580
rect 7500 1540 7540 1580
rect 7580 1570 7670 1580
rect 7580 1540 7590 1570
rect 7450 1520 7590 1540
rect 1300 1440 1380 1500
rect 1300 1400 1320 1440
rect 1360 1400 1380 1440
rect 1300 1380 1380 1400
rect 10 1279 9470 1320
rect 10 1256 1506 1279
rect 10 1222 1410 1256
rect 1444 1245 1506 1256
rect 1540 1245 1596 1279
rect 1630 1245 1686 1279
rect 1720 1245 1776 1279
rect 1810 1245 1866 1279
rect 1900 1245 1956 1279
rect 1990 1245 2046 1279
rect 2080 1245 2136 1279
rect 2170 1245 2226 1279
rect 2260 1245 2316 1279
rect 2350 1245 2406 1279
rect 2440 1245 2496 1279
rect 2530 1256 2866 1279
rect 2530 1245 2597 1256
rect 1444 1222 2597 1245
rect 2631 1222 2770 1256
rect 2804 1245 2866 1256
rect 2900 1245 2956 1279
rect 2990 1245 3046 1279
rect 3080 1245 3136 1279
rect 3170 1245 3226 1279
rect 3260 1245 3316 1279
rect 3350 1245 3406 1279
rect 3440 1245 3496 1279
rect 3530 1245 3586 1279
rect 3620 1245 3676 1279
rect 3710 1245 3766 1279
rect 3800 1245 3856 1279
rect 3890 1256 4226 1279
rect 3890 1245 3957 1256
rect 2804 1222 3957 1245
rect 3991 1222 4130 1256
rect 4164 1245 4226 1256
rect 4260 1245 4316 1279
rect 4350 1245 4406 1279
rect 4440 1245 4496 1279
rect 4530 1245 4586 1279
rect 4620 1245 4676 1279
rect 4710 1245 4766 1279
rect 4800 1245 4856 1279
rect 4890 1245 4946 1279
rect 4980 1245 5036 1279
rect 5070 1245 5126 1279
rect 5160 1245 5216 1279
rect 5250 1256 5586 1279
rect 5250 1245 5317 1256
rect 4164 1222 5317 1245
rect 5351 1222 5490 1256
rect 5524 1245 5586 1256
rect 5620 1245 5676 1279
rect 5710 1245 5766 1279
rect 5800 1245 5856 1279
rect 5890 1245 5946 1279
rect 5980 1245 6036 1279
rect 6070 1245 6126 1279
rect 6160 1245 6216 1279
rect 6250 1245 6306 1279
rect 6340 1245 6396 1279
rect 6430 1245 6486 1279
rect 6520 1245 6576 1279
rect 6610 1256 6946 1279
rect 6610 1245 6677 1256
rect 5524 1222 6677 1245
rect 6711 1222 6850 1256
rect 6884 1245 6946 1256
rect 6980 1245 7036 1279
rect 7070 1245 7126 1279
rect 7160 1245 7216 1279
rect 7250 1245 7306 1279
rect 7340 1245 7396 1279
rect 7430 1245 7486 1279
rect 7520 1245 7576 1279
rect 7610 1245 7666 1279
rect 7700 1245 7756 1279
rect 7790 1245 7846 1279
rect 7880 1245 7936 1279
rect 7970 1256 8306 1279
rect 7970 1245 8037 1256
rect 6884 1222 8037 1245
rect 8071 1222 8210 1256
rect 8244 1245 8306 1256
rect 8340 1245 8396 1279
rect 8430 1245 8486 1279
rect 8520 1245 8576 1279
rect 8610 1245 8666 1279
rect 8700 1245 8756 1279
rect 8790 1245 8846 1279
rect 8880 1245 8936 1279
rect 8970 1245 9026 1279
rect 9060 1245 9116 1279
rect 9150 1245 9206 1279
rect 9240 1245 9296 1279
rect 9330 1256 9470 1279
rect 9330 1245 9397 1256
rect 8244 1222 9397 1245
rect 9431 1222 9470 1256
rect 10 1166 9470 1222
rect 10 1132 1410 1166
rect 1444 1132 2597 1166
rect 2631 1132 2770 1166
rect 2804 1132 3957 1166
rect 3991 1132 4130 1166
rect 4164 1132 5317 1166
rect 5351 1132 5490 1166
rect 5524 1132 6677 1166
rect 6711 1132 6850 1166
rect 6884 1132 8037 1166
rect 8071 1132 8210 1166
rect 8244 1132 9397 1166
rect 9431 1132 9470 1166
rect 10 1098 1670 1132
rect 1704 1098 1760 1132
rect 1794 1098 1850 1132
rect 1884 1098 1940 1132
rect 1974 1098 2030 1132
rect 2064 1098 2120 1132
rect 2154 1098 2210 1132
rect 2244 1098 2300 1132
rect 2334 1098 2390 1132
rect 2424 1098 3030 1132
rect 3064 1098 3120 1132
rect 3154 1098 3210 1132
rect 3244 1098 3300 1132
rect 3334 1098 3390 1132
rect 3424 1098 3480 1132
rect 3514 1098 3570 1132
rect 3604 1098 3660 1132
rect 3694 1098 3750 1132
rect 3784 1098 4390 1132
rect 4424 1098 4480 1132
rect 4514 1098 4570 1132
rect 4604 1098 4660 1132
rect 4694 1098 4750 1132
rect 4784 1098 4840 1132
rect 4874 1098 4930 1132
rect 4964 1098 5020 1132
rect 5054 1098 5110 1132
rect 5144 1098 5750 1132
rect 5784 1098 5840 1132
rect 5874 1098 5930 1132
rect 5964 1098 6020 1132
rect 6054 1098 6110 1132
rect 6144 1098 6200 1132
rect 6234 1098 6290 1132
rect 6324 1098 6380 1132
rect 6414 1098 6470 1132
rect 6504 1098 7110 1132
rect 7144 1098 7200 1132
rect 7234 1098 7290 1132
rect 7324 1098 7380 1132
rect 7414 1098 7470 1132
rect 7504 1098 7560 1132
rect 7594 1098 7650 1132
rect 7684 1098 7740 1132
rect 7774 1098 7830 1132
rect 7864 1098 8470 1132
rect 8504 1098 8560 1132
rect 8594 1098 8650 1132
rect 8684 1098 8740 1132
rect 8774 1098 8830 1132
rect 8864 1098 8920 1132
rect 8954 1098 9010 1132
rect 9044 1098 9100 1132
rect 9134 1098 9190 1132
rect 9224 1098 9470 1132
rect 10 1076 9470 1098
rect 10 1070 1410 1076
rect 10 270 260 1070
rect 1060 1042 1410 1070
rect 1444 1075 2597 1076
rect 1444 1042 1558 1075
rect 1060 1041 1558 1042
rect 1592 1070 2597 1075
rect 1592 1041 1620 1070
rect 1060 986 1620 1041
rect 2420 1056 2597 1070
rect 2420 1022 2448 1056
rect 2482 1042 2597 1056
rect 2631 1042 2770 1076
rect 2804 1075 3957 1076
rect 2804 1042 2918 1075
rect 2482 1041 2918 1042
rect 2952 1070 3957 1075
rect 2952 1041 2980 1070
rect 2482 1022 2980 1041
rect 1060 952 1410 986
rect 1444 985 1620 986
rect 1444 952 1558 985
rect 1060 951 1558 952
rect 1592 951 1620 985
rect 1060 896 1620 951
rect 1060 862 1410 896
rect 1444 895 1620 896
rect 1444 862 1558 895
rect 1060 861 1558 862
rect 1592 861 1620 895
rect 1060 806 1620 861
rect 1060 772 1410 806
rect 1444 805 1620 806
rect 1444 772 1558 805
rect 1060 771 1558 772
rect 1592 771 1620 805
rect 1060 716 1620 771
rect 1060 682 1410 716
rect 1444 715 1620 716
rect 1444 682 1558 715
rect 1060 681 1558 682
rect 1592 681 1620 715
rect 1060 626 1620 681
rect 1060 592 1410 626
rect 1444 625 1620 626
rect 1444 592 1558 625
rect 1060 591 1558 592
rect 1592 591 1620 625
rect 1060 536 1620 591
rect 1060 502 1410 536
rect 1444 535 1620 536
rect 1444 502 1558 535
rect 1060 501 1558 502
rect 1592 501 1620 535
rect 1060 446 1620 501
rect 1060 412 1410 446
rect 1444 445 1620 446
rect 1444 412 1558 445
rect 1060 411 1558 412
rect 1592 411 1620 445
rect 1060 356 1620 411
rect 1060 322 1410 356
rect 1444 355 1620 356
rect 1444 322 1558 355
rect 1060 321 1558 322
rect 1592 321 1620 355
rect 1673 958 2367 1017
rect 1673 924 1734 958
rect 1768 930 1824 958
rect 1858 930 1914 958
rect 1948 930 2004 958
rect 1780 924 1824 930
rect 1880 924 1914 930
rect 1980 924 2004 930
rect 2038 930 2094 958
rect 2038 924 2046 930
rect 1673 896 1746 924
rect 1780 896 1846 924
rect 1880 896 1946 924
rect 1980 896 2046 924
rect 2080 924 2094 930
rect 2128 930 2184 958
rect 2128 924 2146 930
rect 2080 896 2146 924
rect 2180 924 2184 930
rect 2218 930 2274 958
rect 2218 924 2246 930
rect 2308 924 2367 958
rect 2180 896 2246 924
rect 2280 896 2367 924
rect 1673 868 2367 896
rect 1673 834 1734 868
rect 1768 834 1824 868
rect 1858 834 1914 868
rect 1948 834 2004 868
rect 2038 834 2094 868
rect 2128 834 2184 868
rect 2218 834 2274 868
rect 2308 834 2367 868
rect 1673 830 2367 834
rect 1673 796 1746 830
rect 1780 796 1846 830
rect 1880 796 1946 830
rect 1980 796 2046 830
rect 2080 796 2146 830
rect 2180 796 2246 830
rect 2280 796 2367 830
rect 1673 778 2367 796
rect 1673 744 1734 778
rect 1768 744 1824 778
rect 1858 744 1914 778
rect 1948 744 2004 778
rect 2038 744 2094 778
rect 2128 744 2184 778
rect 2218 744 2274 778
rect 2308 744 2367 778
rect 1673 730 2367 744
rect 1673 696 1746 730
rect 1780 696 1846 730
rect 1880 696 1946 730
rect 1980 696 2046 730
rect 2080 696 2146 730
rect 2180 696 2246 730
rect 2280 696 2367 730
rect 1673 688 2367 696
rect 1673 654 1734 688
rect 1768 654 1824 688
rect 1858 654 1914 688
rect 1948 654 2004 688
rect 2038 654 2094 688
rect 2128 654 2184 688
rect 2218 654 2274 688
rect 2308 654 2367 688
rect 1673 630 2367 654
rect 1673 598 1746 630
rect 1780 598 1846 630
rect 1880 598 1946 630
rect 1980 598 2046 630
rect 1673 564 1734 598
rect 1780 596 1824 598
rect 1880 596 1914 598
rect 1980 596 2004 598
rect 1768 564 1824 596
rect 1858 564 1914 596
rect 1948 564 2004 596
rect 2038 596 2046 598
rect 2080 598 2146 630
rect 2080 596 2094 598
rect 2038 564 2094 596
rect 2128 596 2146 598
rect 2180 598 2246 630
rect 2280 598 2367 630
rect 2180 596 2184 598
rect 2128 564 2184 596
rect 2218 596 2246 598
rect 2218 564 2274 596
rect 2308 564 2367 598
rect 1673 530 2367 564
rect 1673 508 1746 530
rect 1780 508 1846 530
rect 1880 508 1946 530
rect 1980 508 2046 530
rect 1673 474 1734 508
rect 1780 496 1824 508
rect 1880 496 1914 508
rect 1980 496 2004 508
rect 1768 474 1824 496
rect 1858 474 1914 496
rect 1948 474 2004 496
rect 2038 496 2046 508
rect 2080 508 2146 530
rect 2080 496 2094 508
rect 2038 474 2094 496
rect 2128 496 2146 508
rect 2180 508 2246 530
rect 2280 508 2367 530
rect 2180 496 2184 508
rect 2128 474 2184 496
rect 2218 496 2246 508
rect 2218 474 2274 496
rect 2308 474 2367 508
rect 1673 430 2367 474
rect 1673 418 1746 430
rect 1780 418 1846 430
rect 1880 418 1946 430
rect 1980 418 2046 430
rect 1673 384 1734 418
rect 1780 396 1824 418
rect 1880 396 1914 418
rect 1980 396 2004 418
rect 1768 384 1824 396
rect 1858 384 1914 396
rect 1948 384 2004 396
rect 2038 396 2046 418
rect 2080 418 2146 430
rect 2080 396 2094 418
rect 2038 384 2094 396
rect 2128 396 2146 418
rect 2180 418 2246 430
rect 2280 418 2367 430
rect 2180 396 2184 418
rect 2128 384 2184 396
rect 2218 396 2246 418
rect 2218 384 2274 396
rect 2308 384 2367 418
rect 1673 323 2367 384
rect 2420 986 2980 1022
rect 3780 1056 3957 1070
rect 3780 1022 3808 1056
rect 3842 1042 3957 1056
rect 3991 1042 4130 1076
rect 4164 1075 5317 1076
rect 4164 1042 4278 1075
rect 3842 1041 4278 1042
rect 4312 1070 5317 1075
rect 4312 1041 4340 1070
rect 3842 1022 4340 1041
rect 2420 966 2597 986
rect 2420 932 2448 966
rect 2482 952 2597 966
rect 2631 952 2770 986
rect 2804 985 2980 986
rect 2804 952 2918 985
rect 2482 951 2918 952
rect 2952 951 2980 985
rect 2482 932 2980 951
rect 2420 896 2980 932
rect 2420 876 2597 896
rect 2420 842 2448 876
rect 2482 862 2597 876
rect 2631 862 2770 896
rect 2804 895 2980 896
rect 2804 862 2918 895
rect 2482 861 2918 862
rect 2952 861 2980 895
rect 2482 842 2980 861
rect 2420 806 2980 842
rect 2420 786 2597 806
rect 2420 752 2448 786
rect 2482 772 2597 786
rect 2631 772 2770 806
rect 2804 805 2980 806
rect 2804 772 2918 805
rect 2482 771 2918 772
rect 2952 771 2980 805
rect 2482 752 2980 771
rect 2420 716 2980 752
rect 2420 696 2597 716
rect 2420 662 2448 696
rect 2482 682 2597 696
rect 2631 682 2770 716
rect 2804 715 2980 716
rect 2804 682 2918 715
rect 2482 681 2918 682
rect 2952 681 2980 715
rect 2482 662 2980 681
rect 2420 626 2980 662
rect 2420 606 2597 626
rect 2420 572 2448 606
rect 2482 592 2597 606
rect 2631 592 2770 626
rect 2804 625 2980 626
rect 2804 592 2918 625
rect 2482 591 2918 592
rect 2952 591 2980 625
rect 2482 572 2980 591
rect 2420 536 2980 572
rect 2420 516 2597 536
rect 2420 482 2448 516
rect 2482 502 2597 516
rect 2631 502 2770 536
rect 2804 535 2980 536
rect 2804 502 2918 535
rect 2482 501 2918 502
rect 2952 501 2980 535
rect 2482 482 2980 501
rect 2420 446 2980 482
rect 2420 426 2597 446
rect 2420 392 2448 426
rect 2482 412 2597 426
rect 2631 412 2770 446
rect 2804 445 2980 446
rect 2804 412 2918 445
rect 2482 411 2918 412
rect 2952 411 2980 445
rect 2482 392 2980 411
rect 2420 356 2980 392
rect 2420 336 2597 356
rect 1060 270 1620 321
rect 2420 302 2448 336
rect 2482 322 2597 336
rect 2631 322 2770 356
rect 2804 355 2980 356
rect 2804 322 2918 355
rect 2482 321 2918 322
rect 2952 321 2980 355
rect 3033 958 3727 1017
rect 3033 924 3094 958
rect 3128 930 3184 958
rect 3218 930 3274 958
rect 3308 930 3364 958
rect 3140 924 3184 930
rect 3240 924 3274 930
rect 3340 924 3364 930
rect 3398 930 3454 958
rect 3398 924 3406 930
rect 3033 896 3106 924
rect 3140 896 3206 924
rect 3240 896 3306 924
rect 3340 896 3406 924
rect 3440 924 3454 930
rect 3488 930 3544 958
rect 3488 924 3506 930
rect 3440 896 3506 924
rect 3540 924 3544 930
rect 3578 930 3634 958
rect 3578 924 3606 930
rect 3668 924 3727 958
rect 3540 896 3606 924
rect 3640 896 3727 924
rect 3033 868 3727 896
rect 3033 834 3094 868
rect 3128 834 3184 868
rect 3218 834 3274 868
rect 3308 834 3364 868
rect 3398 834 3454 868
rect 3488 834 3544 868
rect 3578 834 3634 868
rect 3668 834 3727 868
rect 3033 830 3727 834
rect 3033 796 3106 830
rect 3140 796 3206 830
rect 3240 796 3306 830
rect 3340 796 3406 830
rect 3440 796 3506 830
rect 3540 796 3606 830
rect 3640 796 3727 830
rect 3033 778 3727 796
rect 3033 744 3094 778
rect 3128 744 3184 778
rect 3218 744 3274 778
rect 3308 744 3364 778
rect 3398 744 3454 778
rect 3488 744 3544 778
rect 3578 744 3634 778
rect 3668 744 3727 778
rect 3033 730 3727 744
rect 3033 696 3106 730
rect 3140 696 3206 730
rect 3240 696 3306 730
rect 3340 696 3406 730
rect 3440 696 3506 730
rect 3540 696 3606 730
rect 3640 696 3727 730
rect 3033 688 3727 696
rect 3033 654 3094 688
rect 3128 654 3184 688
rect 3218 654 3274 688
rect 3308 654 3364 688
rect 3398 654 3454 688
rect 3488 654 3544 688
rect 3578 654 3634 688
rect 3668 654 3727 688
rect 3033 630 3727 654
rect 3033 598 3106 630
rect 3140 598 3206 630
rect 3240 598 3306 630
rect 3340 598 3406 630
rect 3033 564 3094 598
rect 3140 596 3184 598
rect 3240 596 3274 598
rect 3340 596 3364 598
rect 3128 564 3184 596
rect 3218 564 3274 596
rect 3308 564 3364 596
rect 3398 596 3406 598
rect 3440 598 3506 630
rect 3440 596 3454 598
rect 3398 564 3454 596
rect 3488 596 3506 598
rect 3540 598 3606 630
rect 3640 598 3727 630
rect 3540 596 3544 598
rect 3488 564 3544 596
rect 3578 596 3606 598
rect 3578 564 3634 596
rect 3668 564 3727 598
rect 3033 530 3727 564
rect 3033 508 3106 530
rect 3140 508 3206 530
rect 3240 508 3306 530
rect 3340 508 3406 530
rect 3033 474 3094 508
rect 3140 496 3184 508
rect 3240 496 3274 508
rect 3340 496 3364 508
rect 3128 474 3184 496
rect 3218 474 3274 496
rect 3308 474 3364 496
rect 3398 496 3406 508
rect 3440 508 3506 530
rect 3440 496 3454 508
rect 3398 474 3454 496
rect 3488 496 3506 508
rect 3540 508 3606 530
rect 3640 508 3727 530
rect 3540 496 3544 508
rect 3488 474 3544 496
rect 3578 496 3606 508
rect 3578 474 3634 496
rect 3668 474 3727 508
rect 3033 430 3727 474
rect 3033 418 3106 430
rect 3140 418 3206 430
rect 3240 418 3306 430
rect 3340 418 3406 430
rect 3033 384 3094 418
rect 3140 396 3184 418
rect 3240 396 3274 418
rect 3340 396 3364 418
rect 3128 384 3184 396
rect 3218 384 3274 396
rect 3308 384 3364 396
rect 3398 396 3406 418
rect 3440 418 3506 430
rect 3440 396 3454 418
rect 3398 384 3454 396
rect 3488 396 3506 418
rect 3540 418 3606 430
rect 3640 418 3727 430
rect 3540 396 3544 418
rect 3488 384 3544 396
rect 3578 396 3606 418
rect 3578 384 3634 396
rect 3668 384 3727 418
rect 3033 323 3727 384
rect 3780 986 4340 1022
rect 5140 1056 5317 1070
rect 5140 1022 5168 1056
rect 5202 1042 5317 1056
rect 5351 1042 5490 1076
rect 5524 1075 6677 1076
rect 5524 1042 5638 1075
rect 5202 1041 5638 1042
rect 5672 1070 6677 1075
rect 5672 1041 5700 1070
rect 5202 1022 5700 1041
rect 3780 966 3957 986
rect 3780 932 3808 966
rect 3842 952 3957 966
rect 3991 952 4130 986
rect 4164 985 4340 986
rect 4164 952 4278 985
rect 3842 951 4278 952
rect 4312 951 4340 985
rect 3842 932 4340 951
rect 3780 896 4340 932
rect 3780 876 3957 896
rect 3780 842 3808 876
rect 3842 862 3957 876
rect 3991 862 4130 896
rect 4164 895 4340 896
rect 4164 862 4278 895
rect 3842 861 4278 862
rect 4312 861 4340 895
rect 3842 842 4340 861
rect 3780 806 4340 842
rect 3780 786 3957 806
rect 3780 752 3808 786
rect 3842 772 3957 786
rect 3991 772 4130 806
rect 4164 805 4340 806
rect 4164 772 4278 805
rect 3842 771 4278 772
rect 4312 771 4340 805
rect 3842 752 4340 771
rect 3780 716 4340 752
rect 3780 696 3957 716
rect 3780 662 3808 696
rect 3842 682 3957 696
rect 3991 682 4130 716
rect 4164 715 4340 716
rect 4164 682 4278 715
rect 3842 681 4278 682
rect 4312 681 4340 715
rect 3842 662 4340 681
rect 3780 626 4340 662
rect 3780 606 3957 626
rect 3780 572 3808 606
rect 3842 592 3957 606
rect 3991 592 4130 626
rect 4164 625 4340 626
rect 4164 592 4278 625
rect 3842 591 4278 592
rect 4312 591 4340 625
rect 3842 572 4340 591
rect 3780 536 4340 572
rect 3780 516 3957 536
rect 3780 482 3808 516
rect 3842 502 3957 516
rect 3991 502 4130 536
rect 4164 535 4340 536
rect 4164 502 4278 535
rect 3842 501 4278 502
rect 4312 501 4340 535
rect 3842 482 4340 501
rect 3780 446 4340 482
rect 3780 426 3957 446
rect 3780 392 3808 426
rect 3842 412 3957 426
rect 3991 412 4130 446
rect 4164 445 4340 446
rect 4164 412 4278 445
rect 3842 411 4278 412
rect 4312 411 4340 445
rect 3842 392 4340 411
rect 3780 356 4340 392
rect 3780 336 3957 356
rect 2482 302 2980 321
rect 2420 270 2980 302
rect 3780 302 3808 336
rect 3842 322 3957 336
rect 3991 322 4130 356
rect 4164 355 4340 356
rect 4164 322 4278 355
rect 3842 321 4278 322
rect 4312 321 4340 355
rect 4393 958 5087 1017
rect 4393 924 4454 958
rect 4488 930 4544 958
rect 4578 930 4634 958
rect 4668 930 4724 958
rect 4500 924 4544 930
rect 4600 924 4634 930
rect 4700 924 4724 930
rect 4758 930 4814 958
rect 4758 924 4766 930
rect 4393 896 4466 924
rect 4500 896 4566 924
rect 4600 896 4666 924
rect 4700 896 4766 924
rect 4800 924 4814 930
rect 4848 930 4904 958
rect 4848 924 4866 930
rect 4800 896 4866 924
rect 4900 924 4904 930
rect 4938 930 4994 958
rect 4938 924 4966 930
rect 5028 924 5087 958
rect 4900 896 4966 924
rect 5000 896 5087 924
rect 4393 868 5087 896
rect 4393 834 4454 868
rect 4488 834 4544 868
rect 4578 834 4634 868
rect 4668 834 4724 868
rect 4758 834 4814 868
rect 4848 834 4904 868
rect 4938 834 4994 868
rect 5028 834 5087 868
rect 4393 830 5087 834
rect 4393 796 4466 830
rect 4500 796 4566 830
rect 4600 796 4666 830
rect 4700 796 4766 830
rect 4800 796 4866 830
rect 4900 796 4966 830
rect 5000 796 5087 830
rect 4393 778 5087 796
rect 4393 744 4454 778
rect 4488 744 4544 778
rect 4578 744 4634 778
rect 4668 744 4724 778
rect 4758 744 4814 778
rect 4848 744 4904 778
rect 4938 744 4994 778
rect 5028 744 5087 778
rect 4393 730 5087 744
rect 4393 696 4466 730
rect 4500 696 4566 730
rect 4600 696 4666 730
rect 4700 696 4766 730
rect 4800 696 4866 730
rect 4900 696 4966 730
rect 5000 696 5087 730
rect 4393 688 5087 696
rect 4393 654 4454 688
rect 4488 654 4544 688
rect 4578 654 4634 688
rect 4668 654 4724 688
rect 4758 654 4814 688
rect 4848 654 4904 688
rect 4938 654 4994 688
rect 5028 654 5087 688
rect 4393 630 5087 654
rect 4393 598 4466 630
rect 4500 598 4566 630
rect 4600 598 4666 630
rect 4700 598 4766 630
rect 4393 564 4454 598
rect 4500 596 4544 598
rect 4600 596 4634 598
rect 4700 596 4724 598
rect 4488 564 4544 596
rect 4578 564 4634 596
rect 4668 564 4724 596
rect 4758 596 4766 598
rect 4800 598 4866 630
rect 4800 596 4814 598
rect 4758 564 4814 596
rect 4848 596 4866 598
rect 4900 598 4966 630
rect 5000 598 5087 630
rect 4900 596 4904 598
rect 4848 564 4904 596
rect 4938 596 4966 598
rect 4938 564 4994 596
rect 5028 564 5087 598
rect 4393 530 5087 564
rect 4393 508 4466 530
rect 4500 508 4566 530
rect 4600 508 4666 530
rect 4700 508 4766 530
rect 4393 474 4454 508
rect 4500 496 4544 508
rect 4600 496 4634 508
rect 4700 496 4724 508
rect 4488 474 4544 496
rect 4578 474 4634 496
rect 4668 474 4724 496
rect 4758 496 4766 508
rect 4800 508 4866 530
rect 4800 496 4814 508
rect 4758 474 4814 496
rect 4848 496 4866 508
rect 4900 508 4966 530
rect 5000 508 5087 530
rect 4900 496 4904 508
rect 4848 474 4904 496
rect 4938 496 4966 508
rect 4938 474 4994 496
rect 5028 474 5087 508
rect 4393 430 5087 474
rect 4393 418 4466 430
rect 4500 418 4566 430
rect 4600 418 4666 430
rect 4700 418 4766 430
rect 4393 384 4454 418
rect 4500 396 4544 418
rect 4600 396 4634 418
rect 4700 396 4724 418
rect 4488 384 4544 396
rect 4578 384 4634 396
rect 4668 384 4724 396
rect 4758 396 4766 418
rect 4800 418 4866 430
rect 4800 396 4814 418
rect 4758 384 4814 396
rect 4848 396 4866 418
rect 4900 418 4966 430
rect 5000 418 5087 430
rect 4900 396 4904 418
rect 4848 384 4904 396
rect 4938 396 4966 418
rect 4938 384 4994 396
rect 5028 384 5087 418
rect 4393 323 5087 384
rect 5140 986 5700 1022
rect 6500 1056 6677 1070
rect 6500 1022 6528 1056
rect 6562 1042 6677 1056
rect 6711 1042 6850 1076
rect 6884 1075 8037 1076
rect 6884 1042 6998 1075
rect 6562 1041 6998 1042
rect 7032 1070 8037 1075
rect 7032 1041 7060 1070
rect 6562 1022 7060 1041
rect 5140 966 5317 986
rect 5140 932 5168 966
rect 5202 952 5317 966
rect 5351 952 5490 986
rect 5524 985 5700 986
rect 5524 952 5638 985
rect 5202 951 5638 952
rect 5672 951 5700 985
rect 5202 932 5700 951
rect 5140 896 5700 932
rect 5140 876 5317 896
rect 5140 842 5168 876
rect 5202 862 5317 876
rect 5351 862 5490 896
rect 5524 895 5700 896
rect 5524 862 5638 895
rect 5202 861 5638 862
rect 5672 861 5700 895
rect 5202 842 5700 861
rect 5140 806 5700 842
rect 5140 786 5317 806
rect 5140 752 5168 786
rect 5202 772 5317 786
rect 5351 772 5490 806
rect 5524 805 5700 806
rect 5524 772 5638 805
rect 5202 771 5638 772
rect 5672 771 5700 805
rect 5202 752 5700 771
rect 5140 716 5700 752
rect 5140 696 5317 716
rect 5140 662 5168 696
rect 5202 682 5317 696
rect 5351 682 5490 716
rect 5524 715 5700 716
rect 5524 682 5638 715
rect 5202 681 5638 682
rect 5672 681 5700 715
rect 5202 662 5700 681
rect 5140 626 5700 662
rect 5140 606 5317 626
rect 5140 572 5168 606
rect 5202 592 5317 606
rect 5351 592 5490 626
rect 5524 625 5700 626
rect 5524 592 5638 625
rect 5202 591 5638 592
rect 5672 591 5700 625
rect 5202 572 5700 591
rect 5140 536 5700 572
rect 5140 516 5317 536
rect 5140 482 5168 516
rect 5202 502 5317 516
rect 5351 502 5490 536
rect 5524 535 5700 536
rect 5524 502 5638 535
rect 5202 501 5638 502
rect 5672 501 5700 535
rect 5202 482 5700 501
rect 5140 446 5700 482
rect 5140 426 5317 446
rect 5140 392 5168 426
rect 5202 412 5317 426
rect 5351 412 5490 446
rect 5524 445 5700 446
rect 5524 412 5638 445
rect 5202 411 5638 412
rect 5672 411 5700 445
rect 5202 392 5700 411
rect 5140 356 5700 392
rect 5140 336 5317 356
rect 3842 302 4340 321
rect 3780 270 4340 302
rect 5140 302 5168 336
rect 5202 322 5317 336
rect 5351 322 5490 356
rect 5524 355 5700 356
rect 5524 322 5638 355
rect 5202 321 5638 322
rect 5672 321 5700 355
rect 5753 958 6447 1017
rect 5753 924 5814 958
rect 5848 930 5904 958
rect 5938 930 5994 958
rect 6028 930 6084 958
rect 5860 924 5904 930
rect 5960 924 5994 930
rect 6060 924 6084 930
rect 6118 930 6174 958
rect 6118 924 6126 930
rect 5753 896 5826 924
rect 5860 896 5926 924
rect 5960 896 6026 924
rect 6060 896 6126 924
rect 6160 924 6174 930
rect 6208 930 6264 958
rect 6208 924 6226 930
rect 6160 896 6226 924
rect 6260 924 6264 930
rect 6298 930 6354 958
rect 6298 924 6326 930
rect 6388 924 6447 958
rect 6260 896 6326 924
rect 6360 896 6447 924
rect 5753 868 6447 896
rect 5753 834 5814 868
rect 5848 834 5904 868
rect 5938 834 5994 868
rect 6028 834 6084 868
rect 6118 834 6174 868
rect 6208 834 6264 868
rect 6298 834 6354 868
rect 6388 834 6447 868
rect 5753 830 6447 834
rect 5753 796 5826 830
rect 5860 796 5926 830
rect 5960 796 6026 830
rect 6060 796 6126 830
rect 6160 796 6226 830
rect 6260 796 6326 830
rect 6360 796 6447 830
rect 5753 778 6447 796
rect 5753 744 5814 778
rect 5848 744 5904 778
rect 5938 744 5994 778
rect 6028 744 6084 778
rect 6118 744 6174 778
rect 6208 744 6264 778
rect 6298 744 6354 778
rect 6388 744 6447 778
rect 5753 730 6447 744
rect 5753 696 5826 730
rect 5860 696 5926 730
rect 5960 696 6026 730
rect 6060 696 6126 730
rect 6160 696 6226 730
rect 6260 696 6326 730
rect 6360 696 6447 730
rect 5753 688 6447 696
rect 5753 654 5814 688
rect 5848 654 5904 688
rect 5938 654 5994 688
rect 6028 654 6084 688
rect 6118 654 6174 688
rect 6208 654 6264 688
rect 6298 654 6354 688
rect 6388 654 6447 688
rect 5753 630 6447 654
rect 5753 598 5826 630
rect 5860 598 5926 630
rect 5960 598 6026 630
rect 6060 598 6126 630
rect 5753 564 5814 598
rect 5860 596 5904 598
rect 5960 596 5994 598
rect 6060 596 6084 598
rect 5848 564 5904 596
rect 5938 564 5994 596
rect 6028 564 6084 596
rect 6118 596 6126 598
rect 6160 598 6226 630
rect 6160 596 6174 598
rect 6118 564 6174 596
rect 6208 596 6226 598
rect 6260 598 6326 630
rect 6360 598 6447 630
rect 6260 596 6264 598
rect 6208 564 6264 596
rect 6298 596 6326 598
rect 6298 564 6354 596
rect 6388 564 6447 598
rect 5753 530 6447 564
rect 5753 508 5826 530
rect 5860 508 5926 530
rect 5960 508 6026 530
rect 6060 508 6126 530
rect 5753 474 5814 508
rect 5860 496 5904 508
rect 5960 496 5994 508
rect 6060 496 6084 508
rect 5848 474 5904 496
rect 5938 474 5994 496
rect 6028 474 6084 496
rect 6118 496 6126 508
rect 6160 508 6226 530
rect 6160 496 6174 508
rect 6118 474 6174 496
rect 6208 496 6226 508
rect 6260 508 6326 530
rect 6360 508 6447 530
rect 6260 496 6264 508
rect 6208 474 6264 496
rect 6298 496 6326 508
rect 6298 474 6354 496
rect 6388 474 6447 508
rect 5753 430 6447 474
rect 5753 418 5826 430
rect 5860 418 5926 430
rect 5960 418 6026 430
rect 6060 418 6126 430
rect 5753 384 5814 418
rect 5860 396 5904 418
rect 5960 396 5994 418
rect 6060 396 6084 418
rect 5848 384 5904 396
rect 5938 384 5994 396
rect 6028 384 6084 396
rect 6118 396 6126 418
rect 6160 418 6226 430
rect 6160 396 6174 418
rect 6118 384 6174 396
rect 6208 396 6226 418
rect 6260 418 6326 430
rect 6360 418 6447 430
rect 6260 396 6264 418
rect 6208 384 6264 396
rect 6298 396 6326 418
rect 6298 384 6354 396
rect 6388 384 6447 418
rect 5753 323 6447 384
rect 6500 986 7060 1022
rect 7860 1056 8037 1070
rect 7860 1022 7888 1056
rect 7922 1042 8037 1056
rect 8071 1042 8210 1076
rect 8244 1075 9397 1076
rect 8244 1042 8358 1075
rect 7922 1041 8358 1042
rect 8392 1070 9397 1075
rect 8392 1041 8420 1070
rect 7922 1022 8420 1041
rect 6500 966 6677 986
rect 6500 932 6528 966
rect 6562 952 6677 966
rect 6711 952 6850 986
rect 6884 985 7060 986
rect 6884 952 6998 985
rect 6562 951 6998 952
rect 7032 951 7060 985
rect 6562 932 7060 951
rect 6500 896 7060 932
rect 6500 876 6677 896
rect 6500 842 6528 876
rect 6562 862 6677 876
rect 6711 862 6850 896
rect 6884 895 7060 896
rect 6884 862 6998 895
rect 6562 861 6998 862
rect 7032 861 7060 895
rect 6562 842 7060 861
rect 6500 806 7060 842
rect 6500 786 6677 806
rect 6500 752 6528 786
rect 6562 772 6677 786
rect 6711 772 6850 806
rect 6884 805 7060 806
rect 6884 772 6998 805
rect 6562 771 6998 772
rect 7032 771 7060 805
rect 6562 752 7060 771
rect 6500 716 7060 752
rect 6500 696 6677 716
rect 6500 662 6528 696
rect 6562 682 6677 696
rect 6711 682 6850 716
rect 6884 715 7060 716
rect 6884 682 6998 715
rect 6562 681 6998 682
rect 7032 681 7060 715
rect 6562 662 7060 681
rect 6500 626 7060 662
rect 6500 606 6677 626
rect 6500 572 6528 606
rect 6562 592 6677 606
rect 6711 592 6850 626
rect 6884 625 7060 626
rect 6884 592 6998 625
rect 6562 591 6998 592
rect 7032 591 7060 625
rect 6562 572 7060 591
rect 6500 536 7060 572
rect 6500 516 6677 536
rect 6500 482 6528 516
rect 6562 502 6677 516
rect 6711 502 6850 536
rect 6884 535 7060 536
rect 6884 502 6998 535
rect 6562 501 6998 502
rect 7032 501 7060 535
rect 6562 482 7060 501
rect 6500 446 7060 482
rect 6500 426 6677 446
rect 6500 392 6528 426
rect 6562 412 6677 426
rect 6711 412 6850 446
rect 6884 445 7060 446
rect 6884 412 6998 445
rect 6562 411 6998 412
rect 7032 411 7060 445
rect 6562 392 7060 411
rect 6500 356 7060 392
rect 6500 336 6677 356
rect 5202 302 5700 321
rect 5140 270 5700 302
rect 6500 302 6528 336
rect 6562 322 6677 336
rect 6711 322 6850 356
rect 6884 355 7060 356
rect 6884 322 6998 355
rect 6562 321 6998 322
rect 7032 321 7060 355
rect 7113 958 7807 1017
rect 7113 924 7174 958
rect 7208 930 7264 958
rect 7298 930 7354 958
rect 7388 930 7444 958
rect 7220 924 7264 930
rect 7320 924 7354 930
rect 7420 924 7444 930
rect 7478 930 7534 958
rect 7478 924 7486 930
rect 7113 896 7186 924
rect 7220 896 7286 924
rect 7320 896 7386 924
rect 7420 896 7486 924
rect 7520 924 7534 930
rect 7568 930 7624 958
rect 7568 924 7586 930
rect 7520 896 7586 924
rect 7620 924 7624 930
rect 7658 930 7714 958
rect 7658 924 7686 930
rect 7748 924 7807 958
rect 7620 896 7686 924
rect 7720 896 7807 924
rect 7113 868 7807 896
rect 7113 834 7174 868
rect 7208 834 7264 868
rect 7298 834 7354 868
rect 7388 834 7444 868
rect 7478 834 7534 868
rect 7568 834 7624 868
rect 7658 834 7714 868
rect 7748 834 7807 868
rect 7113 830 7807 834
rect 7113 796 7186 830
rect 7220 796 7286 830
rect 7320 796 7386 830
rect 7420 796 7486 830
rect 7520 796 7586 830
rect 7620 796 7686 830
rect 7720 796 7807 830
rect 7113 778 7807 796
rect 7113 744 7174 778
rect 7208 744 7264 778
rect 7298 744 7354 778
rect 7388 744 7444 778
rect 7478 744 7534 778
rect 7568 744 7624 778
rect 7658 744 7714 778
rect 7748 744 7807 778
rect 7113 730 7807 744
rect 7113 696 7186 730
rect 7220 696 7286 730
rect 7320 696 7386 730
rect 7420 696 7486 730
rect 7520 696 7586 730
rect 7620 696 7686 730
rect 7720 696 7807 730
rect 7113 688 7807 696
rect 7113 654 7174 688
rect 7208 654 7264 688
rect 7298 654 7354 688
rect 7388 654 7444 688
rect 7478 654 7534 688
rect 7568 654 7624 688
rect 7658 654 7714 688
rect 7748 654 7807 688
rect 7113 630 7807 654
rect 7113 598 7186 630
rect 7220 598 7286 630
rect 7320 598 7386 630
rect 7420 598 7486 630
rect 7113 564 7174 598
rect 7220 596 7264 598
rect 7320 596 7354 598
rect 7420 596 7444 598
rect 7208 564 7264 596
rect 7298 564 7354 596
rect 7388 564 7444 596
rect 7478 596 7486 598
rect 7520 598 7586 630
rect 7520 596 7534 598
rect 7478 564 7534 596
rect 7568 596 7586 598
rect 7620 598 7686 630
rect 7720 598 7807 630
rect 7620 596 7624 598
rect 7568 564 7624 596
rect 7658 596 7686 598
rect 7658 564 7714 596
rect 7748 564 7807 598
rect 7113 530 7807 564
rect 7113 508 7186 530
rect 7220 508 7286 530
rect 7320 508 7386 530
rect 7420 508 7486 530
rect 7113 474 7174 508
rect 7220 496 7264 508
rect 7320 496 7354 508
rect 7420 496 7444 508
rect 7208 474 7264 496
rect 7298 474 7354 496
rect 7388 474 7444 496
rect 7478 496 7486 508
rect 7520 508 7586 530
rect 7520 496 7534 508
rect 7478 474 7534 496
rect 7568 496 7586 508
rect 7620 508 7686 530
rect 7720 508 7807 530
rect 7620 496 7624 508
rect 7568 474 7624 496
rect 7658 496 7686 508
rect 7658 474 7714 496
rect 7748 474 7807 508
rect 7113 430 7807 474
rect 7113 418 7186 430
rect 7220 418 7286 430
rect 7320 418 7386 430
rect 7420 418 7486 430
rect 7113 384 7174 418
rect 7220 396 7264 418
rect 7320 396 7354 418
rect 7420 396 7444 418
rect 7208 384 7264 396
rect 7298 384 7354 396
rect 7388 384 7444 396
rect 7478 396 7486 418
rect 7520 418 7586 430
rect 7520 396 7534 418
rect 7478 384 7534 396
rect 7568 396 7586 418
rect 7620 418 7686 430
rect 7720 418 7807 430
rect 7620 396 7624 418
rect 7568 384 7624 396
rect 7658 396 7686 418
rect 7658 384 7714 396
rect 7748 384 7807 418
rect 7113 323 7807 384
rect 7860 986 8420 1022
rect 9220 1056 9397 1070
rect 9220 1022 9248 1056
rect 9282 1042 9397 1056
rect 9431 1042 9470 1076
rect 9282 1022 9470 1042
rect 7860 966 8037 986
rect 7860 932 7888 966
rect 7922 952 8037 966
rect 8071 952 8210 986
rect 8244 985 8420 986
rect 8244 952 8358 985
rect 7922 951 8358 952
rect 8392 951 8420 985
rect 7922 932 8420 951
rect 7860 896 8420 932
rect 7860 876 8037 896
rect 7860 842 7888 876
rect 7922 862 8037 876
rect 8071 862 8210 896
rect 8244 895 8420 896
rect 8244 862 8358 895
rect 7922 861 8358 862
rect 8392 861 8420 895
rect 7922 842 8420 861
rect 7860 806 8420 842
rect 7860 786 8037 806
rect 7860 752 7888 786
rect 7922 772 8037 786
rect 8071 772 8210 806
rect 8244 805 8420 806
rect 8244 772 8358 805
rect 7922 771 8358 772
rect 8392 771 8420 805
rect 7922 752 8420 771
rect 7860 716 8420 752
rect 7860 696 8037 716
rect 7860 662 7888 696
rect 7922 682 8037 696
rect 8071 682 8210 716
rect 8244 715 8420 716
rect 8244 682 8358 715
rect 7922 681 8358 682
rect 8392 681 8420 715
rect 7922 662 8420 681
rect 7860 626 8420 662
rect 7860 606 8037 626
rect 7860 572 7888 606
rect 7922 592 8037 606
rect 8071 592 8210 626
rect 8244 625 8420 626
rect 8244 592 8358 625
rect 7922 591 8358 592
rect 8392 591 8420 625
rect 7922 572 8420 591
rect 7860 536 8420 572
rect 7860 516 8037 536
rect 7860 482 7888 516
rect 7922 502 8037 516
rect 8071 502 8210 536
rect 8244 535 8420 536
rect 8244 502 8358 535
rect 7922 501 8358 502
rect 8392 501 8420 535
rect 7922 482 8420 501
rect 7860 446 8420 482
rect 7860 426 8037 446
rect 7860 392 7888 426
rect 7922 412 8037 426
rect 8071 412 8210 446
rect 8244 445 8420 446
rect 8244 412 8358 445
rect 7922 411 8358 412
rect 8392 411 8420 445
rect 7922 392 8420 411
rect 7860 356 8420 392
rect 7860 336 8037 356
rect 6562 302 7060 321
rect 6500 270 7060 302
rect 7860 302 7888 336
rect 7922 322 8037 336
rect 8071 322 8210 356
rect 8244 355 8420 356
rect 8244 322 8358 355
rect 7922 321 8358 322
rect 8392 321 8420 355
rect 8473 958 9167 1017
rect 8473 924 8534 958
rect 8568 930 8624 958
rect 8658 930 8714 958
rect 8748 930 8804 958
rect 8580 924 8624 930
rect 8680 924 8714 930
rect 8780 924 8804 930
rect 8838 930 8894 958
rect 8838 924 8846 930
rect 8473 896 8546 924
rect 8580 896 8646 924
rect 8680 896 8746 924
rect 8780 896 8846 924
rect 8880 924 8894 930
rect 8928 930 8984 958
rect 8928 924 8946 930
rect 8880 896 8946 924
rect 8980 924 8984 930
rect 9018 930 9074 958
rect 9018 924 9046 930
rect 9108 924 9167 958
rect 8980 896 9046 924
rect 9080 896 9167 924
rect 8473 868 9167 896
rect 8473 834 8534 868
rect 8568 834 8624 868
rect 8658 834 8714 868
rect 8748 834 8804 868
rect 8838 834 8894 868
rect 8928 834 8984 868
rect 9018 834 9074 868
rect 9108 834 9167 868
rect 8473 830 9167 834
rect 8473 796 8546 830
rect 8580 796 8646 830
rect 8680 796 8746 830
rect 8780 796 8846 830
rect 8880 796 8946 830
rect 8980 796 9046 830
rect 9080 796 9167 830
rect 8473 778 9167 796
rect 8473 744 8534 778
rect 8568 744 8624 778
rect 8658 744 8714 778
rect 8748 744 8804 778
rect 8838 744 8894 778
rect 8928 744 8984 778
rect 9018 744 9074 778
rect 9108 744 9167 778
rect 8473 730 9167 744
rect 8473 696 8546 730
rect 8580 696 8646 730
rect 8680 696 8746 730
rect 8780 696 8846 730
rect 8880 696 8946 730
rect 8980 696 9046 730
rect 9080 696 9167 730
rect 8473 688 9167 696
rect 8473 654 8534 688
rect 8568 654 8624 688
rect 8658 654 8714 688
rect 8748 654 8804 688
rect 8838 654 8894 688
rect 8928 654 8984 688
rect 9018 654 9074 688
rect 9108 654 9167 688
rect 8473 630 9167 654
rect 8473 598 8546 630
rect 8580 598 8646 630
rect 8680 598 8746 630
rect 8780 598 8846 630
rect 8473 564 8534 598
rect 8580 596 8624 598
rect 8680 596 8714 598
rect 8780 596 8804 598
rect 8568 564 8624 596
rect 8658 564 8714 596
rect 8748 564 8804 596
rect 8838 596 8846 598
rect 8880 598 8946 630
rect 8880 596 8894 598
rect 8838 564 8894 596
rect 8928 596 8946 598
rect 8980 598 9046 630
rect 9080 598 9167 630
rect 8980 596 8984 598
rect 8928 564 8984 596
rect 9018 596 9046 598
rect 9018 564 9074 596
rect 9108 564 9167 598
rect 8473 530 9167 564
rect 8473 508 8546 530
rect 8580 508 8646 530
rect 8680 508 8746 530
rect 8780 508 8846 530
rect 8473 474 8534 508
rect 8580 496 8624 508
rect 8680 496 8714 508
rect 8780 496 8804 508
rect 8568 474 8624 496
rect 8658 474 8714 496
rect 8748 474 8804 496
rect 8838 496 8846 508
rect 8880 508 8946 530
rect 8880 496 8894 508
rect 8838 474 8894 496
rect 8928 496 8946 508
rect 8980 508 9046 530
rect 9080 508 9167 530
rect 8980 496 8984 508
rect 8928 474 8984 496
rect 9018 496 9046 508
rect 9018 474 9074 496
rect 9108 474 9167 508
rect 8473 430 9167 474
rect 8473 418 8546 430
rect 8580 418 8646 430
rect 8680 418 8746 430
rect 8780 418 8846 430
rect 8473 384 8534 418
rect 8580 396 8624 418
rect 8680 396 8714 418
rect 8780 396 8804 418
rect 8568 384 8624 396
rect 8658 384 8714 396
rect 8748 384 8804 396
rect 8838 396 8846 418
rect 8880 418 8946 430
rect 8880 396 8894 418
rect 8838 384 8894 396
rect 8928 396 8946 418
rect 8980 418 9046 430
rect 9080 418 9167 430
rect 8980 396 8984 418
rect 8928 384 8984 396
rect 9018 396 9046 418
rect 9018 384 9074 396
rect 9108 384 9167 418
rect 8473 323 9167 384
rect 9220 986 9470 1022
rect 9220 966 9397 986
rect 9220 932 9248 966
rect 9282 952 9397 966
rect 9431 952 9470 986
rect 9282 932 9470 952
rect 9220 896 9470 932
rect 9220 876 9397 896
rect 9220 842 9248 876
rect 9282 862 9397 876
rect 9431 862 9470 896
rect 9282 842 9470 862
rect 9220 806 9470 842
rect 9220 786 9397 806
rect 9220 752 9248 786
rect 9282 772 9397 786
rect 9431 772 9470 806
rect 9282 752 9470 772
rect 9220 716 9470 752
rect 9220 696 9397 716
rect 9220 662 9248 696
rect 9282 682 9397 696
rect 9431 682 9470 716
rect 9282 662 9470 682
rect 9220 626 9470 662
rect 9220 606 9397 626
rect 9220 572 9248 606
rect 9282 592 9397 606
rect 9431 592 9470 626
rect 9282 572 9470 592
rect 9220 536 9470 572
rect 9220 516 9397 536
rect 9220 482 9248 516
rect 9282 502 9397 516
rect 9431 502 9470 536
rect 9282 482 9470 502
rect 9220 446 9470 482
rect 9220 426 9397 446
rect 9220 392 9248 426
rect 9282 412 9397 426
rect 9431 412 9470 446
rect 9282 392 9470 412
rect 9220 356 9470 392
rect 9220 336 9397 356
rect 7922 302 8420 321
rect 7860 270 8420 302
rect 9220 302 9248 336
rect 9282 322 9397 336
rect 9431 322 9470 356
rect 9282 302 9470 322
rect 9220 270 9470 302
rect 10 266 9470 270
rect 10 232 1410 266
rect 1444 242 2597 266
rect 1444 232 1636 242
rect 10 208 1636 232
rect 1670 208 1726 242
rect 1760 208 1816 242
rect 1850 208 1906 242
rect 1940 208 1996 242
rect 2030 208 2086 242
rect 2120 208 2176 242
rect 2210 208 2266 242
rect 2300 208 2356 242
rect 2390 232 2597 242
rect 2631 232 2770 266
rect 2804 242 3957 266
rect 2804 232 2996 242
rect 2390 208 2996 232
rect 3030 208 3086 242
rect 3120 208 3176 242
rect 3210 208 3266 242
rect 3300 208 3356 242
rect 3390 208 3446 242
rect 3480 208 3536 242
rect 3570 208 3626 242
rect 3660 208 3716 242
rect 3750 232 3957 242
rect 3991 232 4130 266
rect 4164 242 5317 266
rect 4164 232 4356 242
rect 3750 208 4356 232
rect 4390 208 4446 242
rect 4480 208 4536 242
rect 4570 208 4626 242
rect 4660 208 4716 242
rect 4750 208 4806 242
rect 4840 208 4896 242
rect 4930 208 4986 242
rect 5020 208 5076 242
rect 5110 232 5317 242
rect 5351 232 5490 266
rect 5524 242 6677 266
rect 5524 232 5716 242
rect 5110 208 5716 232
rect 5750 208 5806 242
rect 5840 208 5896 242
rect 5930 208 5986 242
rect 6020 208 6076 242
rect 6110 208 6166 242
rect 6200 208 6256 242
rect 6290 208 6346 242
rect 6380 208 6436 242
rect 6470 232 6677 242
rect 6711 232 6850 266
rect 6884 242 8037 266
rect 6884 232 7076 242
rect 6470 208 7076 232
rect 7110 208 7166 242
rect 7200 208 7256 242
rect 7290 208 7346 242
rect 7380 208 7436 242
rect 7470 208 7526 242
rect 7560 208 7616 242
rect 7650 208 7706 242
rect 7740 208 7796 242
rect 7830 232 8037 242
rect 8071 232 8210 266
rect 8244 242 9397 266
rect 8244 232 8436 242
rect 7830 208 8436 232
rect 8470 208 8526 242
rect 8560 208 8616 242
rect 8650 208 8706 242
rect 8740 208 8796 242
rect 8830 208 8886 242
rect 8920 208 8976 242
rect 9010 208 9066 242
rect 9100 208 9156 242
rect 9190 232 9397 242
rect 9431 232 9470 266
rect 9190 208 9470 232
rect 10 176 9470 208
rect 10 142 1410 176
rect 1444 142 2597 176
rect 2631 142 2770 176
rect 2804 142 3957 176
rect 3991 142 4130 176
rect 4164 142 5317 176
rect 5351 142 5490 176
rect 5524 142 6677 176
rect 6711 142 6850 176
rect 6884 142 8037 176
rect 8071 142 8210 176
rect 8244 142 9397 176
rect 9431 142 9470 176
rect 10 92 9470 142
rect 10 90 1506 92
rect 1540 90 1596 92
rect 1630 90 1686 92
rect 1720 90 1776 92
rect 1810 90 1866 92
rect 1900 90 1956 92
rect 1990 90 2046 92
rect 2080 90 2136 92
rect 2170 90 2226 92
rect 2260 90 2316 92
rect 2350 90 2406 92
rect 2440 90 2496 92
rect 2530 90 2866 92
rect 2900 90 2956 92
rect 2990 90 3046 92
rect 3080 90 3136 92
rect 3170 90 3226 92
rect 3260 90 3316 92
rect 3350 90 3406 92
rect 3440 90 3496 92
rect 3530 90 3586 92
rect 3620 90 3676 92
rect 3710 90 3766 92
rect 3800 90 3856 92
rect 3890 90 4226 92
rect 4260 90 4316 92
rect 4350 90 4406 92
rect 4440 90 4496 92
rect 4530 90 4586 92
rect 4620 90 4676 92
rect 4710 90 4766 92
rect 4800 90 4856 92
rect 4890 90 4946 92
rect 4980 90 5036 92
rect 5070 90 5126 92
rect 5160 90 5216 92
rect 5250 90 5586 92
rect 5620 90 5676 92
rect 5710 90 5766 92
rect 5800 90 5856 92
rect 5890 90 5946 92
rect 5980 90 6036 92
rect 6070 90 6126 92
rect 6160 90 6216 92
rect 6250 90 6306 92
rect 6340 90 6396 92
rect 6430 90 6486 92
rect 6520 90 6576 92
rect 6610 90 6946 92
rect 6980 90 7036 92
rect 7070 90 7126 92
rect 7160 90 7216 92
rect 7250 90 7306 92
rect 7340 90 7396 92
rect 7430 90 7486 92
rect 7520 90 7576 92
rect 7610 90 7666 92
rect 7700 90 7756 92
rect 7790 90 7846 92
rect 7880 90 7936 92
rect 7970 90 8306 92
rect 8340 90 8396 92
rect 8430 90 8486 92
rect 8520 90 8576 92
rect 8610 90 8666 92
rect 8700 90 8756 92
rect 8790 90 8846 92
rect 8880 90 8936 92
rect 8970 90 9026 92
rect 9060 90 9116 92
rect 9150 90 9206 92
rect 9240 90 9296 92
rect 9330 90 9470 92
rect 10 50 40 90
rect 80 50 140 90
rect 180 50 240 90
rect 280 50 330 90
rect 370 50 410 90
rect 450 50 500 90
rect 540 50 590 90
rect 630 50 680 90
rect 720 50 770 90
rect 810 50 860 90
rect 900 50 950 90
rect 990 50 1040 90
rect 1080 50 1130 90
rect 1170 50 1230 90
rect 1270 50 1320 90
rect 1360 50 1420 90
rect 1460 50 1500 90
rect 1540 50 1590 90
rect 1630 50 1680 90
rect 1720 50 1770 90
rect 1810 50 1860 90
rect 1900 50 1950 90
rect 1990 50 2040 90
rect 2080 50 2130 90
rect 2170 50 2220 90
rect 2260 50 2310 90
rect 2350 50 2400 90
rect 2440 50 2490 90
rect 2530 50 2590 90
rect 2630 50 2680 90
rect 2720 50 2770 90
rect 2810 50 2860 90
rect 2900 50 2950 90
rect 2990 50 3040 90
rect 3080 50 3130 90
rect 3170 50 3220 90
rect 3260 50 3310 90
rect 3350 50 3400 90
rect 3440 50 3490 90
rect 3530 50 3580 90
rect 3620 50 3670 90
rect 3710 50 3760 90
rect 3800 50 3850 90
rect 3890 50 3950 90
rect 3990 50 4040 90
rect 4080 50 4130 90
rect 4170 50 4220 90
rect 4260 50 4310 90
rect 4350 50 4400 90
rect 4440 50 4490 90
rect 4530 50 4580 90
rect 4620 50 4670 90
rect 4710 50 4760 90
rect 4800 50 4850 90
rect 4890 50 4940 90
rect 4980 50 5030 90
rect 5070 50 5120 90
rect 5160 50 5210 90
rect 5250 50 5310 90
rect 5350 50 5400 90
rect 5440 50 5490 90
rect 5530 50 5580 90
rect 5620 50 5670 90
rect 5710 50 5760 90
rect 5800 50 5850 90
rect 5890 50 5940 90
rect 5980 50 6030 90
rect 6070 50 6120 90
rect 6160 50 6210 90
rect 6250 50 6300 90
rect 6340 50 6390 90
rect 6430 50 6480 90
rect 6520 50 6570 90
rect 6610 50 6660 90
rect 6700 50 6760 90
rect 6800 50 6850 90
rect 6890 50 6940 90
rect 6980 50 7030 90
rect 7070 50 7120 90
rect 7160 50 7210 90
rect 7250 50 7300 90
rect 7340 50 7390 90
rect 7430 50 7480 90
rect 7520 50 7570 90
rect 7610 50 7660 90
rect 7700 50 7750 90
rect 7790 50 7840 90
rect 7880 50 7930 90
rect 7970 50 8020 90
rect 8060 50 8120 90
rect 8160 50 8210 90
rect 8250 50 8300 90
rect 8340 50 8390 90
rect 8430 50 8480 90
rect 8520 50 8570 90
rect 8610 50 8660 90
rect 8700 50 8750 90
rect 8790 50 8840 90
rect 8880 50 8930 90
rect 8970 50 9020 90
rect 9060 50 9110 90
rect 9150 50 9200 90
rect 9240 50 9290 90
rect 9330 50 9390 90
rect 9430 50 9470 90
rect 10 20 9470 50
<< viali >>
rect 4640 5510 4680 5550
rect 5040 5510 5080 5550
rect 5440 5510 5480 5550
rect 5840 5510 5880 5550
rect 6240 5510 6280 5550
rect 6440 5510 6480 5550
rect 6640 5510 6680 5550
rect 7040 5510 7080 5550
rect 7440 5510 7480 5550
rect 7840 5510 7880 5550
rect 8240 5510 8280 5550
rect 1910 4990 1950 5030
rect 4840 4570 4880 4610
rect 5240 4480 5280 4520
rect 6240 4570 6280 4610
rect 6040 4480 6080 4520
rect 6640 4570 6680 4610
rect 6840 4570 6880 4610
rect 7640 4570 7680 4610
rect 8160 4570 8200 4610
rect 8040 4480 8080 4520
rect 3810 4400 3850 4440
rect 3900 4400 3940 4440
rect 3990 4400 4030 4440
rect 4080 4400 4120 4440
rect 4170 4400 4210 4440
rect 5640 4390 5680 4430
rect 6440 4390 6480 4430
rect 7240 4390 7280 4430
rect 8770 4370 8810 4410
rect 5240 4270 5280 4310
rect 5640 4270 5680 4310
rect 6040 4270 6080 4310
rect 6240 4270 6280 4310
rect 6440 4270 6480 4310
rect 6640 4270 6680 4310
rect 6840 4270 6880 4310
rect 7240 4270 7280 4310
rect 7640 4270 7680 4310
rect 9190 4270 9230 4310
rect 1910 3970 1950 4010
rect 5840 3730 5880 3770
rect 6480 3730 6520 3770
rect 7040 3730 7080 3770
rect 5440 3640 5480 3680
rect 6350 3640 6390 3680
rect 7440 3640 7480 3680
rect 6480 3550 6520 3590
rect 5840 3460 5880 3500
rect 7040 3460 7080 3500
rect 3810 3380 3850 3420
rect 3900 3380 3940 3420
rect 3990 3380 4030 3420
rect 4080 3380 4120 3420
rect 4170 3380 4210 3420
rect 6120 3370 6160 3410
rect 6240 3370 6280 3410
rect 6640 3370 6680 3410
rect 6760 3370 6800 3410
rect 8990 3700 9030 3740
rect 8880 3370 8920 3410
rect 1910 3020 1950 3060
rect 3810 3020 3850 3060
rect 3900 3020 3940 3060
rect 3990 3020 4030 3060
rect 4080 3020 4120 3060
rect 4170 3020 4210 3060
rect 5840 3030 5880 3070
rect 7040 3030 7080 3070
rect 5640 2940 5680 2980
rect 6040 2940 6080 2980
rect 6440 2940 6480 2980
rect 6840 2940 6880 2980
rect 7240 2940 7280 2980
rect 7400 2820 7440 2860
rect 1910 2430 1950 2470
rect 6360 1880 6400 1920
rect 6440 1880 6480 1920
rect 6520 1880 6560 1920
rect 7460 1760 7500 1800
rect 1320 1600 1360 1640
rect 7610 1590 7650 1630
rect 1746 924 1768 930
rect 1768 924 1780 930
rect 1846 924 1858 930
rect 1858 924 1880 930
rect 1946 924 1948 930
rect 1948 924 1980 930
rect 1746 896 1780 924
rect 1846 896 1880 924
rect 1946 896 1980 924
rect 2046 896 2080 930
rect 2146 896 2180 930
rect 2246 924 2274 930
rect 2274 924 2280 930
rect 2246 896 2280 924
rect 1746 796 1780 830
rect 1846 796 1880 830
rect 1946 796 1980 830
rect 2046 796 2080 830
rect 2146 796 2180 830
rect 2246 796 2280 830
rect 1746 696 1780 730
rect 1846 696 1880 730
rect 1946 696 1980 730
rect 2046 696 2080 730
rect 2146 696 2180 730
rect 2246 696 2280 730
rect 1746 598 1780 630
rect 1846 598 1880 630
rect 1946 598 1980 630
rect 1746 596 1768 598
rect 1768 596 1780 598
rect 1846 596 1858 598
rect 1858 596 1880 598
rect 1946 596 1948 598
rect 1948 596 1980 598
rect 2046 596 2080 630
rect 2146 596 2180 630
rect 2246 598 2280 630
rect 2246 596 2274 598
rect 2274 596 2280 598
rect 1746 508 1780 530
rect 1846 508 1880 530
rect 1946 508 1980 530
rect 1746 496 1768 508
rect 1768 496 1780 508
rect 1846 496 1858 508
rect 1858 496 1880 508
rect 1946 496 1948 508
rect 1948 496 1980 508
rect 2046 496 2080 530
rect 2146 496 2180 530
rect 2246 508 2280 530
rect 2246 496 2274 508
rect 2274 496 2280 508
rect 1746 418 1780 430
rect 1846 418 1880 430
rect 1946 418 1980 430
rect 1746 396 1768 418
rect 1768 396 1780 418
rect 1846 396 1858 418
rect 1858 396 1880 418
rect 1946 396 1948 418
rect 1948 396 1980 418
rect 2046 396 2080 430
rect 2146 396 2180 430
rect 2246 418 2280 430
rect 2246 396 2274 418
rect 2274 396 2280 418
rect 3106 924 3128 930
rect 3128 924 3140 930
rect 3206 924 3218 930
rect 3218 924 3240 930
rect 3306 924 3308 930
rect 3308 924 3340 930
rect 3106 896 3140 924
rect 3206 896 3240 924
rect 3306 896 3340 924
rect 3406 896 3440 930
rect 3506 896 3540 930
rect 3606 924 3634 930
rect 3634 924 3640 930
rect 3606 896 3640 924
rect 3106 796 3140 830
rect 3206 796 3240 830
rect 3306 796 3340 830
rect 3406 796 3440 830
rect 3506 796 3540 830
rect 3606 796 3640 830
rect 3106 696 3140 730
rect 3206 696 3240 730
rect 3306 696 3340 730
rect 3406 696 3440 730
rect 3506 696 3540 730
rect 3606 696 3640 730
rect 3106 598 3140 630
rect 3206 598 3240 630
rect 3306 598 3340 630
rect 3106 596 3128 598
rect 3128 596 3140 598
rect 3206 596 3218 598
rect 3218 596 3240 598
rect 3306 596 3308 598
rect 3308 596 3340 598
rect 3406 596 3440 630
rect 3506 596 3540 630
rect 3606 598 3640 630
rect 3606 596 3634 598
rect 3634 596 3640 598
rect 3106 508 3140 530
rect 3206 508 3240 530
rect 3306 508 3340 530
rect 3106 496 3128 508
rect 3128 496 3140 508
rect 3206 496 3218 508
rect 3218 496 3240 508
rect 3306 496 3308 508
rect 3308 496 3340 508
rect 3406 496 3440 530
rect 3506 496 3540 530
rect 3606 508 3640 530
rect 3606 496 3634 508
rect 3634 496 3640 508
rect 3106 418 3140 430
rect 3206 418 3240 430
rect 3306 418 3340 430
rect 3106 396 3128 418
rect 3128 396 3140 418
rect 3206 396 3218 418
rect 3218 396 3240 418
rect 3306 396 3308 418
rect 3308 396 3340 418
rect 3406 396 3440 430
rect 3506 396 3540 430
rect 3606 418 3640 430
rect 3606 396 3634 418
rect 3634 396 3640 418
rect 4466 924 4488 930
rect 4488 924 4500 930
rect 4566 924 4578 930
rect 4578 924 4600 930
rect 4666 924 4668 930
rect 4668 924 4700 930
rect 4466 896 4500 924
rect 4566 896 4600 924
rect 4666 896 4700 924
rect 4766 896 4800 930
rect 4866 896 4900 930
rect 4966 924 4994 930
rect 4994 924 5000 930
rect 4966 896 5000 924
rect 4466 796 4500 830
rect 4566 796 4600 830
rect 4666 796 4700 830
rect 4766 796 4800 830
rect 4866 796 4900 830
rect 4966 796 5000 830
rect 4466 696 4500 730
rect 4566 696 4600 730
rect 4666 696 4700 730
rect 4766 696 4800 730
rect 4866 696 4900 730
rect 4966 696 5000 730
rect 4466 598 4500 630
rect 4566 598 4600 630
rect 4666 598 4700 630
rect 4466 596 4488 598
rect 4488 596 4500 598
rect 4566 596 4578 598
rect 4578 596 4600 598
rect 4666 596 4668 598
rect 4668 596 4700 598
rect 4766 596 4800 630
rect 4866 596 4900 630
rect 4966 598 5000 630
rect 4966 596 4994 598
rect 4994 596 5000 598
rect 4466 508 4500 530
rect 4566 508 4600 530
rect 4666 508 4700 530
rect 4466 496 4488 508
rect 4488 496 4500 508
rect 4566 496 4578 508
rect 4578 496 4600 508
rect 4666 496 4668 508
rect 4668 496 4700 508
rect 4766 496 4800 530
rect 4866 496 4900 530
rect 4966 508 5000 530
rect 4966 496 4994 508
rect 4994 496 5000 508
rect 4466 418 4500 430
rect 4566 418 4600 430
rect 4666 418 4700 430
rect 4466 396 4488 418
rect 4488 396 4500 418
rect 4566 396 4578 418
rect 4578 396 4600 418
rect 4666 396 4668 418
rect 4668 396 4700 418
rect 4766 396 4800 430
rect 4866 396 4900 430
rect 4966 418 5000 430
rect 4966 396 4994 418
rect 4994 396 5000 418
rect 5826 924 5848 930
rect 5848 924 5860 930
rect 5926 924 5938 930
rect 5938 924 5960 930
rect 6026 924 6028 930
rect 6028 924 6060 930
rect 5826 896 5860 924
rect 5926 896 5960 924
rect 6026 896 6060 924
rect 6126 896 6160 930
rect 6226 896 6260 930
rect 6326 924 6354 930
rect 6354 924 6360 930
rect 6326 896 6360 924
rect 5826 796 5860 830
rect 5926 796 5960 830
rect 6026 796 6060 830
rect 6126 796 6160 830
rect 6226 796 6260 830
rect 6326 796 6360 830
rect 5826 696 5860 730
rect 5926 696 5960 730
rect 6026 696 6060 730
rect 6126 696 6160 730
rect 6226 696 6260 730
rect 6326 696 6360 730
rect 5826 598 5860 630
rect 5926 598 5960 630
rect 6026 598 6060 630
rect 5826 596 5848 598
rect 5848 596 5860 598
rect 5926 596 5938 598
rect 5938 596 5960 598
rect 6026 596 6028 598
rect 6028 596 6060 598
rect 6126 596 6160 630
rect 6226 596 6260 630
rect 6326 598 6360 630
rect 6326 596 6354 598
rect 6354 596 6360 598
rect 5826 508 5860 530
rect 5926 508 5960 530
rect 6026 508 6060 530
rect 5826 496 5848 508
rect 5848 496 5860 508
rect 5926 496 5938 508
rect 5938 496 5960 508
rect 6026 496 6028 508
rect 6028 496 6060 508
rect 6126 496 6160 530
rect 6226 496 6260 530
rect 6326 508 6360 530
rect 6326 496 6354 508
rect 6354 496 6360 508
rect 5826 418 5860 430
rect 5926 418 5960 430
rect 6026 418 6060 430
rect 5826 396 5848 418
rect 5848 396 5860 418
rect 5926 396 5938 418
rect 5938 396 5960 418
rect 6026 396 6028 418
rect 6028 396 6060 418
rect 6126 396 6160 430
rect 6226 396 6260 430
rect 6326 418 6360 430
rect 6326 396 6354 418
rect 6354 396 6360 418
rect 7186 924 7208 930
rect 7208 924 7220 930
rect 7286 924 7298 930
rect 7298 924 7320 930
rect 7386 924 7388 930
rect 7388 924 7420 930
rect 7186 896 7220 924
rect 7286 896 7320 924
rect 7386 896 7420 924
rect 7486 896 7520 930
rect 7586 896 7620 930
rect 7686 924 7714 930
rect 7714 924 7720 930
rect 7686 896 7720 924
rect 7186 796 7220 830
rect 7286 796 7320 830
rect 7386 796 7420 830
rect 7486 796 7520 830
rect 7586 796 7620 830
rect 7686 796 7720 830
rect 7186 696 7220 730
rect 7286 696 7320 730
rect 7386 696 7420 730
rect 7486 696 7520 730
rect 7586 696 7620 730
rect 7686 696 7720 730
rect 7186 598 7220 630
rect 7286 598 7320 630
rect 7386 598 7420 630
rect 7186 596 7208 598
rect 7208 596 7220 598
rect 7286 596 7298 598
rect 7298 596 7320 598
rect 7386 596 7388 598
rect 7388 596 7420 598
rect 7486 596 7520 630
rect 7586 596 7620 630
rect 7686 598 7720 630
rect 7686 596 7714 598
rect 7714 596 7720 598
rect 7186 508 7220 530
rect 7286 508 7320 530
rect 7386 508 7420 530
rect 7186 496 7208 508
rect 7208 496 7220 508
rect 7286 496 7298 508
rect 7298 496 7320 508
rect 7386 496 7388 508
rect 7388 496 7420 508
rect 7486 496 7520 530
rect 7586 496 7620 530
rect 7686 508 7720 530
rect 7686 496 7714 508
rect 7714 496 7720 508
rect 7186 418 7220 430
rect 7286 418 7320 430
rect 7386 418 7420 430
rect 7186 396 7208 418
rect 7208 396 7220 418
rect 7286 396 7298 418
rect 7298 396 7320 418
rect 7386 396 7388 418
rect 7388 396 7420 418
rect 7486 396 7520 430
rect 7586 396 7620 430
rect 7686 418 7720 430
rect 7686 396 7714 418
rect 7714 396 7720 418
rect 8546 924 8568 930
rect 8568 924 8580 930
rect 8646 924 8658 930
rect 8658 924 8680 930
rect 8746 924 8748 930
rect 8748 924 8780 930
rect 8546 896 8580 924
rect 8646 896 8680 924
rect 8746 896 8780 924
rect 8846 896 8880 930
rect 8946 896 8980 930
rect 9046 924 9074 930
rect 9074 924 9080 930
rect 9046 896 9080 924
rect 8546 796 8580 830
rect 8646 796 8680 830
rect 8746 796 8780 830
rect 8846 796 8880 830
rect 8946 796 8980 830
rect 9046 796 9080 830
rect 8546 696 8580 730
rect 8646 696 8680 730
rect 8746 696 8780 730
rect 8846 696 8880 730
rect 8946 696 8980 730
rect 9046 696 9080 730
rect 8546 598 8580 630
rect 8646 598 8680 630
rect 8746 598 8780 630
rect 8546 596 8568 598
rect 8568 596 8580 598
rect 8646 596 8658 598
rect 8658 596 8680 598
rect 8746 596 8748 598
rect 8748 596 8780 598
rect 8846 596 8880 630
rect 8946 596 8980 630
rect 9046 598 9080 630
rect 9046 596 9074 598
rect 9074 596 9080 598
rect 8546 508 8580 530
rect 8646 508 8680 530
rect 8746 508 8780 530
rect 8546 496 8568 508
rect 8568 496 8580 508
rect 8646 496 8658 508
rect 8658 496 8680 508
rect 8746 496 8748 508
rect 8748 496 8780 508
rect 8846 496 8880 530
rect 8946 496 8980 530
rect 9046 508 9080 530
rect 9046 496 9074 508
rect 9074 496 9080 508
rect 8546 418 8580 430
rect 8646 418 8680 430
rect 8746 418 8780 430
rect 8546 396 8568 418
rect 8568 396 8580 418
rect 8646 396 8658 418
rect 8658 396 8680 418
rect 8746 396 8748 418
rect 8748 396 8780 418
rect 8846 396 8880 430
rect 8946 396 8980 430
rect 9046 418 9080 430
rect 9046 396 9074 418
rect 9074 396 9080 418
rect 40 50 80 90
rect 140 50 180 90
rect 240 50 280 90
rect 330 50 370 90
rect 410 50 450 90
rect 500 50 540 90
rect 590 50 630 90
rect 680 50 720 90
rect 770 50 810 90
rect 860 50 900 90
rect 950 50 990 90
rect 1040 50 1080 90
rect 1130 50 1170 90
rect 1230 50 1270 90
rect 1320 50 1360 90
rect 1420 50 1460 90
rect 1500 58 1506 90
rect 1506 58 1540 90
rect 1500 50 1540 58
rect 1590 58 1596 90
rect 1596 58 1630 90
rect 1590 50 1630 58
rect 1680 58 1686 90
rect 1686 58 1720 90
rect 1680 50 1720 58
rect 1770 58 1776 90
rect 1776 58 1810 90
rect 1770 50 1810 58
rect 1860 58 1866 90
rect 1866 58 1900 90
rect 1860 50 1900 58
rect 1950 58 1956 90
rect 1956 58 1990 90
rect 1950 50 1990 58
rect 2040 58 2046 90
rect 2046 58 2080 90
rect 2040 50 2080 58
rect 2130 58 2136 90
rect 2136 58 2170 90
rect 2130 50 2170 58
rect 2220 58 2226 90
rect 2226 58 2260 90
rect 2220 50 2260 58
rect 2310 58 2316 90
rect 2316 58 2350 90
rect 2310 50 2350 58
rect 2400 58 2406 90
rect 2406 58 2440 90
rect 2400 50 2440 58
rect 2490 58 2496 90
rect 2496 58 2530 90
rect 2490 50 2530 58
rect 2590 50 2630 90
rect 2680 50 2720 90
rect 2770 50 2810 90
rect 2860 58 2866 90
rect 2866 58 2900 90
rect 2860 50 2900 58
rect 2950 58 2956 90
rect 2956 58 2990 90
rect 2950 50 2990 58
rect 3040 58 3046 90
rect 3046 58 3080 90
rect 3040 50 3080 58
rect 3130 58 3136 90
rect 3136 58 3170 90
rect 3130 50 3170 58
rect 3220 58 3226 90
rect 3226 58 3260 90
rect 3220 50 3260 58
rect 3310 58 3316 90
rect 3316 58 3350 90
rect 3310 50 3350 58
rect 3400 58 3406 90
rect 3406 58 3440 90
rect 3400 50 3440 58
rect 3490 58 3496 90
rect 3496 58 3530 90
rect 3490 50 3530 58
rect 3580 58 3586 90
rect 3586 58 3620 90
rect 3580 50 3620 58
rect 3670 58 3676 90
rect 3676 58 3710 90
rect 3670 50 3710 58
rect 3760 58 3766 90
rect 3766 58 3800 90
rect 3760 50 3800 58
rect 3850 58 3856 90
rect 3856 58 3890 90
rect 3850 50 3890 58
rect 3950 50 3990 90
rect 4040 50 4080 90
rect 4130 50 4170 90
rect 4220 58 4226 90
rect 4226 58 4260 90
rect 4220 50 4260 58
rect 4310 58 4316 90
rect 4316 58 4350 90
rect 4310 50 4350 58
rect 4400 58 4406 90
rect 4406 58 4440 90
rect 4400 50 4440 58
rect 4490 58 4496 90
rect 4496 58 4530 90
rect 4490 50 4530 58
rect 4580 58 4586 90
rect 4586 58 4620 90
rect 4580 50 4620 58
rect 4670 58 4676 90
rect 4676 58 4710 90
rect 4670 50 4710 58
rect 4760 58 4766 90
rect 4766 58 4800 90
rect 4760 50 4800 58
rect 4850 58 4856 90
rect 4856 58 4890 90
rect 4850 50 4890 58
rect 4940 58 4946 90
rect 4946 58 4980 90
rect 4940 50 4980 58
rect 5030 58 5036 90
rect 5036 58 5070 90
rect 5030 50 5070 58
rect 5120 58 5126 90
rect 5126 58 5160 90
rect 5120 50 5160 58
rect 5210 58 5216 90
rect 5216 58 5250 90
rect 5210 50 5250 58
rect 5310 50 5350 90
rect 5400 50 5440 90
rect 5490 50 5530 90
rect 5580 58 5586 90
rect 5586 58 5620 90
rect 5580 50 5620 58
rect 5670 58 5676 90
rect 5676 58 5710 90
rect 5670 50 5710 58
rect 5760 58 5766 90
rect 5766 58 5800 90
rect 5760 50 5800 58
rect 5850 58 5856 90
rect 5856 58 5890 90
rect 5850 50 5890 58
rect 5940 58 5946 90
rect 5946 58 5980 90
rect 5940 50 5980 58
rect 6030 58 6036 90
rect 6036 58 6070 90
rect 6030 50 6070 58
rect 6120 58 6126 90
rect 6126 58 6160 90
rect 6120 50 6160 58
rect 6210 58 6216 90
rect 6216 58 6250 90
rect 6210 50 6250 58
rect 6300 58 6306 90
rect 6306 58 6340 90
rect 6300 50 6340 58
rect 6390 58 6396 90
rect 6396 58 6430 90
rect 6390 50 6430 58
rect 6480 58 6486 90
rect 6486 58 6520 90
rect 6480 50 6520 58
rect 6570 58 6576 90
rect 6576 58 6610 90
rect 6570 50 6610 58
rect 6660 50 6700 90
rect 6760 50 6800 90
rect 6850 50 6890 90
rect 6940 58 6946 90
rect 6946 58 6980 90
rect 6940 50 6980 58
rect 7030 58 7036 90
rect 7036 58 7070 90
rect 7030 50 7070 58
rect 7120 58 7126 90
rect 7126 58 7160 90
rect 7120 50 7160 58
rect 7210 58 7216 90
rect 7216 58 7250 90
rect 7210 50 7250 58
rect 7300 58 7306 90
rect 7306 58 7340 90
rect 7300 50 7340 58
rect 7390 58 7396 90
rect 7396 58 7430 90
rect 7390 50 7430 58
rect 7480 58 7486 90
rect 7486 58 7520 90
rect 7480 50 7520 58
rect 7570 58 7576 90
rect 7576 58 7610 90
rect 7570 50 7610 58
rect 7660 58 7666 90
rect 7666 58 7700 90
rect 7660 50 7700 58
rect 7750 58 7756 90
rect 7756 58 7790 90
rect 7750 50 7790 58
rect 7840 58 7846 90
rect 7846 58 7880 90
rect 7840 50 7880 58
rect 7930 58 7936 90
rect 7936 58 7970 90
rect 7930 50 7970 58
rect 8020 50 8060 90
rect 8120 50 8160 90
rect 8210 50 8250 90
rect 8300 58 8306 90
rect 8306 58 8340 90
rect 8300 50 8340 58
rect 8390 58 8396 90
rect 8396 58 8430 90
rect 8390 50 8430 58
rect 8480 58 8486 90
rect 8486 58 8520 90
rect 8480 50 8520 58
rect 8570 58 8576 90
rect 8576 58 8610 90
rect 8570 50 8610 58
rect 8660 58 8666 90
rect 8666 58 8700 90
rect 8660 50 8700 58
rect 8750 58 8756 90
rect 8756 58 8790 90
rect 8750 50 8790 58
rect 8840 58 8846 90
rect 8846 58 8880 90
rect 8840 50 8880 58
rect 8930 58 8936 90
rect 8936 58 8970 90
rect 8930 50 8970 58
rect 9020 58 9026 90
rect 9026 58 9060 90
rect 9020 50 9060 58
rect 9110 58 9116 90
rect 9116 58 9150 90
rect 9110 50 9150 58
rect 9200 58 9206 90
rect 9206 58 9240 90
rect 9200 50 9240 58
rect 9290 58 9296 90
rect 9296 58 9330 90
rect 9290 50 9330 58
rect 9390 50 9430 90
<< metal1 >>
rect 6440 5570 6480 6300
rect 4620 5560 4700 5570
rect 4620 5500 4630 5560
rect 4690 5500 4700 5560
rect 4620 5490 4700 5500
rect 5020 5560 5100 5570
rect 5020 5500 5030 5560
rect 5090 5500 5100 5560
rect 5020 5490 5100 5500
rect 5420 5560 5500 5570
rect 5420 5500 5430 5560
rect 5490 5500 5500 5560
rect 5420 5490 5500 5500
rect 5820 5560 5900 5570
rect 5820 5500 5830 5560
rect 5890 5500 5900 5560
rect 5820 5490 5900 5500
rect 6220 5560 6300 5570
rect 6220 5500 6230 5560
rect 6290 5500 6300 5560
rect 6220 5490 6300 5500
rect 6420 5550 6500 5570
rect 6420 5510 6440 5550
rect 6480 5510 6500 5550
rect 6420 5490 6500 5510
rect 6620 5560 6700 5570
rect 6620 5500 6630 5560
rect 6690 5500 6700 5560
rect 6620 5490 6700 5500
rect 7020 5560 7100 5570
rect 7020 5500 7030 5560
rect 7090 5500 7100 5560
rect 7020 5490 7100 5500
rect 7420 5560 7500 5570
rect 7420 5500 7430 5560
rect 7490 5500 7500 5560
rect 7420 5490 7500 5500
rect 7820 5560 7900 5570
rect 7820 5500 7830 5560
rect 7890 5500 7900 5560
rect 7820 5490 7900 5500
rect 8220 5560 8300 5570
rect 8220 5500 8230 5560
rect 8290 5500 8300 5560
rect 8220 5490 8300 5500
rect 1890 5040 1970 5050
rect 1890 4980 1900 5040
rect 1960 4980 1970 5040
rect 1890 4970 1970 4980
rect 4300 4620 4380 4630
rect 4300 4560 4310 4620
rect 4370 4560 4380 4620
rect 4300 4550 4380 4560
rect 4820 4620 4900 4630
rect 4820 4560 4830 4620
rect 4890 4560 4900 4620
rect 4820 4550 4900 4560
rect 6220 4610 6300 4630
rect 6220 4570 6240 4610
rect 6280 4570 6300 4610
rect 6220 4550 6300 4570
rect 6620 4610 6700 4630
rect 6620 4570 6640 4610
rect 6680 4570 6700 4610
rect 6620 4550 6700 4570
rect 6820 4620 6900 4630
rect 6820 4560 6830 4620
rect 6890 4560 6900 4620
rect 6820 4550 6900 4560
rect 7620 4620 7700 4630
rect 7620 4560 7630 4620
rect 7690 4560 7700 4620
rect 7620 4550 7700 4560
rect 8140 4620 8220 4630
rect 8140 4560 8150 4620
rect 8210 4560 8220 4620
rect 8140 4550 8220 4560
rect 8750 4620 8830 4630
rect 8750 4560 8760 4620
rect 8820 4560 8830 4620
rect 8750 4550 8830 4560
rect 3790 4450 4230 4460
rect 3790 4390 3800 4450
rect 4220 4390 4230 4450
rect 3790 4380 4230 4390
rect 1890 4020 1970 4030
rect 1890 3960 1900 4020
rect 1960 3960 1970 4020
rect 1890 3950 1970 3960
rect 4320 3440 4360 4550
rect 5220 4530 5300 4540
rect 5220 4470 5230 4530
rect 5290 4470 5300 4530
rect 5220 4460 5300 4470
rect 6020 4530 6100 4540
rect 6020 4470 6030 4530
rect 6090 4470 6100 4530
rect 6020 4460 6100 4470
rect 5620 4440 5700 4450
rect 5620 4380 5630 4440
rect 5690 4380 5700 4440
rect 5620 4370 5700 4380
rect 6240 4330 6280 4550
rect 6420 4440 6500 4450
rect 6420 4380 6430 4440
rect 6490 4380 6500 4440
rect 6420 4370 6500 4380
rect 6640 4330 6680 4550
rect 8020 4530 8100 4540
rect 8020 4470 8030 4530
rect 8090 4470 8100 4530
rect 8020 4460 8100 4470
rect 8630 4530 8710 4540
rect 8630 4470 8640 4530
rect 8700 4470 8710 4530
rect 8630 4460 8710 4470
rect 7220 4440 7300 4450
rect 7220 4380 7230 4440
rect 7290 4380 7300 4440
rect 7220 4370 7300 4380
rect 5220 4320 5300 4330
rect 5220 4260 5230 4320
rect 5290 4260 5300 4320
rect 5220 4250 5300 4260
rect 5620 4320 5700 4330
rect 5620 4260 5630 4320
rect 5690 4260 5700 4320
rect 5620 4250 5700 4260
rect 6020 4320 6100 4330
rect 6020 4260 6030 4320
rect 6090 4260 6100 4320
rect 6020 4250 6100 4260
rect 6220 4310 6300 4330
rect 6220 4270 6240 4310
rect 6280 4270 6300 4310
rect 6220 4250 6300 4270
rect 6420 4320 6500 4330
rect 6420 4260 6430 4320
rect 6490 4260 6500 4320
rect 6420 4250 6500 4260
rect 6620 4310 6700 4330
rect 6620 4270 6640 4310
rect 6680 4270 6700 4310
rect 6620 4250 6700 4270
rect 6820 4320 6900 4330
rect 6820 4260 6830 4320
rect 6890 4260 6900 4320
rect 6820 4250 6900 4260
rect 7220 4320 7300 4330
rect 7220 4260 7230 4320
rect 7290 4260 7300 4320
rect 7220 4250 7300 4260
rect 7620 4320 7700 4330
rect 7620 4260 7630 4320
rect 7690 4260 7700 4320
rect 7620 4250 7700 4260
rect 5820 3780 5900 3790
rect 5820 3720 5830 3780
rect 5890 3720 5900 3780
rect 5820 3710 5900 3720
rect 6220 3780 6300 3790
rect 6220 3720 6230 3780
rect 6290 3720 6300 3780
rect 6220 3710 6300 3720
rect 6460 3770 6540 3790
rect 6460 3730 6480 3770
rect 6520 3730 6540 3770
rect 6460 3710 6540 3730
rect 6620 3780 6700 3790
rect 6620 3720 6630 3780
rect 6690 3720 6700 3780
rect 6620 3710 6700 3720
rect 7020 3780 7100 3790
rect 7020 3720 7030 3780
rect 7090 3720 7100 3780
rect 7020 3710 7100 3720
rect 5420 3690 5500 3700
rect 5420 3630 5430 3690
rect 5490 3630 5500 3690
rect 5420 3620 5500 3630
rect 5980 3690 6060 3700
rect 5980 3630 5990 3690
rect 6050 3630 6060 3690
rect 5980 3620 6060 3630
rect 6000 3520 6040 3620
rect 5820 3510 5900 3520
rect 5820 3450 5830 3510
rect 5890 3450 5900 3510
rect 5820 3440 5900 3450
rect 5980 3510 6060 3520
rect 5980 3450 5990 3510
rect 6050 3450 6060 3510
rect 5980 3440 6060 3450
rect 880 3430 960 3440
rect 880 3370 890 3430
rect 950 3370 960 3430
rect 880 1450 960 3370
rect 3790 3430 4230 3440
rect 3790 3370 3800 3430
rect 4220 3370 4230 3430
rect 3790 3360 4230 3370
rect 4300 3420 4380 3440
rect 6240 3430 6280 3710
rect 6330 3690 6410 3700
rect 6330 3630 6340 3690
rect 6400 3630 6410 3690
rect 6330 3620 6410 3630
rect 6480 3610 6520 3710
rect 6460 3600 6540 3610
rect 6460 3540 6470 3600
rect 6530 3540 6540 3600
rect 6460 3530 6540 3540
rect 6640 3430 6680 3710
rect 6860 3690 6940 3700
rect 6860 3630 6870 3690
rect 6930 3630 6940 3690
rect 6860 3620 6940 3630
rect 7420 3690 7500 3700
rect 7420 3630 7430 3690
rect 7490 3630 7500 3690
rect 7420 3620 7500 3630
rect 6880 3520 6920 3620
rect 8440 3600 8520 3610
rect 8440 3540 8450 3600
rect 8510 3540 8520 3600
rect 8440 3530 8520 3540
rect 6860 3510 6940 3520
rect 6860 3450 6870 3510
rect 6930 3450 6940 3510
rect 6860 3440 6940 3450
rect 7020 3510 7100 3520
rect 7020 3450 7030 3510
rect 7090 3450 7100 3510
rect 7020 3440 7100 3450
rect 4300 3360 4310 3420
rect 4370 3360 4380 3420
rect 4300 3350 4380 3360
rect 6100 3420 6180 3430
rect 6100 3360 6110 3420
rect 6170 3360 6180 3420
rect 6100 3350 6180 3360
rect 6220 3410 6300 3430
rect 6220 3370 6240 3410
rect 6280 3370 6300 3410
rect 6220 3350 6300 3370
rect 6620 3410 6700 3430
rect 6620 3370 6640 3410
rect 6680 3370 6700 3410
rect 6620 3350 6700 3370
rect 6740 3420 6820 3430
rect 6740 3360 6750 3420
rect 6810 3360 6820 3420
rect 6740 3350 6820 3360
rect 5820 3080 5900 3090
rect 1720 3070 1800 3080
rect 1720 3010 1730 3070
rect 1790 3010 1800 3070
rect 1300 1650 1380 1660
rect 1300 1590 1310 1650
rect 1370 1590 1380 1650
rect 1300 1580 1380 1590
rect 360 370 960 1450
rect 1720 1460 1800 3010
rect 1890 3070 1970 3080
rect 1890 3010 1900 3070
rect 1960 3010 1970 3070
rect 1890 3000 1970 3010
rect 3790 3070 4230 3080
rect 3790 3010 3800 3070
rect 4220 3010 4230 3070
rect 5820 3020 5830 3080
rect 5890 3020 5900 3080
rect 5820 3010 5900 3020
rect 7020 3080 7100 3090
rect 7020 3020 7030 3080
rect 7090 3020 7100 3080
rect 7020 3010 7100 3020
rect 3790 3000 4230 3010
rect 5620 2990 5700 3000
rect 5620 2930 5630 2990
rect 5690 2930 5700 2990
rect 5620 2920 5700 2930
rect 6020 2990 6100 3000
rect 6020 2930 6030 2990
rect 6090 2930 6100 2990
rect 6020 2920 6100 2930
rect 6420 2990 6500 3000
rect 6420 2930 6430 2990
rect 6490 2930 6500 2990
rect 6420 2920 6500 2930
rect 6820 2990 6900 3000
rect 6820 2930 6830 2990
rect 6890 2930 6900 2990
rect 6820 2920 6900 2930
rect 7220 2990 7300 3000
rect 7220 2930 7230 2990
rect 7290 2930 7300 2990
rect 7220 2920 7300 2930
rect 8460 2880 8500 3530
rect 8650 3090 8690 4460
rect 8770 4420 8810 4550
rect 8750 4410 8830 4420
rect 8750 4370 8770 4410
rect 8810 4370 8830 4410
rect 8750 4350 8830 4370
rect 9170 4320 9250 4330
rect 9170 4260 9180 4320
rect 9240 4260 9250 4320
rect 9170 4250 9250 4260
rect 8970 3740 9050 3760
rect 8970 3700 8990 3740
rect 9030 3700 9050 3740
rect 8970 3680 9050 3700
rect 8860 3420 8940 3430
rect 8860 3360 8870 3420
rect 8930 3360 8940 3420
rect 8860 3350 8940 3360
rect 8630 3080 8710 3090
rect 8630 3020 8640 3080
rect 8700 3020 8710 3080
rect 8630 3010 8710 3020
rect 7380 2870 7460 2880
rect 7380 2810 7390 2870
rect 7450 2810 7460 2870
rect 7380 2800 7460 2810
rect 8440 2870 8520 2880
rect 8440 2810 8450 2870
rect 8510 2810 8520 2870
rect 8440 2800 8520 2810
rect 1890 2480 1970 2490
rect 1890 2420 1900 2480
rect 1960 2420 1970 2480
rect 1890 2410 1970 2420
rect 6340 1930 6580 1940
rect 6340 1870 6350 1930
rect 6410 1870 6430 1930
rect 6490 1870 6510 1930
rect 6570 1870 6580 1930
rect 6340 1860 6580 1870
rect 9010 1820 9050 3680
rect 7440 1810 7520 1820
rect 7440 1750 7450 1810
rect 7510 1750 7520 1810
rect 7440 1740 7520 1750
rect 8990 1810 9070 1820
rect 8990 1750 9000 1810
rect 9060 1750 9070 1810
rect 8990 1740 9070 1750
rect 7590 1640 7670 1650
rect 7590 1580 7600 1640
rect 7660 1580 7670 1640
rect 7590 1570 7670 1580
rect 1720 1380 9120 1460
rect 1720 975 2320 1380
rect 3080 975 3680 1380
rect 4440 975 5040 1380
rect 5800 975 6400 1380
rect 7160 975 7760 1380
rect 8520 975 9120 1380
rect 1715 930 2325 975
rect 1715 896 1746 930
rect 1780 896 1846 930
rect 1880 896 1946 930
rect 1980 896 2046 930
rect 2080 896 2146 930
rect 2180 896 2246 930
rect 2280 896 2325 930
rect 1715 830 2325 896
rect 1715 796 1746 830
rect 1780 796 1846 830
rect 1880 796 1946 830
rect 1980 796 2046 830
rect 2080 796 2146 830
rect 2180 796 2246 830
rect 2280 796 2325 830
rect 1715 730 2325 796
rect 1715 696 1746 730
rect 1780 696 1846 730
rect 1880 696 1946 730
rect 1980 696 2046 730
rect 2080 696 2146 730
rect 2180 696 2246 730
rect 2280 696 2325 730
rect 1715 630 2325 696
rect 1715 596 1746 630
rect 1780 596 1846 630
rect 1880 596 1946 630
rect 1980 596 2046 630
rect 2080 596 2146 630
rect 2180 596 2246 630
rect 2280 596 2325 630
rect 1715 530 2325 596
rect 1715 496 1746 530
rect 1780 496 1846 530
rect 1880 496 1946 530
rect 1980 496 2046 530
rect 2080 496 2146 530
rect 2180 496 2246 530
rect 2280 496 2325 530
rect 1715 430 2325 496
rect 1715 396 1746 430
rect 1780 396 1846 430
rect 1880 396 1946 430
rect 1980 396 2046 430
rect 2080 396 2146 430
rect 2180 396 2246 430
rect 2280 396 2325 430
rect 1715 365 2325 396
rect 3075 930 3685 975
rect 3075 896 3106 930
rect 3140 896 3206 930
rect 3240 896 3306 930
rect 3340 896 3406 930
rect 3440 896 3506 930
rect 3540 896 3606 930
rect 3640 896 3685 930
rect 3075 830 3685 896
rect 3075 796 3106 830
rect 3140 796 3206 830
rect 3240 796 3306 830
rect 3340 796 3406 830
rect 3440 796 3506 830
rect 3540 796 3606 830
rect 3640 796 3685 830
rect 3075 730 3685 796
rect 3075 696 3106 730
rect 3140 696 3206 730
rect 3240 696 3306 730
rect 3340 696 3406 730
rect 3440 696 3506 730
rect 3540 696 3606 730
rect 3640 696 3685 730
rect 3075 630 3685 696
rect 3075 596 3106 630
rect 3140 596 3206 630
rect 3240 596 3306 630
rect 3340 596 3406 630
rect 3440 596 3506 630
rect 3540 596 3606 630
rect 3640 596 3685 630
rect 3075 530 3685 596
rect 3075 496 3106 530
rect 3140 496 3206 530
rect 3240 496 3306 530
rect 3340 496 3406 530
rect 3440 496 3506 530
rect 3540 496 3606 530
rect 3640 496 3685 530
rect 3075 430 3685 496
rect 3075 396 3106 430
rect 3140 396 3206 430
rect 3240 396 3306 430
rect 3340 396 3406 430
rect 3440 396 3506 430
rect 3540 396 3606 430
rect 3640 396 3685 430
rect 3075 365 3685 396
rect 4435 930 5045 975
rect 4435 896 4466 930
rect 4500 896 4566 930
rect 4600 896 4666 930
rect 4700 896 4766 930
rect 4800 896 4866 930
rect 4900 896 4966 930
rect 5000 896 5045 930
rect 4435 830 5045 896
rect 4435 796 4466 830
rect 4500 796 4566 830
rect 4600 796 4666 830
rect 4700 796 4766 830
rect 4800 796 4866 830
rect 4900 796 4966 830
rect 5000 796 5045 830
rect 4435 730 5045 796
rect 4435 696 4466 730
rect 4500 696 4566 730
rect 4600 696 4666 730
rect 4700 696 4766 730
rect 4800 696 4866 730
rect 4900 696 4966 730
rect 5000 696 5045 730
rect 4435 630 5045 696
rect 4435 596 4466 630
rect 4500 596 4566 630
rect 4600 596 4666 630
rect 4700 596 4766 630
rect 4800 596 4866 630
rect 4900 596 4966 630
rect 5000 596 5045 630
rect 4435 530 5045 596
rect 4435 496 4466 530
rect 4500 496 4566 530
rect 4600 496 4666 530
rect 4700 496 4766 530
rect 4800 496 4866 530
rect 4900 496 4966 530
rect 5000 496 5045 530
rect 4435 430 5045 496
rect 4435 396 4466 430
rect 4500 396 4566 430
rect 4600 396 4666 430
rect 4700 396 4766 430
rect 4800 396 4866 430
rect 4900 396 4966 430
rect 5000 396 5045 430
rect 4435 365 5045 396
rect 5795 930 6405 975
rect 5795 896 5826 930
rect 5860 896 5926 930
rect 5960 896 6026 930
rect 6060 896 6126 930
rect 6160 896 6226 930
rect 6260 896 6326 930
rect 6360 896 6405 930
rect 5795 830 6405 896
rect 5795 796 5826 830
rect 5860 796 5926 830
rect 5960 796 6026 830
rect 6060 796 6126 830
rect 6160 796 6226 830
rect 6260 796 6326 830
rect 6360 796 6405 830
rect 5795 730 6405 796
rect 5795 696 5826 730
rect 5860 696 5926 730
rect 5960 696 6026 730
rect 6060 696 6126 730
rect 6160 696 6226 730
rect 6260 696 6326 730
rect 6360 696 6405 730
rect 5795 630 6405 696
rect 5795 596 5826 630
rect 5860 596 5926 630
rect 5960 596 6026 630
rect 6060 596 6126 630
rect 6160 596 6226 630
rect 6260 596 6326 630
rect 6360 596 6405 630
rect 5795 530 6405 596
rect 5795 496 5826 530
rect 5860 496 5926 530
rect 5960 496 6026 530
rect 6060 496 6126 530
rect 6160 496 6226 530
rect 6260 496 6326 530
rect 6360 496 6405 530
rect 5795 430 6405 496
rect 5795 396 5826 430
rect 5860 396 5926 430
rect 5960 396 6026 430
rect 6060 396 6126 430
rect 6160 396 6226 430
rect 6260 396 6326 430
rect 6360 396 6405 430
rect 5795 365 6405 396
rect 7155 930 7765 975
rect 7155 896 7186 930
rect 7220 896 7286 930
rect 7320 896 7386 930
rect 7420 896 7486 930
rect 7520 896 7586 930
rect 7620 896 7686 930
rect 7720 896 7765 930
rect 7155 830 7765 896
rect 7155 796 7186 830
rect 7220 796 7286 830
rect 7320 796 7386 830
rect 7420 796 7486 830
rect 7520 796 7586 830
rect 7620 796 7686 830
rect 7720 796 7765 830
rect 7155 730 7765 796
rect 7155 696 7186 730
rect 7220 696 7286 730
rect 7320 696 7386 730
rect 7420 696 7486 730
rect 7520 696 7586 730
rect 7620 696 7686 730
rect 7720 696 7765 730
rect 7155 630 7765 696
rect 7155 596 7186 630
rect 7220 596 7286 630
rect 7320 596 7386 630
rect 7420 596 7486 630
rect 7520 596 7586 630
rect 7620 596 7686 630
rect 7720 596 7765 630
rect 7155 530 7765 596
rect 7155 496 7186 530
rect 7220 496 7286 530
rect 7320 496 7386 530
rect 7420 496 7486 530
rect 7520 496 7586 530
rect 7620 496 7686 530
rect 7720 496 7765 530
rect 7155 430 7765 496
rect 7155 396 7186 430
rect 7220 396 7286 430
rect 7320 396 7386 430
rect 7420 396 7486 430
rect 7520 396 7586 430
rect 7620 396 7686 430
rect 7720 396 7765 430
rect 7155 365 7765 396
rect 8515 930 9125 975
rect 8515 896 8546 930
rect 8580 896 8646 930
rect 8680 896 8746 930
rect 8780 896 8846 930
rect 8880 896 8946 930
rect 8980 896 9046 930
rect 9080 896 9125 930
rect 8515 830 9125 896
rect 8515 796 8546 830
rect 8580 796 8646 830
rect 8680 796 8746 830
rect 8780 796 8846 830
rect 8880 796 8946 830
rect 8980 796 9046 830
rect 9080 796 9125 830
rect 8515 730 9125 796
rect 8515 696 8546 730
rect 8580 696 8646 730
rect 8680 696 8746 730
rect 8780 696 8846 730
rect 8880 696 8946 730
rect 8980 696 9046 730
rect 9080 696 9125 730
rect 8515 630 9125 696
rect 8515 596 8546 630
rect 8580 596 8646 630
rect 8680 596 8746 630
rect 8780 596 8846 630
rect 8880 596 8946 630
rect 8980 596 9046 630
rect 9080 596 9125 630
rect 8515 530 9125 596
rect 8515 496 8546 530
rect 8580 496 8646 530
rect 8680 496 8746 530
rect 8780 496 8846 530
rect 8880 496 8946 530
rect 8980 496 9046 530
rect 9080 496 9125 530
rect 8515 430 9125 496
rect 8515 396 8546 430
rect 8580 396 8646 430
rect 8680 396 8746 430
rect 8780 396 8846 430
rect 8880 396 8946 430
rect 8980 396 9046 430
rect 9080 396 9125 430
rect 8515 365 9125 396
rect 10 100 9460 120
rect 10 40 30 100
rect 90 40 130 100
rect 190 40 230 100
rect 290 40 320 100
rect 380 40 400 100
rect 460 40 490 100
rect 550 40 580 100
rect 640 40 670 100
rect 730 40 760 100
rect 820 40 850 100
rect 910 40 940 100
rect 1000 40 1030 100
rect 1090 40 1120 100
rect 1180 40 1220 100
rect 1280 40 1310 100
rect 1370 40 1410 100
rect 1470 40 1490 100
rect 1550 40 1580 100
rect 1640 40 1670 100
rect 1730 40 1760 100
rect 1820 40 1850 100
rect 1910 40 1940 100
rect 2000 40 2030 100
rect 2090 40 2120 100
rect 2180 40 2210 100
rect 2270 40 2300 100
rect 2360 40 2390 100
rect 2450 40 2480 100
rect 2540 40 2580 100
rect 2640 40 2670 100
rect 2730 40 2760 100
rect 2820 40 2850 100
rect 2910 40 2940 100
rect 3000 40 3030 100
rect 3090 40 3120 100
rect 3180 40 3210 100
rect 3270 40 3300 100
rect 3360 40 3390 100
rect 3450 40 3480 100
rect 3540 40 3570 100
rect 3630 40 3660 100
rect 3720 40 3750 100
rect 3810 40 3840 100
rect 3900 40 3940 100
rect 4000 40 4030 100
rect 4090 40 4120 100
rect 4180 40 4210 100
rect 4270 40 4300 100
rect 4360 40 4390 100
rect 4450 40 4480 100
rect 4540 40 4570 100
rect 4630 40 4660 100
rect 4720 40 4750 100
rect 4810 40 4840 100
rect 4900 40 4930 100
rect 4990 40 5020 100
rect 5080 40 5110 100
rect 5170 40 5200 100
rect 5260 40 5300 100
rect 5360 40 5390 100
rect 5450 40 5480 100
rect 5540 40 5570 100
rect 5630 40 5660 100
rect 5720 40 5750 100
rect 5810 40 5840 100
rect 5900 40 5930 100
rect 5990 40 6020 100
rect 6080 40 6110 100
rect 6170 40 6200 100
rect 6260 40 6290 100
rect 6350 40 6380 100
rect 6440 40 6470 100
rect 6530 40 6560 100
rect 6620 40 6650 100
rect 6710 40 6750 100
rect 6810 40 6840 100
rect 6900 40 6930 100
rect 6990 40 7020 100
rect 7080 40 7110 100
rect 7170 40 7200 100
rect 7260 40 7290 100
rect 7350 40 7380 100
rect 7440 40 7470 100
rect 7530 40 7560 100
rect 7620 40 7650 100
rect 7710 40 7740 100
rect 7800 40 7830 100
rect 7890 40 7920 100
rect 7980 40 8010 100
rect 8070 40 8110 100
rect 8170 40 8200 100
rect 8260 40 8290 100
rect 8350 40 8380 100
rect 8440 40 8470 100
rect 8530 40 8560 100
rect 8620 40 8650 100
rect 8710 40 8740 100
rect 8800 40 8830 100
rect 8890 40 8920 100
rect 8980 40 9010 100
rect 9070 40 9100 100
rect 9160 40 9190 100
rect 9250 40 9280 100
rect 9340 40 9380 100
rect 9440 40 9460 100
rect 10 20 9460 40
<< via1 >>
rect 4630 5550 4690 5560
rect 4630 5510 4640 5550
rect 4640 5510 4680 5550
rect 4680 5510 4690 5550
rect 4630 5500 4690 5510
rect 5030 5550 5090 5560
rect 5030 5510 5040 5550
rect 5040 5510 5080 5550
rect 5080 5510 5090 5550
rect 5030 5500 5090 5510
rect 5430 5550 5490 5560
rect 5430 5510 5440 5550
rect 5440 5510 5480 5550
rect 5480 5510 5490 5550
rect 5430 5500 5490 5510
rect 5830 5550 5890 5560
rect 5830 5510 5840 5550
rect 5840 5510 5880 5550
rect 5880 5510 5890 5550
rect 5830 5500 5890 5510
rect 6230 5550 6290 5560
rect 6230 5510 6240 5550
rect 6240 5510 6280 5550
rect 6280 5510 6290 5550
rect 6230 5500 6290 5510
rect 6630 5550 6690 5560
rect 6630 5510 6640 5550
rect 6640 5510 6680 5550
rect 6680 5510 6690 5550
rect 6630 5500 6690 5510
rect 7030 5550 7090 5560
rect 7030 5510 7040 5550
rect 7040 5510 7080 5550
rect 7080 5510 7090 5550
rect 7030 5500 7090 5510
rect 7430 5550 7490 5560
rect 7430 5510 7440 5550
rect 7440 5510 7480 5550
rect 7480 5510 7490 5550
rect 7430 5500 7490 5510
rect 7830 5550 7890 5560
rect 7830 5510 7840 5550
rect 7840 5510 7880 5550
rect 7880 5510 7890 5550
rect 7830 5500 7890 5510
rect 8230 5550 8290 5560
rect 8230 5510 8240 5550
rect 8240 5510 8280 5550
rect 8280 5510 8290 5550
rect 8230 5500 8290 5510
rect 1900 5030 1960 5040
rect 1900 4990 1910 5030
rect 1910 4990 1950 5030
rect 1950 4990 1960 5030
rect 1900 4980 1960 4990
rect 4310 4560 4370 4620
rect 4830 4610 4890 4620
rect 4830 4570 4840 4610
rect 4840 4570 4880 4610
rect 4880 4570 4890 4610
rect 4830 4560 4890 4570
rect 6830 4610 6890 4620
rect 6830 4570 6840 4610
rect 6840 4570 6880 4610
rect 6880 4570 6890 4610
rect 6830 4560 6890 4570
rect 7630 4610 7690 4620
rect 7630 4570 7640 4610
rect 7640 4570 7680 4610
rect 7680 4570 7690 4610
rect 7630 4560 7690 4570
rect 8150 4610 8210 4620
rect 8150 4570 8160 4610
rect 8160 4570 8200 4610
rect 8200 4570 8210 4610
rect 8150 4560 8210 4570
rect 8760 4560 8820 4620
rect 3800 4440 4220 4450
rect 3800 4400 3810 4440
rect 3810 4400 3850 4440
rect 3850 4400 3900 4440
rect 3900 4400 3940 4440
rect 3940 4400 3990 4440
rect 3990 4400 4030 4440
rect 4030 4400 4080 4440
rect 4080 4400 4120 4440
rect 4120 4400 4170 4440
rect 4170 4400 4210 4440
rect 4210 4400 4220 4440
rect 3800 4390 4220 4400
rect 1900 4010 1960 4020
rect 1900 3970 1910 4010
rect 1910 3970 1950 4010
rect 1950 3970 1960 4010
rect 1900 3960 1960 3970
rect 5230 4520 5290 4530
rect 5230 4480 5240 4520
rect 5240 4480 5280 4520
rect 5280 4480 5290 4520
rect 5230 4470 5290 4480
rect 6030 4520 6090 4530
rect 6030 4480 6040 4520
rect 6040 4480 6080 4520
rect 6080 4480 6090 4520
rect 6030 4470 6090 4480
rect 5630 4430 5690 4440
rect 5630 4390 5640 4430
rect 5640 4390 5680 4430
rect 5680 4390 5690 4430
rect 5630 4380 5690 4390
rect 6430 4430 6490 4440
rect 6430 4390 6440 4430
rect 6440 4390 6480 4430
rect 6480 4390 6490 4430
rect 6430 4380 6490 4390
rect 8030 4520 8090 4530
rect 8030 4480 8040 4520
rect 8040 4480 8080 4520
rect 8080 4480 8090 4520
rect 8030 4470 8090 4480
rect 8640 4470 8700 4530
rect 7230 4430 7290 4440
rect 7230 4390 7240 4430
rect 7240 4390 7280 4430
rect 7280 4390 7290 4430
rect 7230 4380 7290 4390
rect 5230 4310 5290 4320
rect 5230 4270 5240 4310
rect 5240 4270 5280 4310
rect 5280 4270 5290 4310
rect 5230 4260 5290 4270
rect 5630 4310 5690 4320
rect 5630 4270 5640 4310
rect 5640 4270 5680 4310
rect 5680 4270 5690 4310
rect 5630 4260 5690 4270
rect 6030 4310 6090 4320
rect 6030 4270 6040 4310
rect 6040 4270 6080 4310
rect 6080 4270 6090 4310
rect 6030 4260 6090 4270
rect 6430 4310 6490 4320
rect 6430 4270 6440 4310
rect 6440 4270 6480 4310
rect 6480 4270 6490 4310
rect 6430 4260 6490 4270
rect 6830 4310 6890 4320
rect 6830 4270 6840 4310
rect 6840 4270 6880 4310
rect 6880 4270 6890 4310
rect 6830 4260 6890 4270
rect 7230 4310 7290 4320
rect 7230 4270 7240 4310
rect 7240 4270 7280 4310
rect 7280 4270 7290 4310
rect 7230 4260 7290 4270
rect 7630 4310 7690 4320
rect 7630 4270 7640 4310
rect 7640 4270 7680 4310
rect 7680 4270 7690 4310
rect 7630 4260 7690 4270
rect 5830 3770 5890 3780
rect 5830 3730 5840 3770
rect 5840 3730 5880 3770
rect 5880 3730 5890 3770
rect 5830 3720 5890 3730
rect 6230 3720 6290 3780
rect 6630 3720 6690 3780
rect 7030 3770 7090 3780
rect 7030 3730 7040 3770
rect 7040 3730 7080 3770
rect 7080 3730 7090 3770
rect 7030 3720 7090 3730
rect 5430 3680 5490 3690
rect 5430 3640 5440 3680
rect 5440 3640 5480 3680
rect 5480 3640 5490 3680
rect 5430 3630 5490 3640
rect 5990 3630 6050 3690
rect 5830 3500 5890 3510
rect 5830 3460 5840 3500
rect 5840 3460 5880 3500
rect 5880 3460 5890 3500
rect 5830 3450 5890 3460
rect 5990 3450 6050 3510
rect 890 3370 950 3430
rect 3800 3420 4220 3430
rect 3800 3380 3810 3420
rect 3810 3380 3850 3420
rect 3850 3380 3900 3420
rect 3900 3380 3940 3420
rect 3940 3380 3990 3420
rect 3990 3380 4030 3420
rect 4030 3380 4080 3420
rect 4080 3380 4120 3420
rect 4120 3380 4170 3420
rect 4170 3380 4210 3420
rect 4210 3380 4220 3420
rect 3800 3370 4220 3380
rect 6340 3680 6400 3690
rect 6340 3640 6350 3680
rect 6350 3640 6390 3680
rect 6390 3640 6400 3680
rect 6340 3630 6400 3640
rect 6470 3590 6530 3600
rect 6470 3550 6480 3590
rect 6480 3550 6520 3590
rect 6520 3550 6530 3590
rect 6470 3540 6530 3550
rect 6870 3630 6930 3690
rect 7430 3680 7490 3690
rect 7430 3640 7440 3680
rect 7440 3640 7480 3680
rect 7480 3640 7490 3680
rect 7430 3630 7490 3640
rect 8450 3540 8510 3600
rect 6870 3450 6930 3510
rect 7030 3500 7090 3510
rect 7030 3460 7040 3500
rect 7040 3460 7080 3500
rect 7080 3460 7090 3500
rect 7030 3450 7090 3460
rect 4310 3360 4370 3420
rect 6110 3410 6170 3420
rect 6110 3370 6120 3410
rect 6120 3370 6160 3410
rect 6160 3370 6170 3410
rect 6110 3360 6170 3370
rect 6750 3410 6810 3420
rect 6750 3370 6760 3410
rect 6760 3370 6800 3410
rect 6800 3370 6810 3410
rect 6750 3360 6810 3370
rect 1730 3010 1790 3070
rect 1310 1640 1370 1650
rect 1310 1600 1320 1640
rect 1320 1600 1360 1640
rect 1360 1600 1370 1640
rect 1310 1590 1370 1600
rect 1900 3060 1960 3070
rect 1900 3020 1910 3060
rect 1910 3020 1950 3060
rect 1950 3020 1960 3060
rect 1900 3010 1960 3020
rect 3800 3060 4220 3070
rect 3800 3020 3810 3060
rect 3810 3020 3850 3060
rect 3850 3020 3900 3060
rect 3900 3020 3940 3060
rect 3940 3020 3990 3060
rect 3990 3020 4030 3060
rect 4030 3020 4080 3060
rect 4080 3020 4120 3060
rect 4120 3020 4170 3060
rect 4170 3020 4210 3060
rect 4210 3020 4220 3060
rect 3800 3010 4220 3020
rect 5830 3070 5890 3080
rect 5830 3030 5840 3070
rect 5840 3030 5880 3070
rect 5880 3030 5890 3070
rect 5830 3020 5890 3030
rect 7030 3070 7090 3080
rect 7030 3030 7040 3070
rect 7040 3030 7080 3070
rect 7080 3030 7090 3070
rect 7030 3020 7090 3030
rect 5630 2980 5690 2990
rect 5630 2940 5640 2980
rect 5640 2940 5680 2980
rect 5680 2940 5690 2980
rect 5630 2930 5690 2940
rect 6030 2980 6090 2990
rect 6030 2940 6040 2980
rect 6040 2940 6080 2980
rect 6080 2940 6090 2980
rect 6030 2930 6090 2940
rect 6430 2980 6490 2990
rect 6430 2940 6440 2980
rect 6440 2940 6480 2980
rect 6480 2940 6490 2980
rect 6430 2930 6490 2940
rect 6830 2980 6890 2990
rect 6830 2940 6840 2980
rect 6840 2940 6880 2980
rect 6880 2940 6890 2980
rect 6830 2930 6890 2940
rect 7230 2980 7290 2990
rect 7230 2940 7240 2980
rect 7240 2940 7280 2980
rect 7280 2940 7290 2980
rect 7230 2930 7290 2940
rect 9180 4310 9240 4320
rect 9180 4270 9190 4310
rect 9190 4270 9230 4310
rect 9230 4270 9240 4310
rect 9180 4260 9240 4270
rect 8870 3410 8930 3420
rect 8870 3370 8880 3410
rect 8880 3370 8920 3410
rect 8920 3370 8930 3410
rect 8870 3360 8930 3370
rect 8640 3020 8700 3080
rect 7390 2860 7450 2870
rect 7390 2820 7400 2860
rect 7400 2820 7440 2860
rect 7440 2820 7450 2860
rect 7390 2810 7450 2820
rect 8450 2810 8510 2870
rect 1900 2470 1960 2480
rect 1900 2430 1910 2470
rect 1910 2430 1950 2470
rect 1950 2430 1960 2470
rect 1900 2420 1960 2430
rect 6350 1920 6410 1930
rect 6350 1880 6360 1920
rect 6360 1880 6400 1920
rect 6400 1880 6410 1920
rect 6350 1870 6410 1880
rect 6430 1920 6490 1930
rect 6430 1880 6440 1920
rect 6440 1880 6480 1920
rect 6480 1880 6490 1920
rect 6430 1870 6490 1880
rect 6510 1920 6570 1930
rect 6510 1880 6520 1920
rect 6520 1880 6560 1920
rect 6560 1880 6570 1920
rect 6510 1870 6570 1880
rect 7450 1800 7510 1810
rect 7450 1760 7460 1800
rect 7460 1760 7500 1800
rect 7500 1760 7510 1800
rect 7450 1750 7510 1760
rect 9000 1750 9060 1810
rect 7600 1630 7660 1640
rect 7600 1590 7610 1630
rect 7610 1590 7650 1630
rect 7650 1590 7660 1630
rect 7600 1580 7660 1590
rect 30 90 90 100
rect 30 50 40 90
rect 40 50 80 90
rect 80 50 90 90
rect 30 40 90 50
rect 130 90 190 100
rect 130 50 140 90
rect 140 50 180 90
rect 180 50 190 90
rect 130 40 190 50
rect 230 90 290 100
rect 230 50 240 90
rect 240 50 280 90
rect 280 50 290 90
rect 230 40 290 50
rect 320 90 380 100
rect 320 50 330 90
rect 330 50 370 90
rect 370 50 380 90
rect 320 40 380 50
rect 400 90 460 100
rect 400 50 410 90
rect 410 50 450 90
rect 450 50 460 90
rect 400 40 460 50
rect 490 90 550 100
rect 490 50 500 90
rect 500 50 540 90
rect 540 50 550 90
rect 490 40 550 50
rect 580 90 640 100
rect 580 50 590 90
rect 590 50 630 90
rect 630 50 640 90
rect 580 40 640 50
rect 670 90 730 100
rect 670 50 680 90
rect 680 50 720 90
rect 720 50 730 90
rect 670 40 730 50
rect 760 90 820 100
rect 760 50 770 90
rect 770 50 810 90
rect 810 50 820 90
rect 760 40 820 50
rect 850 90 910 100
rect 850 50 860 90
rect 860 50 900 90
rect 900 50 910 90
rect 850 40 910 50
rect 940 90 1000 100
rect 940 50 950 90
rect 950 50 990 90
rect 990 50 1000 90
rect 940 40 1000 50
rect 1030 90 1090 100
rect 1030 50 1040 90
rect 1040 50 1080 90
rect 1080 50 1090 90
rect 1030 40 1090 50
rect 1120 90 1180 100
rect 1120 50 1130 90
rect 1130 50 1170 90
rect 1170 50 1180 90
rect 1120 40 1180 50
rect 1220 90 1280 100
rect 1220 50 1230 90
rect 1230 50 1270 90
rect 1270 50 1280 90
rect 1220 40 1280 50
rect 1310 90 1370 100
rect 1310 50 1320 90
rect 1320 50 1360 90
rect 1360 50 1370 90
rect 1310 40 1370 50
rect 1410 90 1470 100
rect 1410 50 1420 90
rect 1420 50 1460 90
rect 1460 50 1470 90
rect 1410 40 1470 50
rect 1490 90 1550 100
rect 1490 50 1500 90
rect 1500 50 1540 90
rect 1540 50 1550 90
rect 1490 40 1550 50
rect 1580 90 1640 100
rect 1580 50 1590 90
rect 1590 50 1630 90
rect 1630 50 1640 90
rect 1580 40 1640 50
rect 1670 90 1730 100
rect 1670 50 1680 90
rect 1680 50 1720 90
rect 1720 50 1730 90
rect 1670 40 1730 50
rect 1760 90 1820 100
rect 1760 50 1770 90
rect 1770 50 1810 90
rect 1810 50 1820 90
rect 1760 40 1820 50
rect 1850 90 1910 100
rect 1850 50 1860 90
rect 1860 50 1900 90
rect 1900 50 1910 90
rect 1850 40 1910 50
rect 1940 90 2000 100
rect 1940 50 1950 90
rect 1950 50 1990 90
rect 1990 50 2000 90
rect 1940 40 2000 50
rect 2030 90 2090 100
rect 2030 50 2040 90
rect 2040 50 2080 90
rect 2080 50 2090 90
rect 2030 40 2090 50
rect 2120 90 2180 100
rect 2120 50 2130 90
rect 2130 50 2170 90
rect 2170 50 2180 90
rect 2120 40 2180 50
rect 2210 90 2270 100
rect 2210 50 2220 90
rect 2220 50 2260 90
rect 2260 50 2270 90
rect 2210 40 2270 50
rect 2300 90 2360 100
rect 2300 50 2310 90
rect 2310 50 2350 90
rect 2350 50 2360 90
rect 2300 40 2360 50
rect 2390 90 2450 100
rect 2390 50 2400 90
rect 2400 50 2440 90
rect 2440 50 2450 90
rect 2390 40 2450 50
rect 2480 90 2540 100
rect 2480 50 2490 90
rect 2490 50 2530 90
rect 2530 50 2540 90
rect 2480 40 2540 50
rect 2580 90 2640 100
rect 2580 50 2590 90
rect 2590 50 2630 90
rect 2630 50 2640 90
rect 2580 40 2640 50
rect 2670 90 2730 100
rect 2670 50 2680 90
rect 2680 50 2720 90
rect 2720 50 2730 90
rect 2670 40 2730 50
rect 2760 90 2820 100
rect 2760 50 2770 90
rect 2770 50 2810 90
rect 2810 50 2820 90
rect 2760 40 2820 50
rect 2850 90 2910 100
rect 2850 50 2860 90
rect 2860 50 2900 90
rect 2900 50 2910 90
rect 2850 40 2910 50
rect 2940 90 3000 100
rect 2940 50 2950 90
rect 2950 50 2990 90
rect 2990 50 3000 90
rect 2940 40 3000 50
rect 3030 90 3090 100
rect 3030 50 3040 90
rect 3040 50 3080 90
rect 3080 50 3090 90
rect 3030 40 3090 50
rect 3120 90 3180 100
rect 3120 50 3130 90
rect 3130 50 3170 90
rect 3170 50 3180 90
rect 3120 40 3180 50
rect 3210 90 3270 100
rect 3210 50 3220 90
rect 3220 50 3260 90
rect 3260 50 3270 90
rect 3210 40 3270 50
rect 3300 90 3360 100
rect 3300 50 3310 90
rect 3310 50 3350 90
rect 3350 50 3360 90
rect 3300 40 3360 50
rect 3390 90 3450 100
rect 3390 50 3400 90
rect 3400 50 3440 90
rect 3440 50 3450 90
rect 3390 40 3450 50
rect 3480 90 3540 100
rect 3480 50 3490 90
rect 3490 50 3530 90
rect 3530 50 3540 90
rect 3480 40 3540 50
rect 3570 90 3630 100
rect 3570 50 3580 90
rect 3580 50 3620 90
rect 3620 50 3630 90
rect 3570 40 3630 50
rect 3660 90 3720 100
rect 3660 50 3670 90
rect 3670 50 3710 90
rect 3710 50 3720 90
rect 3660 40 3720 50
rect 3750 90 3810 100
rect 3750 50 3760 90
rect 3760 50 3800 90
rect 3800 50 3810 90
rect 3750 40 3810 50
rect 3840 90 3900 100
rect 3840 50 3850 90
rect 3850 50 3890 90
rect 3890 50 3900 90
rect 3840 40 3900 50
rect 3940 90 4000 100
rect 3940 50 3950 90
rect 3950 50 3990 90
rect 3990 50 4000 90
rect 3940 40 4000 50
rect 4030 90 4090 100
rect 4030 50 4040 90
rect 4040 50 4080 90
rect 4080 50 4090 90
rect 4030 40 4090 50
rect 4120 90 4180 100
rect 4120 50 4130 90
rect 4130 50 4170 90
rect 4170 50 4180 90
rect 4120 40 4180 50
rect 4210 90 4270 100
rect 4210 50 4220 90
rect 4220 50 4260 90
rect 4260 50 4270 90
rect 4210 40 4270 50
rect 4300 90 4360 100
rect 4300 50 4310 90
rect 4310 50 4350 90
rect 4350 50 4360 90
rect 4300 40 4360 50
rect 4390 90 4450 100
rect 4390 50 4400 90
rect 4400 50 4440 90
rect 4440 50 4450 90
rect 4390 40 4450 50
rect 4480 90 4540 100
rect 4480 50 4490 90
rect 4490 50 4530 90
rect 4530 50 4540 90
rect 4480 40 4540 50
rect 4570 90 4630 100
rect 4570 50 4580 90
rect 4580 50 4620 90
rect 4620 50 4630 90
rect 4570 40 4630 50
rect 4660 90 4720 100
rect 4660 50 4670 90
rect 4670 50 4710 90
rect 4710 50 4720 90
rect 4660 40 4720 50
rect 4750 90 4810 100
rect 4750 50 4760 90
rect 4760 50 4800 90
rect 4800 50 4810 90
rect 4750 40 4810 50
rect 4840 90 4900 100
rect 4840 50 4850 90
rect 4850 50 4890 90
rect 4890 50 4900 90
rect 4840 40 4900 50
rect 4930 90 4990 100
rect 4930 50 4940 90
rect 4940 50 4980 90
rect 4980 50 4990 90
rect 4930 40 4990 50
rect 5020 90 5080 100
rect 5020 50 5030 90
rect 5030 50 5070 90
rect 5070 50 5080 90
rect 5020 40 5080 50
rect 5110 90 5170 100
rect 5110 50 5120 90
rect 5120 50 5160 90
rect 5160 50 5170 90
rect 5110 40 5170 50
rect 5200 90 5260 100
rect 5200 50 5210 90
rect 5210 50 5250 90
rect 5250 50 5260 90
rect 5200 40 5260 50
rect 5300 90 5360 100
rect 5300 50 5310 90
rect 5310 50 5350 90
rect 5350 50 5360 90
rect 5300 40 5360 50
rect 5390 90 5450 100
rect 5390 50 5400 90
rect 5400 50 5440 90
rect 5440 50 5450 90
rect 5390 40 5450 50
rect 5480 90 5540 100
rect 5480 50 5490 90
rect 5490 50 5530 90
rect 5530 50 5540 90
rect 5480 40 5540 50
rect 5570 90 5630 100
rect 5570 50 5580 90
rect 5580 50 5620 90
rect 5620 50 5630 90
rect 5570 40 5630 50
rect 5660 90 5720 100
rect 5660 50 5670 90
rect 5670 50 5710 90
rect 5710 50 5720 90
rect 5660 40 5720 50
rect 5750 90 5810 100
rect 5750 50 5760 90
rect 5760 50 5800 90
rect 5800 50 5810 90
rect 5750 40 5810 50
rect 5840 90 5900 100
rect 5840 50 5850 90
rect 5850 50 5890 90
rect 5890 50 5900 90
rect 5840 40 5900 50
rect 5930 90 5990 100
rect 5930 50 5940 90
rect 5940 50 5980 90
rect 5980 50 5990 90
rect 5930 40 5990 50
rect 6020 90 6080 100
rect 6020 50 6030 90
rect 6030 50 6070 90
rect 6070 50 6080 90
rect 6020 40 6080 50
rect 6110 90 6170 100
rect 6110 50 6120 90
rect 6120 50 6160 90
rect 6160 50 6170 90
rect 6110 40 6170 50
rect 6200 90 6260 100
rect 6200 50 6210 90
rect 6210 50 6250 90
rect 6250 50 6260 90
rect 6200 40 6260 50
rect 6290 90 6350 100
rect 6290 50 6300 90
rect 6300 50 6340 90
rect 6340 50 6350 90
rect 6290 40 6350 50
rect 6380 90 6440 100
rect 6380 50 6390 90
rect 6390 50 6430 90
rect 6430 50 6440 90
rect 6380 40 6440 50
rect 6470 90 6530 100
rect 6470 50 6480 90
rect 6480 50 6520 90
rect 6520 50 6530 90
rect 6470 40 6530 50
rect 6560 90 6620 100
rect 6560 50 6570 90
rect 6570 50 6610 90
rect 6610 50 6620 90
rect 6560 40 6620 50
rect 6650 90 6710 100
rect 6650 50 6660 90
rect 6660 50 6700 90
rect 6700 50 6710 90
rect 6650 40 6710 50
rect 6750 90 6810 100
rect 6750 50 6760 90
rect 6760 50 6800 90
rect 6800 50 6810 90
rect 6750 40 6810 50
rect 6840 90 6900 100
rect 6840 50 6850 90
rect 6850 50 6890 90
rect 6890 50 6900 90
rect 6840 40 6900 50
rect 6930 90 6990 100
rect 6930 50 6940 90
rect 6940 50 6980 90
rect 6980 50 6990 90
rect 6930 40 6990 50
rect 7020 90 7080 100
rect 7020 50 7030 90
rect 7030 50 7070 90
rect 7070 50 7080 90
rect 7020 40 7080 50
rect 7110 90 7170 100
rect 7110 50 7120 90
rect 7120 50 7160 90
rect 7160 50 7170 90
rect 7110 40 7170 50
rect 7200 90 7260 100
rect 7200 50 7210 90
rect 7210 50 7250 90
rect 7250 50 7260 90
rect 7200 40 7260 50
rect 7290 90 7350 100
rect 7290 50 7300 90
rect 7300 50 7340 90
rect 7340 50 7350 90
rect 7290 40 7350 50
rect 7380 90 7440 100
rect 7380 50 7390 90
rect 7390 50 7430 90
rect 7430 50 7440 90
rect 7380 40 7440 50
rect 7470 90 7530 100
rect 7470 50 7480 90
rect 7480 50 7520 90
rect 7520 50 7530 90
rect 7470 40 7530 50
rect 7560 90 7620 100
rect 7560 50 7570 90
rect 7570 50 7610 90
rect 7610 50 7620 90
rect 7560 40 7620 50
rect 7650 90 7710 100
rect 7650 50 7660 90
rect 7660 50 7700 90
rect 7700 50 7710 90
rect 7650 40 7710 50
rect 7740 90 7800 100
rect 7740 50 7750 90
rect 7750 50 7790 90
rect 7790 50 7800 90
rect 7740 40 7800 50
rect 7830 90 7890 100
rect 7830 50 7840 90
rect 7840 50 7880 90
rect 7880 50 7890 90
rect 7830 40 7890 50
rect 7920 90 7980 100
rect 7920 50 7930 90
rect 7930 50 7970 90
rect 7970 50 7980 90
rect 7920 40 7980 50
rect 8010 90 8070 100
rect 8010 50 8020 90
rect 8020 50 8060 90
rect 8060 50 8070 90
rect 8010 40 8070 50
rect 8110 90 8170 100
rect 8110 50 8120 90
rect 8120 50 8160 90
rect 8160 50 8170 90
rect 8110 40 8170 50
rect 8200 90 8260 100
rect 8200 50 8210 90
rect 8210 50 8250 90
rect 8250 50 8260 90
rect 8200 40 8260 50
rect 8290 90 8350 100
rect 8290 50 8300 90
rect 8300 50 8340 90
rect 8340 50 8350 90
rect 8290 40 8350 50
rect 8380 90 8440 100
rect 8380 50 8390 90
rect 8390 50 8430 90
rect 8430 50 8440 90
rect 8380 40 8440 50
rect 8470 90 8530 100
rect 8470 50 8480 90
rect 8480 50 8520 90
rect 8520 50 8530 90
rect 8470 40 8530 50
rect 8560 90 8620 100
rect 8560 50 8570 90
rect 8570 50 8610 90
rect 8610 50 8620 90
rect 8560 40 8620 50
rect 8650 90 8710 100
rect 8650 50 8660 90
rect 8660 50 8700 90
rect 8700 50 8710 90
rect 8650 40 8710 50
rect 8740 90 8800 100
rect 8740 50 8750 90
rect 8750 50 8790 90
rect 8790 50 8800 90
rect 8740 40 8800 50
rect 8830 90 8890 100
rect 8830 50 8840 90
rect 8840 50 8880 90
rect 8880 50 8890 90
rect 8830 40 8890 50
rect 8920 90 8980 100
rect 8920 50 8930 90
rect 8930 50 8970 90
rect 8970 50 8980 90
rect 8920 40 8980 50
rect 9010 90 9070 100
rect 9010 50 9020 90
rect 9020 50 9060 90
rect 9060 50 9070 90
rect 9010 40 9070 50
rect 9100 90 9160 100
rect 9100 50 9110 90
rect 9110 50 9150 90
rect 9150 50 9160 90
rect 9100 40 9160 50
rect 9190 90 9250 100
rect 9190 50 9200 90
rect 9200 50 9240 90
rect 9240 50 9250 90
rect 9190 40 9250 50
rect 9280 90 9340 100
rect 9280 50 9290 90
rect 9290 50 9330 90
rect 9330 50 9340 90
rect 9280 40 9340 50
rect 9380 90 9440 100
rect 9380 50 9390 90
rect 9390 50 9430 90
rect 9430 50 9440 90
rect 9380 40 9440 50
<< metal2 >>
rect -260 5810 -180 5820
rect -260 5750 -250 5810
rect -190 5750 -180 5810
rect -260 5740 -180 5750
rect 9660 5810 9740 5820
rect 9660 5750 9670 5810
rect 9730 5750 9740 5810
rect 9660 5740 9740 5750
rect -260 5560 -180 5570
rect -260 5500 -250 5560
rect -190 5550 -180 5560
rect 4620 5560 4700 5570
rect 4620 5550 4630 5560
rect -190 5510 4630 5550
rect -190 5500 -180 5510
rect -260 5490 -180 5500
rect 4620 5500 4630 5510
rect 4690 5550 4700 5560
rect 5020 5560 5100 5570
rect 5020 5550 5030 5560
rect 4690 5510 5030 5550
rect 4690 5500 4700 5510
rect 4620 5490 4700 5500
rect 5020 5500 5030 5510
rect 5090 5550 5100 5560
rect 5420 5560 5500 5570
rect 5420 5550 5430 5560
rect 5090 5510 5430 5550
rect 5090 5500 5100 5510
rect 5020 5490 5100 5500
rect 5420 5500 5430 5510
rect 5490 5550 5500 5560
rect 5820 5560 5900 5570
rect 5820 5550 5830 5560
rect 5490 5510 5830 5550
rect 5490 5500 5500 5510
rect 5420 5490 5500 5500
rect 5820 5500 5830 5510
rect 5890 5550 5900 5560
rect 6220 5560 6300 5570
rect 6220 5550 6230 5560
rect 5890 5510 6230 5550
rect 5890 5500 5900 5510
rect 5820 5490 5900 5500
rect 6220 5500 6230 5510
rect 6290 5550 6300 5560
rect 6620 5560 6700 5570
rect 6620 5550 6630 5560
rect 6290 5510 6630 5550
rect 6290 5500 6300 5510
rect 6220 5490 6300 5500
rect 6620 5500 6630 5510
rect 6690 5550 6700 5560
rect 7020 5560 7100 5570
rect 7020 5550 7030 5560
rect 6690 5510 7030 5550
rect 6690 5500 6700 5510
rect 6620 5490 6700 5500
rect 7020 5500 7030 5510
rect 7090 5550 7100 5560
rect 7420 5560 7500 5570
rect 7420 5550 7430 5560
rect 7090 5510 7430 5550
rect 7090 5500 7100 5510
rect 7020 5490 7100 5500
rect 7420 5500 7430 5510
rect 7490 5550 7500 5560
rect 7820 5560 7900 5570
rect 7820 5550 7830 5560
rect 7490 5510 7830 5550
rect 7490 5500 7500 5510
rect 7420 5490 7500 5500
rect 7820 5500 7830 5510
rect 7890 5550 7900 5560
rect 8220 5560 8300 5570
rect 8220 5550 8230 5560
rect 7890 5510 8230 5550
rect 7890 5500 7900 5510
rect 7820 5490 7900 5500
rect 8220 5500 8230 5510
rect 8290 5550 8300 5560
rect 9660 5560 9740 5570
rect 9660 5550 9670 5560
rect 8290 5510 9670 5550
rect 8290 5500 8300 5510
rect 8220 5490 8300 5500
rect 9660 5500 9670 5510
rect 9730 5500 9740 5560
rect 9660 5490 9740 5500
rect -110 5040 1970 5050
rect -110 4980 -100 5040
rect -40 4980 1900 5040
rect 1960 4980 1970 5040
rect -110 4970 1970 4980
rect 4300 4620 4380 4630
rect 4300 4560 4310 4620
rect 4370 4610 4380 4620
rect 4820 4620 4900 4630
rect 4820 4610 4830 4620
rect 4370 4570 4830 4610
rect 4370 4560 4380 4570
rect 4300 4550 4380 4560
rect 4820 4560 4830 4570
rect 4890 4610 4900 4620
rect 6820 4620 6900 4630
rect 6820 4610 6830 4620
rect 4890 4570 6830 4610
rect 4890 4560 4900 4570
rect 4820 4550 4900 4560
rect 6820 4560 6830 4570
rect 6890 4610 6900 4620
rect 7620 4620 7700 4630
rect 7620 4610 7630 4620
rect 6890 4570 7630 4610
rect 6890 4560 6900 4570
rect 6820 4550 6900 4560
rect 7620 4560 7630 4570
rect 7690 4560 7700 4620
rect 7620 4550 7700 4560
rect 8140 4620 8220 4630
rect 8140 4560 8150 4620
rect 8210 4610 8220 4620
rect 8750 4620 8830 4630
rect 8750 4610 8760 4620
rect 8210 4570 8760 4610
rect 8210 4560 8220 4570
rect 8140 4550 8220 4560
rect 8750 4560 8760 4570
rect 8820 4560 8830 4620
rect 8750 4550 8830 4560
rect 5220 4530 5300 4540
rect 5220 4470 5230 4530
rect 5290 4520 5300 4530
rect 6020 4530 6100 4540
rect 6020 4520 6030 4530
rect 5290 4480 6030 4520
rect 5290 4470 5300 4480
rect 5220 4460 5300 4470
rect 6020 4470 6030 4480
rect 6090 4520 6100 4530
rect 8020 4530 8100 4540
rect 8020 4520 8030 4530
rect 6090 4480 8030 4520
rect 6090 4470 6100 4480
rect 6020 4460 6100 4470
rect 8020 4470 8030 4480
rect 8090 4520 8100 4530
rect 8630 4530 8710 4540
rect 8630 4520 8640 4530
rect 8090 4480 8640 4520
rect 8090 4470 8100 4480
rect 8020 4460 8100 4470
rect 8630 4470 8640 4480
rect 8700 4470 8710 4530
rect 8630 4460 8710 4470
rect 3790 4450 4230 4460
rect 3790 4390 3800 4450
rect 4220 4430 4230 4450
rect 5620 4440 5700 4450
rect 5620 4430 5630 4440
rect 4220 4390 5630 4430
rect 3790 4380 4230 4390
rect 5620 4380 5630 4390
rect 5690 4430 5700 4440
rect 6420 4440 6500 4450
rect 6420 4430 6430 4440
rect 5690 4390 6430 4430
rect 5690 4380 5700 4390
rect 5620 4370 5700 4380
rect 6420 4380 6430 4390
rect 6490 4430 6500 4440
rect 7220 4440 7300 4450
rect 7220 4430 7230 4440
rect 6490 4390 7230 4430
rect 6490 4380 6500 4390
rect 6420 4370 6500 4380
rect 7220 4380 7230 4390
rect 7290 4380 7300 4440
rect 7220 4370 7300 4380
rect -260 4320 -180 4330
rect -260 4260 -250 4320
rect -190 4310 -180 4320
rect 5220 4320 5300 4330
rect 5220 4310 5230 4320
rect -190 4270 5230 4310
rect -190 4260 -180 4270
rect -260 4250 -180 4260
rect 5220 4260 5230 4270
rect 5290 4310 5300 4320
rect 5620 4320 5700 4330
rect 5620 4310 5630 4320
rect 5290 4270 5630 4310
rect 5290 4260 5300 4270
rect 5220 4250 5300 4260
rect 5620 4260 5630 4270
rect 5690 4310 5700 4320
rect 6020 4320 6100 4330
rect 6020 4310 6030 4320
rect 5690 4270 6030 4310
rect 5690 4260 5700 4270
rect 5620 4250 5700 4260
rect 6020 4260 6030 4270
rect 6090 4310 6100 4320
rect 6420 4320 6500 4330
rect 6420 4310 6430 4320
rect 6090 4270 6430 4310
rect 6090 4260 6100 4270
rect 6020 4250 6100 4260
rect 6420 4260 6430 4270
rect 6490 4310 6500 4320
rect 6820 4320 6900 4330
rect 6820 4310 6830 4320
rect 6490 4270 6830 4310
rect 6490 4260 6500 4270
rect 6420 4250 6500 4260
rect 6820 4260 6830 4270
rect 6890 4310 6900 4320
rect 7220 4320 7300 4330
rect 7220 4310 7230 4320
rect 6890 4270 7230 4310
rect 6890 4260 6900 4270
rect 6820 4250 6900 4260
rect 7220 4260 7230 4270
rect 7290 4310 7300 4320
rect 7620 4320 7700 4330
rect 7620 4310 7630 4320
rect 7290 4270 7630 4310
rect 7290 4260 7300 4270
rect 7220 4250 7300 4260
rect 7620 4260 7630 4270
rect 7690 4310 7700 4320
rect 9170 4320 9250 4330
rect 9170 4310 9180 4320
rect 7690 4270 9180 4310
rect 7690 4260 7700 4270
rect 7620 4250 7700 4260
rect 9170 4260 9180 4270
rect 9240 4310 9250 4320
rect 9660 4320 9740 4330
rect 9660 4310 9670 4320
rect 9240 4270 9670 4310
rect 9240 4260 9250 4270
rect 9170 4250 9250 4260
rect 9660 4260 9670 4270
rect 9730 4260 9740 4320
rect 9660 4250 9740 4260
rect -110 4020 1970 4030
rect -110 3960 -100 4020
rect -40 3960 1900 4020
rect 1960 3960 1970 4020
rect -110 3950 1970 3960
rect 5820 3780 5900 3790
rect 5820 3720 5830 3780
rect 5890 3770 5900 3780
rect 6220 3780 6300 3790
rect 6220 3770 6230 3780
rect 5890 3730 6230 3770
rect 5890 3720 5900 3730
rect 5820 3710 5900 3720
rect 6220 3720 6230 3730
rect 6290 3770 6300 3780
rect 6620 3780 6700 3790
rect 6620 3770 6630 3780
rect 6290 3730 6630 3770
rect 6290 3720 6300 3730
rect 6220 3710 6300 3720
rect 6620 3720 6630 3730
rect 6690 3770 6700 3780
rect 7020 3780 7100 3790
rect 7020 3770 7030 3780
rect 6690 3730 7030 3770
rect 6690 3720 6700 3730
rect 6620 3710 6700 3720
rect 7020 3720 7030 3730
rect 7090 3720 7100 3780
rect 7020 3710 7100 3720
rect 5420 3690 5500 3700
rect 5420 3630 5430 3690
rect 5490 3680 5500 3690
rect 5980 3690 6060 3700
rect 5980 3680 5990 3690
rect 5490 3640 5990 3680
rect 5490 3630 5500 3640
rect 5420 3620 5500 3630
rect 5980 3630 5990 3640
rect 6050 3680 6060 3690
rect 6330 3690 6410 3700
rect 6330 3680 6340 3690
rect 6050 3640 6340 3680
rect 6050 3630 6060 3640
rect 5980 3620 6060 3630
rect 6330 3630 6340 3640
rect 6400 3680 6410 3690
rect 6860 3690 6940 3700
rect 6860 3680 6870 3690
rect 6400 3640 6870 3680
rect 6400 3630 6410 3640
rect 6330 3620 6410 3630
rect 6860 3630 6870 3640
rect 6930 3680 6940 3690
rect 7420 3690 7500 3700
rect 7420 3680 7430 3690
rect 6930 3640 7430 3680
rect 6930 3630 6940 3640
rect 6860 3620 6940 3630
rect 7420 3630 7430 3640
rect 7490 3630 7500 3690
rect 7420 3620 7500 3630
rect 6460 3600 6540 3610
rect 6460 3540 6470 3600
rect 6530 3590 6540 3600
rect 8440 3600 8520 3610
rect 8440 3590 8450 3600
rect 6530 3550 8450 3590
rect 6530 3540 6540 3550
rect 6460 3530 6540 3540
rect 8440 3540 8450 3550
rect 8510 3540 8520 3600
rect 8440 3530 8520 3540
rect 5820 3510 5900 3520
rect 5820 3450 5830 3510
rect 5890 3500 5900 3510
rect 5980 3510 6060 3520
rect 5980 3500 5990 3510
rect 5890 3460 5990 3500
rect 5890 3450 5900 3460
rect 5820 3440 5900 3450
rect 5980 3450 5990 3460
rect 6050 3500 6060 3510
rect 6860 3510 6940 3520
rect 6860 3500 6870 3510
rect 6050 3460 6870 3500
rect 6050 3450 6060 3460
rect 5980 3440 6060 3450
rect 6860 3450 6870 3460
rect 6930 3500 6940 3510
rect 7020 3510 7100 3520
rect 7020 3500 7030 3510
rect 6930 3460 7030 3500
rect 6930 3450 6940 3460
rect 6860 3440 6940 3450
rect 7020 3450 7030 3460
rect 7090 3450 7100 3510
rect 7020 3440 7100 3450
rect 880 3430 4230 3440
rect 880 3370 890 3430
rect 950 3370 3800 3430
rect 4220 3410 4230 3430
rect 4300 3420 4380 3440
rect 4300 3410 4310 3420
rect 4220 3370 4310 3410
rect 880 3360 4230 3370
rect 4300 3360 4310 3370
rect 4370 3410 4380 3420
rect 6100 3420 6180 3430
rect 6100 3410 6110 3420
rect 4370 3370 6110 3410
rect 4370 3360 4380 3370
rect 4300 3350 4380 3360
rect 6100 3360 6110 3370
rect 6170 3410 6180 3420
rect 6740 3420 6820 3430
rect 6740 3410 6750 3420
rect 6170 3370 6750 3410
rect 6170 3360 6180 3370
rect 6100 3350 6180 3360
rect 6740 3360 6750 3370
rect 6810 3410 6820 3420
rect 8860 3420 8940 3430
rect 8860 3410 8870 3420
rect 6810 3370 8870 3410
rect 6810 3360 6820 3370
rect 6740 3350 6820 3360
rect 8860 3360 8870 3370
rect 8930 3360 8940 3420
rect 8860 3350 8940 3360
rect 5820 3080 5900 3090
rect 1720 3070 1970 3080
rect 1720 3010 1730 3070
rect 1790 3010 1900 3070
rect 1960 3010 1970 3070
rect 1720 3000 1970 3010
rect 3790 3070 4230 3080
rect 5820 3070 5830 3080
rect 3790 3010 3800 3070
rect 4220 3030 5830 3070
rect 4220 3010 4230 3030
rect 5820 3020 5830 3030
rect 5890 3070 5900 3080
rect 7020 3080 7100 3090
rect 7020 3070 7030 3080
rect 5890 3030 7030 3070
rect 5890 3020 5900 3030
rect 5820 3010 5900 3020
rect 7020 3020 7030 3030
rect 7090 3070 7100 3080
rect 8630 3080 8710 3090
rect 8630 3070 8640 3080
rect 7090 3030 8640 3070
rect 7090 3020 7100 3030
rect 7020 3010 7100 3020
rect 8630 3020 8640 3030
rect 8700 3020 8710 3080
rect 8630 3010 8710 3020
rect 3790 3000 4230 3010
rect 5620 2990 5700 3000
rect 5620 2930 5630 2990
rect 5690 2980 5700 2990
rect 6020 2990 6100 3000
rect 6020 2980 6030 2990
rect 5690 2940 6030 2980
rect 5690 2930 5700 2940
rect 5620 2920 5700 2930
rect 6020 2930 6030 2940
rect 6090 2980 6100 2990
rect 6420 2990 6500 3000
rect 6420 2980 6430 2990
rect 6090 2940 6430 2980
rect 6090 2930 6100 2940
rect 6020 2920 6100 2930
rect 6420 2930 6430 2940
rect 6490 2980 6500 2990
rect 6820 2990 6900 3000
rect 6820 2980 6830 2990
rect 6490 2940 6830 2980
rect 6490 2930 6500 2940
rect 6420 2920 6500 2930
rect 6820 2930 6830 2940
rect 6890 2980 6900 2990
rect 7220 2990 7300 3000
rect 7220 2980 7230 2990
rect 6890 2940 7230 2980
rect 6890 2930 6900 2940
rect 6820 2920 6900 2930
rect 7220 2930 7230 2940
rect 7290 2930 7300 2990
rect 7220 2920 7300 2930
rect 7380 2870 7460 2880
rect 7380 2810 7390 2870
rect 7450 2860 7460 2870
rect 8440 2870 8520 2880
rect 8440 2860 8450 2870
rect 7450 2820 8450 2860
rect 7450 2810 7460 2820
rect 7380 2800 7460 2810
rect 8440 2810 8450 2820
rect 8510 2810 8520 2870
rect 8440 2800 8520 2810
rect -110 2480 1970 2490
rect -110 2420 -100 2480
rect -40 2420 1900 2480
rect 1960 2420 1970 2480
rect -110 2410 1970 2420
rect -110 1930 -30 1940
rect -110 1870 -100 1930
rect -40 1920 -30 1930
rect 6340 1930 6580 1940
rect 6340 1920 6350 1930
rect -40 1880 6350 1920
rect -40 1870 -30 1880
rect -110 1860 -30 1870
rect 6340 1870 6350 1880
rect 6410 1870 6430 1930
rect 6490 1870 6510 1930
rect 6570 1920 6580 1930
rect 9510 1930 9590 1940
rect 9510 1920 9520 1930
rect 6570 1880 9520 1920
rect 6570 1870 6580 1880
rect 6340 1860 6580 1870
rect 9510 1870 9520 1880
rect 9580 1870 9590 1930
rect 9510 1860 9590 1870
rect 7440 1810 7520 1820
rect 7440 1750 7450 1810
rect 7510 1800 7520 1810
rect 8990 1810 9070 1820
rect 8990 1800 9000 1810
rect 7510 1760 9000 1800
rect 7510 1750 7520 1760
rect 7440 1740 7520 1750
rect 8990 1750 9000 1760
rect 9060 1750 9070 1810
rect 8990 1740 9070 1750
rect -110 1650 -30 1660
rect -110 1590 -100 1650
rect -40 1640 -30 1650
rect 1300 1650 1380 1660
rect 1300 1640 1310 1650
rect -40 1600 1310 1640
rect -40 1590 -30 1600
rect -110 1580 -30 1590
rect 1300 1590 1310 1600
rect 1370 1590 1380 1650
rect 1300 1580 1380 1590
rect 7590 1640 7670 1650
rect 7590 1580 7600 1640
rect 7660 1630 7670 1640
rect 9510 1640 9590 1650
rect 9510 1630 9520 1640
rect 7660 1590 9520 1630
rect 7660 1580 7670 1590
rect 7590 1570 7670 1580
rect 9510 1580 9520 1590
rect 9580 1580 9590 1640
rect 9510 1570 9590 1580
rect -110 100 9590 110
rect -110 40 -100 100
rect -40 40 30 100
rect 90 40 130 100
rect 190 40 230 100
rect 290 40 320 100
rect 380 40 400 100
rect 460 40 490 100
rect 550 40 580 100
rect 640 40 670 100
rect 730 40 760 100
rect 820 40 850 100
rect 910 40 940 100
rect 1000 40 1030 100
rect 1090 40 1120 100
rect 1180 40 1220 100
rect 1280 40 1310 100
rect 1370 40 1410 100
rect 1470 40 1490 100
rect 1550 40 1580 100
rect 1640 40 1670 100
rect 1730 40 1760 100
rect 1820 40 1850 100
rect 1910 40 1940 100
rect 2000 40 2030 100
rect 2090 40 2120 100
rect 2180 40 2210 100
rect 2270 40 2300 100
rect 2360 40 2390 100
rect 2450 40 2480 100
rect 2540 40 2580 100
rect 2640 40 2670 100
rect 2730 40 2760 100
rect 2820 40 2850 100
rect 2910 40 2940 100
rect 3000 40 3030 100
rect 3090 40 3120 100
rect 3180 40 3210 100
rect 3270 40 3300 100
rect 3360 40 3390 100
rect 3450 40 3480 100
rect 3540 40 3570 100
rect 3630 40 3660 100
rect 3720 40 3750 100
rect 3810 40 3840 100
rect 3900 40 3940 100
rect 4000 40 4030 100
rect 4090 40 4120 100
rect 4180 40 4210 100
rect 4270 40 4300 100
rect 4360 40 4390 100
rect 4450 40 4480 100
rect 4540 40 4570 100
rect 4630 40 4660 100
rect 4720 40 4750 100
rect 4810 40 4840 100
rect 4900 40 4930 100
rect 4990 40 5020 100
rect 5080 40 5110 100
rect 5170 40 5200 100
rect 5260 40 5300 100
rect 5360 40 5390 100
rect 5450 40 5480 100
rect 5540 40 5570 100
rect 5630 40 5660 100
rect 5720 40 5750 100
rect 5810 40 5840 100
rect 5900 40 5930 100
rect 5990 40 6020 100
rect 6080 40 6110 100
rect 6170 40 6200 100
rect 6260 40 6290 100
rect 6350 40 6380 100
rect 6440 40 6470 100
rect 6530 40 6560 100
rect 6620 40 6650 100
rect 6710 40 6750 100
rect 6810 40 6840 100
rect 6900 40 6930 100
rect 6990 40 7020 100
rect 7080 40 7110 100
rect 7170 40 7200 100
rect 7260 40 7290 100
rect 7350 40 7380 100
rect 7440 40 7470 100
rect 7530 40 7560 100
rect 7620 40 7650 100
rect 7710 40 7740 100
rect 7800 40 7830 100
rect 7890 40 7920 100
rect 7980 40 8010 100
rect 8070 40 8110 100
rect 8170 40 8200 100
rect 8260 40 8290 100
rect 8350 40 8380 100
rect 8440 40 8470 100
rect 8530 40 8560 100
rect 8620 40 8650 100
rect 8710 40 8740 100
rect 8800 40 8830 100
rect 8890 40 8920 100
rect 8980 40 9010 100
rect 9070 40 9100 100
rect 9160 40 9190 100
rect 9250 40 9280 100
rect 9340 40 9380 100
rect 9440 40 9520 100
rect 9580 40 9590 100
rect -110 30 9590 40
rect -260 -180 -180 -170
rect -260 -240 -250 -180
rect -190 -240 -180 -180
rect -260 -250 -180 -240
<< via2 >>
rect -250 5750 -190 5810
rect 9670 5750 9730 5810
rect -250 5500 -190 5560
rect 9670 5500 9730 5560
rect -100 4980 -40 5040
rect -250 4260 -190 4320
rect 9670 4260 9730 4320
rect -100 3960 -40 4020
rect -100 2420 -40 2480
rect -100 1870 -40 1930
rect 9520 1870 9580 1930
rect -100 1590 -40 1650
rect 9520 1580 9580 1640
rect -100 40 -40 100
rect 9520 40 9580 100
rect -250 -240 -190 -180
<< metal3 >>
rect -270 5820 -170 5830
rect -270 5740 -260 5820
rect -180 5740 -170 5820
rect -270 5730 -170 5740
rect 9650 5820 9750 5830
rect 9650 5740 9660 5820
rect 9740 5740 9750 5820
rect 9650 5730 9750 5740
rect -260 5560 -180 5730
rect -120 5670 -20 5680
rect -120 5590 -110 5670
rect -30 5590 -20 5670
rect -120 5580 -20 5590
rect 9500 5670 9600 5680
rect 9500 5590 9510 5670
rect 9590 5590 9600 5670
rect 9500 5580 9600 5590
rect -260 5500 -250 5560
rect -190 5500 -180 5560
rect -260 4320 -180 5500
rect -260 4260 -250 4320
rect -190 4260 -180 4320
rect -260 -160 -180 4260
rect -110 5040 -30 5580
rect -110 4980 -100 5040
rect -40 4980 -30 5040
rect -110 4020 -30 4980
rect -110 3960 -100 4020
rect -40 3960 -30 4020
rect -110 2480 -30 3960
rect -110 2420 -100 2480
rect -40 2420 -30 2480
rect -110 1930 -30 2420
rect -110 1870 -100 1930
rect -40 1870 -30 1930
rect -110 1650 -30 1870
rect -110 1590 -100 1650
rect -40 1590 -30 1650
rect -110 100 -30 1590
rect -110 40 -100 100
rect -40 40 -30 100
rect -110 -10 -30 40
rect 9510 1930 9590 5580
rect 9510 1870 9520 1930
rect 9580 1870 9590 1930
rect 9510 1640 9590 1870
rect 9510 1580 9520 1640
rect 9580 1580 9590 1640
rect 9510 100 9590 1580
rect 9510 40 9520 100
rect 9580 40 9590 100
rect 9510 -10 9590 40
rect 9660 5560 9740 5730
rect 9660 5500 9670 5560
rect 9730 5500 9740 5560
rect 9660 4320 9740 5500
rect 9660 4260 9670 4320
rect 9730 4260 9740 4320
rect -120 -20 -20 -10
rect -120 -100 -110 -20
rect -30 -100 -20 -20
rect -120 -110 -20 -100
rect 9500 -20 9600 -10
rect 9500 -100 9510 -20
rect 9590 -100 9600 -20
rect 9500 -110 9600 -100
rect 9660 -160 9740 4260
rect -270 -170 -170 -160
rect -270 -250 -260 -170
rect -180 -250 -170 -170
rect -270 -260 -170 -250
rect 9650 -170 9750 -160
rect 9650 -250 9660 -170
rect 9740 -250 9750 -170
rect 9650 -260 9750 -250
<< via3 >>
rect -260 5810 -180 5820
rect -260 5750 -250 5810
rect -250 5750 -190 5810
rect -190 5750 -180 5810
rect -260 5740 -180 5750
rect 9660 5810 9740 5820
rect 9660 5750 9670 5810
rect 9670 5750 9730 5810
rect 9730 5750 9740 5810
rect 9660 5740 9740 5750
rect -110 5590 -30 5670
rect 9510 5590 9590 5670
rect -110 -100 -30 -20
rect 9510 -100 9590 -20
rect -260 -180 -180 -170
rect -260 -240 -250 -180
rect -250 -240 -190 -180
rect -190 -240 -180 -180
rect -260 -250 -180 -240
rect 9660 -250 9740 -170
<< metal4 >>
rect -270 5820 -170 5830
rect 9650 5820 9750 5830
rect -270 5740 -260 5820
rect -180 5740 9660 5820
rect 9740 5740 9750 5820
rect -270 5730 -170 5740
rect 9650 5730 9750 5740
rect -120 5670 -20 5680
rect 9500 5670 9600 5680
rect -120 5590 -110 5670
rect -30 5590 9510 5670
rect 9590 5590 9600 5670
rect -120 5580 -20 5590
rect 9500 5580 9600 5590
rect -120 -20 -20 -10
rect 9500 -20 9600 -10
rect -120 -100 -110 -20
rect -30 -100 9510 -20
rect 9590 -100 9600 -20
rect -120 -110 -20 -100
rect 9500 -110 9600 -100
rect -270 -170 -170 -160
rect 9650 -170 9750 -160
rect -270 -250 -260 -170
rect -180 -250 9660 -170
rect 9740 -250 9750 -170
rect -270 -260 -170 -250
rect 9650 -260 9750 -250
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0 $PDKPATH/libs.ref/sky130_fd_pr/mag
timestamp 1723858470
transform 1 0 2710 0 1 0
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_1
timestamp 1723858470
transform 1 0 -10 0 1 0
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_2
timestamp 1723858470
transform 1 0 1350 0 1 0
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_3
timestamp 1723858470
transform 1 0 2710 0 1 0
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_4
timestamp 1723858470
transform 1 0 4070 0 1 0
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5
timestamp 1723858470
transform 1 0 5430 0 1 0
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_6
timestamp 1723858470
transform 1 0 6790 0 1 0
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_7
timestamp 1723858470
transform 1 0 4070 0 1 0
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8
timestamp 1723858470
transform 1 0 5430 0 1 0
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_9
timestamp 1723858470
transform 1 0 6790 0 1 0
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_10
timestamp 1723858470
transform 1 0 8150 0 1 0
box 0 0 1340 1340
<< labels >>
flabel locali s 8740 1102 8858 1142 0 FreeSans 400 0 0 0 Base
port 4 nsew
flabel locali s 8763 1252 8864 1301 0 FreeSans 400 0 0 0 Collector
port 3 nsew
flabel locali s 8704 626 8952 730 0 FreeSans 400 0 0 0 Emitter
port 2 nsew
flabel locali s 7380 1102 7498 1142 0 FreeSans 400 0 0 0 Base
port 4 nsew
flabel locali s 7403 1252 7504 1301 0 FreeSans 400 0 0 0 Collector
port 3 nsew
flabel locali s 7344 626 7592 730 0 FreeSans 400 0 0 0 Emitter
port 2 nsew
flabel locali s 6020 1102 6138 1142 0 FreeSans 400 0 0 0 Base
port 4 nsew
flabel locali s 6043 1252 6144 1301 0 FreeSans 400 0 0 0 Collector
port 3 nsew
flabel locali s 5984 626 6232 730 0 FreeSans 400 0 0 0 Emitter
port 2 nsew
flabel locali s 4660 1102 4778 1142 0 FreeSans 400 0 0 0 Base
port 4 nsew
flabel locali s 4683 1252 4784 1301 0 FreeSans 400 0 0 0 Collector
port 3 nsew
flabel locali s 4624 626 4872 730 0 FreeSans 400 0 0 0 Emitter
port 2 nsew
flabel locali s 3300 1102 3418 1142 0 FreeSans 400 0 0 0 Base
port 4 nsew
flabel locali s 3323 1252 3424 1301 0 FreeSans 400 0 0 0 Collector
port 3 nsew
flabel locali s 3264 626 3512 730 0 FreeSans 400 0 0 0 Emitter
port 2 nsew
flabel locali s 1940 1102 2058 1142 0 FreeSans 400 0 0 0 Base
port 4 nsew
flabel locali s 1963 1252 2064 1301 0 FreeSans 400 0 0 0 Collector
port 3 nsew
flabel locali s 1904 626 2152 730 0 FreeSans 400 0 0 0 Emitter
port 2 nsew
flabel metal3 9740 2800 9740 2800 3 FreeSans 1600 0 160 0 VDDA
port 1 e
flabel metal3 9590 2350 9590 2350 3 FreeSans 1600 0 160 0 GNDA
port 6 e
flabel metal1 6460 6300 6460 6300 1 FreeSans 1600 0 0 800 V_out
port 5 n
flabel metal1 1800 2080 1800 2080 3 FreeSans 800 0 160 0 Vbe2
flabel metal1 9050 3230 9050 3230 3 FreeSans 800 0 160 0 start_up
flabel locali 5640 2900 5640 2900 7 FreeSans 800 0 -160 0 V_p
flabel metal2 4570 3370 4570 3370 5 FreeSans 800 0 0 -160 Vin-
flabel metal2 4570 3030 4570 3030 5 FreeSans 800 0 0 -160 Vin+
flabel metal1 8830 4590 8830 4590 3 FreeSans 800 0 160 0 V_TOP
flabel metal2 7500 3660 7500 3660 3 FreeSans 800 0 160 0 1st_Vout
flabel metal1 6240 3580 6240 3580 7 FreeSans 800 0 -160 0 V_mirror
<< end >>
