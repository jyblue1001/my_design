magic
tech sky130A
timestamp 1738167617
<< nwell >>
rect 480 190 865 430
<< pwell >>
rect 565 -10 865 115
rect 575 -15 865 -10
<< nmos >>
rect 700 0 715 100
<< pmos >>
rect 700 210 715 410
<< ndiff >>
rect 650 85 700 100
rect 650 15 665 85
rect 685 15 700 85
rect 650 0 700 15
rect 715 85 765 100
rect 715 15 730 85
rect 750 15 765 85
rect 715 0 765 15
<< pdiff >>
rect 650 395 700 410
rect 650 225 665 395
rect 685 225 700 395
rect 650 210 700 225
rect 715 395 765 410
rect 715 225 730 395
rect 750 225 765 395
rect 715 210 765 225
<< ndiffc >>
rect 665 15 685 85
rect 730 15 750 85
<< pdiffc >>
rect 665 225 685 395
rect 730 225 750 395
<< psubdiff >>
rect 570 85 620 100
rect 570 15 585 85
rect 605 15 620 85
rect 570 0 620 15
<< nsubdiff >>
rect 795 395 845 410
rect 795 225 810 395
rect 830 225 845 395
rect 795 210 845 225
<< psubdiffcont >>
rect 585 15 605 85
<< nsubdiffcont >>
rect 810 225 830 395
<< poly >>
rect 685 455 725 465
rect 685 435 695 455
rect 715 435 725 455
rect 685 425 725 435
rect 700 410 715 425
rect 565 370 605 380
rect 565 350 575 370
rect 595 350 605 370
rect 565 340 605 350
rect 700 195 715 210
rect 700 100 715 115
rect 810 30 850 40
rect 810 10 820 30
rect 840 10 850 30
rect 810 0 850 10
rect 700 -15 715 0
rect 685 -25 725 -15
rect 685 -45 695 -25
rect 715 -45 725 -25
rect 685 -55 725 -45
<< polycont >>
rect 695 435 715 455
rect 575 350 595 370
rect 820 10 840 30
rect 695 -45 715 -25
<< locali >>
rect 685 455 725 465
rect 685 435 695 455
rect 715 435 725 455
rect 685 425 725 435
rect 655 395 695 405
rect 565 370 605 380
rect 565 350 575 370
rect 595 350 605 370
rect 565 340 605 350
rect 585 95 605 340
rect 655 225 665 395
rect 685 225 695 395
rect 655 215 695 225
rect 720 395 765 405
rect 720 225 730 395
rect 750 225 765 395
rect 720 215 765 225
rect 795 395 840 405
rect 795 225 810 395
rect 830 225 840 395
rect 795 215 840 225
rect 665 195 685 215
rect 660 175 685 195
rect 665 95 685 175
rect 730 135 750 215
rect 730 115 755 135
rect 730 95 750 115
rect 575 85 620 95
rect 575 15 585 85
rect 605 15 620 85
rect 575 5 620 15
rect 650 85 695 95
rect 650 15 665 85
rect 685 15 695 85
rect 650 5 695 15
rect 720 85 760 95
rect 720 15 730 85
rect 750 15 760 85
rect 720 5 760 15
rect 810 40 830 215
rect 810 30 850 40
rect 810 10 820 30
rect 840 10 850 30
rect 810 0 850 10
rect 685 -25 725 -15
rect 685 -45 695 -25
rect 715 -45 725 -25
rect 685 -55 725 -45
<< viali >>
rect 695 435 715 455
rect 575 350 595 370
rect 820 10 840 30
rect 695 -45 715 -25
<< metal1 >>
rect 480 455 850 465
rect 480 435 695 455
rect 715 435 850 455
rect 480 370 850 435
rect 480 350 575 370
rect 595 350 850 370
rect 480 210 850 350
rect 480 30 850 100
rect 480 10 820 30
rect 840 10 850 30
rect 480 -25 850 10
rect 480 -45 695 -25
rect 715 -45 850 -25
rect 480 -55 850 -45
<< labels >>
flabel metal1 480 315 480 320 7 FreeSans 400 0 -80 0 VDDA
flabel metal1 480 20 480 25 7 FreeSans 400 0 -80 0 GNDA
flabel locali 660 185 660 185 7 FreeSans 400 0 -80 0 A
flabel locali 755 125 755 125 3 FreeSans 400 0 80 0 B
<< end >>
