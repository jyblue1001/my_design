magic
tech sky130A
timestamp 1752750078
<< error_p >>
rect 810 205 880 214
rect 810 191 880 200
rect 1845 -335 1859 -326
rect 1831 -349 1845 -340
rect 845 -1290 855 -1281
rect 845 -1295 849 -1290
rect 845 -1304 855 -1295
<< nwell >>
rect -30 2305 310 2695
rect 440 2305 780 2525
rect 910 2305 1250 2695
rect 1380 2305 1720 2695
rect -1225 1730 -345 2120
rect -100 1730 780 2120
rect 910 1730 1790 2120
rect 2035 1730 2915 2120
rect -1195 815 -375 1455
rect 395 1215 1295 1505
rect 2065 815 2885 1455
rect -1195 400 -375 640
rect 2065 400 2885 640
<< nmos >>
rect -65 700 -50 850
rect -10 700 5 850
rect 45 700 60 850
rect 100 700 115 850
rect 155 700 170 850
rect 210 700 225 850
rect 265 700 280 850
rect 320 700 335 850
rect 375 700 390 850
rect 430 700 445 850
rect 485 700 500 850
rect 540 700 555 850
rect 755 625 770 875
rect 810 625 825 875
rect 865 625 880 875
rect 920 625 935 875
rect 1135 700 1150 850
rect 1190 700 1205 850
rect 1245 700 1260 850
rect 1300 700 1315 850
rect 1355 700 1370 850
rect 1410 700 1425 850
rect 1465 700 1480 850
rect 1520 700 1535 850
rect 1575 700 1590 850
rect 1630 700 1645 850
rect 1685 700 1700 850
rect 1740 700 1755 850
rect -65 280 -50 430
rect -10 280 5 430
rect 45 280 60 430
rect 100 280 115 430
rect 155 280 170 430
rect 210 280 225 430
rect 265 280 280 430
rect 320 280 335 430
rect 375 280 390 430
rect 430 280 445 430
rect 485 280 500 430
rect 540 280 555 430
rect 755 280 770 430
rect 810 280 825 430
rect 865 280 880 430
rect 920 280 935 430
rect 1135 280 1150 430
rect 1190 280 1205 430
rect 1245 280 1260 430
rect 1300 280 1315 430
rect 1355 280 1370 430
rect 1410 280 1425 430
rect 1465 280 1480 430
rect 1520 280 1535 430
rect 1575 280 1590 430
rect 1630 280 1645 430
rect 1685 280 1700 430
rect 1740 280 1755 430
rect -1095 -70 -1080 230
rect -1040 -70 -1025 230
rect -985 -70 -970 230
rect -930 -70 -915 230
rect -875 -70 -860 230
rect -820 -70 -805 230
rect -765 -70 -750 230
rect -710 -70 -695 230
rect -655 -70 -640 230
rect -600 -70 -585 230
rect -545 -70 -530 230
rect -490 -70 -475 230
rect 755 -315 770 -65
rect 810 -315 825 -65
rect 865 -315 880 -65
rect 920 -315 935 -65
rect 2165 -70 2180 230
rect 2220 -70 2235 230
rect 2275 -70 2290 230
rect 2330 -70 2345 230
rect 2385 -70 2400 230
rect 2440 -70 2455 230
rect 2495 -70 2510 230
rect 2550 -70 2565 230
rect 2605 -70 2620 230
rect 2660 -70 2675 230
rect 2715 -70 2730 230
rect 2770 -70 2785 230
rect -1065 -1055 -1005 -355
rect -965 -1055 -905 -355
rect -865 -1055 -805 -355
rect -765 -1055 -705 -355
rect -665 -1055 -605 -355
rect -565 -1055 -505 -355
rect 315 -785 330 -535
rect 370 -785 385 -535
rect 425 -785 440 -535
rect 480 -785 495 -535
rect 535 -785 550 -535
rect 590 -785 605 -535
rect 645 -785 660 -535
rect 700 -785 715 -535
rect 755 -785 770 -535
rect 810 -785 825 -535
rect 865 -785 880 -535
rect 920 -785 935 -535
rect 975 -785 990 -535
rect 1030 -785 1045 -535
rect 1085 -785 1100 -535
rect 1140 -785 1155 -535
rect 1195 -785 1210 -535
rect 1250 -785 1265 -535
rect 1305 -785 1320 -535
rect 1360 -785 1375 -535
rect 1415 -785 1430 -535
rect 525 -1160 540 -1010
rect 580 -1160 595 -1010
rect 635 -1160 650 -1010
rect 690 -1160 705 -1010
rect 745 -1160 760 -1010
rect 800 -1160 815 -1010
rect 965 -1160 1265 -1010
rect 2195 -1055 2255 -355
rect 2295 -1055 2355 -355
rect 2395 -1055 2455 -355
rect 2495 -1055 2555 -355
rect 2595 -1055 2655 -355
rect 2695 -1055 2755 -355
<< pmos >>
rect 70 2325 90 2675
rect 130 2325 150 2675
rect 190 2325 210 2675
rect 540 2325 560 2505
rect 600 2325 620 2505
rect 660 2325 680 2505
rect 1010 2325 1030 2675
rect 1070 2325 1090 2675
rect 1130 2325 1150 2675
rect 1480 2325 1500 2675
rect 1540 2325 1560 2675
rect 1600 2325 1620 2675
rect -1125 1750 -1105 2100
rect -1065 1750 -1045 2100
rect -1005 1750 -985 2100
rect -945 1750 -925 2100
rect -885 1750 -865 2100
rect -825 1750 -805 2100
rect -765 1750 -745 2100
rect -705 1750 -685 2100
rect -645 1750 -625 2100
rect -585 1750 -565 2100
rect -525 1750 -505 2100
rect -465 1750 -445 2100
rect 0 1750 20 2100
rect 60 1750 80 2100
rect 120 1750 140 2100
rect 180 1750 200 2100
rect 240 1750 260 2100
rect 300 1750 320 2100
rect 360 1750 380 2100
rect 420 1750 440 2100
rect 480 1750 500 2100
rect 540 1750 560 2100
rect 600 1750 620 2100
rect 660 1750 680 2100
rect 1010 1750 1030 2100
rect 1070 1750 1090 2100
rect 1130 1750 1150 2100
rect 1190 1750 1210 2100
rect 1250 1750 1270 2100
rect 1310 1750 1330 2100
rect 1370 1750 1390 2100
rect 1430 1750 1450 2100
rect 1490 1750 1510 2100
rect 1550 1750 1570 2100
rect 1610 1750 1630 2100
rect 1670 1750 1690 2100
rect 2135 1750 2155 2100
rect 2195 1750 2215 2100
rect 2255 1750 2275 2100
rect 2315 1750 2335 2100
rect 2375 1750 2395 2100
rect 2435 1750 2455 2100
rect 2495 1750 2515 2100
rect 2555 1750 2575 2100
rect 2615 1750 2635 2100
rect 2675 1750 2695 2100
rect 2735 1750 2755 2100
rect 2795 1750 2815 2100
rect -1095 835 -1080 1435
rect -1040 835 -1025 1435
rect -985 835 -970 1435
rect -930 835 -915 1435
rect -875 835 -860 1435
rect -820 835 -805 1435
rect -765 835 -750 1435
rect -710 835 -695 1435
rect -655 835 -640 1435
rect -600 835 -585 1435
rect -545 835 -530 1435
rect -490 835 -475 1435
rect 495 1235 510 1485
rect 550 1235 565 1485
rect 605 1235 620 1485
rect 660 1235 675 1485
rect 715 1235 730 1485
rect 770 1235 785 1485
rect 905 1235 920 1485
rect 960 1235 975 1485
rect 1015 1235 1030 1485
rect 1070 1235 1085 1485
rect 1125 1235 1140 1485
rect 1180 1235 1195 1485
rect 2165 835 2180 1435
rect 2220 835 2235 1435
rect 2275 835 2290 1435
rect 2330 835 2345 1435
rect 2385 835 2400 1435
rect 2440 835 2455 1435
rect 2495 835 2510 1435
rect 2550 835 2565 1435
rect 2605 835 2620 1435
rect 2660 835 2675 1435
rect 2715 835 2730 1435
rect 2770 835 2785 1435
rect -1095 420 -1080 620
rect -1040 420 -1025 620
rect -985 420 -970 620
rect -930 420 -915 620
rect -875 420 -860 620
rect -820 420 -805 620
rect -765 420 -750 620
rect -710 420 -695 620
rect -655 420 -640 620
rect -600 420 -585 620
rect -545 420 -530 620
rect -490 420 -475 620
rect 2165 420 2180 620
rect 2220 420 2235 620
rect 2275 420 2290 620
rect 2330 420 2345 620
rect 2385 420 2400 620
rect 2440 420 2455 620
rect 2495 420 2510 620
rect 2550 420 2565 620
rect 2605 420 2620 620
rect 2660 420 2675 620
rect 2715 420 2730 620
rect 2770 420 2785 620
<< ndiff >>
rect 715 860 755 875
rect -105 835 -65 850
rect -105 715 -95 835
rect -75 715 -65 835
rect -105 700 -65 715
rect -50 835 -10 850
rect -50 715 -40 835
rect -20 715 -10 835
rect -50 700 -10 715
rect 5 835 45 850
rect 5 715 15 835
rect 35 715 45 835
rect 5 700 45 715
rect 60 835 100 850
rect 60 715 70 835
rect 90 715 100 835
rect 60 700 100 715
rect 115 835 155 850
rect 115 715 125 835
rect 145 715 155 835
rect 115 700 155 715
rect 170 835 210 850
rect 170 715 180 835
rect 200 715 210 835
rect 170 700 210 715
rect 225 835 265 850
rect 225 715 235 835
rect 255 715 265 835
rect 225 700 265 715
rect 280 835 320 850
rect 280 715 290 835
rect 310 715 320 835
rect 280 700 320 715
rect 335 835 375 850
rect 335 715 345 835
rect 365 715 375 835
rect 335 700 375 715
rect 390 835 430 850
rect 390 715 400 835
rect 420 715 430 835
rect 390 700 430 715
rect 445 835 485 850
rect 445 715 455 835
rect 475 715 485 835
rect 445 700 485 715
rect 500 835 540 850
rect 500 715 510 835
rect 530 715 540 835
rect 500 700 540 715
rect 555 835 595 850
rect 555 715 565 835
rect 585 715 595 835
rect 555 700 595 715
rect 715 640 725 860
rect 745 640 755 860
rect 715 625 755 640
rect 770 860 810 875
rect 770 640 780 860
rect 800 640 810 860
rect 770 625 810 640
rect 825 860 865 875
rect 825 640 835 860
rect 855 640 865 860
rect 825 625 865 640
rect 880 860 920 875
rect 880 640 890 860
rect 910 640 920 860
rect 880 625 920 640
rect 935 860 975 875
rect 935 640 945 860
rect 965 640 975 860
rect 1095 835 1135 850
rect 1095 715 1105 835
rect 1125 715 1135 835
rect 1095 700 1135 715
rect 1150 835 1190 850
rect 1150 715 1160 835
rect 1180 715 1190 835
rect 1150 700 1190 715
rect 1205 835 1245 850
rect 1205 715 1215 835
rect 1235 715 1245 835
rect 1205 700 1245 715
rect 1260 835 1300 850
rect 1260 715 1270 835
rect 1290 715 1300 835
rect 1260 700 1300 715
rect 1315 835 1355 850
rect 1315 715 1325 835
rect 1345 715 1355 835
rect 1315 700 1355 715
rect 1370 835 1410 850
rect 1370 715 1380 835
rect 1400 715 1410 835
rect 1370 700 1410 715
rect 1425 835 1465 850
rect 1425 715 1435 835
rect 1455 715 1465 835
rect 1425 700 1465 715
rect 1480 835 1520 850
rect 1480 715 1490 835
rect 1510 715 1520 835
rect 1480 700 1520 715
rect 1535 835 1575 850
rect 1535 715 1545 835
rect 1565 715 1575 835
rect 1535 700 1575 715
rect 1590 835 1630 850
rect 1590 715 1600 835
rect 1620 715 1630 835
rect 1590 700 1630 715
rect 1645 835 1685 850
rect 1645 715 1655 835
rect 1675 715 1685 835
rect 1645 700 1685 715
rect 1700 835 1740 850
rect 1700 715 1710 835
rect 1730 715 1740 835
rect 1700 700 1740 715
rect 1755 835 1795 850
rect 1755 715 1765 835
rect 1785 715 1795 835
rect 1755 700 1795 715
rect 935 625 975 640
rect -105 415 -65 430
rect -105 295 -95 415
rect -75 295 -65 415
rect -105 280 -65 295
rect -50 415 -10 430
rect -50 295 -40 415
rect -20 295 -10 415
rect -50 280 -10 295
rect 5 415 45 430
rect 5 295 15 415
rect 35 295 45 415
rect 5 280 45 295
rect 60 415 100 430
rect 60 295 70 415
rect 90 295 100 415
rect 60 280 100 295
rect 115 415 155 430
rect 115 295 125 415
rect 145 295 155 415
rect 115 280 155 295
rect 170 415 210 430
rect 170 295 180 415
rect 200 295 210 415
rect 170 280 210 295
rect 225 415 265 430
rect 225 295 235 415
rect 255 295 265 415
rect 225 280 265 295
rect 280 415 320 430
rect 280 295 290 415
rect 310 295 320 415
rect 280 280 320 295
rect 335 415 375 430
rect 335 295 345 415
rect 365 295 375 415
rect 335 280 375 295
rect 390 415 430 430
rect 390 295 400 415
rect 420 295 430 415
rect 390 280 430 295
rect 445 415 485 430
rect 445 295 455 415
rect 475 295 485 415
rect 445 280 485 295
rect 500 415 540 430
rect 500 295 510 415
rect 530 295 540 415
rect 500 280 540 295
rect 555 415 595 430
rect 555 295 565 415
rect 585 295 595 415
rect 555 280 595 295
rect 715 415 755 430
rect 715 295 725 415
rect 745 295 755 415
rect 715 280 755 295
rect 770 415 810 430
rect 770 295 780 415
rect 800 295 810 415
rect 770 280 810 295
rect 825 415 865 430
rect 825 295 835 415
rect 855 295 865 415
rect 825 280 865 295
rect 880 415 920 430
rect 880 295 890 415
rect 910 295 920 415
rect 880 280 920 295
rect 935 415 975 430
rect 935 295 945 415
rect 965 295 975 415
rect 935 280 975 295
rect 1095 415 1135 430
rect 1095 295 1105 415
rect 1125 295 1135 415
rect 1095 280 1135 295
rect 1150 415 1190 430
rect 1150 295 1160 415
rect 1180 295 1190 415
rect 1150 280 1190 295
rect 1205 415 1245 430
rect 1205 295 1215 415
rect 1235 295 1245 415
rect 1205 280 1245 295
rect 1260 415 1300 430
rect 1260 295 1270 415
rect 1290 295 1300 415
rect 1260 280 1300 295
rect 1315 415 1355 430
rect 1315 295 1325 415
rect 1345 295 1355 415
rect 1315 280 1355 295
rect 1370 415 1410 430
rect 1370 295 1380 415
rect 1400 295 1410 415
rect 1370 280 1410 295
rect 1425 415 1465 430
rect 1425 295 1435 415
rect 1455 295 1465 415
rect 1425 280 1465 295
rect 1480 415 1520 430
rect 1480 295 1490 415
rect 1510 295 1520 415
rect 1480 280 1520 295
rect 1535 415 1575 430
rect 1535 295 1545 415
rect 1565 295 1575 415
rect 1535 280 1575 295
rect 1590 415 1630 430
rect 1590 295 1600 415
rect 1620 295 1630 415
rect 1590 280 1630 295
rect 1645 415 1685 430
rect 1645 295 1655 415
rect 1675 295 1685 415
rect 1645 280 1685 295
rect 1700 415 1740 430
rect 1700 295 1710 415
rect 1730 295 1740 415
rect 1700 280 1740 295
rect 1755 415 1795 430
rect 1755 295 1765 415
rect 1785 295 1795 415
rect 1755 280 1795 295
rect -1135 215 -1095 230
rect -1135 -55 -1125 215
rect -1105 -55 -1095 215
rect -1135 -70 -1095 -55
rect -1080 215 -1040 230
rect -1080 -55 -1070 215
rect -1050 -55 -1040 215
rect -1080 -70 -1040 -55
rect -1025 215 -985 230
rect -1025 -55 -1015 215
rect -995 -55 -985 215
rect -1025 -70 -985 -55
rect -970 215 -930 230
rect -970 -55 -960 215
rect -940 -55 -930 215
rect -970 -70 -930 -55
rect -915 215 -875 230
rect -915 -55 -905 215
rect -885 -55 -875 215
rect -915 -70 -875 -55
rect -860 215 -820 230
rect -860 -55 -850 215
rect -830 -55 -820 215
rect -860 -70 -820 -55
rect -805 215 -765 230
rect -805 -55 -795 215
rect -775 -55 -765 215
rect -805 -70 -765 -55
rect -750 215 -710 230
rect -750 -55 -740 215
rect -720 -55 -710 215
rect -750 -70 -710 -55
rect -695 215 -655 230
rect -695 -55 -685 215
rect -665 -55 -655 215
rect -695 -70 -655 -55
rect -640 215 -600 230
rect -640 -55 -630 215
rect -610 -55 -600 215
rect -640 -70 -600 -55
rect -585 215 -545 230
rect -585 -55 -575 215
rect -555 -55 -545 215
rect -585 -70 -545 -55
rect -530 215 -490 230
rect -530 -55 -520 215
rect -500 -55 -490 215
rect -530 -70 -490 -55
rect -475 215 -435 230
rect -475 -55 -465 215
rect -445 -55 -435 215
rect 2125 215 2165 230
rect -475 -70 -435 -55
rect 2125 -55 2135 215
rect 2155 -55 2165 215
rect 715 -80 755 -65
rect 715 -300 725 -80
rect 745 -300 755 -80
rect 715 -315 755 -300
rect 770 -80 810 -65
rect 770 -300 780 -80
rect 800 -300 810 -80
rect 770 -315 810 -300
rect 825 -80 865 -65
rect 825 -300 835 -80
rect 855 -300 865 -80
rect 825 -315 865 -300
rect 880 -80 920 -65
rect 880 -300 890 -80
rect 910 -300 920 -80
rect 880 -315 920 -300
rect 935 -80 975 -65
rect 2125 -70 2165 -55
rect 2180 215 2220 230
rect 2180 -55 2190 215
rect 2210 -55 2220 215
rect 2180 -70 2220 -55
rect 2235 215 2275 230
rect 2235 -55 2245 215
rect 2265 -55 2275 215
rect 2235 -70 2275 -55
rect 2290 215 2330 230
rect 2290 -55 2300 215
rect 2320 -55 2330 215
rect 2290 -70 2330 -55
rect 2345 215 2385 230
rect 2345 -55 2355 215
rect 2375 -55 2385 215
rect 2345 -70 2385 -55
rect 2400 215 2440 230
rect 2400 -55 2410 215
rect 2430 -55 2440 215
rect 2400 -70 2440 -55
rect 2455 215 2495 230
rect 2455 -55 2465 215
rect 2485 -55 2495 215
rect 2455 -70 2495 -55
rect 2510 215 2550 230
rect 2510 -55 2520 215
rect 2540 -55 2550 215
rect 2510 -70 2550 -55
rect 2565 215 2605 230
rect 2565 -55 2575 215
rect 2595 -55 2605 215
rect 2565 -70 2605 -55
rect 2620 215 2660 230
rect 2620 -55 2630 215
rect 2650 -55 2660 215
rect 2620 -70 2660 -55
rect 2675 215 2715 230
rect 2675 -55 2685 215
rect 2705 -55 2715 215
rect 2675 -70 2715 -55
rect 2730 215 2770 230
rect 2730 -55 2740 215
rect 2760 -55 2770 215
rect 2730 -70 2770 -55
rect 2785 215 2825 230
rect 2785 -55 2795 215
rect 2815 -55 2825 215
rect 2785 -70 2825 -55
rect 935 -300 945 -80
rect 965 -300 975 -80
rect 935 -315 975 -300
rect -1105 -370 -1065 -355
rect -1105 -1040 -1095 -370
rect -1075 -1040 -1065 -370
rect -1105 -1055 -1065 -1040
rect -1005 -370 -965 -355
rect -1005 -1040 -995 -370
rect -975 -1040 -965 -370
rect -1005 -1055 -965 -1040
rect -905 -370 -865 -355
rect -905 -1040 -895 -370
rect -875 -1040 -865 -370
rect -905 -1055 -865 -1040
rect -805 -370 -765 -355
rect -805 -1040 -795 -370
rect -775 -1040 -765 -370
rect -805 -1055 -765 -1040
rect -705 -370 -665 -355
rect -705 -1040 -695 -370
rect -675 -1040 -665 -370
rect -705 -1055 -665 -1040
rect -605 -370 -565 -355
rect -605 -1040 -595 -370
rect -575 -1040 -565 -370
rect -605 -1055 -565 -1040
rect -505 -370 -465 -355
rect 2155 -370 2195 -355
rect -505 -1040 -495 -370
rect -475 -1040 -465 -370
rect 275 -550 315 -535
rect 275 -770 285 -550
rect 305 -770 315 -550
rect 275 -785 315 -770
rect 330 -550 370 -535
rect 330 -770 340 -550
rect 360 -770 370 -550
rect 330 -785 370 -770
rect 385 -550 425 -535
rect 385 -770 395 -550
rect 415 -770 425 -550
rect 385 -785 425 -770
rect 440 -550 480 -535
rect 440 -770 450 -550
rect 470 -770 480 -550
rect 440 -785 480 -770
rect 495 -550 535 -535
rect 495 -770 505 -550
rect 525 -770 535 -550
rect 495 -785 535 -770
rect 550 -550 590 -535
rect 550 -770 560 -550
rect 580 -770 590 -550
rect 550 -785 590 -770
rect 605 -550 645 -535
rect 605 -770 615 -550
rect 635 -770 645 -550
rect 605 -785 645 -770
rect 660 -550 700 -535
rect 660 -770 670 -550
rect 690 -770 700 -550
rect 660 -785 700 -770
rect 715 -550 755 -535
rect 715 -770 725 -550
rect 745 -770 755 -550
rect 715 -785 755 -770
rect 770 -550 810 -535
rect 770 -770 780 -550
rect 800 -770 810 -550
rect 770 -785 810 -770
rect 825 -550 865 -535
rect 825 -770 835 -550
rect 855 -770 865 -550
rect 825 -785 865 -770
rect 880 -550 920 -535
rect 880 -770 890 -550
rect 910 -770 920 -550
rect 880 -785 920 -770
rect 935 -550 975 -535
rect 935 -770 945 -550
rect 965 -770 975 -550
rect 935 -785 975 -770
rect 990 -550 1030 -535
rect 990 -770 1000 -550
rect 1020 -770 1030 -550
rect 990 -785 1030 -770
rect 1045 -550 1085 -535
rect 1045 -770 1055 -550
rect 1075 -770 1085 -550
rect 1045 -785 1085 -770
rect 1100 -550 1140 -535
rect 1100 -770 1110 -550
rect 1130 -770 1140 -550
rect 1100 -785 1140 -770
rect 1155 -550 1195 -535
rect 1155 -770 1165 -550
rect 1185 -770 1195 -550
rect 1155 -785 1195 -770
rect 1210 -550 1250 -535
rect 1210 -770 1220 -550
rect 1240 -770 1250 -550
rect 1210 -785 1250 -770
rect 1265 -550 1305 -535
rect 1265 -770 1275 -550
rect 1295 -770 1305 -550
rect 1265 -785 1305 -770
rect 1320 -550 1360 -535
rect 1320 -770 1330 -550
rect 1350 -770 1360 -550
rect 1320 -785 1360 -770
rect 1375 -550 1415 -535
rect 1375 -770 1385 -550
rect 1405 -770 1415 -550
rect 1375 -785 1415 -770
rect 1430 -550 1470 -535
rect 1430 -770 1440 -550
rect 1460 -770 1470 -550
rect 1430 -785 1470 -770
rect -505 -1055 -465 -1040
rect 485 -1025 525 -1010
rect 485 -1145 495 -1025
rect 515 -1145 525 -1025
rect 485 -1160 525 -1145
rect 540 -1025 580 -1010
rect 540 -1145 550 -1025
rect 570 -1145 580 -1025
rect 540 -1160 580 -1145
rect 595 -1025 635 -1010
rect 595 -1145 605 -1025
rect 625 -1145 635 -1025
rect 595 -1160 635 -1145
rect 650 -1025 690 -1010
rect 650 -1145 660 -1025
rect 680 -1145 690 -1025
rect 650 -1160 690 -1145
rect 705 -1025 745 -1010
rect 705 -1145 715 -1025
rect 735 -1145 745 -1025
rect 705 -1160 745 -1145
rect 760 -1025 800 -1010
rect 760 -1145 770 -1025
rect 790 -1145 800 -1025
rect 760 -1160 800 -1145
rect 815 -1025 855 -1010
rect 815 -1145 825 -1025
rect 845 -1145 855 -1025
rect 815 -1160 855 -1145
rect 925 -1025 965 -1010
rect 925 -1145 935 -1025
rect 955 -1145 965 -1025
rect 925 -1160 965 -1145
rect 1265 -1025 1305 -1010
rect 1265 -1145 1275 -1025
rect 1295 -1145 1305 -1025
rect 2155 -1040 2165 -370
rect 2185 -1040 2195 -370
rect 2155 -1055 2195 -1040
rect 2255 -370 2295 -355
rect 2255 -1040 2265 -370
rect 2285 -1040 2295 -370
rect 2255 -1055 2295 -1040
rect 2355 -370 2395 -355
rect 2355 -1040 2365 -370
rect 2385 -1040 2395 -370
rect 2355 -1055 2395 -1040
rect 2455 -370 2495 -355
rect 2455 -1040 2465 -370
rect 2485 -1040 2495 -370
rect 2455 -1055 2495 -1040
rect 2555 -370 2595 -355
rect 2555 -1040 2565 -370
rect 2585 -1040 2595 -370
rect 2555 -1055 2595 -1040
rect 2655 -370 2695 -355
rect 2655 -1040 2665 -370
rect 2685 -1040 2695 -370
rect 2655 -1055 2695 -1040
rect 2755 -370 2795 -355
rect 2755 -1040 2765 -370
rect 2785 -1040 2795 -370
rect 2755 -1055 2795 -1040
rect 1265 -1160 1305 -1145
<< pdiff >>
rect 30 2660 70 2675
rect 30 2340 40 2660
rect 60 2340 70 2660
rect 30 2325 70 2340
rect 90 2660 130 2675
rect 90 2340 100 2660
rect 120 2340 130 2660
rect 90 2325 130 2340
rect 150 2660 190 2675
rect 150 2340 160 2660
rect 180 2340 190 2660
rect 150 2325 190 2340
rect 210 2660 250 2675
rect 210 2340 220 2660
rect 240 2340 250 2660
rect 970 2660 1010 2675
rect 210 2325 250 2340
rect 500 2490 540 2505
rect 500 2340 510 2490
rect 530 2340 540 2490
rect 500 2325 540 2340
rect 560 2490 600 2505
rect 560 2340 570 2490
rect 590 2340 600 2490
rect 560 2325 600 2340
rect 620 2490 660 2505
rect 620 2340 630 2490
rect 650 2340 660 2490
rect 620 2325 660 2340
rect 680 2490 720 2505
rect 680 2340 690 2490
rect 710 2340 720 2490
rect 680 2325 720 2340
rect 970 2340 980 2660
rect 1000 2340 1010 2660
rect 970 2325 1010 2340
rect 1030 2660 1070 2675
rect 1030 2340 1040 2660
rect 1060 2340 1070 2660
rect 1030 2325 1070 2340
rect 1090 2660 1130 2675
rect 1090 2340 1100 2660
rect 1120 2340 1130 2660
rect 1090 2325 1130 2340
rect 1150 2660 1190 2675
rect 1150 2340 1160 2660
rect 1180 2340 1190 2660
rect 1150 2325 1190 2340
rect 1440 2660 1480 2675
rect 1440 2340 1450 2660
rect 1470 2340 1480 2660
rect 1440 2325 1480 2340
rect 1500 2660 1540 2675
rect 1500 2340 1510 2660
rect 1530 2340 1540 2660
rect 1500 2325 1540 2340
rect 1560 2660 1600 2675
rect 1560 2340 1570 2660
rect 1590 2340 1600 2660
rect 1560 2325 1600 2340
rect 1620 2660 1660 2675
rect 1620 2340 1630 2660
rect 1650 2340 1660 2660
rect 1620 2325 1660 2340
rect -1165 2085 -1125 2100
rect -1165 1765 -1155 2085
rect -1135 1765 -1125 2085
rect -1165 1750 -1125 1765
rect -1105 2085 -1065 2100
rect -1105 1765 -1095 2085
rect -1075 1765 -1065 2085
rect -1105 1750 -1065 1765
rect -1045 2085 -1005 2100
rect -1045 1765 -1035 2085
rect -1015 1765 -1005 2085
rect -1045 1750 -1005 1765
rect -985 2085 -945 2100
rect -985 1765 -975 2085
rect -955 1765 -945 2085
rect -985 1750 -945 1765
rect -925 2085 -885 2100
rect -925 1765 -915 2085
rect -895 1765 -885 2085
rect -925 1750 -885 1765
rect -865 2085 -825 2100
rect -865 1765 -855 2085
rect -835 1765 -825 2085
rect -865 1750 -825 1765
rect -805 2085 -765 2100
rect -805 1765 -795 2085
rect -775 1765 -765 2085
rect -805 1750 -765 1765
rect -745 2085 -705 2100
rect -745 1765 -735 2085
rect -715 1765 -705 2085
rect -745 1750 -705 1765
rect -685 2085 -645 2100
rect -685 1765 -675 2085
rect -655 1765 -645 2085
rect -685 1750 -645 1765
rect -625 2085 -585 2100
rect -625 1765 -615 2085
rect -595 1765 -585 2085
rect -625 1750 -585 1765
rect -565 2085 -525 2100
rect -565 1765 -555 2085
rect -535 1765 -525 2085
rect -565 1750 -525 1765
rect -505 2085 -465 2100
rect -505 1765 -495 2085
rect -475 1765 -465 2085
rect -505 1750 -465 1765
rect -445 2085 -405 2100
rect -445 1765 -435 2085
rect -415 1765 -405 2085
rect -445 1750 -405 1765
rect -40 2085 0 2100
rect -40 1765 -30 2085
rect -10 1765 0 2085
rect -40 1750 0 1765
rect 20 2085 60 2100
rect 20 1765 30 2085
rect 50 1765 60 2085
rect 20 1750 60 1765
rect 80 2085 120 2100
rect 80 1765 90 2085
rect 110 1765 120 2085
rect 80 1750 120 1765
rect 140 2085 180 2100
rect 140 1765 150 2085
rect 170 1765 180 2085
rect 140 1750 180 1765
rect 200 2085 240 2100
rect 200 1765 210 2085
rect 230 1765 240 2085
rect 200 1750 240 1765
rect 260 2085 300 2100
rect 260 1765 270 2085
rect 290 1765 300 2085
rect 260 1750 300 1765
rect 320 2085 360 2100
rect 320 1765 330 2085
rect 350 1765 360 2085
rect 320 1750 360 1765
rect 380 2085 420 2100
rect 380 1765 390 2085
rect 410 1765 420 2085
rect 380 1750 420 1765
rect 440 2085 480 2100
rect 440 1765 450 2085
rect 470 1765 480 2085
rect 440 1750 480 1765
rect 500 2085 540 2100
rect 500 1765 510 2085
rect 530 1765 540 2085
rect 500 1750 540 1765
rect 560 2085 600 2100
rect 560 1765 570 2085
rect 590 1765 600 2085
rect 560 1750 600 1765
rect 620 2085 660 2100
rect 620 1765 630 2085
rect 650 1765 660 2085
rect 620 1750 660 1765
rect 680 2085 720 2100
rect 680 1765 690 2085
rect 710 1765 720 2085
rect 680 1750 720 1765
rect 970 2085 1010 2100
rect 970 1765 980 2085
rect 1000 1765 1010 2085
rect 970 1750 1010 1765
rect 1030 2085 1070 2100
rect 1030 1765 1040 2085
rect 1060 1765 1070 2085
rect 1030 1750 1070 1765
rect 1090 2085 1130 2100
rect 1090 1765 1100 2085
rect 1120 1765 1130 2085
rect 1090 1750 1130 1765
rect 1150 2085 1190 2100
rect 1150 1765 1160 2085
rect 1180 1765 1190 2085
rect 1150 1750 1190 1765
rect 1210 2085 1250 2100
rect 1210 1765 1220 2085
rect 1240 1765 1250 2085
rect 1210 1750 1250 1765
rect 1270 2085 1310 2100
rect 1270 1765 1280 2085
rect 1300 1765 1310 2085
rect 1270 1750 1310 1765
rect 1330 2085 1370 2100
rect 1330 1765 1340 2085
rect 1360 1765 1370 2085
rect 1330 1750 1370 1765
rect 1390 2085 1430 2100
rect 1390 1765 1400 2085
rect 1420 1765 1430 2085
rect 1390 1750 1430 1765
rect 1450 2085 1490 2100
rect 1450 1765 1460 2085
rect 1480 1765 1490 2085
rect 1450 1750 1490 1765
rect 1510 2085 1550 2100
rect 1510 1765 1520 2085
rect 1540 1765 1550 2085
rect 1510 1750 1550 1765
rect 1570 2085 1610 2100
rect 1570 1765 1580 2085
rect 1600 1765 1610 2085
rect 1570 1750 1610 1765
rect 1630 2085 1670 2100
rect 1630 1765 1640 2085
rect 1660 1765 1670 2085
rect 1630 1750 1670 1765
rect 1690 2085 1730 2100
rect 1690 1765 1700 2085
rect 1720 1765 1730 2085
rect 1690 1750 1730 1765
rect 2095 2085 2135 2100
rect 2095 1765 2105 2085
rect 2125 1765 2135 2085
rect 2095 1750 2135 1765
rect 2155 2085 2195 2100
rect 2155 1765 2165 2085
rect 2185 1765 2195 2085
rect 2155 1750 2195 1765
rect 2215 2085 2255 2100
rect 2215 1765 2225 2085
rect 2245 1765 2255 2085
rect 2215 1750 2255 1765
rect 2275 2085 2315 2100
rect 2275 1765 2285 2085
rect 2305 1765 2315 2085
rect 2275 1750 2315 1765
rect 2335 2085 2375 2100
rect 2335 1765 2345 2085
rect 2365 1765 2375 2085
rect 2335 1750 2375 1765
rect 2395 2085 2435 2100
rect 2395 1765 2405 2085
rect 2425 1765 2435 2085
rect 2395 1750 2435 1765
rect 2455 2085 2495 2100
rect 2455 1765 2465 2085
rect 2485 1765 2495 2085
rect 2455 1750 2495 1765
rect 2515 2085 2555 2100
rect 2515 1765 2525 2085
rect 2545 1765 2555 2085
rect 2515 1750 2555 1765
rect 2575 2085 2615 2100
rect 2575 1765 2585 2085
rect 2605 1765 2615 2085
rect 2575 1750 2615 1765
rect 2635 2085 2675 2100
rect 2635 1765 2645 2085
rect 2665 1765 2675 2085
rect 2635 1750 2675 1765
rect 2695 2085 2735 2100
rect 2695 1765 2705 2085
rect 2725 1765 2735 2085
rect 2695 1750 2735 1765
rect 2755 2085 2795 2100
rect 2755 1765 2765 2085
rect 2785 1765 2795 2085
rect 2755 1750 2795 1765
rect 2815 2085 2855 2100
rect 2815 1765 2825 2085
rect 2845 1765 2855 2085
rect 2815 1750 2855 1765
rect 455 1470 495 1485
rect -1135 1420 -1095 1435
rect -1135 850 -1125 1420
rect -1105 850 -1095 1420
rect -1135 835 -1095 850
rect -1080 1420 -1040 1435
rect -1080 850 -1070 1420
rect -1050 850 -1040 1420
rect -1080 835 -1040 850
rect -1025 1420 -985 1435
rect -1025 850 -1015 1420
rect -995 850 -985 1420
rect -1025 835 -985 850
rect -970 1420 -930 1435
rect -970 850 -960 1420
rect -940 850 -930 1420
rect -970 835 -930 850
rect -915 1420 -875 1435
rect -915 850 -905 1420
rect -885 850 -875 1420
rect -915 835 -875 850
rect -860 1420 -820 1435
rect -860 850 -850 1420
rect -830 850 -820 1420
rect -860 835 -820 850
rect -805 1420 -765 1435
rect -805 850 -795 1420
rect -775 850 -765 1420
rect -805 835 -765 850
rect -750 1420 -710 1435
rect -750 850 -740 1420
rect -720 850 -710 1420
rect -750 835 -710 850
rect -695 1420 -655 1435
rect -695 850 -685 1420
rect -665 850 -655 1420
rect -695 835 -655 850
rect -640 1420 -600 1435
rect -640 850 -630 1420
rect -610 850 -600 1420
rect -640 835 -600 850
rect -585 1420 -545 1435
rect -585 850 -575 1420
rect -555 850 -545 1420
rect -585 835 -545 850
rect -530 1420 -490 1435
rect -530 850 -520 1420
rect -500 850 -490 1420
rect -530 835 -490 850
rect -475 1420 -435 1435
rect -475 850 -465 1420
rect -445 850 -435 1420
rect 455 1250 465 1470
rect 485 1250 495 1470
rect 455 1235 495 1250
rect 510 1470 550 1485
rect 510 1250 520 1470
rect 540 1250 550 1470
rect 510 1235 550 1250
rect 565 1470 605 1485
rect 565 1250 575 1470
rect 595 1250 605 1470
rect 565 1235 605 1250
rect 620 1470 660 1485
rect 620 1250 630 1470
rect 650 1250 660 1470
rect 620 1235 660 1250
rect 675 1470 715 1485
rect 675 1250 685 1470
rect 705 1250 715 1470
rect 675 1235 715 1250
rect 730 1470 770 1485
rect 730 1250 740 1470
rect 760 1250 770 1470
rect 730 1235 770 1250
rect 785 1470 825 1485
rect 865 1470 905 1485
rect 785 1250 795 1470
rect 815 1250 825 1470
rect 865 1250 875 1470
rect 895 1250 905 1470
rect 785 1235 825 1250
rect 865 1235 905 1250
rect 920 1470 960 1485
rect 920 1250 930 1470
rect 950 1250 960 1470
rect 920 1235 960 1250
rect 975 1470 1015 1485
rect 975 1250 985 1470
rect 1005 1250 1015 1470
rect 975 1235 1015 1250
rect 1030 1470 1070 1485
rect 1030 1250 1040 1470
rect 1060 1250 1070 1470
rect 1030 1235 1070 1250
rect 1085 1470 1125 1485
rect 1085 1250 1095 1470
rect 1115 1250 1125 1470
rect 1085 1235 1125 1250
rect 1140 1470 1180 1485
rect 1140 1250 1150 1470
rect 1170 1250 1180 1470
rect 1140 1235 1180 1250
rect 1195 1470 1235 1485
rect 1195 1250 1205 1470
rect 1225 1250 1235 1470
rect 1195 1235 1235 1250
rect 2125 1420 2165 1435
rect -475 835 -435 850
rect 2125 850 2135 1420
rect 2155 850 2165 1420
rect 2125 835 2165 850
rect 2180 1420 2220 1435
rect 2180 850 2190 1420
rect 2210 850 2220 1420
rect 2180 835 2220 850
rect 2235 1420 2275 1435
rect 2235 850 2245 1420
rect 2265 850 2275 1420
rect 2235 835 2275 850
rect 2290 1420 2330 1435
rect 2290 850 2300 1420
rect 2320 850 2330 1420
rect 2290 835 2330 850
rect 2345 1420 2385 1435
rect 2345 850 2355 1420
rect 2375 850 2385 1420
rect 2345 835 2385 850
rect 2400 1420 2440 1435
rect 2400 850 2410 1420
rect 2430 850 2440 1420
rect 2400 835 2440 850
rect 2455 1420 2495 1435
rect 2455 850 2465 1420
rect 2485 850 2495 1420
rect 2455 835 2495 850
rect 2510 1420 2550 1435
rect 2510 850 2520 1420
rect 2540 850 2550 1420
rect 2510 835 2550 850
rect 2565 1420 2605 1435
rect 2565 850 2575 1420
rect 2595 850 2605 1420
rect 2565 835 2605 850
rect 2620 1420 2660 1435
rect 2620 850 2630 1420
rect 2650 850 2660 1420
rect 2620 835 2660 850
rect 2675 1420 2715 1435
rect 2675 850 2685 1420
rect 2705 850 2715 1420
rect 2675 835 2715 850
rect 2730 1420 2770 1435
rect 2730 850 2740 1420
rect 2760 850 2770 1420
rect 2730 835 2770 850
rect 2785 1420 2825 1435
rect 2785 850 2795 1420
rect 2815 850 2825 1420
rect 2785 835 2825 850
rect -1135 605 -1095 620
rect -1135 435 -1125 605
rect -1105 435 -1095 605
rect -1135 420 -1095 435
rect -1080 605 -1040 620
rect -1080 435 -1070 605
rect -1050 435 -1040 605
rect -1080 420 -1040 435
rect -1025 605 -985 620
rect -1025 435 -1015 605
rect -995 435 -985 605
rect -1025 420 -985 435
rect -970 605 -930 620
rect -970 435 -960 605
rect -940 435 -930 605
rect -970 420 -930 435
rect -915 605 -875 620
rect -915 435 -905 605
rect -885 435 -875 605
rect -915 420 -875 435
rect -860 605 -820 620
rect -860 435 -850 605
rect -830 435 -820 605
rect -860 420 -820 435
rect -805 605 -765 620
rect -805 435 -795 605
rect -775 435 -765 605
rect -805 420 -765 435
rect -750 605 -710 620
rect -750 435 -740 605
rect -720 435 -710 605
rect -750 420 -710 435
rect -695 605 -655 620
rect -695 435 -685 605
rect -665 435 -655 605
rect -695 420 -655 435
rect -640 605 -600 620
rect -640 435 -630 605
rect -610 435 -600 605
rect -640 420 -600 435
rect -585 605 -545 620
rect -585 435 -575 605
rect -555 435 -545 605
rect -585 420 -545 435
rect -530 605 -490 620
rect -530 435 -520 605
rect -500 435 -490 605
rect -530 420 -490 435
rect -475 605 -435 620
rect -475 435 -465 605
rect -445 435 -435 605
rect 2125 605 2165 620
rect -475 420 -435 435
rect 2125 435 2135 605
rect 2155 435 2165 605
rect 2125 420 2165 435
rect 2180 605 2220 620
rect 2180 435 2190 605
rect 2210 435 2220 605
rect 2180 420 2220 435
rect 2235 605 2275 620
rect 2235 435 2245 605
rect 2265 435 2275 605
rect 2235 420 2275 435
rect 2290 605 2330 620
rect 2290 435 2300 605
rect 2320 435 2330 605
rect 2290 420 2330 435
rect 2345 605 2385 620
rect 2345 435 2355 605
rect 2375 435 2385 605
rect 2345 420 2385 435
rect 2400 605 2440 620
rect 2400 435 2410 605
rect 2430 435 2440 605
rect 2400 420 2440 435
rect 2455 605 2495 620
rect 2455 435 2465 605
rect 2485 435 2495 605
rect 2455 420 2495 435
rect 2510 605 2550 620
rect 2510 435 2520 605
rect 2540 435 2550 605
rect 2510 420 2550 435
rect 2565 605 2605 620
rect 2565 435 2575 605
rect 2595 435 2605 605
rect 2565 420 2605 435
rect 2620 605 2660 620
rect 2620 435 2630 605
rect 2650 435 2660 605
rect 2620 420 2660 435
rect 2675 605 2715 620
rect 2675 435 2685 605
rect 2705 435 2715 605
rect 2675 420 2715 435
rect 2730 605 2770 620
rect 2730 435 2740 605
rect 2760 435 2770 605
rect 2730 420 2770 435
rect 2785 605 2825 620
rect 2785 435 2795 605
rect 2815 435 2825 605
rect 2785 420 2825 435
<< ndiffc >>
rect -95 715 -75 835
rect -40 715 -20 835
rect 15 715 35 835
rect 70 715 90 835
rect 125 715 145 835
rect 180 715 200 835
rect 235 715 255 835
rect 290 715 310 835
rect 345 715 365 835
rect 400 715 420 835
rect 455 715 475 835
rect 510 715 530 835
rect 565 715 585 835
rect 725 640 745 860
rect 780 640 800 860
rect 835 640 855 860
rect 890 640 910 860
rect 945 640 965 860
rect 1105 715 1125 835
rect 1160 715 1180 835
rect 1215 715 1235 835
rect 1270 715 1290 835
rect 1325 715 1345 835
rect 1380 715 1400 835
rect 1435 715 1455 835
rect 1490 715 1510 835
rect 1545 715 1565 835
rect 1600 715 1620 835
rect 1655 715 1675 835
rect 1710 715 1730 835
rect 1765 715 1785 835
rect -95 295 -75 415
rect -40 295 -20 415
rect 15 295 35 415
rect 70 295 90 415
rect 125 295 145 415
rect 180 295 200 415
rect 235 295 255 415
rect 290 295 310 415
rect 345 295 365 415
rect 400 295 420 415
rect 455 295 475 415
rect 510 295 530 415
rect 565 295 585 415
rect 725 295 745 415
rect 780 295 800 415
rect 835 295 855 415
rect 890 295 910 415
rect 945 295 965 415
rect 1105 295 1125 415
rect 1160 295 1180 415
rect 1215 295 1235 415
rect 1270 295 1290 415
rect 1325 295 1345 415
rect 1380 295 1400 415
rect 1435 295 1455 415
rect 1490 295 1510 415
rect 1545 295 1565 415
rect 1600 295 1620 415
rect 1655 295 1675 415
rect 1710 295 1730 415
rect 1765 295 1785 415
rect -1125 -55 -1105 215
rect -1070 -55 -1050 215
rect -1015 -55 -995 215
rect -960 -55 -940 215
rect -905 -55 -885 215
rect -850 -55 -830 215
rect -795 -55 -775 215
rect -740 -55 -720 215
rect -685 -55 -665 215
rect -630 -55 -610 215
rect -575 -55 -555 215
rect -520 -55 -500 215
rect -465 -55 -445 215
rect 2135 -55 2155 215
rect 725 -300 745 -80
rect 780 -300 800 -80
rect 835 -300 855 -80
rect 890 -300 910 -80
rect 2190 -55 2210 215
rect 2245 -55 2265 215
rect 2300 -55 2320 215
rect 2355 -55 2375 215
rect 2410 -55 2430 215
rect 2465 -55 2485 215
rect 2520 -55 2540 215
rect 2575 -55 2595 215
rect 2630 -55 2650 215
rect 2685 -55 2705 215
rect 2740 -55 2760 215
rect 2795 -55 2815 215
rect 945 -300 965 -80
rect -1095 -1040 -1075 -370
rect -995 -1040 -975 -370
rect -895 -1040 -875 -370
rect -795 -1040 -775 -370
rect -695 -1040 -675 -370
rect -595 -1040 -575 -370
rect -495 -1040 -475 -370
rect 285 -770 305 -550
rect 340 -770 360 -550
rect 395 -770 415 -550
rect 450 -770 470 -550
rect 505 -770 525 -550
rect 560 -770 580 -550
rect 615 -770 635 -550
rect 670 -770 690 -550
rect 725 -770 745 -550
rect 780 -770 800 -550
rect 835 -770 855 -550
rect 890 -770 910 -550
rect 945 -770 965 -550
rect 1000 -770 1020 -550
rect 1055 -770 1075 -550
rect 1110 -770 1130 -550
rect 1165 -770 1185 -550
rect 1220 -770 1240 -550
rect 1275 -770 1295 -550
rect 1330 -770 1350 -550
rect 1385 -770 1405 -550
rect 1440 -770 1460 -550
rect 495 -1145 515 -1025
rect 550 -1145 570 -1025
rect 605 -1145 625 -1025
rect 660 -1145 680 -1025
rect 715 -1145 735 -1025
rect 770 -1145 790 -1025
rect 825 -1145 845 -1025
rect 935 -1145 955 -1025
rect 1275 -1145 1295 -1025
rect 2165 -1040 2185 -370
rect 2265 -1040 2285 -370
rect 2365 -1040 2385 -370
rect 2465 -1040 2485 -370
rect 2565 -1040 2585 -370
rect 2665 -1040 2685 -370
rect 2765 -1040 2785 -370
<< pdiffc >>
rect 40 2340 60 2660
rect 100 2340 120 2660
rect 160 2340 180 2660
rect 220 2340 240 2660
rect 510 2340 530 2490
rect 570 2340 590 2490
rect 630 2340 650 2490
rect 690 2340 710 2490
rect 980 2340 1000 2660
rect 1040 2340 1060 2660
rect 1100 2340 1120 2660
rect 1160 2340 1180 2660
rect 1450 2340 1470 2660
rect 1510 2340 1530 2660
rect 1570 2340 1590 2660
rect 1630 2340 1650 2660
rect -1155 1765 -1135 2085
rect -1095 1765 -1075 2085
rect -1035 1765 -1015 2085
rect -975 1765 -955 2085
rect -915 1765 -895 2085
rect -855 1765 -835 2085
rect -795 1765 -775 2085
rect -735 1765 -715 2085
rect -675 1765 -655 2085
rect -615 1765 -595 2085
rect -555 1765 -535 2085
rect -495 1765 -475 2085
rect -435 1765 -415 2085
rect -30 1765 -10 2085
rect 30 1765 50 2085
rect 90 1765 110 2085
rect 150 1765 170 2085
rect 210 1765 230 2085
rect 270 1765 290 2085
rect 330 1765 350 2085
rect 390 1765 410 2085
rect 450 1765 470 2085
rect 510 1765 530 2085
rect 570 1765 590 2085
rect 630 1765 650 2085
rect 690 1765 710 2085
rect 980 1765 1000 2085
rect 1040 1765 1060 2085
rect 1100 1765 1120 2085
rect 1160 1765 1180 2085
rect 1220 1765 1240 2085
rect 1280 1765 1300 2085
rect 1340 1765 1360 2085
rect 1400 1765 1420 2085
rect 1460 1765 1480 2085
rect 1520 1765 1540 2085
rect 1580 1765 1600 2085
rect 1640 1765 1660 2085
rect 1700 1765 1720 2085
rect 2105 1765 2125 2085
rect 2165 1765 2185 2085
rect 2225 1765 2245 2085
rect 2285 1765 2305 2085
rect 2345 1765 2365 2085
rect 2405 1765 2425 2085
rect 2465 1765 2485 2085
rect 2525 1765 2545 2085
rect 2585 1765 2605 2085
rect 2645 1765 2665 2085
rect 2705 1765 2725 2085
rect 2765 1765 2785 2085
rect 2825 1765 2845 2085
rect -1125 850 -1105 1420
rect -1070 850 -1050 1420
rect -1015 850 -995 1420
rect -960 850 -940 1420
rect -905 850 -885 1420
rect -850 850 -830 1420
rect -795 850 -775 1420
rect -740 850 -720 1420
rect -685 850 -665 1420
rect -630 850 -610 1420
rect -575 850 -555 1420
rect -520 850 -500 1420
rect -465 850 -445 1420
rect 465 1250 485 1470
rect 520 1250 540 1470
rect 575 1250 595 1470
rect 630 1250 650 1470
rect 685 1250 705 1470
rect 740 1250 760 1470
rect 795 1250 815 1470
rect 875 1250 895 1470
rect 930 1250 950 1470
rect 985 1250 1005 1470
rect 1040 1250 1060 1470
rect 1095 1250 1115 1470
rect 1150 1250 1170 1470
rect 1205 1250 1225 1470
rect 2135 850 2155 1420
rect 2190 850 2210 1420
rect 2245 850 2265 1420
rect 2300 850 2320 1420
rect 2355 850 2375 1420
rect 2410 850 2430 1420
rect 2465 850 2485 1420
rect 2520 850 2540 1420
rect 2575 850 2595 1420
rect 2630 850 2650 1420
rect 2685 850 2705 1420
rect 2740 850 2760 1420
rect 2795 850 2815 1420
rect -1125 435 -1105 605
rect -1070 435 -1050 605
rect -1015 435 -995 605
rect -960 435 -940 605
rect -905 435 -885 605
rect -850 435 -830 605
rect -795 435 -775 605
rect -740 435 -720 605
rect -685 435 -665 605
rect -630 435 -610 605
rect -575 435 -555 605
rect -520 435 -500 605
rect -465 435 -445 605
rect 2135 435 2155 605
rect 2190 435 2210 605
rect 2245 435 2265 605
rect 2300 435 2320 605
rect 2355 435 2375 605
rect 2410 435 2430 605
rect 2465 435 2485 605
rect 2520 435 2540 605
rect 2575 435 2595 605
rect 2630 435 2650 605
rect 2685 435 2705 605
rect 2740 435 2760 605
rect 2795 435 2815 605
<< psubdiff >>
rect 675 860 715 875
rect -145 835 -105 850
rect -145 715 -135 835
rect -115 715 -105 835
rect -145 700 -105 715
rect 595 835 635 850
rect 595 715 605 835
rect 625 715 635 835
rect 595 700 635 715
rect 675 640 685 860
rect 705 640 715 860
rect 675 625 715 640
rect 975 860 1015 875
rect 975 640 985 860
rect 1005 640 1015 860
rect 1055 835 1095 850
rect 1055 715 1065 835
rect 1085 715 1095 835
rect 1055 700 1095 715
rect 1795 835 1835 850
rect 1795 715 1805 835
rect 1825 715 1835 835
rect 1795 700 1835 715
rect 975 625 1015 640
rect -145 415 -105 430
rect -145 295 -135 415
rect -115 295 -105 415
rect -145 280 -105 295
rect 595 415 635 430
rect 595 295 605 415
rect 625 295 635 415
rect 595 280 635 295
rect 675 415 715 430
rect 675 295 685 415
rect 705 295 715 415
rect 675 280 715 295
rect 975 415 1015 430
rect 975 295 985 415
rect 1005 295 1015 415
rect 975 280 1015 295
rect 1055 415 1095 430
rect 1055 295 1065 415
rect 1085 295 1095 415
rect 1055 280 1095 295
rect 1795 415 1835 430
rect 1795 295 1805 415
rect 1825 295 1835 415
rect 1795 280 1835 295
rect -1175 215 -1135 230
rect -1175 -55 -1165 215
rect -1145 -55 -1135 215
rect -1175 -70 -1135 -55
rect -435 215 -395 230
rect -435 -55 -425 215
rect -405 -55 -395 215
rect 2085 215 2125 230
rect -435 -70 -395 -55
rect 2085 -55 2095 215
rect 2115 -55 2125 215
rect 675 -80 715 -65
rect 675 -300 685 -80
rect 705 -300 715 -80
rect 675 -315 715 -300
rect 975 -80 1015 -65
rect 2085 -70 2125 -55
rect 2825 215 2865 230
rect 2825 -55 2835 215
rect 2855 -55 2865 215
rect 2825 -70 2865 -55
rect 975 -300 985 -80
rect 1005 -300 1015 -80
rect 975 -315 1015 -300
rect -1145 -370 -1105 -355
rect -1145 -1040 -1135 -370
rect -1115 -1040 -1105 -370
rect -1145 -1055 -1105 -1040
rect -465 -370 -425 -355
rect 2115 -370 2155 -355
rect -465 -1040 -455 -370
rect -435 -1040 -425 -370
rect 235 -550 275 -535
rect 235 -770 245 -550
rect 265 -770 275 -550
rect 235 -785 275 -770
rect 1470 -550 1510 -535
rect 1470 -770 1480 -550
rect 1500 -770 1510 -550
rect 1470 -785 1510 -770
rect -465 -1055 -425 -1040
rect 445 -1025 485 -1010
rect 445 -1145 455 -1025
rect 475 -1145 485 -1025
rect 445 -1160 485 -1145
rect 855 -1025 895 -1010
rect 855 -1145 865 -1025
rect 885 -1145 895 -1025
rect 855 -1160 895 -1145
rect 2115 -1040 2125 -370
rect 2145 -1040 2155 -370
rect 2115 -1055 2155 -1040
rect 2795 -370 2835 -355
rect 2795 -1040 2805 -370
rect 2825 -1040 2835 -370
rect 2795 -1055 2835 -1040
<< nsubdiff >>
rect -10 2660 30 2675
rect -10 2340 0 2660
rect 20 2340 30 2660
rect -10 2325 30 2340
rect 250 2660 290 2675
rect 250 2340 260 2660
rect 280 2340 290 2660
rect 930 2660 970 2675
rect 250 2325 290 2340
rect 460 2490 500 2505
rect 460 2340 470 2490
rect 490 2340 500 2490
rect 460 2325 500 2340
rect 720 2490 760 2505
rect 720 2340 730 2490
rect 750 2340 760 2490
rect 720 2325 760 2340
rect 930 2340 940 2660
rect 960 2340 970 2660
rect 930 2325 970 2340
rect 1190 2660 1230 2675
rect 1190 2340 1200 2660
rect 1220 2340 1230 2660
rect 1190 2325 1230 2340
rect 1400 2660 1440 2675
rect 1400 2340 1410 2660
rect 1430 2340 1440 2660
rect 1400 2325 1440 2340
rect 1660 2660 1700 2675
rect 1660 2340 1670 2660
rect 1690 2340 1700 2660
rect 1660 2325 1700 2340
rect -1205 2085 -1165 2100
rect -1205 1765 -1195 2085
rect -1175 1765 -1165 2085
rect -1205 1750 -1165 1765
rect -405 2085 -365 2100
rect -405 1765 -395 2085
rect -375 1765 -365 2085
rect -405 1750 -365 1765
rect -80 2085 -40 2100
rect -80 1765 -70 2085
rect -50 1765 -40 2085
rect -80 1750 -40 1765
rect 720 2085 760 2100
rect 720 1765 730 2085
rect 750 1765 760 2085
rect 720 1750 760 1765
rect 930 2085 970 2100
rect 930 1765 940 2085
rect 960 1765 970 2085
rect 930 1750 970 1765
rect 1730 2085 1770 2100
rect 1730 1765 1740 2085
rect 1760 1765 1770 2085
rect 1730 1750 1770 1765
rect 2055 2085 2095 2100
rect 2055 1765 2065 2085
rect 2085 1765 2095 2085
rect 2055 1750 2095 1765
rect 2855 2085 2895 2100
rect 2855 1765 2865 2085
rect 2885 1765 2895 2085
rect 2855 1750 2895 1765
rect 415 1470 455 1485
rect -1175 1420 -1135 1435
rect -1175 850 -1165 1420
rect -1145 850 -1135 1420
rect -1175 835 -1135 850
rect -435 1420 -395 1435
rect -435 850 -425 1420
rect -405 850 -395 1420
rect 415 1250 425 1470
rect 445 1250 455 1470
rect 415 1235 455 1250
rect 825 1470 865 1485
rect 825 1250 835 1470
rect 855 1250 865 1470
rect 825 1235 865 1250
rect 1235 1470 1275 1485
rect 1235 1250 1245 1470
rect 1265 1250 1275 1470
rect 1235 1235 1275 1250
rect 2085 1420 2125 1435
rect -435 835 -395 850
rect 2085 850 2095 1420
rect 2115 850 2125 1420
rect 2085 835 2125 850
rect 2825 1420 2865 1435
rect 2825 850 2835 1420
rect 2855 850 2865 1420
rect 2825 835 2865 850
rect -1175 605 -1135 620
rect -1175 435 -1165 605
rect -1145 435 -1135 605
rect -1175 420 -1135 435
rect -435 605 -395 620
rect -435 435 -425 605
rect -405 435 -395 605
rect 2085 605 2125 620
rect -435 420 -395 435
rect 2085 435 2095 605
rect 2115 435 2125 605
rect 2085 420 2125 435
rect 2825 605 2865 620
rect 2825 435 2835 605
rect 2855 435 2865 605
rect 2825 420 2865 435
<< psubdiffcont >>
rect -135 715 -115 835
rect 605 715 625 835
rect 685 640 705 860
rect 985 640 1005 860
rect 1065 715 1085 835
rect 1805 715 1825 835
rect -135 295 -115 415
rect 605 295 625 415
rect 685 295 705 415
rect 985 295 1005 415
rect 1065 295 1085 415
rect 1805 295 1825 415
rect -1165 -55 -1145 215
rect -425 -55 -405 215
rect 2095 -55 2115 215
rect 685 -300 705 -80
rect 2835 -55 2855 215
rect 985 -300 1005 -80
rect -1135 -1040 -1115 -370
rect -455 -1040 -435 -370
rect 245 -770 265 -550
rect 1480 -770 1500 -550
rect 455 -1145 475 -1025
rect 865 -1145 885 -1025
rect 2125 -1040 2145 -370
rect 2805 -1040 2825 -370
<< nsubdiffcont >>
rect 0 2340 20 2660
rect 260 2340 280 2660
rect 470 2340 490 2490
rect 730 2340 750 2490
rect 940 2340 960 2660
rect 1200 2340 1220 2660
rect 1410 2340 1430 2660
rect 1670 2340 1690 2660
rect -1195 1765 -1175 2085
rect -395 1765 -375 2085
rect -70 1765 -50 2085
rect 730 1765 750 2085
rect 940 1765 960 2085
rect 1740 1765 1760 2085
rect 2065 1765 2085 2085
rect 2865 1765 2885 2085
rect -1165 850 -1145 1420
rect -425 850 -405 1420
rect 425 1250 445 1470
rect 835 1250 855 1470
rect 1245 1250 1265 1470
rect 2095 850 2115 1420
rect 2835 850 2855 1420
rect -1165 435 -1145 605
rect -425 435 -405 605
rect 2095 435 2115 605
rect 2835 435 2855 605
<< poly >>
rect 30 2720 70 2730
rect 30 2700 40 2720
rect 60 2705 70 2720
rect 210 2720 250 2730
rect 210 2705 220 2720
rect 60 2700 90 2705
rect 30 2690 90 2700
rect 190 2700 220 2705
rect 240 2700 250 2720
rect 190 2690 250 2700
rect 970 2720 1010 2730
rect 970 2700 980 2720
rect 1000 2705 1010 2720
rect 1150 2720 1190 2730
rect 1150 2705 1160 2720
rect 1000 2700 1030 2705
rect 970 2690 1030 2700
rect 1130 2700 1160 2705
rect 1180 2700 1190 2720
rect 1130 2690 1190 2700
rect 1440 2720 1480 2730
rect 1440 2700 1450 2720
rect 1470 2705 1480 2720
rect 1620 2720 1660 2730
rect 1620 2705 1630 2720
rect 1470 2700 1500 2705
rect 1440 2690 1500 2700
rect 1600 2700 1630 2705
rect 1650 2700 1660 2720
rect 1600 2690 1660 2700
rect 70 2675 90 2690
rect 130 2675 150 2690
rect 190 2675 210 2690
rect 1010 2675 1030 2690
rect 1070 2675 1090 2690
rect 1130 2675 1150 2690
rect 1480 2675 1500 2690
rect 1540 2675 1560 2690
rect 1600 2675 1620 2690
rect 500 2550 540 2560
rect 500 2530 510 2550
rect 530 2535 540 2550
rect 680 2550 720 2560
rect 680 2535 690 2550
rect 530 2530 560 2535
rect 500 2520 560 2530
rect 660 2530 690 2535
rect 710 2530 720 2550
rect 660 2520 720 2530
rect 540 2505 560 2520
rect 600 2505 620 2520
rect 660 2505 680 2520
rect 70 2310 90 2325
rect 130 2310 150 2325
rect 190 2310 210 2325
rect 540 2310 560 2325
rect 600 2310 620 2325
rect 660 2310 680 2325
rect 1010 2310 1030 2325
rect 1070 2310 1090 2325
rect 1130 2310 1150 2325
rect 1480 2310 1500 2325
rect 1540 2310 1560 2325
rect 1600 2310 1620 2325
rect 130 2300 169 2310
rect 130 2295 144 2300
rect 139 2280 144 2295
rect 164 2280 169 2300
rect 600 2300 639 2310
rect 600 2295 614 2300
rect 139 2270 169 2280
rect 609 2280 614 2295
rect 634 2280 639 2300
rect 609 2270 639 2280
rect 1051 2300 1090 2310
rect 1051 2280 1056 2300
rect 1076 2295 1090 2300
rect 1521 2300 1560 2310
rect 1076 2280 1081 2295
rect 1051 2270 1081 2280
rect 1521 2280 1526 2300
rect 1546 2295 1560 2300
rect 1546 2280 1551 2295
rect 1521 2270 1551 2280
rect -1165 2145 -1125 2155
rect -1165 2125 -1155 2145
rect -1135 2130 -1125 2145
rect -445 2145 -405 2155
rect -445 2130 -435 2145
rect -1135 2125 -1105 2130
rect -1165 2115 -1105 2125
rect -465 2125 -435 2130
rect -415 2125 -405 2145
rect -465 2115 -405 2125
rect -40 2145 0 2155
rect -40 2125 -30 2145
rect -10 2130 0 2145
rect 680 2145 720 2155
rect 680 2130 690 2145
rect -10 2125 20 2130
rect -40 2115 20 2125
rect 660 2125 690 2130
rect 710 2125 720 2145
rect 660 2115 720 2125
rect 970 2145 1010 2155
rect 970 2125 980 2145
rect 1000 2130 1010 2145
rect 1690 2145 1730 2155
rect 1690 2130 1700 2145
rect 1000 2125 1030 2130
rect 970 2115 1030 2125
rect 1670 2125 1700 2130
rect 1720 2125 1730 2145
rect 1670 2115 1730 2125
rect 2095 2145 2135 2155
rect 2095 2125 2105 2145
rect 2125 2130 2135 2145
rect 2815 2145 2855 2155
rect 2815 2130 2825 2145
rect 2125 2125 2155 2130
rect 2095 2115 2155 2125
rect 2795 2125 2825 2130
rect 2845 2125 2855 2145
rect 2795 2115 2855 2125
rect -1125 2100 -1105 2115
rect -1065 2100 -1045 2115
rect -1005 2100 -985 2115
rect -945 2100 -925 2115
rect -885 2100 -865 2115
rect -825 2100 -805 2115
rect -765 2100 -745 2115
rect -705 2100 -685 2115
rect -645 2100 -625 2115
rect -585 2100 -565 2115
rect -525 2100 -505 2115
rect -465 2100 -445 2115
rect 0 2100 20 2115
rect 60 2100 80 2115
rect 120 2100 140 2115
rect 180 2100 200 2115
rect 240 2100 260 2115
rect 300 2100 320 2115
rect 360 2100 380 2115
rect 420 2100 440 2115
rect 480 2100 500 2115
rect 540 2100 560 2115
rect 600 2100 620 2115
rect 660 2100 680 2115
rect 1010 2100 1030 2115
rect 1070 2100 1090 2115
rect 1130 2100 1150 2115
rect 1190 2100 1210 2115
rect 1250 2100 1270 2115
rect 1310 2100 1330 2115
rect 1370 2100 1390 2115
rect 1430 2100 1450 2115
rect 1490 2100 1510 2115
rect 1550 2100 1570 2115
rect 1610 2100 1630 2115
rect 1670 2100 1690 2115
rect 2135 2100 2155 2115
rect 2195 2100 2215 2115
rect 2255 2100 2275 2115
rect 2315 2100 2335 2115
rect 2375 2100 2395 2115
rect 2435 2100 2455 2115
rect 2495 2100 2515 2115
rect 2555 2100 2575 2115
rect 2615 2100 2635 2115
rect 2675 2100 2695 2115
rect 2735 2100 2755 2115
rect 2795 2100 2815 2115
rect -1125 1735 -1105 1750
rect -1065 1740 -1045 1750
rect -1005 1740 -985 1750
rect -945 1740 -925 1750
rect -885 1740 -865 1750
rect -825 1740 -805 1750
rect -765 1740 -745 1750
rect -705 1740 -685 1750
rect -645 1740 -625 1750
rect -585 1740 -565 1750
rect -525 1740 -505 1750
rect -1065 1725 -505 1740
rect -465 1735 -445 1750
rect 0 1735 20 1750
rect 60 1740 80 1750
rect 120 1740 140 1750
rect 180 1740 200 1750
rect 240 1740 260 1750
rect 300 1740 320 1750
rect 360 1740 380 1750
rect 420 1740 440 1750
rect 480 1740 500 1750
rect 540 1740 560 1750
rect 600 1740 620 1750
rect 60 1725 620 1740
rect 660 1735 680 1750
rect 1010 1735 1030 1750
rect 1070 1740 1090 1750
rect 1130 1740 1150 1750
rect 1190 1740 1210 1750
rect 1250 1740 1270 1750
rect 1310 1740 1330 1750
rect 1370 1740 1390 1750
rect 1430 1740 1450 1750
rect 1490 1740 1510 1750
rect 1550 1740 1570 1750
rect 1610 1740 1630 1750
rect 1070 1725 1630 1740
rect 1670 1735 1690 1750
rect 2135 1735 2155 1750
rect 2195 1740 2215 1750
rect 2255 1740 2275 1750
rect 2315 1740 2335 1750
rect 2375 1740 2395 1750
rect 2435 1740 2455 1750
rect 2495 1740 2515 1750
rect 2555 1740 2575 1750
rect 2615 1740 2635 1750
rect 2675 1740 2695 1750
rect 2735 1740 2755 1750
rect 2195 1725 2755 1740
rect 2795 1735 2815 1750
rect -705 1630 -685 1725
rect 420 1675 440 1725
rect 1250 1675 1270 1725
rect 410 1665 450 1675
rect 410 1645 420 1665
rect 440 1645 450 1665
rect 410 1635 450 1645
rect 1240 1665 1280 1675
rect 1240 1645 1250 1665
rect 1270 1645 1280 1665
rect 1240 1635 1280 1645
rect 2375 1630 2395 1725
rect -715 1620 -675 1630
rect -715 1600 -705 1620
rect -685 1600 -675 1620
rect -715 1590 -675 1600
rect 2365 1620 2405 1630
rect 2365 1600 2375 1620
rect 2395 1600 2405 1620
rect 2365 1590 2405 1600
rect 455 1560 495 1570
rect 455 1540 465 1560
rect 485 1545 495 1560
rect 785 1560 825 1570
rect 785 1545 795 1560
rect 485 1540 510 1545
rect 455 1530 510 1540
rect -1135 1480 -1095 1490
rect -1135 1460 -1125 1480
rect -1105 1465 -1095 1480
rect -475 1480 -435 1490
rect 495 1485 510 1530
rect 770 1540 795 1545
rect 815 1540 825 1560
rect 770 1530 825 1540
rect 865 1560 905 1570
rect 865 1540 875 1560
rect 895 1545 905 1560
rect 1195 1560 1235 1570
rect 1195 1545 1205 1560
rect 895 1540 920 1545
rect 865 1530 920 1540
rect 550 1485 565 1500
rect 605 1485 620 1500
rect 660 1485 675 1500
rect 715 1485 730 1500
rect 770 1485 785 1530
rect 905 1485 920 1530
rect 1180 1540 1205 1545
rect 1225 1540 1235 1560
rect 1180 1530 1235 1540
rect 960 1485 975 1500
rect 1015 1485 1030 1500
rect 1070 1485 1085 1500
rect 1125 1485 1140 1500
rect 1180 1485 1195 1530
rect -475 1465 -465 1480
rect -1105 1460 -1080 1465
rect -1135 1450 -1080 1460
rect -490 1460 -465 1465
rect -445 1460 -435 1480
rect -490 1450 -435 1460
rect -1095 1435 -1080 1450
rect -1040 1435 -1025 1450
rect -985 1435 -970 1450
rect -930 1435 -915 1450
rect -875 1435 -860 1450
rect -820 1435 -805 1450
rect -765 1435 -750 1450
rect -710 1435 -695 1450
rect -655 1435 -640 1450
rect -600 1435 -585 1450
rect -545 1435 -530 1450
rect -490 1435 -475 1450
rect 2125 1480 2165 1490
rect 2125 1460 2135 1480
rect 2155 1465 2165 1480
rect 2785 1480 2825 1490
rect 2785 1465 2795 1480
rect 2155 1460 2180 1465
rect 2125 1450 2180 1460
rect 2770 1460 2795 1465
rect 2815 1460 2825 1480
rect 2770 1450 2825 1460
rect 2165 1435 2180 1450
rect 2220 1435 2235 1450
rect 2275 1435 2290 1450
rect 2330 1435 2345 1450
rect 2385 1435 2400 1450
rect 2440 1435 2455 1450
rect 2495 1435 2510 1450
rect 2550 1435 2565 1450
rect 2605 1435 2620 1450
rect 2660 1435 2675 1450
rect 2715 1435 2730 1450
rect 2770 1435 2785 1450
rect 495 1220 510 1235
rect 550 1220 565 1235
rect 605 1225 620 1235
rect 660 1225 675 1235
rect 550 1210 580 1220
rect 605 1210 675 1225
rect 715 1220 730 1235
rect 770 1220 785 1235
rect 905 1220 920 1235
rect 960 1220 975 1235
rect 1015 1225 1030 1235
rect 1070 1225 1085 1235
rect 700 1210 730 1220
rect 550 1190 555 1210
rect 575 1190 580 1210
rect 550 1180 580 1190
rect 620 1190 630 1210
rect 650 1190 660 1210
rect 620 1180 660 1190
rect 700 1190 705 1210
rect 725 1190 730 1210
rect 700 1180 730 1190
rect 960 1210 990 1220
rect 1015 1210 1085 1225
rect 1125 1220 1140 1235
rect 1180 1220 1195 1235
rect 1110 1210 1140 1220
rect 960 1190 965 1210
rect 985 1190 990 1210
rect 960 1180 990 1190
rect 1030 1190 1040 1210
rect 1060 1190 1070 1210
rect 1030 1180 1070 1190
rect 1110 1190 1115 1210
rect 1135 1190 1140 1210
rect 1110 1180 1140 1190
rect 120 945 150 955
rect 120 925 125 945
rect 145 925 150 945
rect 1540 945 1570 955
rect 120 915 150 925
rect 795 920 835 930
rect 130 875 145 915
rect 795 900 805 920
rect 825 900 835 920
rect 1540 925 1545 945
rect 1565 925 1570 945
rect 1540 915 1570 925
rect 795 890 880 900
rect 755 875 770 890
rect 810 885 880 890
rect 810 875 825 885
rect 865 875 880 885
rect 920 875 935 890
rect 1545 875 1560 915
rect -65 850 -50 865
rect -10 860 500 875
rect -10 850 5 860
rect 45 850 60 860
rect 100 850 115 860
rect 155 850 170 860
rect 210 850 225 860
rect 265 850 280 860
rect 320 850 335 860
rect 375 850 390 860
rect 430 850 445 860
rect 485 850 500 860
rect 540 850 555 865
rect -1095 820 -1080 835
rect -1040 825 -1025 835
rect -985 825 -970 835
rect -930 825 -915 835
rect -875 825 -860 835
rect -820 825 -805 835
rect -765 825 -750 835
rect -710 825 -695 835
rect -655 825 -640 835
rect -600 825 -585 835
rect -545 825 -530 835
rect -1040 810 -530 825
rect -490 820 -475 835
rect -795 720 -775 810
rect -805 710 -765 720
rect -805 690 -795 710
rect -775 690 -765 710
rect -805 680 -765 690
rect -65 685 -50 700
rect -10 685 5 700
rect 45 685 60 700
rect 100 685 115 700
rect 155 685 170 700
rect 210 685 225 700
rect 265 685 280 700
rect 320 685 335 700
rect 375 685 390 700
rect 430 685 445 700
rect 485 685 500 700
rect 540 685 555 700
rect -100 675 -50 685
rect -1135 665 -1095 675
rect -1135 645 -1125 665
rect -1105 650 -1095 665
rect -475 665 -435 675
rect -475 650 -465 665
rect -1105 645 -1080 650
rect -1135 635 -1080 645
rect -490 645 -465 650
rect -445 645 -435 665
rect -100 655 -95 675
rect -75 670 -50 675
rect 540 675 590 685
rect 540 670 565 675
rect -75 655 -70 670
rect -100 645 -70 655
rect 560 655 565 670
rect 585 655 590 675
rect 560 645 590 655
rect -490 635 -435 645
rect -1095 620 -1080 635
rect -1040 620 -1025 635
rect -985 620 -970 635
rect -930 620 -915 635
rect -875 620 -860 635
rect -820 620 -805 635
rect -765 620 -750 635
rect -710 620 -695 635
rect -655 620 -640 635
rect -600 620 -585 635
rect -545 620 -530 635
rect -490 620 -475 635
rect 1135 850 1150 865
rect 1190 860 1700 875
rect 1190 850 1205 860
rect 1245 850 1260 860
rect 1300 850 1315 860
rect 1355 850 1370 860
rect 1410 850 1425 860
rect 1465 850 1480 860
rect 1520 850 1535 860
rect 1575 850 1590 860
rect 1630 850 1645 860
rect 1685 850 1700 860
rect 1740 850 1755 865
rect 2165 820 2180 835
rect 2220 825 2235 835
rect 2275 825 2290 835
rect 2330 825 2345 835
rect 2385 825 2400 835
rect 2440 825 2455 835
rect 2495 825 2510 835
rect 2550 825 2565 835
rect 2605 825 2620 835
rect 2660 825 2675 835
rect 2715 825 2730 835
rect 2220 810 2730 825
rect 2770 820 2785 835
rect 2465 720 2485 810
rect 2455 710 2495 720
rect 1135 685 1150 700
rect 1190 685 1205 700
rect 1245 685 1260 700
rect 1300 685 1315 700
rect 1355 685 1370 700
rect 1410 685 1425 700
rect 1465 685 1480 700
rect 1520 685 1535 700
rect 1575 685 1590 700
rect 1630 685 1645 700
rect 1685 685 1700 700
rect 1740 685 1755 700
rect 2455 690 2465 710
rect 2485 690 2495 710
rect 1100 675 1150 685
rect 1100 655 1105 675
rect 1125 670 1150 675
rect 1740 675 1790 685
rect 2455 680 2495 690
rect 1740 670 1765 675
rect 1125 655 1130 670
rect 1100 645 1130 655
rect 1760 655 1765 670
rect 1785 655 1790 675
rect 1760 645 1790 655
rect 2125 665 2165 675
rect 2125 645 2135 665
rect 2155 650 2165 665
rect 2785 665 2825 675
rect 2785 650 2795 665
rect 2155 645 2180 650
rect 2125 635 2180 645
rect 2770 645 2795 650
rect 2815 645 2825 665
rect 2770 635 2825 645
rect 755 610 770 625
rect 810 610 825 625
rect 865 610 880 625
rect 920 610 935 625
rect 2165 620 2180 635
rect 2220 620 2235 635
rect 2275 620 2290 635
rect 2330 620 2345 635
rect 2385 620 2400 635
rect 2440 620 2455 635
rect 2495 620 2510 635
rect 2550 620 2565 635
rect 2605 620 2620 635
rect 2660 620 2675 635
rect 2715 620 2730 635
rect 2770 620 2785 635
rect 715 600 770 610
rect 715 580 725 600
rect 745 595 770 600
rect 920 600 975 610
rect 920 595 945 600
rect 745 580 755 595
rect 715 570 755 580
rect 935 580 945 595
rect 965 580 975 600
rect 935 570 975 580
rect 145 545 175 555
rect 145 525 150 545
rect 170 525 175 545
rect 145 515 175 525
rect 795 545 825 555
rect 795 525 800 545
rect 820 525 825 545
rect 795 515 825 525
rect 155 455 170 515
rect 715 475 755 485
rect 715 455 725 475
rect 745 460 755 475
rect 745 455 770 460
rect -65 430 -50 445
rect -10 440 500 455
rect 715 445 770 455
rect -10 430 5 440
rect 45 430 60 440
rect 100 430 115 440
rect 155 430 170 440
rect 210 430 225 440
rect 265 430 280 440
rect 320 430 335 440
rect 375 430 390 440
rect 430 430 445 440
rect 485 430 500 440
rect 540 430 555 445
rect 755 430 770 445
rect 810 430 825 515
rect 865 545 895 555
rect 865 525 870 545
rect 890 525 895 545
rect 865 515 895 525
rect 1515 545 1545 555
rect 1515 525 1520 545
rect 1540 525 1545 545
rect 1515 515 1545 525
rect 865 430 880 515
rect 935 475 975 485
rect 935 460 945 475
rect 920 455 945 460
rect 965 455 975 475
rect 1520 455 1535 515
rect 920 445 975 455
rect 920 430 935 445
rect 1135 430 1150 445
rect 1190 440 1700 455
rect 1190 430 1205 440
rect 1245 430 1260 440
rect 1300 430 1315 440
rect 1355 430 1370 440
rect 1410 430 1425 440
rect 1465 430 1480 440
rect 1520 430 1535 440
rect 1575 430 1590 440
rect 1630 430 1645 440
rect 1685 430 1700 440
rect 1740 430 1755 445
rect -1095 405 -1080 420
rect -1040 410 -1025 420
rect -985 410 -970 420
rect -930 410 -915 420
rect -875 410 -860 420
rect -820 410 -805 420
rect -765 410 -750 420
rect -710 410 -695 420
rect -655 410 -640 420
rect -600 410 -585 420
rect -545 410 -530 420
rect -1040 395 -530 410
rect -490 405 -475 420
rect -740 345 -720 395
rect -750 335 -710 345
rect -750 315 -740 335
rect -720 315 -710 335
rect -750 305 -710 315
rect -740 255 -720 305
rect 2165 405 2180 420
rect 2220 410 2235 420
rect 2275 410 2290 420
rect 2330 410 2345 420
rect 2385 410 2400 420
rect 2440 410 2455 420
rect 2495 410 2510 420
rect 2550 410 2565 420
rect 2605 410 2620 420
rect 2660 410 2675 420
rect 2715 410 2730 420
rect 2220 395 2730 410
rect 2770 405 2785 420
rect 2410 345 2430 395
rect 2400 335 2440 345
rect 2400 315 2410 335
rect 2430 315 2440 335
rect 2400 305 2440 315
rect -65 265 -50 280
rect -10 265 5 280
rect 45 265 60 280
rect 100 265 115 280
rect 155 265 170 280
rect 210 265 225 280
rect 265 265 280 280
rect 320 265 335 280
rect 375 265 390 280
rect 430 265 445 280
rect 485 265 500 280
rect 540 265 555 280
rect 755 265 770 280
rect 810 265 825 280
rect 865 265 880 280
rect 920 265 935 280
rect 1135 265 1150 280
rect 1190 265 1205 280
rect 1245 265 1260 280
rect 1300 265 1315 280
rect 1355 265 1370 280
rect 1410 265 1425 280
rect 1465 265 1480 280
rect 1520 265 1535 280
rect 1575 265 1590 280
rect 1630 265 1645 280
rect 1685 265 1700 280
rect 1740 265 1755 280
rect -100 255 -50 265
rect -1095 230 -1080 245
rect -1040 240 -530 255
rect -1040 230 -1025 240
rect -985 230 -970 240
rect -930 230 -915 240
rect -875 230 -860 240
rect -820 230 -805 240
rect -765 230 -750 240
rect -710 230 -695 240
rect -655 230 -640 240
rect -600 230 -585 240
rect -545 230 -530 240
rect -490 230 -475 245
rect -100 235 -95 255
rect -75 250 -50 255
rect 540 255 590 265
rect 540 250 565 255
rect -75 235 -70 250
rect -100 225 -70 235
rect 560 235 565 250
rect 585 235 590 255
rect 560 225 590 235
rect 1100 255 1150 265
rect 1100 235 1105 255
rect 1125 250 1150 255
rect 1740 255 1790 265
rect 2410 255 2430 305
rect 1740 250 1765 255
rect 1125 235 1130 250
rect 1100 225 1130 235
rect 1760 235 1765 250
rect 1785 235 1790 255
rect 1760 225 1790 235
rect 2165 230 2180 245
rect 2220 240 2730 255
rect 2220 230 2235 240
rect 2275 230 2290 240
rect 2330 230 2345 240
rect 2385 230 2400 240
rect 2440 230 2455 240
rect 2495 230 2510 240
rect 2550 230 2565 240
rect 2605 230 2620 240
rect 2660 230 2675 240
rect 2715 230 2730 240
rect 2770 230 2785 245
rect 830 -15 860 -5
rect 830 -35 835 -15
rect 855 -35 860 -15
rect 830 -40 860 -35
rect 755 -65 770 -50
rect 810 -55 880 -40
rect 810 -65 825 -55
rect 865 -65 880 -55
rect 920 -65 935 -50
rect -1095 -85 -1080 -70
rect -1040 -85 -1025 -70
rect -985 -85 -970 -70
rect -930 -85 -915 -70
rect -875 -85 -860 -70
rect -820 -85 -805 -70
rect -765 -85 -750 -70
rect -710 -85 -695 -70
rect -655 -85 -640 -70
rect -600 -85 -585 -70
rect -545 -85 -530 -70
rect -490 -85 -475 -70
rect -1135 -95 -1080 -85
rect -1135 -115 -1125 -95
rect -1105 -100 -1080 -95
rect -490 -95 -435 -85
rect -490 -100 -465 -95
rect -1105 -115 -1095 -100
rect -1135 -125 -1095 -115
rect -475 -115 -465 -100
rect -445 -115 -435 -95
rect -475 -125 -435 -115
rect -805 -250 -765 -240
rect -805 -270 -795 -250
rect -775 -270 -765 -250
rect -805 -280 -765 -270
rect -795 -330 -775 -280
rect 2165 -85 2180 -70
rect 2220 -85 2235 -70
rect 2275 -85 2290 -70
rect 2330 -85 2345 -70
rect 2385 -85 2400 -70
rect 2440 -85 2455 -70
rect 2495 -85 2510 -70
rect 2550 -85 2565 -70
rect 2605 -85 2620 -70
rect 2660 -85 2675 -70
rect 2715 -85 2730 -70
rect 2770 -85 2785 -70
rect 2125 -95 2180 -85
rect 2125 -115 2135 -95
rect 2155 -100 2180 -95
rect 2770 -95 2825 -85
rect 2770 -100 2795 -95
rect 2155 -115 2165 -100
rect 2125 -125 2165 -115
rect 2785 -115 2795 -100
rect 2815 -115 2825 -95
rect 2785 -125 2825 -115
rect 2455 -250 2495 -240
rect 2455 -270 2465 -250
rect 2485 -270 2495 -250
rect 2455 -280 2495 -270
rect 755 -330 770 -315
rect 810 -330 825 -315
rect 865 -330 880 -315
rect 920 -330 935 -315
rect 2465 -330 2485 -280
rect -1065 -355 -1005 -340
rect -965 -345 -605 -330
rect 715 -340 770 -330
rect -965 -355 -905 -345
rect -865 -355 -805 -345
rect -765 -355 -705 -345
rect -665 -355 -605 -345
rect -565 -355 -505 -340
rect 715 -360 725 -340
rect 745 -345 770 -340
rect 920 -340 975 -330
rect 920 -345 945 -340
rect 745 -360 755 -345
rect 715 -370 755 -360
rect 935 -360 945 -345
rect 965 -360 975 -340
rect 2195 -355 2255 -340
rect 2295 -345 2655 -330
rect 2295 -355 2355 -345
rect 2395 -355 2455 -345
rect 2495 -355 2555 -345
rect 2595 -355 2655 -345
rect 2695 -355 2755 -340
rect 935 -370 975 -360
rect 445 -440 475 -430
rect 445 -460 450 -440
rect 470 -460 475 -440
rect 445 -470 475 -460
rect 1350 -440 1390 -430
rect 1350 -460 1360 -440
rect 1380 -460 1390 -440
rect 1350 -470 1390 -460
rect 450 -510 470 -470
rect 315 -535 330 -520
rect 370 -525 1320 -510
rect 370 -535 385 -525
rect 425 -535 440 -525
rect 480 -535 495 -525
rect 535 -535 550 -525
rect 590 -535 605 -525
rect 645 -535 660 -525
rect 700 -535 715 -525
rect 755 -535 770 -525
rect 810 -535 825 -525
rect 865 -535 880 -525
rect 920 -535 935 -525
rect 975 -535 990 -525
rect 1030 -535 1045 -525
rect 1085 -535 1100 -525
rect 1140 -535 1155 -525
rect 1195 -535 1210 -525
rect 1250 -535 1265 -525
rect 1305 -535 1320 -525
rect 1360 -535 1375 -470
rect 1415 -535 1430 -520
rect 315 -800 330 -785
rect 370 -800 385 -785
rect 425 -800 440 -785
rect 480 -800 495 -785
rect 535 -800 550 -785
rect 590 -800 605 -785
rect 645 -800 660 -785
rect 700 -800 715 -785
rect 755 -800 770 -785
rect 810 -800 825 -785
rect 865 -800 880 -785
rect 920 -800 935 -785
rect 975 -800 990 -785
rect 1030 -800 1045 -785
rect 1085 -800 1100 -785
rect 1140 -800 1155 -785
rect 1195 -800 1210 -785
rect 1250 -800 1265 -785
rect 1305 -800 1320 -785
rect 1360 -800 1375 -785
rect 1415 -800 1430 -785
rect 275 -810 330 -800
rect 275 -830 285 -810
rect 305 -815 330 -810
rect 1415 -810 1470 -800
rect 1415 -815 1440 -810
rect 305 -830 315 -815
rect 275 -840 315 -830
rect 1430 -830 1440 -815
rect 1460 -830 1470 -810
rect 1430 -840 1470 -830
rect 650 -965 690 -955
rect 650 -985 660 -965
rect 680 -985 690 -965
rect 1095 -965 1135 -955
rect 1095 -985 1105 -965
rect 1125 -985 1135 -965
rect 525 -1010 540 -995
rect 580 -1000 760 -985
rect 1095 -995 1135 -985
rect 580 -1010 595 -1000
rect 635 -1010 650 -1000
rect 690 -1010 705 -1000
rect 745 -1010 760 -1000
rect 800 -1010 815 -995
rect 965 -1010 1265 -995
rect -1065 -1070 -1005 -1055
rect -965 -1070 -905 -1055
rect -865 -1070 -805 -1055
rect -765 -1070 -705 -1055
rect -665 -1070 -605 -1055
rect -565 -1070 -505 -1055
rect -1105 -1080 -1005 -1070
rect -1105 -1100 -1095 -1080
rect -1075 -1085 -1005 -1080
rect -565 -1080 -465 -1070
rect -565 -1085 -495 -1080
rect -1075 -1100 -1065 -1085
rect -1105 -1110 -1065 -1100
rect -505 -1100 -495 -1085
rect -475 -1100 -465 -1080
rect -505 -1110 -465 -1100
rect 2195 -1070 2255 -1055
rect 2295 -1070 2355 -1055
rect 2395 -1070 2455 -1055
rect 2495 -1070 2555 -1055
rect 2595 -1070 2655 -1055
rect 2695 -1070 2755 -1055
rect 2155 -1080 2255 -1070
rect 2155 -1100 2165 -1080
rect 2185 -1085 2255 -1080
rect 2695 -1080 2795 -1070
rect 2695 -1085 2765 -1080
rect 2185 -1100 2195 -1085
rect 2155 -1110 2195 -1100
rect 2755 -1100 2765 -1085
rect 2785 -1100 2795 -1080
rect 2755 -1110 2795 -1100
rect 525 -1175 540 -1160
rect 580 -1175 595 -1160
rect 635 -1175 650 -1160
rect 690 -1175 705 -1160
rect 745 -1175 760 -1160
rect 800 -1175 815 -1160
rect 965 -1175 1265 -1160
rect 490 -1185 540 -1175
rect 490 -1205 495 -1185
rect 515 -1190 540 -1185
rect 800 -1185 850 -1175
rect 800 -1190 825 -1185
rect 515 -1205 520 -1190
rect 490 -1215 520 -1205
rect 820 -1205 825 -1190
rect 845 -1205 850 -1185
rect 820 -1215 850 -1205
<< polycont >>
rect 40 2700 60 2720
rect 220 2700 240 2720
rect 980 2700 1000 2720
rect 1160 2700 1180 2720
rect 1450 2700 1470 2720
rect 1630 2700 1650 2720
rect 510 2530 530 2550
rect 690 2530 710 2550
rect 144 2280 164 2300
rect 614 2280 634 2300
rect 1056 2280 1076 2300
rect 1526 2280 1546 2300
rect -1155 2125 -1135 2145
rect -435 2125 -415 2145
rect -30 2125 -10 2145
rect 690 2125 710 2145
rect 980 2125 1000 2145
rect 1700 2125 1720 2145
rect 2105 2125 2125 2145
rect 2825 2125 2845 2145
rect 420 1645 440 1665
rect 1250 1645 1270 1665
rect -705 1600 -685 1620
rect 2375 1600 2395 1620
rect 465 1540 485 1560
rect -1125 1460 -1105 1480
rect 795 1540 815 1560
rect 875 1540 895 1560
rect 1205 1540 1225 1560
rect -465 1460 -445 1480
rect 2135 1460 2155 1480
rect 2795 1460 2815 1480
rect 555 1190 575 1210
rect 630 1190 650 1210
rect 705 1190 725 1210
rect 965 1190 985 1210
rect 1040 1190 1060 1210
rect 1115 1190 1135 1210
rect 125 925 145 945
rect 805 900 825 920
rect 1545 925 1565 945
rect -795 690 -775 710
rect -1125 645 -1105 665
rect -465 645 -445 665
rect -95 655 -75 675
rect 565 655 585 675
rect 2465 690 2485 710
rect 1105 655 1125 675
rect 1765 655 1785 675
rect 2135 645 2155 665
rect 2795 645 2815 665
rect 725 580 745 600
rect 945 580 965 600
rect 150 525 170 545
rect 800 525 820 545
rect 725 455 745 475
rect 870 525 890 545
rect 1520 525 1540 545
rect 945 455 965 475
rect -740 315 -720 335
rect 2410 315 2430 335
rect -95 235 -75 255
rect 565 235 585 255
rect 1105 235 1125 255
rect 1765 235 1785 255
rect 835 -35 855 -15
rect -1125 -115 -1105 -95
rect -465 -115 -445 -95
rect -795 -270 -775 -250
rect 2135 -115 2155 -95
rect 2795 -115 2815 -95
rect 2465 -270 2485 -250
rect 725 -360 745 -340
rect 945 -360 965 -340
rect 450 -460 470 -440
rect 1360 -460 1380 -440
rect 285 -830 305 -810
rect 1440 -830 1460 -810
rect 660 -985 680 -965
rect 1105 -985 1125 -965
rect -1095 -1100 -1075 -1080
rect -495 -1100 -475 -1080
rect 2165 -1100 2185 -1080
rect 2765 -1100 2785 -1080
rect 495 -1205 515 -1185
rect 825 -1205 845 -1185
<< xpolycontact >>
rect -1501 1170 -1360 1390
rect -1501 825 -1360 1045
rect 3050 1170 3191 1390
rect 3050 825 3191 1045
rect -1490 297 -1455 517
rect -1490 -85 -1455 138
rect -1430 297 -1395 517
rect -1430 -85 -1395 138
rect -1370 297 -1335 517
rect -1370 -85 -1335 138
rect -1310 297 -1275 517
rect -1310 -85 -1275 138
rect 2965 297 3000 517
rect 2965 -85 3000 138
rect 3025 297 3060 517
rect 3025 -85 3060 138
rect 3085 297 3120 517
rect 3085 -85 3120 138
rect 3145 297 3180 517
rect 3145 -85 3180 138
rect -1290 -638 -1255 -415
rect -1290 -1105 -1255 -885
rect -1230 -638 -1195 -415
rect -1230 -1105 -1195 -885
rect 2885 -638 2920 -415
rect 2885 -1105 2920 -885
rect 2945 -638 2980 -415
rect 2945 -1105 2980 -885
<< ppolyres >>
rect -1501 1045 -1360 1170
rect 3050 1045 3191 1170
<< xpolyres >>
rect -1490 138 -1455 297
rect -1430 138 -1395 297
rect -1370 138 -1335 297
rect -1310 138 -1275 297
rect 2965 138 3000 297
rect 3025 138 3060 297
rect 3085 138 3120 297
rect 3145 138 3180 297
rect -1290 -885 -1255 -638
rect -1230 -885 -1195 -638
rect 2885 -885 2920 -638
rect 2945 -885 2980 -638
<< locali >>
rect 30 2720 70 2730
rect 30 2700 40 2720
rect 60 2700 70 2720
rect 30 2690 70 2700
rect 210 2720 250 2730
rect 210 2700 220 2720
rect 240 2700 250 2720
rect 210 2690 250 2700
rect 970 2720 1010 2730
rect 970 2700 980 2720
rect 1000 2700 1010 2720
rect 970 2690 1010 2700
rect 1150 2720 1190 2730
rect 1150 2700 1160 2720
rect 1180 2700 1190 2720
rect 1150 2690 1190 2700
rect 1440 2720 1480 2730
rect 1440 2700 1450 2720
rect 1470 2700 1480 2720
rect 1440 2690 1480 2700
rect 1620 2720 1660 2730
rect 1620 2700 1630 2720
rect 1650 2700 1660 2720
rect 1620 2690 1660 2700
rect -5 2660 65 2670
rect -5 2340 0 2660
rect 20 2340 40 2660
rect 60 2340 65 2660
rect -5 2330 65 2340
rect 95 2660 125 2670
rect 95 2340 100 2660
rect 120 2340 125 2660
rect 95 2330 125 2340
rect 155 2660 185 2670
rect 155 2340 160 2660
rect 180 2340 185 2660
rect 155 2330 185 2340
rect 215 2660 285 2670
rect 215 2340 220 2660
rect 240 2340 260 2660
rect 280 2340 285 2660
rect 935 2660 1005 2670
rect 500 2550 540 2560
rect 500 2530 510 2550
rect 530 2530 540 2550
rect 500 2520 540 2530
rect 560 2550 600 2560
rect 560 2530 570 2550
rect 590 2530 600 2550
rect 560 2520 600 2530
rect 680 2550 720 2560
rect 680 2530 690 2550
rect 710 2530 720 2550
rect 680 2520 720 2530
rect 215 2330 285 2340
rect 465 2490 535 2500
rect 465 2340 470 2490
rect 490 2340 510 2490
rect 530 2340 535 2490
rect 465 2330 535 2340
rect 565 2490 595 2500
rect 565 2340 570 2490
rect 590 2340 595 2490
rect 565 2330 595 2340
rect 625 2490 655 2500
rect 625 2340 630 2490
rect 650 2340 655 2490
rect 625 2330 655 2340
rect 685 2490 755 2500
rect 685 2340 690 2490
rect 710 2340 730 2490
rect 750 2340 755 2490
rect 685 2330 755 2340
rect 935 2340 940 2660
rect 960 2340 980 2660
rect 1000 2340 1005 2660
rect 935 2330 1005 2340
rect 1035 2660 1065 2670
rect 1035 2340 1040 2660
rect 1060 2340 1065 2660
rect 1035 2330 1065 2340
rect 1095 2660 1125 2670
rect 1095 2340 1100 2660
rect 1120 2340 1125 2660
rect 1095 2330 1125 2340
rect 1155 2660 1225 2670
rect 1155 2340 1160 2660
rect 1180 2340 1200 2660
rect 1220 2340 1225 2660
rect 1155 2330 1225 2340
rect 1405 2660 1475 2670
rect 1405 2340 1410 2660
rect 1430 2340 1450 2660
rect 1470 2340 1475 2660
rect 1405 2330 1475 2340
rect 1505 2660 1535 2670
rect 1505 2340 1510 2660
rect 1530 2340 1535 2660
rect 1505 2330 1535 2340
rect 1565 2660 1595 2670
rect 1565 2340 1570 2660
rect 1590 2340 1595 2660
rect 1565 2330 1595 2340
rect 1625 2660 1695 2670
rect 1625 2340 1630 2660
rect 1650 2340 1670 2660
rect 1690 2340 1695 2660
rect 1625 2330 1695 2340
rect 95 2310 115 2330
rect 75 2300 115 2310
rect 75 2280 85 2300
rect 105 2280 115 2300
rect 75 2270 115 2280
rect 139 2300 169 2310
rect 139 2280 144 2300
rect 164 2280 169 2300
rect 139 2270 169 2280
rect 609 2300 639 2310
rect 609 2280 614 2300
rect 634 2280 639 2300
rect 609 2270 639 2280
rect 1051 2300 1081 2310
rect 1051 2280 1056 2300
rect 1076 2280 1081 2300
rect 1051 2270 1081 2280
rect 1521 2300 1551 2310
rect 1521 2280 1526 2300
rect 1546 2280 1551 2300
rect 1521 2270 1551 2280
rect -1165 2145 -1125 2155
rect -1165 2125 -1155 2145
rect -1135 2125 -1125 2145
rect -1165 2115 -1125 2125
rect -445 2145 -405 2155
rect -445 2125 -435 2145
rect -415 2125 -405 2145
rect -445 2115 -405 2125
rect -40 2145 0 2155
rect -40 2125 -30 2145
rect -10 2125 0 2145
rect -40 2115 0 2125
rect 680 2145 720 2155
rect 680 2125 690 2145
rect 710 2125 720 2145
rect 680 2115 720 2125
rect 970 2145 1010 2155
rect 970 2125 980 2145
rect 1000 2125 1010 2145
rect 970 2115 1010 2125
rect 1690 2145 1730 2155
rect 1690 2125 1700 2145
rect 1720 2125 1730 2145
rect 1690 2115 1730 2125
rect 2095 2145 2135 2155
rect 2095 2125 2105 2145
rect 2125 2125 2135 2145
rect 2095 2115 2135 2125
rect 2815 2145 2855 2155
rect 2815 2125 2825 2145
rect 2845 2125 2855 2145
rect 2815 2115 2855 2125
rect -1160 2095 -1130 2115
rect -35 2095 -5 2115
rect 685 2095 715 2115
rect 975 2095 1005 2115
rect 1695 2095 1725 2115
rect 2820 2095 2850 2115
rect -1200 2085 -1130 2095
rect -1200 1765 -1195 2085
rect -1175 1765 -1155 2085
rect -1135 1765 -1130 2085
rect -1200 1755 -1130 1765
rect -1100 2085 -1070 2095
rect -1100 1765 -1095 2085
rect -1075 1765 -1070 2085
rect -1100 1755 -1070 1765
rect -1040 2085 -1010 2095
rect -1040 1765 -1035 2085
rect -1015 1765 -1010 2085
rect -1040 1755 -1010 1765
rect -980 2085 -950 2095
rect -980 1765 -975 2085
rect -955 1765 -950 2085
rect -980 1755 -950 1765
rect -920 2085 -890 2095
rect -920 1765 -915 2085
rect -895 1765 -890 2085
rect -920 1755 -890 1765
rect -860 2085 -830 2095
rect -860 1765 -855 2085
rect -835 1765 -830 2085
rect -860 1755 -830 1765
rect -800 2085 -770 2095
rect -800 1765 -795 2085
rect -775 1765 -770 2085
rect -800 1755 -770 1765
rect -740 2085 -710 2095
rect -740 1765 -735 2085
rect -715 1765 -710 2085
rect -740 1755 -710 1765
rect -680 2085 -650 2095
rect -680 1765 -675 2085
rect -655 1765 -650 2085
rect -680 1755 -650 1765
rect -620 2085 -590 2095
rect -620 1765 -615 2085
rect -595 1765 -590 2085
rect -620 1755 -590 1765
rect -560 2085 -530 2095
rect -560 1765 -555 2085
rect -535 1765 -530 2085
rect -560 1755 -530 1765
rect -500 2085 -470 2095
rect -500 1765 -495 2085
rect -475 1765 -470 2085
rect -500 1755 -470 1765
rect -440 2085 -370 2095
rect -440 1765 -435 2085
rect -415 1765 -395 2085
rect -375 1765 -370 2085
rect -440 1755 -370 1765
rect -75 2085 -5 2095
rect -75 1765 -70 2085
rect -50 1765 -30 2085
rect -10 1765 -5 2085
rect -75 1755 -5 1765
rect 25 2085 55 2095
rect 25 1765 30 2085
rect 50 1765 55 2085
rect 25 1755 55 1765
rect 85 2085 115 2095
rect 85 1765 90 2085
rect 110 1765 115 2085
rect 85 1755 115 1765
rect 145 2085 175 2095
rect 145 1765 150 2085
rect 170 1765 175 2085
rect 145 1755 175 1765
rect 205 2085 235 2095
rect 205 1765 210 2085
rect 230 1765 235 2085
rect 205 1755 235 1765
rect 265 2085 295 2095
rect 265 1765 270 2085
rect 290 1765 295 2085
rect 265 1755 295 1765
rect 325 2085 355 2095
rect 325 1765 330 2085
rect 350 1765 355 2085
rect 325 1755 355 1765
rect 385 2085 415 2095
rect 385 1765 390 2085
rect 410 1765 415 2085
rect 385 1755 415 1765
rect 445 2085 475 2095
rect 445 1765 450 2085
rect 470 1765 475 2085
rect 445 1755 475 1765
rect 505 2085 535 2095
rect 505 1765 510 2085
rect 530 1765 535 2085
rect 505 1755 535 1765
rect 565 2085 595 2095
rect 565 1765 570 2085
rect 590 1765 595 2085
rect 565 1755 595 1765
rect 625 2085 655 2095
rect 625 1765 630 2085
rect 650 1765 655 2085
rect 625 1755 655 1765
rect 685 2085 755 2095
rect 685 1765 690 2085
rect 710 1765 730 2085
rect 750 1765 755 2085
rect 685 1755 755 1765
rect 935 2085 1005 2095
rect 935 1765 940 2085
rect 960 1765 980 2085
rect 1000 1765 1005 2085
rect 935 1755 1005 1765
rect 1035 2085 1065 2095
rect 1035 1765 1040 2085
rect 1060 1765 1065 2085
rect 1035 1755 1065 1765
rect 1095 2085 1125 2095
rect 1095 1765 1100 2085
rect 1120 1765 1125 2085
rect 1095 1755 1125 1765
rect 1155 2085 1185 2095
rect 1155 1765 1160 2085
rect 1180 1765 1185 2085
rect 1155 1755 1185 1765
rect 1215 2085 1245 2095
rect 1215 1765 1220 2085
rect 1240 1765 1245 2085
rect 1215 1755 1245 1765
rect 1275 2085 1305 2095
rect 1275 1765 1280 2085
rect 1300 1765 1305 2085
rect 1275 1755 1305 1765
rect 1335 2085 1365 2095
rect 1335 1765 1340 2085
rect 1360 1765 1365 2085
rect 1335 1755 1365 1765
rect 1395 2085 1425 2095
rect 1395 1765 1400 2085
rect 1420 1765 1425 2085
rect 1395 1755 1425 1765
rect 1455 2085 1485 2095
rect 1455 1765 1460 2085
rect 1480 1765 1485 2085
rect 1455 1755 1485 1765
rect 1515 2085 1545 2095
rect 1515 1765 1520 2085
rect 1540 1765 1545 2085
rect 1515 1755 1545 1765
rect 1575 2085 1605 2095
rect 1575 1765 1580 2085
rect 1600 1765 1605 2085
rect 1575 1755 1605 1765
rect 1635 2085 1665 2095
rect 1635 1765 1640 2085
rect 1660 1765 1665 2085
rect 1635 1755 1665 1765
rect 1695 2085 1765 2095
rect 1695 1765 1700 2085
rect 1720 1765 1740 2085
rect 1760 1765 1765 2085
rect 1695 1755 1765 1765
rect 2060 2085 2130 2095
rect 2060 1765 2065 2085
rect 2085 1765 2105 2085
rect 2125 1765 2130 2085
rect 2060 1755 2130 1765
rect 2160 2085 2190 2095
rect 2160 1765 2165 2085
rect 2185 1765 2190 2085
rect 2160 1755 2190 1765
rect 2220 2085 2250 2095
rect 2220 1765 2225 2085
rect 2245 1765 2250 2085
rect 2220 1755 2250 1765
rect 2280 2085 2310 2095
rect 2280 1765 2285 2085
rect 2305 1765 2310 2085
rect 2280 1755 2310 1765
rect 2340 2085 2370 2095
rect 2340 1765 2345 2085
rect 2365 1765 2370 2085
rect 2340 1755 2370 1765
rect 2400 2085 2430 2095
rect 2400 1765 2405 2085
rect 2425 1765 2430 2085
rect 2400 1755 2430 1765
rect 2460 2085 2490 2095
rect 2460 1765 2465 2085
rect 2485 1765 2490 2085
rect 2460 1755 2490 1765
rect 2520 2085 2550 2095
rect 2520 1765 2525 2085
rect 2545 1765 2550 2085
rect 2520 1755 2550 1765
rect 2580 2085 2610 2095
rect 2580 1765 2585 2085
rect 2605 1765 2610 2085
rect 2580 1755 2610 1765
rect 2640 2085 2670 2095
rect 2640 1765 2645 2085
rect 2665 1765 2670 2085
rect 2640 1755 2670 1765
rect 2700 2085 2730 2095
rect 2700 1765 2705 2085
rect 2725 1765 2730 2085
rect 2700 1755 2730 1765
rect 2760 2085 2790 2095
rect 2760 1765 2765 2085
rect 2785 1765 2790 2085
rect 2760 1755 2790 1765
rect 2820 2085 2890 2095
rect 2820 1765 2825 2085
rect 2845 1765 2865 2085
rect 2885 1765 2890 2085
rect 2820 1755 2890 1765
rect 410 1665 450 1675
rect 410 1645 420 1665
rect 440 1645 450 1665
rect 410 1635 450 1645
rect 1240 1665 1280 1675
rect 1240 1645 1250 1665
rect 1270 1645 1280 1665
rect 1240 1635 1280 1645
rect -715 1620 -675 1630
rect -715 1600 -705 1620
rect -685 1600 -675 1620
rect -715 1590 -675 1600
rect 2365 1620 2405 1630
rect 2365 1600 2375 1620
rect 2395 1600 2405 1620
rect 2365 1590 2405 1600
rect 455 1560 495 1570
rect 455 1540 465 1560
rect 485 1540 495 1560
rect 455 1530 495 1540
rect 785 1560 825 1570
rect 785 1540 795 1560
rect 815 1540 825 1560
rect 785 1530 825 1540
rect 865 1560 905 1570
rect 865 1540 875 1560
rect 895 1540 905 1560
rect 865 1530 905 1540
rect 1195 1560 1235 1570
rect 1195 1540 1205 1560
rect 1225 1540 1235 1560
rect 1195 1530 1235 1540
rect -1135 1480 -1095 1490
rect -1135 1460 -1125 1480
rect -1105 1460 -1095 1480
rect -1135 1450 -1095 1460
rect -475 1480 -435 1490
rect 2125 1480 2165 1490
rect -475 1460 -465 1480
rect -445 1460 -435 1480
rect -475 1450 -435 1460
rect 420 1470 490 1480
rect -1501 1420 -1360 1430
rect -1501 1400 -1495 1420
rect -1475 1400 -1440 1420
rect -1420 1400 -1385 1420
rect -1365 1400 -1360 1420
rect -1501 1390 -1360 1400
rect -1170 1420 -1100 1430
rect -1170 850 -1165 1420
rect -1145 850 -1125 1420
rect -1105 850 -1100 1420
rect -1170 840 -1100 850
rect -1075 1420 -1045 1430
rect -1075 850 -1070 1420
rect -1050 850 -1045 1420
rect -1075 840 -1045 850
rect -1020 1420 -990 1430
rect -1020 850 -1015 1420
rect -995 850 -990 1420
rect -1020 840 -990 850
rect -965 1420 -935 1430
rect -965 850 -960 1420
rect -940 850 -935 1420
rect -965 840 -935 850
rect -910 1420 -880 1430
rect -910 850 -905 1420
rect -885 850 -880 1420
rect -910 840 -880 850
rect -855 1420 -825 1430
rect -855 850 -850 1420
rect -830 850 -825 1420
rect -855 840 -825 850
rect -800 1420 -770 1430
rect -800 850 -795 1420
rect -775 850 -770 1420
rect -800 840 -770 850
rect -745 1420 -715 1430
rect -745 850 -740 1420
rect -720 850 -715 1420
rect -745 840 -715 850
rect -690 1420 -660 1430
rect -690 850 -685 1420
rect -665 850 -660 1420
rect -690 840 -660 850
rect -635 1420 -605 1430
rect -635 850 -630 1420
rect -610 850 -605 1420
rect -635 840 -605 850
rect -580 1420 -550 1430
rect -580 850 -575 1420
rect -555 850 -550 1420
rect -580 840 -550 850
rect -525 1420 -495 1430
rect -525 850 -520 1420
rect -500 850 -495 1420
rect -525 840 -495 850
rect -470 1420 -400 1430
rect -470 850 -465 1420
rect -445 850 -425 1420
rect -405 850 -400 1420
rect 420 1250 425 1470
rect 445 1250 465 1470
rect 485 1250 490 1470
rect 420 1240 490 1250
rect 515 1470 545 1480
rect 515 1250 520 1470
rect 540 1250 545 1470
rect 515 1240 545 1250
rect 570 1470 600 1480
rect 570 1250 575 1470
rect 595 1250 600 1470
rect 570 1240 600 1250
rect 625 1470 655 1480
rect 625 1250 630 1470
rect 650 1250 655 1470
rect 625 1240 655 1250
rect 680 1470 710 1480
rect 680 1250 685 1470
rect 705 1250 710 1470
rect 680 1240 710 1250
rect 735 1470 765 1480
rect 735 1250 740 1470
rect 760 1250 765 1470
rect 735 1240 765 1250
rect 790 1470 900 1480
rect 790 1250 795 1470
rect 815 1250 835 1470
rect 855 1250 875 1470
rect 895 1250 900 1470
rect 790 1240 900 1250
rect 925 1470 955 1480
rect 925 1250 930 1470
rect 950 1250 955 1470
rect 925 1240 955 1250
rect 980 1470 1010 1480
rect 980 1250 985 1470
rect 1005 1250 1010 1470
rect 980 1240 1010 1250
rect 1035 1470 1065 1480
rect 1035 1250 1040 1470
rect 1060 1250 1065 1470
rect 1035 1240 1065 1250
rect 1090 1470 1120 1480
rect 1090 1250 1095 1470
rect 1115 1250 1120 1470
rect 1090 1240 1120 1250
rect 1145 1470 1175 1480
rect 1145 1250 1150 1470
rect 1170 1250 1175 1470
rect 1145 1240 1175 1250
rect 1200 1470 1270 1480
rect 1200 1250 1205 1470
rect 1225 1250 1245 1470
rect 1265 1250 1270 1470
rect 2125 1460 2135 1480
rect 2155 1460 2165 1480
rect 2125 1450 2165 1460
rect 2785 1480 2825 1490
rect 2785 1460 2795 1480
rect 2815 1460 2825 1480
rect 2785 1450 2825 1460
rect 1200 1240 1270 1250
rect 2090 1420 2160 1430
rect 550 1210 580 1220
rect 550 1190 555 1210
rect 575 1190 580 1210
rect 550 1180 580 1190
rect 620 1210 660 1220
rect 620 1190 630 1210
rect 650 1190 660 1210
rect 620 1180 660 1190
rect 700 1210 730 1220
rect 700 1190 705 1210
rect 725 1190 730 1210
rect 700 1180 730 1190
rect 960 1210 990 1220
rect 960 1190 965 1210
rect 985 1190 990 1210
rect 960 1180 990 1190
rect 1030 1210 1070 1220
rect 1030 1190 1040 1210
rect 1060 1190 1070 1210
rect 1030 1180 1070 1190
rect 1110 1210 1140 1220
rect 1110 1190 1115 1210
rect 1135 1190 1140 1210
rect 1110 1180 1140 1190
rect 545 1150 585 1160
rect 545 1130 555 1150
rect 575 1130 585 1150
rect 545 1120 585 1130
rect 120 945 150 955
rect 120 925 125 945
rect 145 925 150 945
rect 1540 945 1570 955
rect 120 915 150 925
rect 795 920 835 930
rect 795 900 805 920
rect 825 900 835 920
rect 795 890 835 900
rect 880 920 920 930
rect 880 900 890 920
rect 910 900 920 920
rect 1540 925 1545 945
rect 1565 925 1570 945
rect 1540 915 1570 925
rect 880 890 920 900
rect -470 840 -400 850
rect 680 860 750 870
rect -1501 815 -1360 825
rect -1501 795 -1495 815
rect -1475 795 -1440 815
rect -1420 795 -1385 815
rect -1365 795 -1360 815
rect -1501 785 -1360 795
rect -140 835 -70 845
rect -805 710 -765 720
rect -805 690 -795 710
rect -775 690 -765 710
rect -140 715 -135 835
rect -115 715 -95 835
rect -75 715 -70 835
rect -140 705 -70 715
rect -45 835 -15 845
rect -45 715 -40 835
rect -20 715 -15 835
rect -45 705 -15 715
rect 10 835 40 845
rect 10 715 15 835
rect 35 715 40 835
rect 10 705 40 715
rect 65 835 95 845
rect 65 715 70 835
rect 90 715 95 835
rect 65 705 95 715
rect 120 835 150 845
rect 120 715 125 835
rect 145 715 150 835
rect 120 705 150 715
rect 175 835 205 845
rect 175 715 180 835
rect 200 715 205 835
rect 175 705 205 715
rect 230 835 260 845
rect 230 715 235 835
rect 255 715 260 835
rect 230 705 260 715
rect 285 835 315 845
rect 285 715 290 835
rect 310 715 315 835
rect 285 705 315 715
rect 340 835 370 845
rect 340 715 345 835
rect 365 715 370 835
rect 340 705 370 715
rect 395 835 425 845
rect 395 715 400 835
rect 420 715 425 835
rect 395 705 425 715
rect 450 835 480 845
rect 450 715 455 835
rect 475 715 480 835
rect 450 705 480 715
rect 505 835 535 845
rect 505 715 510 835
rect 530 715 535 835
rect 505 705 535 715
rect 560 835 630 845
rect 560 715 565 835
rect 585 715 605 835
rect 625 715 630 835
rect 560 705 630 715
rect -805 680 -765 690
rect -100 675 -70 685
rect -1135 665 -1095 675
rect -1135 645 -1125 665
rect -1105 645 -1095 665
rect -1135 635 -1095 645
rect -475 665 -435 675
rect -475 645 -465 665
rect -445 645 -435 665
rect -100 655 -95 675
rect -75 655 -70 675
rect -100 645 -70 655
rect 560 675 590 685
rect 560 655 565 675
rect 585 655 590 675
rect 560 645 590 655
rect -475 635 -435 645
rect 680 640 685 860
rect 705 640 725 860
rect 745 640 750 860
rect 680 630 750 640
rect 775 860 805 870
rect 775 640 780 860
rect 800 640 805 860
rect 775 630 805 640
rect 830 860 860 870
rect 830 640 835 860
rect 855 640 860 860
rect 830 630 860 640
rect 885 860 915 870
rect 885 640 890 860
rect 910 640 915 860
rect 885 630 915 640
rect 940 860 1010 870
rect 940 640 945 860
rect 965 640 985 860
rect 1005 640 1010 860
rect 2090 850 2095 1420
rect 2115 850 2135 1420
rect 2155 850 2160 1420
rect 1060 835 1130 845
rect 1060 715 1065 835
rect 1085 715 1105 835
rect 1125 715 1130 835
rect 1060 705 1130 715
rect 1155 835 1185 845
rect 1155 715 1160 835
rect 1180 715 1185 835
rect 1155 705 1185 715
rect 1210 835 1240 845
rect 1210 715 1215 835
rect 1235 715 1240 835
rect 1210 705 1240 715
rect 1265 835 1295 845
rect 1265 715 1270 835
rect 1290 715 1295 835
rect 1265 705 1295 715
rect 1320 835 1350 845
rect 1320 715 1325 835
rect 1345 715 1350 835
rect 1320 705 1350 715
rect 1375 835 1405 845
rect 1375 715 1380 835
rect 1400 715 1405 835
rect 1375 705 1405 715
rect 1430 835 1460 845
rect 1430 715 1435 835
rect 1455 715 1460 835
rect 1430 705 1460 715
rect 1485 835 1515 845
rect 1485 715 1490 835
rect 1510 715 1515 835
rect 1485 705 1515 715
rect 1540 835 1570 845
rect 1540 715 1545 835
rect 1565 715 1570 835
rect 1540 705 1570 715
rect 1595 835 1625 845
rect 1595 715 1600 835
rect 1620 715 1625 835
rect 1595 705 1625 715
rect 1650 835 1680 845
rect 1650 715 1655 835
rect 1675 715 1680 835
rect 1650 705 1680 715
rect 1705 835 1735 845
rect 1705 715 1710 835
rect 1730 715 1735 835
rect 1705 705 1735 715
rect 1760 835 1830 845
rect 2090 840 2160 850
rect 2185 1420 2215 1430
rect 2185 850 2190 1420
rect 2210 850 2215 1420
rect 2185 840 2215 850
rect 2240 1420 2270 1430
rect 2240 850 2245 1420
rect 2265 850 2270 1420
rect 2240 840 2270 850
rect 2295 1420 2325 1430
rect 2295 850 2300 1420
rect 2320 850 2325 1420
rect 2295 840 2325 850
rect 2350 1420 2380 1430
rect 2350 850 2355 1420
rect 2375 850 2380 1420
rect 2350 840 2380 850
rect 2405 1420 2435 1430
rect 2405 850 2410 1420
rect 2430 850 2435 1420
rect 2405 840 2435 850
rect 2460 1420 2490 1430
rect 2460 850 2465 1420
rect 2485 850 2490 1420
rect 2460 840 2490 850
rect 2515 1420 2545 1430
rect 2515 850 2520 1420
rect 2540 850 2545 1420
rect 2515 840 2545 850
rect 2570 1420 2600 1430
rect 2570 850 2575 1420
rect 2595 850 2600 1420
rect 2570 840 2600 850
rect 2625 1420 2655 1430
rect 2625 850 2630 1420
rect 2650 850 2655 1420
rect 2625 840 2655 850
rect 2680 1420 2710 1430
rect 2680 850 2685 1420
rect 2705 850 2710 1420
rect 2680 840 2710 850
rect 2735 1420 2765 1430
rect 2735 850 2740 1420
rect 2760 850 2765 1420
rect 2735 840 2765 850
rect 2790 1420 2860 1430
rect 2790 850 2795 1420
rect 2815 850 2835 1420
rect 2855 850 2860 1420
rect 3050 1420 3191 1430
rect 3050 1400 3055 1420
rect 3075 1400 3110 1420
rect 3130 1400 3165 1420
rect 3185 1400 3191 1420
rect 3050 1390 3191 1400
rect 2790 840 2860 850
rect 1760 715 1765 835
rect 1785 715 1805 835
rect 1825 715 1830 835
rect 3050 815 3191 825
rect 3050 795 3055 815
rect 3075 795 3110 815
rect 3130 795 3165 815
rect 3185 795 3191 815
rect 3050 785 3191 795
rect 1760 705 1830 715
rect 2455 710 2495 720
rect 2455 690 2465 710
rect 2485 690 2495 710
rect 1100 675 1130 685
rect 1100 655 1105 675
rect 1125 655 1130 675
rect 1100 645 1130 655
rect 1760 675 1790 685
rect 2455 680 2495 690
rect 1760 655 1765 675
rect 1785 655 1790 675
rect 1760 645 1790 655
rect 2125 665 2165 675
rect 2125 645 2135 665
rect 2155 645 2165 665
rect 940 630 1010 640
rect 2125 635 2165 645
rect 2785 665 2825 675
rect 2785 645 2795 665
rect 2815 645 2825 665
rect 2785 635 2825 645
rect -1170 605 -1100 615
rect -1490 537 -1275 572
rect -1490 517 -1455 537
rect -1310 517 -1275 537
rect -1395 467 -1370 517
rect -1170 435 -1165 605
rect -1145 435 -1125 605
rect -1105 435 -1100 605
rect -1170 425 -1100 435
rect -1075 605 -1045 615
rect -1075 435 -1070 605
rect -1050 435 -1045 605
rect -1075 425 -1045 435
rect -1020 605 -990 615
rect -1020 435 -1015 605
rect -995 435 -990 605
rect -1020 425 -990 435
rect -965 605 -935 615
rect -965 435 -960 605
rect -940 435 -935 605
rect -965 425 -935 435
rect -910 605 -880 615
rect -910 435 -905 605
rect -885 435 -880 605
rect -910 425 -880 435
rect -855 605 -825 615
rect -855 435 -850 605
rect -830 435 -825 605
rect -855 425 -825 435
rect -800 605 -770 615
rect -800 435 -795 605
rect -775 435 -770 605
rect -800 425 -770 435
rect -745 605 -715 615
rect -745 435 -740 605
rect -720 435 -715 605
rect -745 425 -715 435
rect -690 605 -660 615
rect -690 435 -685 605
rect -665 435 -660 605
rect -690 425 -660 435
rect -635 605 -605 615
rect -635 435 -630 605
rect -610 435 -605 605
rect -635 425 -605 435
rect -580 605 -550 615
rect -580 435 -575 605
rect -555 435 -550 605
rect -580 425 -550 435
rect -525 605 -495 615
rect -525 435 -520 605
rect -500 435 -495 605
rect -525 425 -495 435
rect -470 605 -400 615
rect -470 435 -465 605
rect -445 435 -425 605
rect -405 435 -400 605
rect 715 600 755 610
rect 715 580 725 600
rect 745 580 755 600
rect 715 570 755 580
rect 935 600 975 610
rect 935 580 945 600
rect 965 580 975 600
rect 935 570 975 580
rect 2090 605 2160 615
rect 145 545 175 555
rect 145 525 150 545
rect 170 525 175 545
rect 145 515 175 525
rect 795 545 825 555
rect 795 525 800 545
rect 820 525 825 545
rect 795 515 825 525
rect 865 545 895 555
rect 865 525 870 545
rect 890 525 895 545
rect 865 515 895 525
rect 1515 545 1545 555
rect 1515 525 1520 545
rect 1540 525 1545 545
rect 1515 515 1545 525
rect 715 475 755 485
rect 715 455 725 475
rect 745 455 755 475
rect 715 445 755 455
rect 935 475 975 485
rect 935 455 945 475
rect 965 455 975 475
rect 935 445 975 455
rect -470 425 -400 435
rect 2090 435 2095 605
rect 2115 435 2135 605
rect 2155 435 2160 605
rect 2090 425 2160 435
rect 2185 605 2215 615
rect 2185 435 2190 605
rect 2210 435 2215 605
rect 2185 425 2215 435
rect 2240 605 2270 615
rect 2240 435 2245 605
rect 2265 435 2270 605
rect 2240 425 2270 435
rect 2295 605 2325 615
rect 2295 435 2300 605
rect 2320 435 2325 605
rect 2295 425 2325 435
rect 2350 605 2380 615
rect 2350 435 2355 605
rect 2375 435 2380 605
rect 2350 425 2380 435
rect 2405 605 2435 615
rect 2405 435 2410 605
rect 2430 435 2435 605
rect 2405 425 2435 435
rect 2460 605 2490 615
rect 2460 435 2465 605
rect 2485 435 2490 605
rect 2460 425 2490 435
rect 2515 605 2545 615
rect 2515 435 2520 605
rect 2540 435 2545 605
rect 2515 425 2545 435
rect 2570 605 2600 615
rect 2570 435 2575 605
rect 2595 435 2600 605
rect 2570 425 2600 435
rect 2625 605 2655 615
rect 2625 435 2630 605
rect 2650 435 2655 605
rect 2625 425 2655 435
rect 2680 605 2710 615
rect 2680 435 2685 605
rect 2705 435 2710 605
rect 2680 425 2710 435
rect 2735 605 2765 615
rect 2735 435 2740 605
rect 2760 435 2765 605
rect 2735 425 2765 435
rect 2790 605 2860 615
rect 2790 435 2795 605
rect 2815 435 2835 605
rect 2855 435 2860 605
rect 2790 425 2860 435
rect 2965 537 3180 572
rect 2965 517 3000 537
rect 3145 517 3180 537
rect -140 415 -70 425
rect -750 335 -710 345
rect -750 315 -740 335
rect -720 315 -710 335
rect -750 305 -710 315
rect -140 295 -135 415
rect -115 295 -95 415
rect -75 295 -70 415
rect -140 285 -70 295
rect -45 415 -15 425
rect -45 295 -40 415
rect -20 295 -15 415
rect -45 285 -15 295
rect 10 415 40 425
rect 10 295 15 415
rect 35 295 40 415
rect 10 285 40 295
rect 65 415 95 425
rect 65 295 70 415
rect 90 295 95 415
rect 65 285 95 295
rect 120 415 150 425
rect 120 295 125 415
rect 145 295 150 415
rect 120 285 150 295
rect 175 415 205 425
rect 175 295 180 415
rect 200 295 205 415
rect 175 285 205 295
rect 230 415 260 425
rect 230 295 235 415
rect 255 295 260 415
rect 230 285 260 295
rect 285 415 315 425
rect 285 295 290 415
rect 310 295 315 415
rect 285 285 315 295
rect 340 415 370 425
rect 340 295 345 415
rect 365 295 370 415
rect 340 285 370 295
rect 395 415 425 425
rect 395 295 400 415
rect 420 295 425 415
rect 395 285 425 295
rect 450 415 480 425
rect 450 295 455 415
rect 475 295 480 415
rect 450 285 480 295
rect 505 415 535 425
rect 505 295 510 415
rect 530 295 535 415
rect 505 285 535 295
rect 560 415 630 425
rect 560 295 565 415
rect 585 295 605 415
rect 625 295 630 415
rect 560 285 630 295
rect 680 415 750 425
rect 680 295 685 415
rect 705 295 725 415
rect 745 295 750 415
rect 680 285 750 295
rect 775 415 805 425
rect 775 295 780 415
rect 800 295 805 415
rect 775 285 805 295
rect 830 415 860 425
rect 830 295 835 415
rect 855 295 860 415
rect 830 285 860 295
rect 885 415 915 425
rect 885 295 890 415
rect 910 295 915 415
rect 885 285 915 295
rect 940 415 1010 425
rect 940 295 945 415
rect 965 295 985 415
rect 1005 295 1010 415
rect 940 285 1010 295
rect 1060 415 1130 425
rect 1060 295 1065 415
rect 1085 295 1105 415
rect 1125 295 1130 415
rect 1060 285 1130 295
rect 1155 415 1185 425
rect 1155 295 1160 415
rect 1180 295 1185 415
rect 1155 285 1185 295
rect 1210 415 1240 425
rect 1210 295 1215 415
rect 1235 295 1240 415
rect 1210 285 1240 295
rect 1265 415 1295 425
rect 1265 295 1270 415
rect 1290 295 1295 415
rect 1265 285 1295 295
rect 1320 415 1350 425
rect 1320 295 1325 415
rect 1345 295 1350 415
rect 1320 285 1350 295
rect 1375 415 1405 425
rect 1375 295 1380 415
rect 1400 295 1405 415
rect 1375 285 1405 295
rect 1430 415 1460 425
rect 1430 295 1435 415
rect 1455 295 1460 415
rect 1430 285 1460 295
rect 1485 415 1515 425
rect 1485 295 1490 415
rect 1510 295 1515 415
rect 1485 285 1515 295
rect 1540 415 1570 425
rect 1540 295 1545 415
rect 1565 295 1570 415
rect 1540 285 1570 295
rect 1595 415 1625 425
rect 1595 295 1600 415
rect 1620 295 1625 415
rect 1595 285 1625 295
rect 1650 415 1680 425
rect 1650 295 1655 415
rect 1675 295 1680 415
rect 1650 285 1680 295
rect 1705 415 1735 425
rect 1705 295 1710 415
rect 1730 295 1735 415
rect 1705 285 1735 295
rect 1760 415 1830 425
rect 1760 295 1765 415
rect 1785 295 1805 415
rect 1825 295 1830 415
rect 2400 335 2440 345
rect 2400 315 2410 335
rect 2430 315 2440 335
rect 2400 305 2440 315
rect 3060 467 3085 517
rect 1760 285 1830 295
rect -100 255 -70 265
rect -100 235 -95 255
rect -75 235 -70 255
rect -100 225 -70 235
rect 560 255 590 265
rect 560 235 565 255
rect 585 235 590 255
rect 560 225 590 235
rect 1100 255 1130 265
rect 1100 235 1105 255
rect 1125 235 1130 255
rect 1100 225 1130 235
rect 1760 255 1790 265
rect 1760 235 1765 255
rect 1785 235 1790 255
rect 1760 225 1790 235
rect -1170 215 -1100 225
rect -1490 -93 -1455 -85
rect -1490 -113 -1485 -93
rect -1460 -113 -1455 -93
rect -1490 -120 -1455 -113
rect -1430 -93 -1395 -85
rect -1430 -113 -1425 -93
rect -1400 -113 -1395 -93
rect -1430 -120 -1395 -113
rect -1370 -93 -1335 -85
rect -1370 -113 -1365 -93
rect -1340 -113 -1335 -93
rect -1370 -120 -1335 -113
rect -1170 -55 -1165 215
rect -1145 -55 -1125 215
rect -1105 -55 -1100 215
rect -1170 -65 -1100 -55
rect -1075 215 -1045 225
rect -1075 -55 -1070 215
rect -1050 -55 -1045 215
rect -1075 -65 -1045 -55
rect -1020 215 -990 225
rect -1020 -55 -1015 215
rect -995 -55 -990 215
rect -1020 -65 -990 -55
rect -965 215 -935 225
rect -965 -55 -960 215
rect -940 -55 -935 215
rect -965 -65 -935 -55
rect -910 215 -880 225
rect -910 -55 -905 215
rect -885 -55 -880 215
rect -910 -65 -880 -55
rect -855 215 -825 225
rect -855 -55 -850 215
rect -830 -55 -825 215
rect -855 -65 -825 -55
rect -800 215 -770 225
rect -800 -55 -795 215
rect -775 -55 -770 215
rect -800 -65 -770 -55
rect -745 215 -715 225
rect -745 -55 -740 215
rect -720 -55 -715 215
rect -745 -65 -715 -55
rect -690 215 -660 225
rect -690 -55 -685 215
rect -665 -55 -660 215
rect -690 -65 -660 -55
rect -635 215 -605 225
rect -635 -55 -630 215
rect -610 -55 -605 215
rect -635 -65 -605 -55
rect -580 215 -550 225
rect -580 -55 -575 215
rect -555 -55 -550 215
rect -580 -65 -550 -55
rect -525 215 -495 225
rect -525 -55 -520 215
rect -500 -55 -495 215
rect -525 -65 -495 -55
rect -470 215 -400 225
rect -470 -55 -465 215
rect -445 -55 -425 215
rect -405 -55 -400 215
rect 2090 215 2160 225
rect 830 -15 860 -5
rect 830 -35 835 -15
rect 855 -35 860 -15
rect 830 -45 860 -35
rect -470 -65 -400 -55
rect 2090 -55 2095 215
rect 2115 -55 2135 215
rect 2155 -55 2160 215
rect 2090 -65 2160 -55
rect 2185 215 2215 225
rect 2185 -55 2190 215
rect 2210 -55 2215 215
rect 2185 -65 2215 -55
rect 2240 215 2270 225
rect 2240 -55 2245 215
rect 2265 -55 2270 215
rect 2240 -65 2270 -55
rect 2295 215 2325 225
rect 2295 -55 2300 215
rect 2320 -55 2325 215
rect 2295 -65 2325 -55
rect 2350 215 2380 225
rect 2350 -55 2355 215
rect 2375 -55 2380 215
rect 2350 -65 2380 -55
rect 2405 215 2435 225
rect 2405 -55 2410 215
rect 2430 -55 2435 215
rect 2405 -65 2435 -55
rect 2460 215 2490 225
rect 2460 -55 2465 215
rect 2485 -55 2490 215
rect 2460 -65 2490 -55
rect 2515 215 2545 225
rect 2515 -55 2520 215
rect 2540 -55 2545 215
rect 2515 -65 2545 -55
rect 2570 215 2600 225
rect 2570 -55 2575 215
rect 2595 -55 2600 215
rect 2570 -65 2600 -55
rect 2625 215 2655 225
rect 2625 -55 2630 215
rect 2650 -55 2655 215
rect 2625 -65 2655 -55
rect 2680 215 2710 225
rect 2680 -55 2685 215
rect 2705 -55 2710 215
rect 2680 -65 2710 -55
rect 2735 215 2765 225
rect 2735 -55 2740 215
rect 2760 -55 2765 215
rect 2735 -65 2765 -55
rect 2790 215 2860 225
rect 2790 -55 2795 215
rect 2815 -55 2835 215
rect 2855 -55 2860 215
rect 2790 -65 2860 -55
rect 680 -80 750 -70
rect -1310 -93 -1275 -85
rect -1310 -113 -1305 -93
rect -1280 -113 -1275 -93
rect -1310 -120 -1275 -113
rect -1135 -95 -1095 -85
rect -1135 -115 -1125 -95
rect -1105 -115 -1095 -95
rect -1135 -125 -1095 -115
rect -475 -95 -435 -85
rect -475 -115 -465 -95
rect -445 -115 -435 -95
rect -475 -125 -435 -115
rect -805 -250 -765 -240
rect -805 -270 -795 -250
rect -775 -270 -765 -250
rect -805 -280 -765 -270
rect 680 -300 685 -80
rect 705 -300 725 -80
rect 745 -300 750 -80
rect 680 -310 750 -300
rect 775 -80 805 -70
rect 775 -300 780 -80
rect 800 -300 805 -80
rect 775 -310 805 -300
rect 830 -80 860 -70
rect 830 -300 835 -80
rect 855 -300 860 -80
rect 830 -310 860 -300
rect 885 -80 915 -70
rect 885 -300 890 -80
rect 910 -300 915 -80
rect 885 -310 915 -300
rect 940 -80 1010 -70
rect 940 -300 945 -80
rect 965 -300 985 -80
rect 1005 -300 1010 -80
rect 2125 -95 2165 -85
rect 2125 -115 2135 -95
rect 2155 -115 2165 -95
rect 2125 -125 2165 -115
rect 2785 -95 2825 -85
rect 2785 -115 2795 -95
rect 2815 -115 2825 -95
rect 2785 -125 2825 -115
rect 2965 -93 3000 -85
rect 2965 -113 2970 -93
rect 2995 -113 3000 -93
rect 2965 -120 3000 -113
rect 3025 -93 3060 -85
rect 3025 -113 3030 -93
rect 3055 -113 3060 -93
rect 3025 -120 3060 -113
rect 3085 -93 3120 -85
rect 3085 -113 3090 -93
rect 3115 -113 3120 -93
rect 3085 -120 3120 -113
rect 3145 -93 3180 -85
rect 3145 -113 3150 -93
rect 3175 -113 3180 -93
rect 3145 -120 3180 -113
rect 2455 -250 2495 -240
rect 2455 -270 2465 -250
rect 2485 -270 2495 -250
rect 2455 -280 2495 -270
rect 940 -310 1010 -300
rect 715 -340 755 -330
rect 715 -360 725 -340
rect 745 -360 755 -340
rect -1140 -370 -1070 -360
rect -1290 -387 -1255 -380
rect -1290 -407 -1285 -387
rect -1260 -407 -1255 -387
rect -1290 -415 -1255 -407
rect -1230 -387 -1195 -380
rect -1230 -407 -1225 -387
rect -1200 -407 -1195 -387
rect -1230 -415 -1195 -407
rect -1255 -1105 -1230 -1055
rect -1140 -1040 -1135 -370
rect -1115 -1040 -1095 -370
rect -1075 -1040 -1070 -370
rect -1140 -1050 -1070 -1040
rect -1000 -370 -970 -360
rect -1000 -1040 -995 -370
rect -975 -1040 -970 -370
rect -1000 -1050 -970 -1040
rect -900 -370 -870 -360
rect -900 -1040 -895 -370
rect -875 -1040 -870 -370
rect -900 -1050 -870 -1040
rect -800 -370 -770 -360
rect -800 -1040 -795 -370
rect -775 -1040 -770 -370
rect -800 -1050 -770 -1040
rect -700 -370 -670 -360
rect -700 -1040 -695 -370
rect -675 -1040 -670 -370
rect -700 -1050 -670 -1040
rect -600 -370 -570 -360
rect -600 -1040 -595 -370
rect -575 -1040 -570 -370
rect -600 -1050 -570 -1040
rect -500 -370 -430 -360
rect 715 -370 755 -360
rect 935 -340 975 -330
rect 935 -360 945 -340
rect 965 -360 975 -340
rect 935 -370 975 -360
rect 2120 -370 2190 -360
rect -500 -1040 -495 -370
rect -475 -1040 -455 -370
rect -435 -1040 -430 -370
rect 445 -440 475 -430
rect 445 -460 450 -440
rect 470 -460 475 -440
rect 445 -470 475 -460
rect 1350 -440 1390 -430
rect 1350 -460 1360 -440
rect 1380 -460 1390 -440
rect 1350 -470 1390 -460
rect 240 -550 310 -540
rect 240 -770 245 -550
rect 265 -770 285 -550
rect 305 -770 310 -550
rect 240 -780 310 -770
rect 335 -550 365 -540
rect 335 -770 340 -550
rect 360 -770 365 -550
rect 335 -780 365 -770
rect 390 -550 420 -540
rect 390 -770 395 -550
rect 415 -770 420 -550
rect 390 -780 420 -770
rect 445 -550 475 -540
rect 445 -770 450 -550
rect 470 -770 475 -550
rect 445 -780 475 -770
rect 500 -550 530 -540
rect 500 -770 505 -550
rect 525 -770 530 -550
rect 500 -780 530 -770
rect 555 -550 585 -540
rect 555 -770 560 -550
rect 580 -770 585 -550
rect 555 -780 585 -770
rect 610 -550 640 -540
rect 610 -770 615 -550
rect 635 -770 640 -550
rect 610 -780 640 -770
rect 665 -550 695 -540
rect 665 -770 670 -550
rect 690 -770 695 -550
rect 665 -780 695 -770
rect 720 -550 750 -540
rect 720 -770 725 -550
rect 745 -770 750 -550
rect 720 -780 750 -770
rect 775 -550 805 -540
rect 775 -770 780 -550
rect 800 -770 805 -550
rect 775 -780 805 -770
rect 830 -550 860 -540
rect 830 -770 835 -550
rect 855 -770 860 -550
rect 830 -780 860 -770
rect 885 -550 915 -540
rect 885 -770 890 -550
rect 910 -770 915 -550
rect 885 -780 915 -770
rect 940 -550 970 -540
rect 940 -770 945 -550
rect 965 -770 970 -550
rect 940 -780 970 -770
rect 995 -550 1025 -540
rect 995 -770 1000 -550
rect 1020 -770 1025 -550
rect 995 -780 1025 -770
rect 1050 -550 1080 -540
rect 1050 -770 1055 -550
rect 1075 -770 1080 -550
rect 1050 -780 1080 -770
rect 1105 -550 1135 -540
rect 1105 -770 1110 -550
rect 1130 -770 1135 -550
rect 1105 -780 1135 -770
rect 1160 -550 1190 -540
rect 1160 -770 1165 -550
rect 1185 -770 1190 -550
rect 1160 -780 1190 -770
rect 1215 -550 1245 -540
rect 1215 -770 1220 -550
rect 1240 -770 1245 -550
rect 1215 -780 1245 -770
rect 1270 -550 1300 -540
rect 1270 -770 1275 -550
rect 1295 -770 1300 -550
rect 1270 -780 1300 -770
rect 1325 -550 1355 -540
rect 1325 -770 1330 -550
rect 1350 -770 1355 -550
rect 1325 -780 1355 -770
rect 1380 -550 1410 -540
rect 1380 -770 1385 -550
rect 1405 -770 1410 -550
rect 1380 -780 1410 -770
rect 1435 -550 1505 -540
rect 1435 -770 1440 -550
rect 1460 -770 1480 -550
rect 1500 -770 1505 -550
rect 1435 -780 1505 -770
rect 275 -810 330 -800
rect 275 -830 285 -810
rect 305 -820 330 -810
rect 1415 -810 1470 -800
rect 1415 -820 1440 -810
rect 305 -830 315 -820
rect 275 -840 315 -830
rect 1430 -830 1440 -820
rect 1460 -830 1470 -810
rect 1430 -840 1470 -830
rect 650 -965 690 -955
rect 650 -985 660 -965
rect 680 -985 690 -965
rect 650 -995 690 -985
rect 1095 -965 1135 -955
rect 1095 -985 1105 -965
rect 1125 -985 1135 -965
rect 1095 -995 1135 -985
rect -500 -1050 -430 -1040
rect 450 -1025 520 -1015
rect -1105 -1080 -1065 -1070
rect -1105 -1100 -1095 -1080
rect -1075 -1100 -1065 -1080
rect -1105 -1110 -1065 -1100
rect -505 -1080 -465 -1070
rect -505 -1100 -495 -1080
rect -475 -1100 -465 -1080
rect -505 -1110 -465 -1100
rect 450 -1145 455 -1025
rect 475 -1145 495 -1025
rect 515 -1145 520 -1025
rect 450 -1155 520 -1145
rect 545 -1025 575 -1015
rect 545 -1145 550 -1025
rect 570 -1145 575 -1025
rect 545 -1155 575 -1145
rect 600 -1025 630 -1015
rect 600 -1145 605 -1025
rect 625 -1145 630 -1025
rect 600 -1155 630 -1145
rect 655 -1025 685 -1015
rect 655 -1145 660 -1025
rect 680 -1145 685 -1025
rect 655 -1155 685 -1145
rect 710 -1025 740 -1015
rect 710 -1145 715 -1025
rect 735 -1145 740 -1025
rect 710 -1155 740 -1145
rect 765 -1025 795 -1015
rect 765 -1145 770 -1025
rect 790 -1145 795 -1025
rect 765 -1155 795 -1145
rect 820 -1025 890 -1015
rect 820 -1145 825 -1025
rect 845 -1145 865 -1025
rect 885 -1145 890 -1025
rect 820 -1155 890 -1145
rect 930 -1025 960 -1015
rect 930 -1145 935 -1025
rect 955 -1145 960 -1025
rect 930 -1155 960 -1145
rect 1270 -1025 1300 -1015
rect 1270 -1145 1275 -1025
rect 1295 -1145 1300 -1025
rect 2120 -1040 2125 -370
rect 2145 -1040 2165 -370
rect 2185 -1040 2190 -370
rect 2120 -1050 2190 -1040
rect 2260 -370 2290 -360
rect 2260 -1040 2265 -370
rect 2285 -1040 2290 -370
rect 2260 -1050 2290 -1040
rect 2360 -370 2390 -360
rect 2360 -1040 2365 -370
rect 2385 -1040 2390 -370
rect 2360 -1050 2390 -1040
rect 2460 -370 2490 -360
rect 2460 -1040 2465 -370
rect 2485 -1040 2490 -370
rect 2460 -1050 2490 -1040
rect 2560 -370 2590 -360
rect 2560 -1040 2565 -370
rect 2585 -1040 2590 -370
rect 2560 -1050 2590 -1040
rect 2660 -370 2690 -360
rect 2660 -1040 2665 -370
rect 2685 -1040 2690 -370
rect 2660 -1050 2690 -1040
rect 2760 -370 2830 -360
rect 2760 -1040 2765 -370
rect 2785 -1040 2805 -370
rect 2825 -1040 2830 -370
rect 2885 -387 2920 -380
rect 2885 -407 2890 -387
rect 2915 -407 2920 -387
rect 2885 -415 2920 -407
rect 2945 -387 2980 -380
rect 2945 -407 2950 -387
rect 2975 -407 2980 -387
rect 2945 -415 2980 -407
rect 2760 -1050 2830 -1040
rect 2155 -1080 2195 -1070
rect 2155 -1100 2165 -1080
rect 2185 -1100 2195 -1080
rect 2155 -1110 2195 -1100
rect 2755 -1080 2795 -1070
rect 2755 -1100 2765 -1080
rect 2785 -1100 2795 -1080
rect 2755 -1110 2795 -1100
rect 2920 -1105 2945 -1055
rect 1270 -1155 1300 -1145
rect 490 -1185 520 -1175
rect 490 -1205 495 -1185
rect 515 -1205 520 -1185
rect 490 -1215 520 -1205
rect 820 -1185 850 -1175
rect 820 -1205 825 -1185
rect 845 -1205 850 -1185
rect 820 -1215 850 -1205
<< viali >>
rect 40 2700 60 2720
rect 220 2700 240 2720
rect 980 2700 1000 2720
rect 1160 2700 1180 2720
rect 1450 2700 1470 2720
rect 1630 2700 1650 2720
rect 40 2340 60 2660
rect 100 2340 120 2660
rect 160 2340 180 2660
rect 220 2340 240 2660
rect 510 2530 530 2550
rect 570 2530 590 2550
rect 690 2530 710 2550
rect 510 2340 530 2490
rect 570 2340 590 2490
rect 630 2340 650 2490
rect 690 2340 710 2490
rect 980 2340 1000 2660
rect 1040 2340 1060 2660
rect 1100 2340 1120 2660
rect 1160 2340 1180 2660
rect 1450 2340 1470 2660
rect 1510 2340 1530 2660
rect 1570 2340 1590 2660
rect 1630 2340 1650 2660
rect 85 2280 105 2300
rect 144 2280 164 2300
rect 614 2280 634 2300
rect 1056 2280 1076 2300
rect 1526 2280 1546 2300
rect -435 2125 -415 2145
rect -30 2125 -10 2145
rect 690 2125 710 2145
rect 980 2125 1000 2145
rect 1700 2125 1720 2145
rect 2105 2125 2125 2145
rect -1155 1765 -1135 2085
rect -1095 1765 -1075 2085
rect -1035 1765 -1015 2085
rect -975 1765 -955 2085
rect -915 1765 -895 2085
rect -855 1765 -835 2085
rect -795 1765 -775 2085
rect -735 1765 -715 2085
rect -675 1765 -655 2085
rect -615 1765 -595 2085
rect -555 1765 -535 2085
rect -495 1765 -475 2085
rect -435 1765 -415 2085
rect -30 1765 -10 2085
rect 30 1765 50 2085
rect 90 1765 110 2085
rect 150 1765 170 2085
rect 210 1765 230 2085
rect 270 1765 290 2085
rect 330 1765 350 2085
rect 390 1765 410 2085
rect 450 1765 470 2085
rect 510 1765 530 2085
rect 570 1765 590 2085
rect 630 1765 650 2085
rect 690 1765 710 2085
rect 980 1765 1000 2085
rect 1040 1765 1060 2085
rect 1100 1765 1120 2085
rect 1160 1765 1180 2085
rect 1220 1765 1240 2085
rect 1280 1765 1300 2085
rect 1340 1765 1360 2085
rect 1400 1765 1420 2085
rect 1460 1765 1480 2085
rect 1520 1765 1540 2085
rect 1580 1765 1600 2085
rect 1640 1765 1660 2085
rect 1700 1765 1720 2085
rect 2105 1765 2125 2085
rect 2165 1765 2185 2085
rect 2225 1765 2245 2085
rect 2285 1765 2305 2085
rect 2345 1765 2365 2085
rect 2405 1765 2425 2085
rect 2465 1765 2485 2085
rect 2525 1765 2545 2085
rect 2585 1765 2605 2085
rect 2645 1765 2665 2085
rect 2705 1765 2725 2085
rect 2765 1765 2785 2085
rect 2825 1765 2845 2085
rect 420 1645 440 1665
rect 1250 1645 1270 1665
rect -705 1600 -685 1620
rect 2375 1600 2395 1620
rect 465 1540 485 1560
rect 795 1540 815 1560
rect 875 1540 895 1560
rect 1205 1540 1225 1560
rect -1125 1460 -1105 1480
rect -465 1460 -445 1480
rect -1495 1400 -1475 1420
rect -1440 1400 -1420 1420
rect -1385 1400 -1365 1420
rect -1125 850 -1105 1420
rect -1070 850 -1050 1420
rect -1015 850 -995 1420
rect -960 850 -940 1420
rect -905 850 -885 1420
rect -850 850 -830 1420
rect -795 850 -775 1420
rect -740 850 -720 1420
rect -685 850 -665 1420
rect -630 850 -610 1420
rect -575 850 -555 1420
rect -520 850 -500 1420
rect -465 850 -445 1420
rect 465 1250 485 1470
rect 520 1250 540 1470
rect 575 1250 595 1470
rect 630 1250 650 1470
rect 685 1250 705 1470
rect 740 1250 760 1470
rect 795 1250 815 1470
rect 875 1250 895 1470
rect 930 1250 950 1470
rect 985 1250 1005 1470
rect 1040 1250 1060 1470
rect 1095 1250 1115 1470
rect 1150 1250 1170 1470
rect 1205 1250 1225 1470
rect 2135 1460 2155 1480
rect 2795 1460 2815 1480
rect 555 1190 575 1210
rect 630 1190 650 1210
rect 705 1190 725 1210
rect 965 1190 985 1210
rect 1040 1190 1060 1210
rect 1115 1190 1135 1210
rect 555 1130 575 1150
rect 125 925 145 945
rect 805 900 825 920
rect 890 900 910 920
rect 1545 925 1565 945
rect -1495 795 -1475 815
rect -1440 795 -1420 815
rect -1385 795 -1365 815
rect -795 690 -775 710
rect -95 715 -75 835
rect -40 715 -20 835
rect 15 715 35 835
rect 70 715 90 835
rect 125 715 145 835
rect 180 715 200 835
rect 235 715 255 835
rect 290 715 310 835
rect 345 715 365 835
rect 400 715 420 835
rect 455 715 475 835
rect 510 715 530 835
rect 565 715 585 835
rect -1125 645 -1105 665
rect -465 645 -445 665
rect -95 655 -75 675
rect 565 655 585 675
rect 725 640 745 860
rect 780 640 800 860
rect 835 640 855 860
rect 890 640 910 860
rect 945 640 965 860
rect 2135 850 2155 1420
rect 1105 715 1125 835
rect 1160 715 1180 835
rect 1215 715 1235 835
rect 1270 715 1290 835
rect 1325 715 1345 835
rect 1380 715 1400 835
rect 1435 715 1455 835
rect 1490 715 1510 835
rect 1545 715 1565 835
rect 1600 715 1620 835
rect 1655 715 1675 835
rect 1710 715 1730 835
rect 2190 850 2210 1420
rect 2245 850 2265 1420
rect 2300 850 2320 1420
rect 2355 850 2375 1420
rect 2410 850 2430 1420
rect 2465 850 2485 1420
rect 2520 850 2540 1420
rect 2575 850 2595 1420
rect 2630 850 2650 1420
rect 2685 850 2705 1420
rect 2740 850 2760 1420
rect 2795 850 2815 1420
rect 3055 1400 3075 1420
rect 3110 1400 3130 1420
rect 3165 1400 3185 1420
rect 1765 715 1785 835
rect 3055 795 3075 815
rect 3110 795 3130 815
rect 3165 795 3185 815
rect 2465 690 2485 710
rect 1105 655 1125 675
rect 1765 655 1785 675
rect 2135 645 2155 665
rect 2795 645 2815 665
rect -1125 435 -1105 605
rect -1070 435 -1050 605
rect -1015 435 -995 605
rect -960 435 -940 605
rect -905 435 -885 605
rect -850 435 -830 605
rect -795 435 -775 605
rect -740 435 -720 605
rect -685 435 -665 605
rect -630 435 -610 605
rect -575 435 -555 605
rect -520 435 -500 605
rect -465 435 -445 605
rect 725 580 745 600
rect 945 580 965 600
rect 150 525 170 545
rect 800 525 820 545
rect 870 525 890 545
rect 1520 525 1540 545
rect 725 455 745 475
rect 945 455 965 475
rect 2135 435 2155 605
rect 2190 435 2210 605
rect 2245 435 2265 605
rect 2300 435 2320 605
rect 2355 435 2375 605
rect 2410 435 2430 605
rect 2465 435 2485 605
rect 2520 435 2540 605
rect 2575 435 2595 605
rect 2630 435 2650 605
rect 2685 435 2705 605
rect 2740 435 2760 605
rect 2795 435 2815 605
rect -740 315 -720 335
rect -95 295 -75 415
rect -40 295 -20 415
rect 15 295 35 415
rect 70 295 90 415
rect 125 295 145 415
rect 180 295 200 415
rect 235 295 255 415
rect 290 295 310 415
rect 345 295 365 415
rect 400 295 420 415
rect 455 295 475 415
rect 510 295 530 415
rect 565 295 585 415
rect 725 295 745 415
rect 780 295 800 415
rect 835 295 855 415
rect 890 295 910 415
rect 945 295 965 415
rect 1105 295 1125 415
rect 1160 295 1180 415
rect 1215 295 1235 415
rect 1270 295 1290 415
rect 1325 295 1345 415
rect 1380 295 1400 415
rect 1435 295 1455 415
rect 1490 295 1510 415
rect 1545 295 1565 415
rect 1600 295 1620 415
rect 1655 295 1675 415
rect 1710 295 1730 415
rect 1765 295 1785 415
rect 2410 315 2430 335
rect -95 235 -75 255
rect 565 235 585 255
rect 1105 235 1125 255
rect 1765 235 1785 255
rect -1485 -113 -1460 -93
rect -1425 -113 -1400 -93
rect -1365 -113 -1340 -93
rect -1125 -55 -1105 215
rect -1070 -55 -1050 215
rect -1015 -55 -995 215
rect -960 -55 -940 215
rect -905 -55 -885 215
rect -850 -55 -830 215
rect -795 -55 -775 215
rect -740 -55 -720 215
rect -685 -55 -665 215
rect -630 -55 -610 215
rect -575 -55 -555 215
rect -520 -55 -500 215
rect -465 -55 -445 215
rect 835 -35 855 -15
rect 2135 -55 2155 215
rect 2190 -55 2210 215
rect 2245 -55 2265 215
rect 2300 -55 2320 215
rect 2355 -55 2375 215
rect 2410 -55 2430 215
rect 2465 -55 2485 215
rect 2520 -55 2540 215
rect 2575 -55 2595 215
rect 2630 -55 2650 215
rect 2685 -55 2705 215
rect 2740 -55 2760 215
rect 2795 -55 2815 215
rect -1305 -113 -1280 -93
rect -1125 -115 -1105 -95
rect -465 -115 -445 -95
rect -795 -270 -775 -250
rect 725 -300 745 -80
rect 780 -300 800 -80
rect 835 -300 855 -80
rect 890 -300 910 -80
rect 945 -300 965 -80
rect 2135 -115 2155 -95
rect 2795 -115 2815 -95
rect 2970 -113 2995 -93
rect 3030 -113 3055 -93
rect 3090 -113 3115 -93
rect 3150 -113 3175 -93
rect 2465 -270 2485 -250
rect 725 -360 745 -340
rect -1285 -407 -1260 -387
rect -1225 -407 -1200 -387
rect -1095 -1040 -1075 -370
rect -995 -1040 -975 -370
rect -895 -1040 -875 -370
rect -795 -1040 -775 -370
rect -695 -1040 -675 -370
rect -595 -1040 -575 -370
rect 945 -360 965 -340
rect -495 -1040 -475 -370
rect 450 -460 470 -440
rect 1360 -460 1380 -440
rect 285 -770 305 -550
rect 340 -770 360 -550
rect 395 -770 415 -550
rect 450 -770 470 -550
rect 505 -770 525 -550
rect 560 -770 580 -550
rect 615 -770 635 -550
rect 670 -770 690 -550
rect 725 -770 745 -550
rect 780 -770 800 -550
rect 835 -770 855 -550
rect 890 -770 910 -550
rect 945 -770 965 -550
rect 1000 -770 1020 -550
rect 1055 -770 1075 -550
rect 1110 -770 1130 -550
rect 1165 -770 1185 -550
rect 1220 -770 1240 -550
rect 1275 -770 1295 -550
rect 1330 -770 1350 -550
rect 1385 -770 1405 -550
rect 1440 -770 1460 -550
rect 285 -830 305 -810
rect 1440 -830 1460 -810
rect 660 -985 680 -965
rect 1105 -985 1125 -965
rect -1095 -1100 -1075 -1080
rect -495 -1100 -475 -1080
rect 495 -1145 515 -1025
rect 550 -1145 570 -1025
rect 605 -1145 625 -1025
rect 660 -1145 680 -1025
rect 715 -1145 735 -1025
rect 770 -1145 790 -1025
rect 825 -1145 845 -1025
rect 935 -1145 955 -1025
rect 1275 -1145 1295 -1025
rect 2165 -1040 2185 -370
rect 2265 -1040 2285 -370
rect 2365 -1040 2385 -370
rect 2465 -1040 2485 -370
rect 2565 -1040 2585 -370
rect 2665 -1040 2685 -370
rect 2765 -1040 2785 -370
rect 2890 -407 2915 -387
rect 2950 -407 2975 -387
rect 2165 -1100 2185 -1080
rect 2765 -1100 2785 -1080
rect 495 -1205 515 -1185
rect 825 -1205 845 -1185
<< metal1 >>
rect 825 4275 865 4280
rect 825 4245 830 4275
rect 860 4245 865 4275
rect 825 4240 865 4245
rect 210 2780 250 2785
rect 210 2750 215 2780
rect 245 2750 250 2780
rect 30 2725 70 2730
rect 30 2695 35 2725
rect 65 2695 70 2725
rect 30 2690 70 2695
rect 150 2725 190 2730
rect 150 2695 155 2725
rect 185 2695 190 2725
rect 150 2690 190 2695
rect 210 2725 250 2750
rect 620 2780 660 2785
rect 620 2750 625 2780
rect 655 2750 660 2780
rect 620 2745 660 2750
rect 210 2695 215 2725
rect 245 2695 250 2725
rect 210 2690 250 2695
rect 35 2660 65 2690
rect 35 2340 40 2660
rect 60 2340 65 2660
rect 35 2330 65 2340
rect 95 2660 125 2670
rect 95 2340 100 2660
rect 120 2340 125 2660
rect 95 2330 125 2340
rect 155 2660 185 2690
rect 155 2340 160 2660
rect 180 2340 185 2660
rect 155 2330 185 2340
rect 215 2660 245 2690
rect 215 2340 220 2660
rect 240 2340 245 2660
rect 500 2555 540 2560
rect 500 2525 505 2555
rect 535 2525 540 2555
rect 500 2520 540 2525
rect 560 2555 600 2560
rect 560 2525 565 2555
rect 595 2525 600 2555
rect 560 2520 600 2525
rect 215 2330 245 2340
rect 505 2490 535 2520
rect 505 2340 510 2490
rect 530 2340 535 2490
rect 505 2330 535 2340
rect 565 2490 595 2520
rect 630 2500 650 2745
rect 835 2730 855 4240
rect 1030 2780 1070 2785
rect 1030 2750 1035 2780
rect 1065 2750 1070 2780
rect 1030 2745 1070 2750
rect 1440 2780 1480 2785
rect 1440 2750 1445 2780
rect 1475 2750 1480 2780
rect 825 2725 865 2730
rect 825 2695 830 2725
rect 860 2695 865 2725
rect 825 2690 865 2695
rect 970 2725 1010 2730
rect 970 2695 975 2725
rect 1005 2695 1010 2725
rect 970 2690 1010 2695
rect 835 2560 855 2690
rect 975 2660 1005 2690
rect 680 2555 720 2560
rect 680 2525 685 2555
rect 715 2525 720 2555
rect 680 2520 720 2525
rect 825 2555 865 2560
rect 825 2525 830 2555
rect 860 2525 865 2555
rect 825 2520 865 2525
rect 565 2340 570 2490
rect 590 2340 595 2490
rect 565 2330 595 2340
rect 625 2490 655 2500
rect 625 2340 630 2490
rect 650 2340 655 2490
rect 625 2330 655 2340
rect 685 2490 715 2500
rect 685 2340 690 2490
rect 710 2340 715 2490
rect 685 2330 715 2340
rect 75 2305 115 2310
rect 75 2275 80 2305
rect 110 2275 115 2305
rect 75 2270 115 2275
rect 139 2305 169 2310
rect 139 2270 169 2275
rect 609 2305 639 2310
rect 609 2270 639 2275
rect 770 2305 810 2310
rect 770 2275 775 2305
rect 805 2275 810 2305
rect 770 2270 810 2275
rect -805 2205 -765 2210
rect -805 2175 -800 2205
rect -770 2175 -765 2205
rect -805 2170 -765 2175
rect -235 2205 -195 2210
rect -235 2175 -230 2205
rect -200 2175 -195 2205
rect -235 2170 -195 2175
rect -800 2155 -770 2170
rect -1165 2150 -1125 2155
rect -1165 2120 -1160 2150
rect -1130 2120 -1125 2150
rect -1165 2115 -1125 2120
rect -1045 2150 -1005 2155
rect -1045 2120 -1040 2150
rect -1010 2120 -1005 2150
rect -1045 2115 -1005 2120
rect -925 2150 -885 2155
rect -925 2120 -920 2150
rect -890 2120 -885 2150
rect -925 2115 -885 2120
rect -805 2150 -765 2155
rect -805 2120 -800 2150
rect -770 2120 -765 2150
rect -805 2115 -765 2120
rect -685 2150 -645 2155
rect -685 2120 -680 2150
rect -650 2120 -645 2150
rect -685 2115 -645 2120
rect -565 2150 -525 2155
rect -565 2120 -560 2150
rect -530 2120 -525 2150
rect -565 2115 -525 2120
rect -445 2150 -405 2155
rect -445 2120 -440 2150
rect -410 2120 -405 2150
rect -445 2115 -405 2120
rect -280 2150 -240 2155
rect -280 2120 -275 2150
rect -245 2120 -240 2150
rect -280 2115 -240 2120
rect -1160 2085 -1130 2115
rect -1160 1765 -1155 2085
rect -1135 1765 -1130 2085
rect -1160 1755 -1130 1765
rect -1100 2085 -1070 2095
rect -1100 1765 -1095 2085
rect -1075 1765 -1070 2085
rect -1100 1735 -1070 1765
rect -1040 2085 -1010 2115
rect -1040 1765 -1035 2085
rect -1015 1765 -1010 2085
rect -1040 1755 -1010 1765
rect -980 2085 -950 2095
rect -980 1765 -975 2085
rect -955 1765 -950 2085
rect -980 1735 -950 1765
rect -920 2085 -890 2115
rect -920 1765 -915 2085
rect -895 1765 -890 2085
rect -920 1755 -890 1765
rect -860 2085 -830 2095
rect -860 1765 -855 2085
rect -835 1765 -830 2085
rect -860 1735 -830 1765
rect -800 2085 -770 2115
rect -800 1765 -795 2085
rect -775 1765 -770 2085
rect -800 1755 -770 1765
rect -740 2085 -710 2095
rect -740 1765 -735 2085
rect -715 1765 -710 2085
rect -740 1735 -710 1765
rect -680 2085 -650 2115
rect -680 1765 -675 2085
rect -655 1765 -650 2085
rect -680 1755 -650 1765
rect -620 2085 -590 2095
rect -620 1765 -615 2085
rect -595 1765 -590 2085
rect -620 1735 -590 1765
rect -560 2085 -530 2115
rect -560 1765 -555 2085
rect -535 1765 -530 2085
rect -560 1755 -530 1765
rect -500 2085 -470 2095
rect -500 1765 -495 2085
rect -475 1765 -470 2085
rect -500 1735 -470 1765
rect -440 2085 -410 2115
rect -440 1765 -435 2085
rect -415 1765 -410 2085
rect -440 1755 -410 1765
rect -270 1735 -250 2115
rect -1105 1730 -1065 1735
rect -1105 1700 -1100 1730
rect -1070 1700 -1065 1730
rect -1105 1695 -1065 1700
rect -985 1730 -945 1735
rect -985 1700 -980 1730
rect -950 1700 -945 1730
rect -985 1695 -945 1700
rect -865 1730 -825 1735
rect -865 1700 -860 1730
rect -830 1700 -825 1730
rect -865 1695 -825 1700
rect -745 1730 -705 1735
rect -745 1700 -740 1730
rect -710 1700 -705 1730
rect -745 1695 -705 1700
rect -625 1730 -585 1735
rect -625 1700 -620 1730
rect -590 1700 -585 1730
rect -625 1695 -585 1700
rect -505 1730 -465 1735
rect -505 1700 -500 1730
rect -470 1700 -465 1730
rect -505 1695 -465 1700
rect -280 1730 -240 1735
rect -280 1700 -275 1730
rect -245 1700 -240 1730
rect -280 1695 -240 1700
rect -370 1670 -330 1675
rect -370 1640 -365 1670
rect -335 1640 -330 1670
rect -370 1635 -330 1640
rect -715 1625 -675 1630
rect -715 1595 -710 1625
rect -680 1595 -675 1625
rect -715 1590 -675 1595
rect -1450 1540 -1410 1545
rect -1450 1510 -1445 1540
rect -1415 1510 -1410 1540
rect -1450 1505 -1410 1510
rect -1440 1430 -1420 1505
rect -1135 1485 -1095 1490
rect -1135 1455 -1130 1485
rect -1100 1455 -1095 1485
rect -1135 1450 -1095 1455
rect -1025 1485 -985 1490
rect -1025 1455 -1020 1485
rect -990 1455 -985 1485
rect -1025 1450 -985 1455
rect -915 1485 -875 1490
rect -915 1455 -910 1485
rect -880 1455 -875 1485
rect -915 1450 -875 1455
rect -805 1485 -765 1490
rect -805 1455 -800 1485
rect -770 1455 -765 1485
rect -805 1450 -765 1455
rect -695 1485 -655 1490
rect -695 1455 -690 1485
rect -660 1455 -655 1485
rect -695 1450 -655 1455
rect -585 1485 -545 1490
rect -585 1455 -580 1485
rect -550 1455 -545 1485
rect -585 1450 -545 1455
rect -475 1485 -435 1490
rect -475 1455 -470 1485
rect -440 1455 -435 1485
rect -475 1450 -435 1455
rect -1501 1420 -1360 1430
rect -1501 1400 -1495 1420
rect -1475 1400 -1440 1420
rect -1420 1400 -1385 1420
rect -1365 1400 -1360 1420
rect -1501 1390 -1360 1400
rect -1130 1420 -1100 1450
rect -1130 850 -1125 1420
rect -1105 850 -1100 1420
rect -1130 840 -1100 850
rect -1075 1420 -1045 1430
rect -1075 850 -1070 1420
rect -1050 850 -1045 1420
rect -1501 815 -1360 825
rect -1075 820 -1045 850
rect -1020 1420 -990 1450
rect -1020 850 -1015 1420
rect -995 850 -990 1420
rect -1020 840 -990 850
rect -965 1420 -935 1430
rect -965 850 -960 1420
rect -940 850 -935 1420
rect -965 820 -935 850
rect -910 1420 -880 1450
rect -910 850 -905 1420
rect -885 850 -880 1420
rect -910 840 -880 850
rect -855 1420 -825 1430
rect -855 850 -850 1420
rect -830 850 -825 1420
rect -855 820 -825 850
rect -800 1420 -770 1450
rect -800 850 -795 1420
rect -775 850 -770 1420
rect -800 840 -770 850
rect -745 1420 -715 1430
rect -745 850 -740 1420
rect -720 850 -715 1420
rect -745 820 -715 850
rect -690 1420 -660 1450
rect -690 850 -685 1420
rect -665 850 -660 1420
rect -690 840 -660 850
rect -635 1420 -605 1430
rect -635 850 -630 1420
rect -610 850 -605 1420
rect -635 820 -605 850
rect -580 1420 -550 1450
rect -580 850 -575 1420
rect -555 850 -550 1420
rect -580 840 -550 850
rect -525 1420 -495 1430
rect -525 850 -520 1420
rect -500 850 -495 1420
rect -525 820 -495 850
rect -470 1420 -440 1450
rect -470 850 -465 1420
rect -445 850 -440 1420
rect -360 905 -340 1635
rect -225 1490 -205 2170
rect -40 2150 0 2155
rect -40 2120 -35 2150
rect -5 2120 0 2150
rect -40 2115 0 2120
rect 80 2150 120 2155
rect 80 2120 85 2150
rect 115 2120 120 2150
rect 80 2115 120 2120
rect 200 2150 240 2155
rect 200 2120 205 2150
rect 235 2120 240 2150
rect 200 2115 240 2120
rect 320 2150 360 2155
rect 320 2120 325 2150
rect 355 2120 360 2150
rect 320 2115 360 2120
rect 440 2150 480 2155
rect 440 2120 445 2150
rect 475 2120 480 2150
rect 440 2115 480 2120
rect 560 2150 600 2155
rect 560 2120 565 2150
rect 595 2120 600 2150
rect 560 2115 600 2120
rect 680 2150 720 2155
rect 680 2120 685 2150
rect 715 2120 720 2150
rect 680 2115 720 2120
rect -35 2085 -5 2095
rect -35 1765 -30 2085
rect -10 1765 -5 2085
rect -35 1755 -5 1765
rect 25 2085 55 2095
rect 25 1765 30 2085
rect 50 1765 55 2085
rect 25 1735 55 1765
rect 85 2085 115 2115
rect 85 1765 90 2085
rect 110 1765 115 2085
rect 85 1755 115 1765
rect 145 2085 175 2095
rect 145 1765 150 2085
rect 170 1765 175 2085
rect 145 1735 175 1765
rect 205 2085 235 2115
rect 205 1765 210 2085
rect 230 1765 235 2085
rect 205 1755 235 1765
rect 265 2085 295 2095
rect 265 1765 270 2085
rect 290 1765 295 2085
rect 265 1735 295 1765
rect 325 2085 355 2115
rect 325 1765 330 2085
rect 350 1765 355 2085
rect 325 1755 355 1765
rect 385 2085 415 2095
rect 385 1765 390 2085
rect 410 1765 415 2085
rect 385 1735 415 1765
rect 445 2085 475 2115
rect 445 1765 450 2085
rect 470 1765 475 2085
rect 445 1755 475 1765
rect 505 2085 535 2095
rect 505 1765 510 2085
rect 530 1765 535 2085
rect 505 1735 535 1765
rect 565 2085 595 2115
rect 565 1765 570 2085
rect 590 1765 595 2085
rect 565 1755 595 1765
rect 625 2085 655 2095
rect 625 1765 630 2085
rect 650 1765 655 2085
rect 625 1735 655 1765
rect 685 2085 715 2095
rect 685 1765 690 2085
rect 710 1765 715 2085
rect 685 1755 715 1765
rect 20 1730 60 1735
rect 20 1700 25 1730
rect 55 1700 60 1730
rect 20 1695 60 1700
rect 140 1730 180 1735
rect 140 1700 145 1730
rect 175 1700 180 1730
rect 140 1695 180 1700
rect 260 1730 300 1735
rect 260 1700 265 1730
rect 295 1700 300 1730
rect 260 1670 300 1700
rect 380 1730 420 1735
rect 380 1700 385 1730
rect 415 1700 420 1730
rect 380 1695 420 1700
rect 500 1730 540 1735
rect 500 1700 505 1730
rect 535 1700 540 1730
rect 500 1695 540 1700
rect 620 1730 660 1735
rect 620 1700 625 1730
rect 655 1700 660 1730
rect 620 1695 660 1700
rect 790 1675 810 2270
rect 835 2210 855 2520
rect 975 2340 980 2660
rect 1000 2340 1005 2660
rect 975 2330 1005 2340
rect 1035 2660 1065 2745
rect 1090 2725 1130 2730
rect 1090 2695 1095 2725
rect 1125 2695 1130 2725
rect 1090 2690 1130 2695
rect 1150 2725 1190 2730
rect 1150 2695 1155 2725
rect 1185 2695 1190 2725
rect 1150 2690 1190 2695
rect 1440 2725 1480 2750
rect 1440 2695 1445 2725
rect 1475 2695 1480 2725
rect 1440 2690 1480 2695
rect 1500 2725 1540 2730
rect 1500 2695 1505 2725
rect 1535 2695 1540 2725
rect 1500 2690 1540 2695
rect 1620 2725 1660 2730
rect 1620 2695 1625 2725
rect 1655 2695 1660 2725
rect 1620 2690 1660 2695
rect 1035 2340 1040 2660
rect 1060 2340 1065 2660
rect 1035 2330 1065 2340
rect 1095 2660 1125 2690
rect 1095 2340 1100 2660
rect 1120 2340 1125 2660
rect 1095 2330 1125 2340
rect 1155 2660 1185 2690
rect 1155 2340 1160 2660
rect 1180 2340 1185 2660
rect 1155 2330 1185 2340
rect 1445 2660 1475 2690
rect 1445 2340 1450 2660
rect 1470 2340 1475 2660
rect 1445 2330 1475 2340
rect 1505 2660 1535 2690
rect 1505 2340 1510 2660
rect 1530 2340 1535 2660
rect 1505 2330 1535 2340
rect 1565 2660 1595 2670
rect 1565 2340 1570 2660
rect 1590 2340 1595 2660
rect 1051 2300 1081 2310
rect 1051 2280 1056 2300
rect 1076 2280 1081 2300
rect 1051 2270 1081 2280
rect 1521 2305 1551 2310
rect 1521 2270 1551 2275
rect 880 2260 920 2265
rect 880 2230 885 2260
rect 915 2230 920 2260
rect 1055 2255 1075 2270
rect 1565 2255 1595 2340
rect 1625 2660 1655 2690
rect 1625 2340 1630 2660
rect 1650 2340 1655 2660
rect 1625 2330 1655 2340
rect 880 2225 920 2230
rect 1045 2250 1085 2255
rect 825 2205 865 2210
rect 825 2175 830 2205
rect 860 2175 865 2205
rect 825 2170 865 2175
rect 260 1640 265 1670
rect 295 1640 300 1670
rect 260 1635 300 1640
rect 410 1670 450 1675
rect 410 1640 415 1670
rect 445 1640 450 1670
rect 410 1635 450 1640
rect 780 1670 820 1675
rect 780 1640 785 1670
rect 815 1640 820 1670
rect 780 1635 820 1640
rect 880 1630 900 2225
rect 1045 2220 1050 2250
rect 1080 2220 1085 2250
rect 1045 2215 1085 2220
rect 1560 2250 1600 2255
rect 1560 2220 1565 2250
rect 1595 2220 1600 2250
rect 1560 2215 1600 2220
rect 1885 2205 1925 2210
rect 1885 2175 1890 2205
rect 1920 2175 1925 2205
rect 1885 2170 1925 2175
rect 2455 2205 2495 2210
rect 2455 2175 2460 2205
rect 2490 2175 2495 2205
rect 2455 2170 2495 2175
rect 970 2150 1010 2155
rect 970 2120 975 2150
rect 1005 2120 1010 2150
rect 970 2115 1010 2120
rect 1090 2150 1130 2155
rect 1090 2120 1095 2150
rect 1125 2120 1130 2150
rect 1090 2115 1130 2120
rect 1210 2150 1250 2155
rect 1210 2120 1215 2150
rect 1245 2120 1250 2150
rect 1210 2115 1250 2120
rect 1330 2150 1370 2155
rect 1330 2120 1335 2150
rect 1365 2120 1370 2150
rect 1330 2115 1370 2120
rect 1450 2150 1490 2155
rect 1450 2120 1455 2150
rect 1485 2120 1490 2150
rect 1450 2115 1490 2120
rect 1570 2150 1610 2155
rect 1570 2120 1575 2150
rect 1605 2120 1610 2150
rect 1570 2115 1610 2120
rect 1690 2150 1730 2155
rect 1690 2120 1695 2150
rect 1725 2120 1730 2150
rect 1690 2115 1730 2120
rect 975 2085 1005 2095
rect 975 1765 980 2085
rect 1000 1765 1005 2085
rect 975 1755 1005 1765
rect 1035 2085 1065 2095
rect 1035 1765 1040 2085
rect 1060 1765 1065 2085
rect 1035 1735 1065 1765
rect 1095 2085 1125 2115
rect 1095 1765 1100 2085
rect 1120 1765 1125 2085
rect 1095 1755 1125 1765
rect 1155 2085 1185 2095
rect 1155 1765 1160 2085
rect 1180 1765 1185 2085
rect 1155 1735 1185 1765
rect 1215 2085 1245 2115
rect 1215 1765 1220 2085
rect 1240 1765 1245 2085
rect 1215 1755 1245 1765
rect 1275 2085 1305 2095
rect 1275 1765 1280 2085
rect 1300 1765 1305 2085
rect 1275 1735 1305 1765
rect 1335 2085 1365 2115
rect 1335 1765 1340 2085
rect 1360 1765 1365 2085
rect 1335 1755 1365 1765
rect 1395 2085 1425 2095
rect 1395 1765 1400 2085
rect 1420 1765 1425 2085
rect 1395 1735 1425 1765
rect 1455 2085 1485 2115
rect 1455 1765 1460 2085
rect 1480 1765 1485 2085
rect 1455 1755 1485 1765
rect 1515 2085 1545 2095
rect 1515 1765 1520 2085
rect 1540 1765 1545 2085
rect 1515 1735 1545 1765
rect 1575 2085 1605 2115
rect 1575 1765 1580 2085
rect 1600 1765 1605 2085
rect 1575 1755 1605 1765
rect 1635 2085 1665 2095
rect 1635 1765 1640 2085
rect 1660 1765 1665 2085
rect 1635 1735 1665 1765
rect 1695 2085 1725 2095
rect 1695 1765 1700 2085
rect 1720 1765 1725 2085
rect 1695 1755 1725 1765
rect 1030 1730 1070 1735
rect 1030 1700 1035 1730
rect 1065 1700 1070 1730
rect 1030 1695 1070 1700
rect 1150 1730 1190 1735
rect 1150 1700 1155 1730
rect 1185 1700 1190 1730
rect 1150 1695 1190 1700
rect 1270 1730 1310 1735
rect 1270 1700 1275 1730
rect 1305 1700 1310 1730
rect 1270 1695 1310 1700
rect 1390 1730 1430 1735
rect 1390 1700 1395 1730
rect 1425 1700 1430 1730
rect 1240 1670 1280 1675
rect 1240 1640 1245 1670
rect 1275 1640 1280 1670
rect 1240 1635 1280 1640
rect 1390 1670 1430 1700
rect 1510 1730 1550 1735
rect 1510 1700 1515 1730
rect 1545 1700 1550 1730
rect 1510 1695 1550 1700
rect 1630 1730 1670 1735
rect 1630 1700 1635 1730
rect 1665 1700 1670 1730
rect 1630 1695 1670 1700
rect 1390 1640 1395 1670
rect 1425 1640 1430 1670
rect 1390 1635 1430 1640
rect 870 1600 875 1630
rect 905 1600 910 1630
rect 1895 1570 1915 2170
rect 2460 2155 2490 2170
rect 1930 2150 1970 2155
rect 1930 2120 1935 2150
rect 1965 2120 1970 2150
rect 1930 2115 1970 2120
rect 2095 2150 2135 2155
rect 2095 2120 2100 2150
rect 2130 2120 2135 2150
rect 2095 2115 2135 2120
rect 2215 2150 2255 2155
rect 2215 2120 2220 2150
rect 2250 2120 2255 2150
rect 2215 2115 2255 2120
rect 2335 2150 2375 2155
rect 2335 2120 2340 2150
rect 2370 2120 2375 2150
rect 2335 2115 2375 2120
rect 2455 2150 2495 2155
rect 2455 2120 2460 2150
rect 2490 2120 2495 2150
rect 2455 2115 2495 2120
rect 2575 2150 2615 2155
rect 2575 2120 2580 2150
rect 2610 2120 2615 2150
rect 2575 2115 2615 2120
rect 2695 2150 2735 2155
rect 2695 2120 2700 2150
rect 2730 2120 2735 2150
rect 2695 2115 2735 2120
rect 2815 2150 2855 2155
rect 2815 2120 2820 2150
rect 2850 2120 2855 2150
rect 2815 2115 2855 2120
rect 1940 1735 1960 2115
rect 2100 2085 2130 2115
rect 2100 1765 2105 2085
rect 2125 1765 2130 2085
rect 2100 1755 2130 1765
rect 2160 2085 2190 2095
rect 2160 1765 2165 2085
rect 2185 1765 2190 2085
rect 2160 1735 2190 1765
rect 2220 2085 2250 2115
rect 2220 1765 2225 2085
rect 2245 1765 2250 2085
rect 2220 1755 2250 1765
rect 2280 2085 2310 2095
rect 2280 1765 2285 2085
rect 2305 1765 2310 2085
rect 2280 1735 2310 1765
rect 2340 2085 2370 2115
rect 2340 1765 2345 2085
rect 2365 1765 2370 2085
rect 2340 1755 2370 1765
rect 2400 2085 2430 2095
rect 2400 1765 2405 2085
rect 2425 1765 2430 2085
rect 2400 1735 2430 1765
rect 2460 2085 2490 2115
rect 2460 1765 2465 2085
rect 2485 1765 2490 2085
rect 2460 1755 2490 1765
rect 2520 2085 2550 2095
rect 2520 1765 2525 2085
rect 2545 1765 2550 2085
rect 2520 1735 2550 1765
rect 2580 2085 2610 2115
rect 2580 1765 2585 2085
rect 2605 1765 2610 2085
rect 2580 1755 2610 1765
rect 2640 2085 2670 2095
rect 2640 1765 2645 2085
rect 2665 1765 2670 2085
rect 2640 1735 2670 1765
rect 2700 2085 2730 2115
rect 2700 1765 2705 2085
rect 2725 1765 2730 2085
rect 2700 1755 2730 1765
rect 2760 2085 2790 2095
rect 2760 1765 2765 2085
rect 2785 1765 2790 2085
rect 2760 1735 2790 1765
rect 2820 2085 2850 2115
rect 2820 1765 2825 2085
rect 2845 1765 2850 2085
rect 2820 1755 2850 1765
rect 1930 1730 1970 1735
rect 1930 1700 1935 1730
rect 1965 1700 1970 1730
rect 1930 1695 1970 1700
rect 2155 1730 2195 1735
rect 2155 1700 2160 1730
rect 2190 1700 2195 1730
rect 2155 1695 2195 1700
rect 2275 1730 2315 1735
rect 2275 1700 2280 1730
rect 2310 1700 2315 1730
rect 2275 1695 2315 1700
rect 2395 1730 2435 1735
rect 2395 1700 2400 1730
rect 2430 1700 2435 1730
rect 2395 1695 2435 1700
rect 2515 1730 2555 1735
rect 2515 1700 2520 1730
rect 2550 1700 2555 1730
rect 2515 1695 2555 1700
rect 2635 1730 2675 1735
rect 2635 1700 2640 1730
rect 2670 1700 2675 1730
rect 2635 1695 2675 1700
rect 2755 1730 2795 1735
rect 2755 1700 2760 1730
rect 2790 1700 2795 1730
rect 2755 1695 2795 1700
rect 2020 1670 2060 1675
rect 2020 1640 2025 1670
rect 2055 1640 2060 1670
rect 2020 1635 2060 1640
rect 455 1565 495 1570
rect 455 1535 460 1565
rect 490 1535 495 1565
rect 455 1530 495 1535
rect 620 1565 660 1570
rect 620 1535 625 1565
rect 655 1535 660 1565
rect 620 1530 660 1535
rect 785 1565 825 1570
rect 785 1535 790 1565
rect 820 1535 825 1565
rect 785 1530 825 1535
rect 865 1565 905 1570
rect 865 1535 870 1565
rect 900 1535 905 1565
rect 865 1530 905 1535
rect 1030 1565 1070 1570
rect 1030 1535 1035 1565
rect 1065 1535 1070 1565
rect 1030 1530 1070 1535
rect 1195 1565 1235 1570
rect 1195 1535 1200 1565
rect 1230 1535 1235 1565
rect 1195 1530 1235 1535
rect 1885 1565 1925 1570
rect 1885 1535 1890 1565
rect 1920 1535 1925 1565
rect 1885 1530 1925 1535
rect -235 1485 -195 1490
rect -235 1455 -230 1485
rect -200 1455 -195 1485
rect -235 1450 -195 1455
rect 460 1470 490 1530
rect 565 1520 605 1525
rect 565 1490 570 1520
rect 600 1490 605 1520
rect 565 1485 605 1490
rect -325 1105 -285 1110
rect -325 1075 -320 1105
rect -290 1075 -285 1105
rect -325 1070 -285 1075
rect -370 900 -330 905
rect -370 870 -365 900
rect -335 870 -330 900
rect -370 865 -330 870
rect -470 840 -440 850
rect -1501 795 -1495 815
rect -1475 795 -1440 815
rect -1420 795 -1385 815
rect -1365 795 -1360 815
rect -1501 785 -1360 795
rect -1080 815 -1040 820
rect -1080 785 -1075 815
rect -1045 785 -1040 815
rect -1540 760 -1500 765
rect -1540 730 -1535 760
rect -1505 730 -1500 760
rect -1540 725 -1500 730
rect -1530 360 -1510 725
rect -1440 720 -1420 785
rect -1080 780 -1040 785
rect -970 815 -930 820
rect -970 785 -965 815
rect -935 785 -930 815
rect -970 780 -930 785
rect -860 815 -820 820
rect -860 785 -855 815
rect -825 785 -820 815
rect -860 780 -820 785
rect -750 815 -710 820
rect -750 785 -745 815
rect -715 785 -710 815
rect -750 780 -710 785
rect -640 815 -600 820
rect -640 785 -635 815
rect -605 785 -600 815
rect -640 780 -600 785
rect -530 815 -490 820
rect -530 785 -525 815
rect -495 785 -490 815
rect -530 780 -490 785
rect -960 765 -940 780
rect -970 760 -930 765
rect -970 730 -965 760
rect -935 730 -930 760
rect -970 725 -930 730
rect -530 760 -490 765
rect -530 730 -525 760
rect -495 730 -490 760
rect -530 725 -490 730
rect -1450 715 -1410 720
rect -1450 685 -1445 715
rect -1415 685 -1410 715
rect -1450 680 -1410 685
rect -805 715 -765 720
rect -805 685 -800 715
rect -770 685 -765 715
rect -805 680 -765 685
rect -520 675 -500 725
rect -360 720 -340 865
rect -370 715 -330 720
rect -370 685 -365 715
rect -335 685 -330 715
rect -370 680 -330 685
rect -1135 670 -1095 675
rect -1135 640 -1130 670
rect -1100 640 -1095 670
rect -1135 635 -1095 640
rect -1080 670 -1040 675
rect -1080 640 -1075 670
rect -1045 640 -1040 670
rect -1080 635 -1040 640
rect -970 670 -930 675
rect -970 640 -965 670
rect -935 640 -930 670
rect -970 635 -930 640
rect -860 670 -820 675
rect -860 640 -855 670
rect -825 640 -820 670
rect -860 635 -820 640
rect -750 670 -710 675
rect -750 640 -745 670
rect -715 640 -710 670
rect -750 635 -710 640
rect -640 670 -600 675
rect -640 640 -635 670
rect -605 640 -600 670
rect -640 635 -600 640
rect -530 670 -490 675
rect -530 640 -525 670
rect -495 640 -490 670
rect -530 635 -490 640
rect -475 670 -435 675
rect -475 640 -470 670
rect -440 640 -435 670
rect -475 635 -435 640
rect -1130 605 -1100 635
rect -1130 435 -1125 605
rect -1105 435 -1100 605
rect -1130 425 -1100 435
rect -1075 605 -1045 635
rect -1075 435 -1070 605
rect -1050 435 -1045 605
rect -1075 425 -1045 435
rect -1020 605 -990 615
rect -1020 435 -1015 605
rect -995 435 -990 605
rect -1020 420 -990 435
rect -965 605 -935 635
rect -965 435 -960 605
rect -940 435 -935 605
rect -965 425 -935 435
rect -910 605 -880 615
rect -910 435 -905 605
rect -885 435 -880 605
rect -910 420 -880 435
rect -855 605 -825 635
rect -855 435 -850 605
rect -830 435 -825 605
rect -855 425 -825 435
rect -800 605 -770 615
rect -800 435 -795 605
rect -775 435 -770 605
rect -800 420 -770 435
rect -745 605 -715 635
rect -745 435 -740 605
rect -720 435 -715 605
rect -745 425 -715 435
rect -690 605 -660 615
rect -690 435 -685 605
rect -665 435 -660 605
rect -690 420 -660 435
rect -635 605 -605 635
rect -635 435 -630 605
rect -610 435 -605 605
rect -635 425 -605 435
rect -580 605 -550 615
rect -580 435 -575 605
rect -555 435 -550 605
rect -580 420 -550 435
rect -525 605 -495 635
rect -525 435 -520 605
rect -500 435 -495 605
rect -525 425 -495 435
rect -470 605 -440 635
rect -470 435 -465 605
rect -445 435 -440 605
rect -470 425 -440 435
rect -1270 415 -1230 420
rect -1270 385 -1265 415
rect -1235 385 -1230 415
rect -1270 380 -1230 385
rect -1025 415 -985 420
rect -1025 385 -1020 415
rect -990 385 -985 415
rect -1025 380 -985 385
rect -915 415 -875 420
rect -915 385 -910 415
rect -880 385 -875 415
rect -915 380 -875 385
rect -805 415 -765 420
rect -805 385 -800 415
rect -770 385 -765 415
rect -805 380 -765 385
rect -695 415 -655 420
rect -695 385 -690 415
rect -660 385 -655 415
rect -695 380 -655 385
rect -585 415 -545 420
rect -585 385 -580 415
rect -550 385 -545 415
rect -585 380 -545 385
rect -1545 350 -1495 360
rect -1545 320 -1535 350
rect -1505 320 -1495 350
rect -1545 310 -1495 320
rect -1530 -300 -1510 310
rect -1490 -120 -1486 -85
rect -1459 -120 -1455 -85
rect -1430 -120 -1426 -85
rect -1399 -120 -1395 -85
rect -1370 -120 -1366 -85
rect -1339 -120 -1335 -85
rect -1310 -120 -1306 -85
rect -1279 -120 -1275 -85
rect -1485 -185 -1460 -120
rect -1370 -145 -1335 -120
rect -1260 -140 -1240 380
rect -360 345 -340 680
rect -750 340 -710 345
rect -750 310 -745 340
rect -715 310 -710 340
rect -750 305 -710 310
rect -370 340 -330 345
rect -370 310 -365 340
rect -335 310 -330 340
rect -370 305 -330 310
rect -1225 265 -1185 270
rect -1225 235 -1220 265
rect -1190 235 -1185 265
rect -1225 230 -1185 235
rect -1025 265 -985 270
rect -1025 235 -1020 265
rect -990 235 -985 265
rect -1025 230 -985 235
rect -915 265 -875 270
rect -915 235 -910 265
rect -880 235 -875 265
rect -915 230 -875 235
rect -805 265 -765 270
rect -805 235 -800 265
rect -770 235 -765 265
rect -805 230 -765 235
rect -695 265 -655 270
rect -695 235 -690 265
rect -660 235 -655 265
rect -695 230 -655 235
rect -585 265 -545 270
rect -585 235 -580 265
rect -550 235 -545 265
rect -585 230 -545 235
rect -1215 -85 -1195 230
rect -1130 215 -1100 225
rect -1130 -55 -1125 215
rect -1105 -55 -1100 215
rect -1130 -85 -1100 -55
rect -1075 215 -1045 225
rect -1075 -55 -1070 215
rect -1050 -55 -1045 215
rect -1075 -85 -1045 -55
rect -1020 215 -990 230
rect -1020 -55 -1015 215
rect -995 -55 -990 215
rect -1020 -65 -990 -55
rect -965 215 -935 225
rect -965 -55 -960 215
rect -940 -55 -935 215
rect -965 -85 -935 -55
rect -910 215 -880 230
rect -910 -55 -905 215
rect -885 -55 -880 215
rect -910 -65 -880 -55
rect -855 215 -825 225
rect -855 -55 -850 215
rect -830 -55 -825 215
rect -855 -85 -825 -55
rect -800 215 -770 230
rect -800 -55 -795 215
rect -775 -55 -770 215
rect -800 -65 -770 -55
rect -745 215 -715 225
rect -745 -55 -740 215
rect -720 -55 -715 215
rect -745 -85 -715 -55
rect -690 215 -660 230
rect -690 -55 -685 215
rect -665 -55 -660 215
rect -690 -65 -660 -55
rect -635 215 -605 225
rect -635 -55 -630 215
rect -610 -55 -605 215
rect -635 -85 -605 -55
rect -580 215 -550 230
rect -580 -55 -575 215
rect -555 -55 -550 215
rect -580 -65 -550 -55
rect -525 215 -495 225
rect -525 -55 -520 215
rect -500 -55 -495 215
rect -525 -85 -495 -55
rect -470 215 -440 225
rect -470 -55 -465 215
rect -445 -55 -440 215
rect -470 -85 -440 -55
rect -1225 -90 -1185 -85
rect -1225 -120 -1220 -90
rect -1190 -120 -1185 -90
rect -1225 -125 -1185 -120
rect -1135 -90 -1095 -85
rect -1135 -120 -1130 -90
rect -1100 -120 -1095 -90
rect -1370 -180 -1335 -175
rect -1270 -145 -1230 -140
rect -1270 -175 -1265 -145
rect -1235 -175 -1230 -145
rect -1270 -180 -1230 -175
rect -1135 -145 -1095 -120
rect -1080 -90 -1040 -85
rect -1080 -120 -1075 -90
rect -1045 -120 -1040 -90
rect -1080 -125 -1040 -120
rect -970 -90 -930 -85
rect -970 -120 -965 -90
rect -935 -120 -930 -90
rect -970 -125 -930 -120
rect -860 -90 -820 -85
rect -860 -120 -855 -90
rect -825 -120 -820 -90
rect -860 -125 -820 -120
rect -750 -90 -710 -85
rect -750 -120 -745 -90
rect -715 -120 -710 -90
rect -750 -125 -710 -120
rect -640 -90 -600 -85
rect -640 -120 -635 -90
rect -605 -120 -600 -90
rect -640 -125 -600 -120
rect -530 -90 -490 -85
rect -530 -120 -525 -90
rect -495 -120 -490 -90
rect -530 -125 -490 -120
rect -475 -95 -435 -85
rect -475 -115 -465 -95
rect -445 -115 -435 -95
rect -1135 -175 -1130 -145
rect -1100 -175 -1095 -145
rect -1135 -180 -1095 -175
rect -475 -145 -435 -115
rect -475 -175 -470 -145
rect -440 -175 -435 -145
rect -475 -180 -435 -175
rect -1490 -190 -1455 -185
rect -315 -190 -295 1070
rect -280 770 -240 775
rect -280 740 -275 770
rect -245 740 -240 770
rect -280 735 -240 740
rect -270 -140 -250 735
rect -225 675 -205 1450
rect 460 1250 465 1470
rect 485 1250 490 1470
rect 460 1240 490 1250
rect 515 1470 545 1480
rect 515 1250 520 1470
rect 540 1250 545 1470
rect 515 1240 545 1250
rect 570 1470 600 1485
rect 570 1250 575 1470
rect 595 1250 600 1470
rect 570 1240 600 1250
rect 625 1470 655 1530
rect 675 1520 715 1525
rect 675 1490 680 1520
rect 710 1490 715 1520
rect 675 1485 715 1490
rect 625 1250 630 1470
rect 650 1250 655 1470
rect 625 1240 655 1250
rect 680 1470 710 1485
rect 680 1250 685 1470
rect 705 1250 710 1470
rect 680 1240 710 1250
rect 735 1470 765 1480
rect 735 1250 740 1470
rect 760 1250 765 1470
rect 735 1240 765 1250
rect 790 1470 820 1530
rect 790 1250 795 1470
rect 815 1250 820 1470
rect 790 1240 820 1250
rect 870 1470 900 1530
rect 975 1520 1015 1525
rect 975 1490 980 1520
rect 1010 1490 1015 1520
rect 975 1485 1015 1490
rect 870 1250 875 1470
rect 895 1250 900 1470
rect 870 1240 900 1250
rect 925 1470 955 1480
rect 925 1250 930 1470
rect 950 1250 955 1470
rect 925 1240 955 1250
rect 980 1470 1010 1485
rect 980 1250 985 1470
rect 1005 1250 1010 1470
rect 980 1240 1010 1250
rect 1035 1470 1065 1530
rect 1085 1520 1125 1525
rect 1085 1490 1090 1520
rect 1120 1490 1125 1520
rect 1085 1485 1125 1490
rect 1035 1250 1040 1470
rect 1060 1250 1065 1470
rect 1035 1240 1065 1250
rect 1090 1470 1120 1485
rect 1090 1250 1095 1470
rect 1115 1250 1120 1470
rect 1090 1240 1120 1250
rect 1145 1470 1175 1480
rect 1145 1250 1150 1470
rect 1170 1250 1175 1470
rect 1145 1240 1175 1250
rect 1200 1470 1230 1530
rect 1895 1490 1915 1530
rect 1200 1250 1205 1470
rect 1225 1250 1230 1470
rect 1885 1485 1925 1490
rect 1885 1455 1890 1485
rect 1920 1455 1925 1485
rect 1885 1450 1925 1455
rect 1200 1240 1230 1250
rect 515 1210 535 1240
rect 495 1205 535 1210
rect 495 1175 500 1205
rect 530 1175 535 1205
rect 550 1210 580 1220
rect 550 1190 555 1210
rect 575 1190 580 1210
rect 550 1180 580 1190
rect 620 1215 660 1220
rect 620 1185 625 1215
rect 655 1185 660 1215
rect 620 1180 660 1185
rect 700 1210 730 1220
rect 700 1190 705 1210
rect 725 1190 730 1210
rect 700 1180 730 1190
rect 745 1210 765 1240
rect 745 1205 785 1210
rect 495 1170 535 1175
rect 555 1160 575 1180
rect 545 1155 585 1160
rect 545 1125 550 1155
rect 580 1125 585 1155
rect 545 1120 585 1125
rect 705 1110 725 1180
rect 745 1175 750 1205
rect 780 1175 785 1205
rect 745 1170 785 1175
rect 690 1105 730 1110
rect 690 1075 695 1105
rect 725 1075 730 1105
rect 690 1070 730 1075
rect 925 1065 945 1240
rect 960 1210 990 1220
rect 960 1190 965 1210
rect 985 1190 990 1210
rect 960 1180 990 1190
rect 1030 1215 1070 1220
rect 1030 1185 1035 1215
rect 1065 1185 1070 1215
rect 1030 1180 1070 1185
rect 1110 1210 1140 1220
rect 1110 1190 1115 1210
rect 1135 1190 1140 1210
rect 1110 1180 1140 1190
rect 965 1110 985 1180
rect 1115 1160 1135 1180
rect 1095 1155 1135 1160
rect 1095 1125 1100 1155
rect 1130 1125 1135 1155
rect 1095 1120 1135 1125
rect 965 1105 1005 1110
rect 965 1075 970 1105
rect 1000 1075 1005 1105
rect 965 1070 1005 1075
rect 795 1060 835 1065
rect 795 1030 800 1060
rect 830 1030 835 1060
rect 795 1025 835 1030
rect 905 1060 945 1065
rect 905 1030 910 1060
rect 940 1030 945 1060
rect 905 1025 945 1030
rect 805 1010 825 1025
rect 1155 1015 1175 1240
rect 1155 1010 1195 1015
rect 795 1005 835 1010
rect 795 975 800 1005
rect 830 975 835 1005
rect 795 970 835 975
rect 880 1005 920 1010
rect 880 975 885 1005
rect 915 975 920 1005
rect 1155 980 1160 1010
rect 1190 980 1195 1010
rect 1155 975 1195 980
rect 1840 1010 1880 1015
rect 1840 980 1845 1010
rect 1875 980 1880 1010
rect 1840 975 1880 980
rect 880 970 920 975
rect -190 950 -150 955
rect -190 920 -185 950
rect -155 920 -150 950
rect -190 915 -150 920
rect 120 950 150 955
rect 805 930 825 970
rect 890 930 910 970
rect 1540 950 1570 955
rect 120 915 150 920
rect 775 920 835 930
rect -235 670 -195 675
rect -235 640 -230 670
rect -200 640 -195 670
rect -235 635 -195 640
rect -225 -85 -205 635
rect -235 -90 -195 -85
rect -235 -120 -230 -90
rect -200 -120 -195 -90
rect -235 -125 -195 -120
rect -280 -145 -240 -140
rect -280 -175 -275 -145
rect -245 -175 -240 -145
rect -1490 -225 -1455 -220
rect -325 -220 -320 -190
rect -290 -220 -285 -190
rect -325 -225 -285 -220
rect -1290 -245 -1255 -240
rect -1290 -280 -1255 -275
rect -805 -245 -765 -240
rect -805 -275 -800 -245
rect -770 -275 -765 -245
rect -805 -280 -765 -275
rect -1540 -305 -1500 -300
rect -1540 -335 -1535 -305
rect -1505 -335 -1500 -305
rect -1540 -340 -1500 -335
rect -1285 -380 -1260 -280
rect -1230 -305 -1195 -300
rect -1230 -340 -1195 -335
rect -1005 -305 -965 -300
rect -1005 -335 -1000 -305
rect -970 -335 -965 -305
rect -1005 -340 -965 -335
rect -805 -305 -765 -300
rect -805 -335 -800 -305
rect -770 -335 -765 -305
rect -805 -340 -765 -335
rect -605 -305 -565 -300
rect -605 -335 -600 -305
rect -570 -335 -565 -305
rect -605 -340 -565 -335
rect -1225 -380 -1200 -340
rect -1100 -370 -1070 -360
rect -1290 -415 -1286 -380
rect -1259 -415 -1255 -380
rect -1230 -415 -1226 -380
rect -1199 -415 -1195 -380
rect -1100 -1040 -1095 -370
rect -1075 -1040 -1070 -370
rect -1100 -1070 -1070 -1040
rect -1000 -370 -970 -340
rect -1000 -1040 -995 -370
rect -975 -1040 -970 -370
rect -1000 -1050 -970 -1040
rect -900 -370 -870 -360
rect -900 -1040 -895 -370
rect -875 -1040 -870 -370
rect -900 -1070 -870 -1040
rect -800 -370 -770 -340
rect -800 -1040 -795 -370
rect -775 -1040 -770 -370
rect -800 -1050 -770 -1040
rect -700 -370 -670 -360
rect -700 -1040 -695 -370
rect -675 -1040 -670 -370
rect -700 -1070 -670 -1040
rect -600 -370 -570 -340
rect -600 -1040 -595 -370
rect -575 -1040 -570 -370
rect -600 -1050 -570 -1040
rect -500 -370 -470 -360
rect -500 -1040 -495 -370
rect -475 -1040 -470 -370
rect -500 -1070 -470 -1040
rect -1105 -1075 -1065 -1070
rect -1105 -1105 -1100 -1075
rect -1070 -1105 -1065 -1075
rect -1105 -1110 -1065 -1105
rect -905 -1075 -865 -1070
rect -905 -1105 -900 -1075
rect -870 -1105 -865 -1075
rect -905 -1110 -865 -1105
rect -705 -1075 -665 -1070
rect -705 -1105 -700 -1075
rect -670 -1105 -665 -1075
rect -705 -1110 -665 -1105
rect -505 -1075 -465 -1070
rect -505 -1105 -500 -1075
rect -470 -1105 -465 -1075
rect -505 -1110 -465 -1105
rect -695 -1250 -675 -1110
rect -270 -1250 -250 -175
rect -235 -245 -195 -240
rect -235 -275 -230 -245
rect -200 -275 -195 -245
rect -235 -280 -195 -275
rect -225 -375 -205 -280
rect -235 -380 -195 -375
rect -235 -410 -230 -380
rect -200 -410 -195 -380
rect -235 -415 -195 -410
rect -180 -955 -160 915
rect -50 900 -10 905
rect -50 870 -45 900
rect -15 870 -10 900
rect -50 865 -10 870
rect 60 900 100 905
rect 60 870 65 900
rect 95 870 100 900
rect 60 865 100 870
rect 170 900 210 905
rect 170 870 175 900
rect 205 870 210 900
rect 170 865 210 870
rect 280 900 320 905
rect 280 870 285 900
rect 315 870 320 900
rect 280 865 320 870
rect 390 900 430 905
rect 390 870 395 900
rect 425 870 430 900
rect 390 865 430 870
rect 500 900 540 905
rect 500 870 505 900
rect 535 870 540 900
rect 775 900 805 920
rect 825 900 835 920
rect 775 890 835 900
rect 880 920 920 930
rect 880 900 890 920
rect 910 900 920 920
rect 1540 915 1570 920
rect 880 890 920 900
rect 1150 900 1190 905
rect 500 865 540 870
rect -100 835 -70 845
rect -100 715 -95 835
rect -75 715 -70 835
rect -100 675 -70 715
rect -100 655 -95 675
rect -75 655 -70 675
rect -100 610 -70 655
rect -45 835 -15 865
rect -45 715 -40 835
rect -20 715 -15 835
rect -45 640 -15 715
rect 10 835 40 845
rect 10 715 15 835
rect 35 715 40 835
rect 10 685 40 715
rect 65 835 95 865
rect 65 715 70 835
rect 90 715 95 835
rect 5 655 10 685
rect 40 655 45 685
rect 65 640 95 715
rect 120 835 150 845
rect 120 715 125 835
rect 145 715 150 835
rect 120 685 150 715
rect 175 835 205 865
rect 175 715 180 835
rect 200 715 205 835
rect 115 655 120 685
rect 150 655 155 685
rect 175 640 205 715
rect 230 835 260 845
rect 230 715 235 835
rect 255 715 260 835
rect 230 685 260 715
rect 285 835 315 865
rect 285 715 290 835
rect 310 715 315 835
rect 225 655 230 685
rect 260 655 265 685
rect -50 610 -45 640
rect -15 610 -10 640
rect 60 610 65 640
rect 95 610 100 640
rect 170 610 175 640
rect 205 610 210 640
rect -105 605 -65 610
rect -105 575 -100 605
rect -70 575 -65 605
rect -105 570 -65 575
rect 145 550 175 555
rect 145 515 175 520
rect 230 475 260 655
rect 285 640 315 715
rect 340 835 370 845
rect 340 715 345 835
rect 365 715 370 835
rect 340 685 370 715
rect 395 835 425 865
rect 395 715 400 835
rect 420 715 425 835
rect 335 655 340 685
rect 370 655 375 685
rect 395 640 425 715
rect 450 835 480 845
rect 450 715 455 835
rect 475 715 480 835
rect 450 685 480 715
rect 505 835 535 865
rect 720 860 750 870
rect 505 715 510 835
rect 530 715 535 835
rect 445 655 450 685
rect 480 655 485 685
rect 505 640 535 715
rect 560 835 590 845
rect 560 715 565 835
rect 585 715 590 835
rect 560 675 590 715
rect 560 655 565 675
rect 585 655 590 675
rect 280 610 285 640
rect 315 610 320 640
rect 390 610 395 640
rect 425 610 430 640
rect 500 610 505 640
rect 535 610 540 640
rect 560 610 590 655
rect 720 640 725 860
rect 745 640 750 860
rect 720 610 750 640
rect 775 860 805 890
rect 775 640 780 860
rect 800 640 805 860
rect 775 630 805 640
rect 830 860 860 870
rect 830 640 835 860
rect 855 640 860 860
rect 830 610 860 640
rect 885 860 915 890
rect 1150 870 1155 900
rect 1185 870 1190 900
rect 885 640 890 860
rect 910 640 915 860
rect 885 630 915 640
rect 940 860 970 870
rect 1150 865 1190 870
rect 1260 900 1300 905
rect 1260 870 1265 900
rect 1295 870 1300 900
rect 1260 865 1300 870
rect 1370 900 1410 905
rect 1370 870 1375 900
rect 1405 870 1410 900
rect 1370 865 1410 870
rect 1480 900 1520 905
rect 1480 870 1485 900
rect 1515 870 1520 900
rect 1480 865 1520 870
rect 1590 900 1630 905
rect 1590 870 1595 900
rect 1625 870 1630 900
rect 1590 865 1630 870
rect 1700 900 1740 905
rect 1700 870 1705 900
rect 1735 870 1740 900
rect 1700 865 1740 870
rect 940 640 945 860
rect 965 640 970 860
rect 940 610 970 640
rect 1100 835 1130 845
rect 1100 715 1105 835
rect 1125 715 1130 835
rect 1100 675 1130 715
rect 1100 655 1105 675
rect 1125 655 1130 675
rect 1100 610 1130 655
rect 1155 835 1185 865
rect 1155 715 1160 835
rect 1180 715 1185 835
rect 1155 640 1185 715
rect 1210 835 1240 845
rect 1210 715 1215 835
rect 1235 715 1240 835
rect 1210 685 1240 715
rect 1265 835 1295 865
rect 1265 715 1270 835
rect 1290 715 1295 835
rect 1205 655 1210 685
rect 1240 655 1245 685
rect 1265 640 1295 715
rect 1320 835 1350 845
rect 1320 715 1325 835
rect 1345 715 1350 835
rect 1320 685 1350 715
rect 1375 835 1405 865
rect 1375 715 1380 835
rect 1400 715 1405 835
rect 1315 655 1320 685
rect 1350 655 1355 685
rect 1375 640 1405 715
rect 1430 835 1460 845
rect 1430 715 1435 835
rect 1455 715 1460 835
rect 1430 685 1460 715
rect 1485 835 1515 865
rect 1485 715 1490 835
rect 1510 715 1515 835
rect 1425 655 1430 685
rect 1460 655 1465 685
rect 1150 610 1155 640
rect 1185 610 1190 640
rect 1260 610 1265 640
rect 1295 610 1300 640
rect 1370 610 1375 640
rect 1405 610 1410 640
rect 555 605 595 610
rect 555 575 560 605
rect 590 575 595 605
rect 555 570 595 575
rect 715 605 755 610
rect 715 575 720 605
rect 750 575 755 605
rect 715 570 755 575
rect 825 605 865 610
rect 825 575 830 605
rect 860 575 865 605
rect 825 570 865 575
rect 935 605 975 610
rect 935 575 940 605
rect 970 575 975 605
rect 935 570 975 575
rect 1095 605 1135 610
rect 1095 575 1100 605
rect 1130 575 1135 605
rect 1095 570 1135 575
rect 725 485 745 570
rect 795 550 825 555
rect 795 515 825 520
rect 865 550 895 555
rect 865 515 895 520
rect 945 485 965 570
rect -50 465 -10 470
rect -50 435 -45 465
rect -15 435 -10 465
rect -50 430 -10 435
rect 60 465 100 470
rect 60 435 65 465
rect 95 435 100 465
rect 60 430 100 435
rect 170 465 210 470
rect 170 435 175 465
rect 205 435 210 465
rect 715 475 755 485
rect 230 440 260 445
rect 280 465 320 470
rect 170 430 210 435
rect 280 435 285 465
rect 315 435 320 465
rect 280 430 320 435
rect 390 465 430 470
rect 390 435 395 465
rect 425 435 430 465
rect 390 430 430 435
rect 500 465 540 470
rect 500 435 505 465
rect 535 435 540 465
rect 715 455 725 475
rect 745 455 755 475
rect 715 445 755 455
rect 935 475 975 485
rect 935 455 945 475
rect 965 455 975 475
rect 1430 475 1460 655
rect 1485 640 1515 715
rect 1540 835 1570 845
rect 1540 715 1545 835
rect 1565 715 1570 835
rect 1540 685 1570 715
rect 1595 835 1625 865
rect 1595 715 1600 835
rect 1620 715 1625 835
rect 1535 655 1540 685
rect 1570 655 1575 685
rect 1595 640 1625 715
rect 1650 835 1680 845
rect 1650 715 1655 835
rect 1675 715 1680 835
rect 1650 685 1680 715
rect 1705 835 1735 865
rect 1705 715 1710 835
rect 1730 715 1735 835
rect 1645 655 1650 685
rect 1680 655 1685 685
rect 1705 640 1735 715
rect 1760 835 1790 845
rect 1760 715 1765 835
rect 1785 715 1790 835
rect 1760 675 1790 715
rect 1760 655 1765 675
rect 1785 655 1790 675
rect 1480 610 1485 640
rect 1515 610 1520 640
rect 1590 610 1595 640
rect 1625 610 1630 640
rect 1700 610 1705 640
rect 1735 610 1740 640
rect 1760 610 1790 655
rect 1755 605 1795 610
rect 1755 575 1760 605
rect 1790 575 1795 605
rect 1755 570 1795 575
rect 1515 550 1545 555
rect 1515 515 1545 520
rect 935 445 975 455
rect 1150 465 1190 470
rect 500 430 540 435
rect -100 415 -70 425
rect -100 295 -95 415
rect -75 295 -70 415
rect -100 255 -70 295
rect -100 235 -95 255
rect -75 235 -70 255
rect -45 415 -15 430
rect -45 295 -40 415
rect -20 295 -15 415
rect -45 235 -15 295
rect 10 415 40 425
rect 10 295 15 415
rect 35 295 40 415
rect 10 280 40 295
rect 65 415 95 430
rect 65 295 70 415
rect 90 295 95 415
rect 5 275 45 280
rect 5 245 10 275
rect 40 245 45 275
rect 5 240 45 245
rect 65 235 95 295
rect 120 415 150 425
rect 120 295 125 415
rect 145 295 150 415
rect 120 280 150 295
rect 175 415 205 430
rect 175 295 180 415
rect 200 295 205 415
rect 115 275 155 280
rect 115 245 120 275
rect 150 245 155 275
rect 115 240 155 245
rect 175 235 205 295
rect 230 415 260 425
rect 230 295 235 415
rect 255 295 260 415
rect 230 280 260 295
rect 285 415 315 430
rect 285 295 290 415
rect 310 295 315 415
rect 225 275 265 280
rect 225 245 230 275
rect 260 245 265 275
rect 225 240 265 245
rect 285 235 315 295
rect 340 415 370 425
rect 340 295 345 415
rect 365 295 370 415
rect 340 280 370 295
rect 395 415 425 430
rect 395 295 400 415
rect 420 295 425 415
rect 335 275 375 280
rect 335 245 340 275
rect 370 245 375 275
rect 335 240 375 245
rect 395 235 425 295
rect 450 415 480 425
rect 450 295 455 415
rect 475 295 480 415
rect 450 280 480 295
rect 505 415 535 430
rect 505 295 510 415
rect 530 295 535 415
rect 445 275 485 280
rect 445 245 450 275
rect 480 245 485 275
rect 445 240 485 245
rect 505 235 535 295
rect 560 415 590 425
rect 560 295 565 415
rect 585 295 590 415
rect 560 255 590 295
rect 720 415 750 445
rect 720 295 725 415
rect 745 295 750 415
rect 720 285 750 295
rect 775 415 805 425
rect 775 295 780 415
rect 800 295 805 415
rect 560 235 565 255
rect 585 235 590 255
rect -100 225 -70 235
rect -50 230 -10 235
rect -95 -330 -75 225
rect -50 200 -45 230
rect -15 200 -10 230
rect -50 195 -10 200
rect 60 230 100 235
rect 60 200 65 230
rect 95 200 100 230
rect 60 195 100 200
rect 170 230 210 235
rect 170 200 175 230
rect 205 200 210 230
rect 170 195 210 200
rect 280 230 320 235
rect 280 200 285 230
rect 315 200 320 230
rect 280 195 320 200
rect 390 230 430 235
rect 390 200 395 230
rect 425 200 430 230
rect 390 195 430 200
rect 500 230 540 235
rect 500 200 505 230
rect 535 200 540 230
rect 560 225 590 235
rect 500 195 540 200
rect 440 -10 480 -5
rect 440 -40 445 -10
rect 475 -40 480 -10
rect 440 -45 480 -40
rect -105 -335 -65 -330
rect -105 -365 -100 -335
rect -70 -365 -65 -335
rect -105 -370 -65 -365
rect 450 -430 470 -45
rect 565 -330 585 225
rect 775 210 805 295
rect 830 415 860 425
rect 830 295 835 415
rect 855 295 860 415
rect 770 205 810 210
rect 770 175 775 205
rect 805 175 810 205
rect 770 170 810 175
rect 775 100 805 170
rect 830 150 860 295
rect 885 415 915 425
rect 885 295 890 415
rect 910 295 915 415
rect 885 210 915 295
rect 940 415 970 445
rect 1150 435 1155 465
rect 1185 435 1190 465
rect 1150 430 1190 435
rect 1260 465 1300 470
rect 1260 435 1265 465
rect 1295 435 1300 465
rect 1260 430 1300 435
rect 1370 465 1410 470
rect 1370 435 1375 465
rect 1405 435 1410 465
rect 1430 440 1460 445
rect 1480 465 1520 470
rect 1370 430 1410 435
rect 1480 435 1485 465
rect 1515 435 1520 465
rect 1480 430 1520 435
rect 1590 465 1630 470
rect 1590 435 1595 465
rect 1625 435 1630 465
rect 1590 430 1630 435
rect 1700 465 1740 470
rect 1700 435 1705 465
rect 1735 435 1740 465
rect 1700 430 1740 435
rect 940 295 945 415
rect 965 295 970 415
rect 940 285 970 295
rect 1100 415 1130 425
rect 1100 295 1105 415
rect 1125 295 1130 415
rect 1100 255 1130 295
rect 1100 235 1105 255
rect 1125 235 1130 255
rect 1155 415 1185 430
rect 1155 295 1160 415
rect 1180 295 1185 415
rect 1155 235 1185 295
rect 1210 415 1240 425
rect 1210 295 1215 415
rect 1235 295 1240 415
rect 1210 280 1240 295
rect 1265 415 1295 430
rect 1265 295 1270 415
rect 1290 295 1295 415
rect 1205 275 1245 280
rect 1205 245 1210 275
rect 1240 245 1245 275
rect 1205 240 1245 245
rect 1265 235 1295 295
rect 1320 415 1350 425
rect 1320 295 1325 415
rect 1345 295 1350 415
rect 1320 280 1350 295
rect 1375 415 1405 430
rect 1375 295 1380 415
rect 1400 295 1405 415
rect 1315 275 1355 280
rect 1315 245 1320 275
rect 1350 245 1355 275
rect 1315 240 1355 245
rect 1375 235 1405 295
rect 1430 415 1460 425
rect 1430 295 1435 415
rect 1455 295 1460 415
rect 1430 280 1460 295
rect 1485 415 1515 430
rect 1485 295 1490 415
rect 1510 295 1515 415
rect 1425 275 1465 280
rect 1425 245 1430 275
rect 1460 245 1465 275
rect 1425 240 1465 245
rect 1485 235 1515 295
rect 1540 415 1570 425
rect 1540 295 1545 415
rect 1565 295 1570 415
rect 1540 280 1570 295
rect 1595 415 1625 430
rect 1595 295 1600 415
rect 1620 295 1625 415
rect 1535 275 1575 280
rect 1535 245 1540 275
rect 1570 245 1575 275
rect 1535 240 1575 245
rect 1595 235 1625 295
rect 1650 415 1680 425
rect 1650 295 1655 415
rect 1675 295 1680 415
rect 1650 280 1680 295
rect 1705 415 1735 430
rect 1705 295 1710 415
rect 1730 295 1735 415
rect 1645 275 1685 280
rect 1645 245 1650 275
rect 1680 245 1685 275
rect 1645 240 1685 245
rect 1705 235 1735 295
rect 1760 415 1790 425
rect 1760 295 1765 415
rect 1785 295 1790 415
rect 1760 255 1790 295
rect 1760 235 1765 255
rect 1785 235 1790 255
rect 1100 225 1130 235
rect 1150 230 1190 235
rect 880 205 920 210
rect 880 175 885 205
rect 915 175 920 205
rect 880 170 920 175
rect 830 115 860 120
rect 880 150 920 155
rect 880 120 885 150
rect 915 120 920 150
rect 880 115 920 120
rect 770 95 810 100
rect 770 65 775 95
rect 805 65 810 95
rect 770 60 810 65
rect 830 95 860 100
rect 830 60 860 65
rect 770 40 810 45
rect 770 10 775 40
rect 805 10 810 40
rect 770 5 810 10
rect 720 -80 750 -70
rect 720 -300 725 -80
rect 745 -300 750 -80
rect 720 -330 750 -300
rect 775 -80 805 5
rect 835 -5 855 60
rect 890 45 910 115
rect 880 40 920 45
rect 880 10 885 40
rect 915 10 920 40
rect 880 5 920 10
rect 830 -10 860 -5
rect 830 -45 860 -40
rect 775 -300 780 -80
rect 800 -300 805 -80
rect 775 -310 805 -300
rect 830 -80 860 -70
rect 830 -300 835 -80
rect 855 -300 860 -80
rect 830 -330 860 -300
rect 885 -80 915 5
rect 885 -300 890 -80
rect 910 -300 915 -80
rect 885 -310 915 -300
rect 940 -80 970 -70
rect 940 -300 945 -80
rect 965 -300 970 -80
rect 940 -330 970 -300
rect 1105 -330 1125 225
rect 1150 200 1155 230
rect 1185 200 1190 230
rect 1150 195 1190 200
rect 1260 230 1300 235
rect 1260 200 1265 230
rect 1295 200 1300 230
rect 1260 195 1300 200
rect 1370 230 1410 235
rect 1370 200 1375 230
rect 1405 200 1410 230
rect 1370 195 1410 200
rect 1480 230 1520 235
rect 1480 200 1485 230
rect 1515 200 1520 230
rect 1480 195 1520 200
rect 1590 230 1630 235
rect 1590 200 1595 230
rect 1625 200 1630 230
rect 1590 195 1630 200
rect 1700 230 1740 235
rect 1700 200 1705 230
rect 1735 200 1740 230
rect 1760 225 1790 235
rect 1700 195 1740 200
rect 555 -335 595 -330
rect 555 -365 560 -335
rect 590 -365 595 -335
rect 555 -370 595 -365
rect 715 -335 755 -330
rect 715 -365 720 -335
rect 750 -365 755 -335
rect 715 -370 755 -365
rect 825 -335 865 -330
rect 825 -365 830 -335
rect 860 -365 865 -335
rect 825 -370 865 -365
rect 935 -335 975 -330
rect 935 -365 940 -335
rect 970 -365 975 -335
rect 935 -370 975 -365
rect 1095 -335 1135 -330
rect 1095 -365 1100 -335
rect 1130 -365 1135 -335
rect 1095 -370 1135 -365
rect 445 -440 475 -430
rect 445 -460 450 -440
rect 470 -460 475 -440
rect 445 -470 475 -460
rect 1245 -485 1265 175
rect 1765 -330 1785 225
rect 1755 -335 1795 -330
rect 1755 -365 1760 -335
rect 1790 -365 1795 -335
rect 1755 -370 1795 -365
rect 1850 -430 1870 975
rect 1895 675 1915 1450
rect 1975 1105 2015 1110
rect 1975 1075 1980 1105
rect 2010 1075 2015 1105
rect 1975 1070 2015 1075
rect 1930 760 1970 765
rect 1930 730 1935 760
rect 1965 730 1970 760
rect 1930 725 1970 730
rect 1885 670 1925 675
rect 1885 640 1890 670
rect 1920 640 1925 670
rect 1885 635 1925 640
rect 1895 -85 1915 635
rect 1940 610 1960 725
rect 1930 605 1970 610
rect 1930 575 1935 605
rect 1965 575 1970 605
rect 1930 570 1970 575
rect 1885 -90 1925 -85
rect 1885 -120 1890 -90
rect 1920 -120 1925 -90
rect 1885 -125 1925 -120
rect 1940 -140 1960 570
rect 1930 -145 1970 -140
rect 1930 -175 1935 -145
rect 1965 -175 1970 -145
rect 1885 -245 1925 -240
rect 1885 -275 1890 -245
rect 1920 -275 1925 -245
rect 1885 -280 1925 -275
rect 1895 -375 1915 -280
rect 1940 -305 1960 -175
rect 1985 -190 2005 1070
rect 2030 905 2050 1635
rect 2365 1625 2405 1630
rect 2365 1595 2370 1625
rect 2400 1595 2405 1625
rect 2365 1590 2405 1595
rect 3100 1490 3140 1495
rect 2125 1485 2165 1490
rect 2125 1455 2130 1485
rect 2160 1455 2165 1485
rect 2125 1450 2165 1455
rect 2235 1485 2275 1490
rect 2235 1455 2240 1485
rect 2270 1455 2275 1485
rect 2235 1450 2275 1455
rect 2345 1485 2385 1490
rect 2345 1455 2350 1485
rect 2380 1455 2385 1485
rect 2345 1450 2385 1455
rect 2455 1485 2495 1490
rect 2455 1455 2460 1485
rect 2490 1455 2495 1485
rect 2455 1450 2495 1455
rect 2565 1485 2605 1490
rect 2565 1455 2570 1485
rect 2600 1455 2605 1485
rect 2565 1450 2605 1455
rect 2675 1485 2715 1490
rect 2675 1455 2680 1485
rect 2710 1455 2715 1485
rect 2675 1450 2715 1455
rect 2785 1485 2825 1490
rect 2785 1455 2790 1485
rect 2820 1455 2825 1485
rect 3100 1460 3105 1490
rect 3135 1460 3140 1490
rect 3100 1455 3140 1460
rect 2785 1450 2825 1455
rect 2130 1420 2160 1450
rect 2020 900 2060 905
rect 2020 870 2025 900
rect 2055 870 2060 900
rect 2020 865 2060 870
rect 2030 720 2050 865
rect 2130 850 2135 1420
rect 2155 850 2160 1420
rect 2130 840 2160 850
rect 2185 1420 2215 1430
rect 2185 850 2190 1420
rect 2210 850 2215 1420
rect 2185 820 2215 850
rect 2240 1420 2270 1450
rect 2240 850 2245 1420
rect 2265 850 2270 1420
rect 2240 840 2270 850
rect 2295 1420 2325 1430
rect 2295 850 2300 1420
rect 2320 850 2325 1420
rect 2295 820 2325 850
rect 2350 1420 2380 1450
rect 2350 850 2355 1420
rect 2375 850 2380 1420
rect 2350 840 2380 850
rect 2405 1420 2435 1430
rect 2405 850 2410 1420
rect 2430 850 2435 1420
rect 2405 820 2435 850
rect 2460 1420 2490 1450
rect 2460 850 2465 1420
rect 2485 850 2490 1420
rect 2460 840 2490 850
rect 2515 1420 2545 1430
rect 2515 850 2520 1420
rect 2540 850 2545 1420
rect 2515 820 2545 850
rect 2570 1420 2600 1450
rect 2570 850 2575 1420
rect 2595 850 2600 1420
rect 2570 840 2600 850
rect 2625 1420 2655 1430
rect 2625 850 2630 1420
rect 2650 850 2655 1420
rect 2625 820 2655 850
rect 2680 1420 2710 1450
rect 2680 850 2685 1420
rect 2705 850 2710 1420
rect 2680 840 2710 850
rect 2735 1420 2765 1430
rect 2735 850 2740 1420
rect 2760 850 2765 1420
rect 2735 820 2765 850
rect 2790 1420 2820 1450
rect 3110 1430 3130 1455
rect 2790 850 2795 1420
rect 2815 850 2820 1420
rect 3050 1420 3191 1430
rect 3050 1400 3055 1420
rect 3075 1400 3110 1420
rect 3130 1400 3165 1420
rect 3185 1400 3191 1420
rect 3050 1390 3191 1400
rect 2790 840 2820 850
rect 2180 815 2220 820
rect 2180 785 2185 815
rect 2215 785 2220 815
rect 2180 780 2220 785
rect 2290 815 2330 820
rect 2290 785 2295 815
rect 2325 785 2330 815
rect 2290 780 2330 785
rect 2400 815 2440 820
rect 2400 785 2405 815
rect 2435 785 2440 815
rect 2400 780 2440 785
rect 2510 815 2550 820
rect 2510 785 2515 815
rect 2545 785 2550 815
rect 2510 780 2550 785
rect 2620 815 2660 820
rect 2620 785 2625 815
rect 2655 785 2660 815
rect 2620 780 2660 785
rect 2730 815 2770 820
rect 2730 785 2735 815
rect 2765 785 2770 815
rect 3050 815 3191 825
rect 3050 795 3055 815
rect 3075 795 3110 815
rect 3130 795 3165 815
rect 3185 795 3191 815
rect 3050 785 3191 795
rect 2730 780 2770 785
rect 2630 765 2650 780
rect 2180 760 2220 765
rect 2180 730 2185 760
rect 2215 730 2220 760
rect 2180 725 2220 730
rect 2620 760 2660 765
rect 2620 730 2625 760
rect 2655 730 2660 760
rect 2620 725 2660 730
rect 2020 715 2060 720
rect 2020 685 2025 715
rect 2055 685 2060 715
rect 2020 680 2060 685
rect 2030 345 2050 680
rect 2190 675 2210 725
rect 3110 720 3130 785
rect 3190 760 3230 765
rect 3190 730 3195 760
rect 3225 730 3230 760
rect 3190 725 3230 730
rect 2455 715 2495 720
rect 2455 685 2460 715
rect 2490 685 2495 715
rect 2455 680 2495 685
rect 3100 715 3140 720
rect 3100 685 3105 715
rect 3135 685 3140 715
rect 3100 680 3140 685
rect 2125 670 2165 675
rect 2125 640 2130 670
rect 2160 640 2165 670
rect 2125 635 2165 640
rect 2180 670 2220 675
rect 2180 640 2185 670
rect 2215 640 2220 670
rect 2180 635 2220 640
rect 2290 670 2330 675
rect 2290 640 2295 670
rect 2325 640 2330 670
rect 2290 635 2330 640
rect 2400 670 2440 675
rect 2400 640 2405 670
rect 2435 640 2440 670
rect 2400 635 2440 640
rect 2510 670 2550 675
rect 2510 640 2515 670
rect 2545 640 2550 670
rect 2510 635 2550 640
rect 2620 670 2660 675
rect 2620 640 2625 670
rect 2655 640 2660 670
rect 2620 635 2660 640
rect 2730 670 2770 675
rect 2730 640 2735 670
rect 2765 640 2770 670
rect 2730 635 2770 640
rect 2785 670 2825 675
rect 2785 640 2790 670
rect 2820 640 2825 670
rect 2785 635 2825 640
rect 2130 605 2160 635
rect 2130 435 2135 605
rect 2155 435 2160 605
rect 2130 425 2160 435
rect 2185 605 2215 635
rect 2185 435 2190 605
rect 2210 435 2215 605
rect 2185 425 2215 435
rect 2240 605 2270 615
rect 2240 435 2245 605
rect 2265 435 2270 605
rect 2240 420 2270 435
rect 2295 605 2325 635
rect 2295 435 2300 605
rect 2320 435 2325 605
rect 2295 425 2325 435
rect 2350 605 2380 615
rect 2350 435 2355 605
rect 2375 435 2380 605
rect 2350 420 2380 435
rect 2405 605 2435 635
rect 2405 435 2410 605
rect 2430 435 2435 605
rect 2405 425 2435 435
rect 2460 605 2490 615
rect 2460 435 2465 605
rect 2485 435 2490 605
rect 2460 420 2490 435
rect 2515 605 2545 635
rect 2515 435 2520 605
rect 2540 435 2545 605
rect 2515 425 2545 435
rect 2570 605 2600 615
rect 2570 435 2575 605
rect 2595 435 2600 605
rect 2570 420 2600 435
rect 2625 605 2655 635
rect 2625 435 2630 605
rect 2650 435 2655 605
rect 2625 425 2655 435
rect 2680 605 2710 615
rect 2680 435 2685 605
rect 2705 435 2710 605
rect 2680 420 2710 435
rect 2735 605 2765 635
rect 2735 435 2740 605
rect 2760 435 2765 605
rect 2735 425 2765 435
rect 2790 605 2820 635
rect 2790 435 2795 605
rect 2815 435 2820 605
rect 2790 425 2820 435
rect 2235 415 2275 420
rect 2235 385 2240 415
rect 2270 385 2275 415
rect 2235 380 2275 385
rect 2345 415 2385 420
rect 2345 385 2350 415
rect 2380 385 2385 415
rect 2345 380 2385 385
rect 2455 415 2495 420
rect 2455 385 2460 415
rect 2490 385 2495 415
rect 2455 380 2495 385
rect 2565 415 2605 420
rect 2565 385 2570 415
rect 2600 385 2605 415
rect 2565 380 2605 385
rect 2675 415 2715 420
rect 2675 385 2680 415
rect 2710 385 2715 415
rect 2675 380 2715 385
rect 2920 415 2960 420
rect 2920 385 2925 415
rect 2955 385 2960 415
rect 2920 380 2960 385
rect 2020 340 2060 345
rect 2020 310 2025 340
rect 2055 310 2060 340
rect 2020 305 2060 310
rect 2400 340 2440 345
rect 2400 310 2405 340
rect 2435 310 2440 340
rect 2400 305 2440 310
rect 2235 265 2275 270
rect 2235 235 2240 265
rect 2270 235 2275 265
rect 2235 230 2275 235
rect 2345 265 2385 270
rect 2345 235 2350 265
rect 2380 235 2385 265
rect 2345 230 2385 235
rect 2455 265 2495 270
rect 2455 235 2460 265
rect 2490 235 2495 265
rect 2455 230 2495 235
rect 2565 265 2605 270
rect 2565 235 2570 265
rect 2600 235 2605 265
rect 2565 230 2605 235
rect 2675 265 2715 270
rect 2675 235 2680 265
rect 2710 235 2715 265
rect 2675 230 2715 235
rect 2875 265 2915 270
rect 2875 235 2880 265
rect 2910 235 2915 265
rect 2875 230 2915 235
rect 2130 215 2160 225
rect 2130 -55 2135 215
rect 2155 -55 2160 215
rect 2130 -85 2160 -55
rect 2185 215 2215 225
rect 2185 -55 2190 215
rect 2210 -55 2215 215
rect 2185 -85 2215 -55
rect 2240 215 2270 230
rect 2240 -55 2245 215
rect 2265 -55 2270 215
rect 2240 -65 2270 -55
rect 2295 215 2325 225
rect 2295 -55 2300 215
rect 2320 -55 2325 215
rect 2295 -85 2325 -55
rect 2350 215 2380 230
rect 2350 -55 2355 215
rect 2375 -55 2380 215
rect 2350 -65 2380 -55
rect 2405 215 2435 225
rect 2405 -55 2410 215
rect 2430 -55 2435 215
rect 2405 -85 2435 -55
rect 2460 215 2490 230
rect 2460 -55 2465 215
rect 2485 -55 2490 215
rect 2460 -65 2490 -55
rect 2515 215 2545 225
rect 2515 -55 2520 215
rect 2540 -55 2545 215
rect 2515 -85 2545 -55
rect 2570 215 2600 230
rect 2570 -55 2575 215
rect 2595 -55 2600 215
rect 2570 -65 2600 -55
rect 2625 215 2655 225
rect 2625 -55 2630 215
rect 2650 -55 2655 215
rect 2625 -85 2655 -55
rect 2680 215 2710 230
rect 2680 -55 2685 215
rect 2705 -55 2710 215
rect 2680 -65 2710 -55
rect 2735 215 2765 225
rect 2735 -55 2740 215
rect 2760 -55 2765 215
rect 2735 -85 2765 -55
rect 2790 215 2820 225
rect 2790 -55 2795 215
rect 2815 -55 2820 215
rect 2790 -85 2820 -55
rect 2885 -85 2905 230
rect 2125 -95 2165 -85
rect 2125 -115 2135 -95
rect 2155 -115 2165 -95
rect 2125 -145 2165 -115
rect 2180 -90 2220 -85
rect 2180 -120 2185 -90
rect 2215 -120 2220 -90
rect 2180 -125 2220 -120
rect 2290 -90 2330 -85
rect 2290 -120 2295 -90
rect 2325 -120 2330 -90
rect 2290 -125 2330 -120
rect 2400 -90 2440 -85
rect 2400 -120 2405 -90
rect 2435 -120 2440 -90
rect 2400 -125 2440 -120
rect 2510 -90 2550 -85
rect 2510 -120 2515 -90
rect 2545 -120 2550 -90
rect 2510 -125 2550 -120
rect 2620 -90 2660 -85
rect 2620 -120 2625 -90
rect 2655 -120 2660 -90
rect 2620 -125 2660 -120
rect 2730 -90 2770 -85
rect 2730 -120 2735 -90
rect 2765 -120 2770 -90
rect 2730 -125 2770 -120
rect 2785 -90 2825 -85
rect 2785 -120 2790 -90
rect 2820 -120 2825 -90
rect 2125 -175 2130 -145
rect 2160 -175 2165 -145
rect 2125 -180 2165 -175
rect 2785 -145 2825 -120
rect 2875 -90 2915 -85
rect 2875 -120 2880 -90
rect 2910 -120 2915 -90
rect 2875 -125 2915 -120
rect 2930 -140 2950 380
rect 3200 360 3220 725
rect 3185 350 3235 360
rect 3185 320 3195 350
rect 3225 320 3235 350
rect 3185 310 3235 320
rect 2965 -120 2969 -85
rect 2996 -120 3000 -85
rect 3025 -120 3029 -85
rect 3056 -120 3060 -85
rect 3085 -120 3089 -85
rect 3116 -120 3120 -85
rect 3145 -120 3149 -85
rect 3176 -120 3180 -85
rect 2785 -175 2790 -145
rect 2820 -175 2825 -145
rect 2785 -180 2825 -175
rect 2920 -145 2960 -140
rect 2920 -175 2925 -145
rect 2955 -175 2960 -145
rect 2920 -180 2960 -175
rect 3025 -145 3060 -120
rect 3025 -180 3060 -175
rect 3150 -185 3175 -120
rect 3145 -190 3180 -185
rect 1975 -220 1980 -190
rect 2010 -220 2015 -190
rect 1975 -225 2015 -220
rect 3145 -225 3180 -220
rect 2455 -245 2495 -240
rect 2455 -275 2460 -245
rect 2490 -275 2495 -245
rect 2455 -280 2495 -275
rect 2945 -245 2980 -240
rect 2945 -280 2980 -275
rect 2255 -305 2295 -300
rect 1930 -310 1970 -305
rect 1930 -340 1935 -310
rect 1965 -340 1970 -310
rect 2255 -335 2260 -305
rect 2290 -335 2295 -305
rect 2255 -340 2295 -335
rect 2455 -305 2495 -300
rect 2455 -335 2460 -305
rect 2490 -335 2495 -305
rect 2455 -340 2495 -335
rect 2655 -305 2695 -300
rect 2655 -335 2660 -305
rect 2690 -335 2695 -305
rect 2655 -340 2695 -335
rect 2885 -305 2920 -300
rect 2885 -340 2920 -335
rect 1930 -345 1970 -340
rect 1885 -380 1925 -375
rect 1885 -410 1890 -380
rect 1920 -410 1925 -380
rect 1885 -415 1925 -410
rect 1350 -435 1390 -430
rect 1350 -465 1355 -435
rect 1385 -465 1390 -435
rect 1350 -470 1390 -465
rect 1840 -435 1880 -430
rect 1840 -465 1845 -435
rect 1875 -465 1880 -435
rect 1840 -470 1880 -465
rect 385 -490 425 -485
rect 385 -520 390 -490
rect 420 -520 425 -490
rect 385 -525 425 -520
rect 495 -490 535 -485
rect 495 -520 500 -490
rect 530 -520 535 -490
rect 495 -525 535 -520
rect 605 -490 645 -485
rect 605 -520 610 -490
rect 640 -520 645 -490
rect 605 -525 645 -520
rect 715 -490 755 -485
rect 715 -520 720 -490
rect 750 -520 755 -490
rect 715 -525 755 -520
rect 825 -490 865 -485
rect 825 -520 830 -490
rect 860 -520 865 -490
rect 825 -525 865 -520
rect 935 -490 975 -485
rect 935 -520 940 -490
rect 970 -520 975 -490
rect 935 -525 975 -520
rect 1045 -490 1085 -485
rect 1045 -520 1050 -490
rect 1080 -520 1085 -490
rect 1045 -525 1085 -520
rect 1155 -490 1195 -485
rect 1155 -520 1160 -490
rect 1190 -520 1195 -490
rect 1155 -525 1195 -520
rect 1245 -490 1305 -485
rect 1245 -520 1270 -490
rect 1300 -520 1305 -490
rect 1245 -525 1305 -520
rect 1375 -490 1415 -485
rect 1375 -520 1380 -490
rect 1410 -520 1415 -490
rect 1375 -525 1415 -520
rect 280 -550 310 -540
rect 280 -770 285 -550
rect 305 -770 310 -550
rect 280 -800 310 -770
rect 335 -550 365 -540
rect 335 -770 340 -550
rect 360 -770 365 -550
rect 335 -800 365 -770
rect 390 -550 420 -525
rect 390 -770 395 -550
rect 415 -770 420 -550
rect 275 -805 315 -800
rect 275 -835 280 -805
rect 310 -835 315 -805
rect 275 -840 315 -835
rect 330 -805 370 -800
rect 330 -835 335 -805
rect 365 -835 370 -805
rect 330 -840 370 -835
rect 390 -845 420 -770
rect 445 -550 475 -540
rect 445 -770 450 -550
rect 470 -770 475 -550
rect 445 -800 475 -770
rect 500 -550 530 -525
rect 500 -770 505 -550
rect 525 -770 530 -550
rect 440 -805 480 -800
rect 440 -835 445 -805
rect 475 -835 480 -805
rect 440 -840 480 -835
rect 500 -845 530 -770
rect 555 -550 585 -540
rect 555 -770 560 -550
rect 580 -770 585 -550
rect 555 -800 585 -770
rect 610 -550 640 -525
rect 610 -770 615 -550
rect 635 -770 640 -550
rect 550 -805 590 -800
rect 550 -835 555 -805
rect 585 -835 590 -805
rect 550 -840 590 -835
rect 610 -845 640 -770
rect 665 -550 695 -540
rect 665 -770 670 -550
rect 690 -770 695 -550
rect 665 -800 695 -770
rect 720 -550 750 -525
rect 720 -770 725 -550
rect 745 -770 750 -550
rect 660 -805 700 -800
rect 660 -835 665 -805
rect 695 -835 700 -805
rect 660 -840 700 -835
rect 720 -845 750 -770
rect 775 -550 805 -540
rect 775 -770 780 -550
rect 800 -770 805 -550
rect 775 -800 805 -770
rect 830 -550 860 -525
rect 830 -770 835 -550
rect 855 -770 860 -550
rect 770 -805 810 -800
rect 770 -835 775 -805
rect 805 -835 810 -805
rect 770 -840 810 -835
rect 830 -845 860 -770
rect 885 -550 915 -540
rect 885 -770 890 -550
rect 910 -770 915 -550
rect 885 -800 915 -770
rect 940 -550 970 -525
rect 940 -770 945 -550
rect 965 -770 970 -550
rect 880 -805 920 -800
rect 880 -835 885 -805
rect 915 -835 920 -805
rect 880 -840 920 -835
rect 940 -845 970 -770
rect 995 -550 1025 -540
rect 995 -770 1000 -550
rect 1020 -770 1025 -550
rect 995 -800 1025 -770
rect 1050 -550 1080 -525
rect 1050 -770 1055 -550
rect 1075 -770 1080 -550
rect 990 -805 1030 -800
rect 990 -835 995 -805
rect 1025 -835 1030 -805
rect 990 -840 1030 -835
rect 1050 -845 1080 -770
rect 1105 -550 1135 -540
rect 1105 -770 1110 -550
rect 1130 -770 1135 -550
rect 1105 -800 1135 -770
rect 1160 -550 1190 -525
rect 1160 -770 1165 -550
rect 1185 -770 1190 -550
rect 1100 -805 1140 -800
rect 1100 -835 1105 -805
rect 1135 -835 1140 -805
rect 1100 -840 1140 -835
rect 1160 -845 1190 -770
rect 1215 -550 1245 -540
rect 1215 -770 1220 -550
rect 1240 -770 1245 -550
rect 1215 -800 1245 -770
rect 1270 -550 1300 -525
rect 1270 -770 1275 -550
rect 1295 -770 1300 -550
rect 1210 -805 1250 -800
rect 1210 -835 1215 -805
rect 1245 -835 1250 -805
rect 1210 -840 1250 -835
rect 1270 -845 1300 -770
rect 1325 -550 1355 -540
rect 1325 -770 1330 -550
rect 1350 -770 1355 -550
rect 1325 -800 1355 -770
rect 1380 -550 1410 -525
rect 1380 -770 1385 -550
rect 1405 -770 1410 -550
rect 1320 -805 1360 -800
rect 1320 -835 1325 -805
rect 1355 -835 1360 -805
rect 1320 -840 1360 -835
rect 1380 -845 1410 -770
rect 1435 -550 1465 -540
rect 1435 -770 1440 -550
rect 1460 -770 1465 -550
rect 1435 -800 1465 -770
rect 1940 -800 1960 -345
rect 2160 -370 2190 -360
rect 1430 -805 1470 -800
rect 1430 -835 1435 -805
rect 1465 -835 1470 -805
rect 1430 -840 1470 -835
rect 1930 -805 1970 -800
rect 1930 -835 1935 -805
rect 1965 -835 1970 -805
rect 1930 -840 1970 -835
rect 385 -850 425 -845
rect 385 -880 390 -850
rect 420 -880 425 -850
rect 385 -885 425 -880
rect 495 -850 535 -845
rect 495 -880 500 -850
rect 530 -880 535 -850
rect 495 -885 535 -880
rect 605 -850 645 -845
rect 605 -880 610 -850
rect 640 -880 645 -850
rect 605 -885 645 -880
rect 715 -850 755 -845
rect 715 -880 720 -850
rect 750 -880 755 -850
rect 715 -885 755 -880
rect 825 -850 865 -845
rect 825 -880 830 -850
rect 860 -880 865 -850
rect 825 -885 865 -880
rect 935 -850 975 -845
rect 935 -880 940 -850
rect 970 -880 975 -850
rect 935 -885 975 -880
rect 1045 -850 1085 -845
rect 1045 -880 1050 -850
rect 1080 -880 1085 -850
rect 1045 -885 1085 -880
rect 1155 -850 1195 -845
rect 1155 -880 1160 -850
rect 1190 -880 1195 -850
rect 1155 -885 1195 -880
rect 1265 -850 1305 -845
rect 1265 -880 1270 -850
rect 1300 -880 1305 -850
rect 1265 -885 1305 -880
rect 1375 -850 1415 -845
rect 1375 -880 1380 -850
rect 1410 -880 1415 -850
rect 1375 -885 1415 -880
rect 595 -915 635 -910
rect 595 -945 600 -915
rect 630 -945 635 -915
rect 595 -950 635 -945
rect 705 -915 745 -910
rect 705 -945 710 -915
rect 740 -945 745 -915
rect 705 -950 745 -945
rect 925 -915 965 -910
rect 925 -945 930 -915
rect 960 -945 965 -915
rect 925 -950 965 -945
rect -190 -960 -150 -955
rect -190 -990 -185 -960
rect -155 -990 -150 -960
rect -190 -995 -150 -990
rect 540 -960 580 -955
rect 540 -990 545 -960
rect 575 -990 580 -960
rect 540 -995 580 -990
rect 490 -1025 520 -1015
rect 490 -1145 495 -1025
rect 515 -1145 520 -1025
rect 490 -1185 520 -1145
rect 490 -1205 495 -1185
rect 515 -1205 520 -1185
rect 545 -1025 575 -995
rect 545 -1145 550 -1025
rect 570 -1145 575 -1025
rect 545 -1205 575 -1145
rect 600 -1025 630 -950
rect 650 -960 690 -955
rect 650 -990 655 -960
rect 685 -990 690 -960
rect 650 -995 690 -990
rect 600 -1145 605 -1025
rect 625 -1145 630 -1025
rect 600 -1160 630 -1145
rect 655 -1025 685 -995
rect 655 -1145 660 -1025
rect 680 -1145 685 -1025
rect 595 -1165 635 -1160
rect 595 -1195 600 -1165
rect 630 -1195 635 -1165
rect 595 -1200 635 -1195
rect 655 -1205 685 -1145
rect 710 -1025 740 -950
rect 760 -960 800 -955
rect 760 -990 765 -960
rect 795 -990 800 -960
rect 760 -995 800 -990
rect 710 -1145 715 -1025
rect 735 -1145 740 -1025
rect 710 -1160 740 -1145
rect 765 -1025 795 -995
rect 765 -1145 770 -1025
rect 790 -1145 795 -1025
rect 705 -1165 745 -1160
rect 705 -1195 710 -1165
rect 740 -1195 745 -1165
rect 705 -1200 745 -1195
rect 765 -1205 795 -1145
rect 820 -1025 850 -1015
rect 820 -1145 825 -1025
rect 845 -1145 850 -1025
rect 820 -1185 850 -1145
rect 930 -1025 960 -950
rect 1270 -955 1300 -885
rect 1095 -960 1135 -955
rect 1095 -990 1100 -960
rect 1130 -990 1135 -960
rect 1095 -995 1135 -990
rect 1265 -960 1305 -955
rect 1265 -990 1270 -960
rect 1300 -990 1305 -960
rect 1265 -995 1305 -990
rect 930 -1145 935 -1025
rect 955 -1145 960 -1025
rect 930 -1160 960 -1145
rect 1270 -1025 1300 -995
rect 1270 -1145 1275 -1025
rect 1295 -1145 1300 -1025
rect 1270 -1155 1300 -1145
rect 820 -1205 825 -1185
rect 845 -1205 850 -1185
rect 925 -1165 965 -1160
rect 925 -1195 930 -1165
rect 960 -1195 965 -1165
rect 925 -1200 965 -1195
rect 490 -1250 520 -1205
rect 540 -1210 580 -1205
rect 540 -1240 545 -1210
rect 575 -1240 580 -1210
rect 540 -1245 580 -1240
rect 650 -1210 690 -1205
rect 650 -1240 655 -1210
rect 685 -1240 690 -1210
rect 650 -1245 690 -1240
rect 760 -1210 800 -1205
rect 760 -1240 765 -1210
rect 795 -1240 800 -1210
rect 760 -1245 800 -1240
rect 820 -1250 850 -1205
rect 1940 -1250 1960 -840
rect 2160 -1040 2165 -370
rect 2185 -1040 2190 -370
rect 2160 -1070 2190 -1040
rect 2260 -370 2290 -340
rect 2260 -1040 2265 -370
rect 2285 -1040 2290 -370
rect 2260 -1050 2290 -1040
rect 2360 -370 2390 -360
rect 2360 -1040 2365 -370
rect 2385 -1040 2390 -370
rect 2360 -1070 2390 -1040
rect 2460 -370 2490 -340
rect 2460 -1040 2465 -370
rect 2485 -1040 2490 -370
rect 2460 -1050 2490 -1040
rect 2560 -370 2590 -360
rect 2560 -1040 2565 -370
rect 2585 -1040 2590 -370
rect 2560 -1070 2590 -1040
rect 2660 -370 2690 -340
rect 2660 -1040 2665 -370
rect 2685 -1040 2690 -370
rect 2660 -1050 2690 -1040
rect 2760 -370 2790 -360
rect 2760 -1040 2765 -370
rect 2785 -1040 2790 -370
rect 2890 -380 2915 -340
rect 2950 -380 2975 -280
rect 3200 -300 3220 310
rect 3190 -305 3230 -300
rect 3190 -335 3195 -305
rect 3225 -335 3230 -305
rect 3190 -340 3230 -335
rect 2885 -415 2889 -380
rect 2916 -415 2920 -380
rect 2945 -415 2949 -380
rect 2976 -415 2980 -380
rect 2760 -1070 2790 -1040
rect 2155 -1075 2195 -1070
rect 2155 -1105 2160 -1075
rect 2190 -1105 2195 -1075
rect 2155 -1110 2195 -1105
rect 2355 -1075 2395 -1070
rect 2355 -1105 2360 -1075
rect 2390 -1105 2395 -1075
rect 2355 -1110 2395 -1105
rect 2555 -1075 2595 -1070
rect 2555 -1105 2560 -1075
rect 2590 -1105 2595 -1075
rect 2555 -1110 2595 -1105
rect 2755 -1075 2795 -1070
rect 2755 -1105 2760 -1075
rect 2790 -1105 2795 -1075
rect 2755 -1110 2795 -1105
rect 2365 -1250 2385 -1110
rect -705 -1255 -665 -1250
rect -705 -1285 -700 -1255
rect -670 -1285 -665 -1255
rect -705 -1290 -665 -1285
rect -280 -1255 -240 -1250
rect -280 -1285 -275 -1255
rect -245 -1285 -240 -1255
rect -280 -1290 -240 -1285
rect 485 -1255 525 -1250
rect 485 -1285 490 -1255
rect 520 -1285 525 -1255
rect 485 -1290 525 -1285
rect 815 -1255 855 -1250
rect 815 -1285 820 -1255
rect 850 -1285 855 -1255
rect 815 -1290 855 -1285
rect 1930 -1255 1970 -1250
rect 1930 -1285 1935 -1255
rect 1965 -1285 1970 -1255
rect 1930 -1290 1970 -1285
rect 2355 -1255 2395 -1250
rect 2355 -1285 2360 -1255
rect 2390 -1285 2395 -1255
rect 2355 -1290 2395 -1285
rect 825 -1295 845 -1290
rect 835 -2420 855 -1295
rect 825 -2425 865 -2420
rect 825 -2455 830 -2425
rect 860 -2455 865 -2425
rect 825 -2460 865 -2455
<< via1 >>
rect 830 4245 860 4275
rect 215 2750 245 2780
rect 35 2720 65 2725
rect 35 2700 40 2720
rect 40 2700 60 2720
rect 60 2700 65 2720
rect 35 2695 65 2700
rect 155 2695 185 2725
rect 625 2750 655 2780
rect 215 2720 245 2725
rect 215 2700 220 2720
rect 220 2700 240 2720
rect 240 2700 245 2720
rect 215 2695 245 2700
rect 505 2550 535 2555
rect 505 2530 510 2550
rect 510 2530 530 2550
rect 530 2530 535 2550
rect 505 2525 535 2530
rect 565 2550 595 2555
rect 565 2530 570 2550
rect 570 2530 590 2550
rect 590 2530 595 2550
rect 565 2525 595 2530
rect 1035 2750 1065 2780
rect 1445 2750 1475 2780
rect 830 2695 860 2725
rect 975 2720 1005 2725
rect 975 2700 980 2720
rect 980 2700 1000 2720
rect 1000 2700 1005 2720
rect 975 2695 1005 2700
rect 685 2550 715 2555
rect 685 2530 690 2550
rect 690 2530 710 2550
rect 710 2530 715 2550
rect 685 2525 715 2530
rect 830 2525 860 2555
rect 80 2300 110 2305
rect 80 2280 85 2300
rect 85 2280 105 2300
rect 105 2280 110 2300
rect 80 2275 110 2280
rect 139 2300 169 2305
rect 139 2280 144 2300
rect 144 2280 164 2300
rect 164 2280 169 2300
rect 139 2275 169 2280
rect 609 2300 639 2305
rect 609 2280 614 2300
rect 614 2280 634 2300
rect 634 2280 639 2300
rect 609 2275 639 2280
rect 775 2275 805 2305
rect -800 2175 -770 2205
rect -230 2175 -200 2205
rect -1160 2120 -1130 2150
rect -1040 2120 -1010 2150
rect -920 2120 -890 2150
rect -800 2120 -770 2150
rect -680 2120 -650 2150
rect -560 2120 -530 2150
rect -440 2145 -410 2150
rect -440 2125 -435 2145
rect -435 2125 -415 2145
rect -415 2125 -410 2145
rect -440 2120 -410 2125
rect -275 2120 -245 2150
rect -1100 1700 -1070 1730
rect -980 1700 -950 1730
rect -860 1700 -830 1730
rect -740 1700 -710 1730
rect -620 1700 -590 1730
rect -500 1700 -470 1730
rect -275 1700 -245 1730
rect -365 1640 -335 1670
rect -710 1620 -680 1625
rect -710 1600 -705 1620
rect -705 1600 -685 1620
rect -685 1600 -680 1620
rect -710 1595 -680 1600
rect -1445 1510 -1415 1540
rect -1130 1480 -1100 1485
rect -1130 1460 -1125 1480
rect -1125 1460 -1105 1480
rect -1105 1460 -1100 1480
rect -1130 1455 -1100 1460
rect -1020 1455 -990 1485
rect -910 1455 -880 1485
rect -800 1455 -770 1485
rect -690 1455 -660 1485
rect -580 1455 -550 1485
rect -470 1480 -440 1485
rect -470 1460 -465 1480
rect -465 1460 -445 1480
rect -445 1460 -440 1480
rect -470 1455 -440 1460
rect -35 2145 -5 2150
rect -35 2125 -30 2145
rect -30 2125 -10 2145
rect -10 2125 -5 2145
rect -35 2120 -5 2125
rect 85 2120 115 2150
rect 205 2120 235 2150
rect 325 2120 355 2150
rect 445 2120 475 2150
rect 565 2120 595 2150
rect 685 2145 715 2150
rect 685 2125 690 2145
rect 690 2125 710 2145
rect 710 2125 715 2145
rect 685 2120 715 2125
rect 25 1700 55 1730
rect 145 1700 175 1730
rect 265 1700 295 1730
rect 385 1700 415 1730
rect 505 1700 535 1730
rect 625 1700 655 1730
rect 1095 2695 1125 2725
rect 1155 2720 1185 2725
rect 1155 2700 1160 2720
rect 1160 2700 1180 2720
rect 1180 2700 1185 2720
rect 1155 2695 1185 2700
rect 1445 2720 1475 2725
rect 1445 2700 1450 2720
rect 1450 2700 1470 2720
rect 1470 2700 1475 2720
rect 1445 2695 1475 2700
rect 1505 2695 1535 2725
rect 1625 2720 1655 2725
rect 1625 2700 1630 2720
rect 1630 2700 1650 2720
rect 1650 2700 1655 2720
rect 1625 2695 1655 2700
rect 1521 2300 1551 2305
rect 1521 2280 1526 2300
rect 1526 2280 1546 2300
rect 1546 2280 1551 2300
rect 1521 2275 1551 2280
rect 885 2230 915 2260
rect 830 2175 860 2205
rect 265 1640 295 1670
rect 415 1665 445 1670
rect 415 1645 420 1665
rect 420 1645 440 1665
rect 440 1645 445 1665
rect 415 1640 445 1645
rect 785 1640 815 1670
rect 1050 2220 1080 2250
rect 1565 2220 1595 2250
rect 1890 2175 1920 2205
rect 2460 2175 2490 2205
rect 975 2145 1005 2150
rect 975 2125 980 2145
rect 980 2125 1000 2145
rect 1000 2125 1005 2145
rect 975 2120 1005 2125
rect 1095 2120 1125 2150
rect 1215 2120 1245 2150
rect 1335 2120 1365 2150
rect 1455 2120 1485 2150
rect 1575 2120 1605 2150
rect 1695 2145 1725 2150
rect 1695 2125 1700 2145
rect 1700 2125 1720 2145
rect 1720 2125 1725 2145
rect 1695 2120 1725 2125
rect 1035 1700 1065 1730
rect 1155 1700 1185 1730
rect 1275 1700 1305 1730
rect 1395 1700 1425 1730
rect 1245 1665 1275 1670
rect 1245 1645 1250 1665
rect 1250 1645 1270 1665
rect 1270 1645 1275 1665
rect 1245 1640 1275 1645
rect 1515 1700 1545 1730
rect 1635 1700 1665 1730
rect 1395 1640 1425 1670
rect 875 1600 905 1630
rect 1935 2120 1965 2150
rect 2100 2145 2130 2150
rect 2100 2125 2105 2145
rect 2105 2125 2125 2145
rect 2125 2125 2130 2145
rect 2100 2120 2130 2125
rect 2220 2120 2250 2150
rect 2340 2120 2370 2150
rect 2460 2120 2490 2150
rect 2580 2120 2610 2150
rect 2700 2120 2730 2150
rect 2820 2120 2850 2150
rect 1935 1700 1965 1730
rect 2160 1700 2190 1730
rect 2280 1700 2310 1730
rect 2400 1700 2430 1730
rect 2520 1700 2550 1730
rect 2640 1700 2670 1730
rect 2760 1700 2790 1730
rect 2025 1640 2055 1670
rect 460 1560 490 1565
rect 460 1540 465 1560
rect 465 1540 485 1560
rect 485 1540 490 1560
rect 460 1535 490 1540
rect 625 1535 655 1565
rect 790 1560 820 1565
rect 790 1540 795 1560
rect 795 1540 815 1560
rect 815 1540 820 1560
rect 790 1535 820 1540
rect 870 1560 900 1565
rect 870 1540 875 1560
rect 875 1540 895 1560
rect 895 1540 900 1560
rect 870 1535 900 1540
rect 1035 1535 1065 1565
rect 1200 1560 1230 1565
rect 1200 1540 1205 1560
rect 1205 1540 1225 1560
rect 1225 1540 1230 1560
rect 1200 1535 1230 1540
rect 1890 1535 1920 1565
rect -230 1455 -200 1485
rect 570 1490 600 1520
rect -320 1075 -290 1105
rect -365 870 -335 900
rect -1075 785 -1045 815
rect -1535 730 -1505 760
rect -965 785 -935 815
rect -855 785 -825 815
rect -745 785 -715 815
rect -635 785 -605 815
rect -525 785 -495 815
rect -965 730 -935 760
rect -525 730 -495 760
rect -1445 685 -1415 715
rect -800 710 -770 715
rect -800 690 -795 710
rect -795 690 -775 710
rect -775 690 -770 710
rect -800 685 -770 690
rect -365 685 -335 715
rect -1130 665 -1100 670
rect -1130 645 -1125 665
rect -1125 645 -1105 665
rect -1105 645 -1100 665
rect -1130 640 -1100 645
rect -1075 640 -1045 670
rect -965 640 -935 670
rect -855 640 -825 670
rect -745 640 -715 670
rect -635 640 -605 670
rect -525 640 -495 670
rect -470 665 -440 670
rect -470 645 -465 665
rect -465 645 -445 665
rect -445 645 -440 665
rect -470 640 -440 645
rect -1265 385 -1235 415
rect -1020 385 -990 415
rect -910 385 -880 415
rect -800 385 -770 415
rect -690 385 -660 415
rect -580 385 -550 415
rect -1535 320 -1505 350
rect -1486 -93 -1459 -85
rect -1486 -113 -1485 -93
rect -1485 -113 -1460 -93
rect -1460 -113 -1459 -93
rect -1486 -120 -1459 -113
rect -1426 -93 -1399 -85
rect -1426 -113 -1425 -93
rect -1425 -113 -1400 -93
rect -1400 -113 -1399 -93
rect -1426 -120 -1399 -113
rect -1366 -93 -1339 -85
rect -1366 -113 -1365 -93
rect -1365 -113 -1340 -93
rect -1340 -113 -1339 -93
rect -1366 -120 -1339 -113
rect -1306 -93 -1279 -85
rect -1306 -113 -1305 -93
rect -1305 -113 -1280 -93
rect -1280 -113 -1279 -93
rect -1306 -120 -1279 -113
rect -745 335 -715 340
rect -745 315 -740 335
rect -740 315 -720 335
rect -720 315 -715 335
rect -745 310 -715 315
rect -365 310 -335 340
rect -1220 235 -1190 265
rect -1020 235 -990 265
rect -910 235 -880 265
rect -800 235 -770 265
rect -690 235 -660 265
rect -580 235 -550 265
rect -1220 -120 -1190 -90
rect -1130 -95 -1100 -90
rect -1130 -115 -1125 -95
rect -1125 -115 -1105 -95
rect -1105 -115 -1100 -95
rect -1130 -120 -1100 -115
rect -1370 -175 -1335 -145
rect -1265 -175 -1235 -145
rect -1075 -120 -1045 -90
rect -965 -120 -935 -90
rect -855 -120 -825 -90
rect -745 -120 -715 -90
rect -635 -120 -605 -90
rect -525 -120 -495 -90
rect -1130 -175 -1100 -145
rect -470 -175 -440 -145
rect -275 740 -245 770
rect 680 1490 710 1520
rect 980 1490 1010 1520
rect 1090 1490 1120 1520
rect 1890 1455 1920 1485
rect 500 1175 530 1205
rect 625 1210 655 1215
rect 625 1190 630 1210
rect 630 1190 650 1210
rect 650 1190 655 1210
rect 625 1185 655 1190
rect 550 1150 580 1155
rect 550 1130 555 1150
rect 555 1130 575 1150
rect 575 1130 580 1150
rect 550 1125 580 1130
rect 750 1175 780 1205
rect 695 1075 725 1105
rect 1035 1210 1065 1215
rect 1035 1190 1040 1210
rect 1040 1190 1060 1210
rect 1060 1190 1065 1210
rect 1035 1185 1065 1190
rect 1100 1125 1130 1155
rect 970 1075 1000 1105
rect 800 1030 830 1060
rect 910 1030 940 1060
rect 800 975 830 1005
rect 885 975 915 1005
rect 1160 980 1190 1010
rect 1845 980 1875 1010
rect -185 920 -155 950
rect 120 945 150 950
rect 120 925 125 945
rect 125 925 145 945
rect 145 925 150 945
rect 1540 945 1570 950
rect 120 920 150 925
rect -230 640 -200 670
rect -230 -120 -200 -90
rect -275 -175 -245 -145
rect -1490 -220 -1455 -190
rect -320 -220 -290 -190
rect -1290 -275 -1255 -245
rect -800 -250 -770 -245
rect -800 -270 -795 -250
rect -795 -270 -775 -250
rect -775 -270 -770 -250
rect -800 -275 -770 -270
rect -1535 -335 -1505 -305
rect -1230 -335 -1195 -305
rect -1000 -335 -970 -305
rect -800 -335 -770 -305
rect -600 -335 -570 -305
rect -1286 -387 -1259 -380
rect -1286 -407 -1285 -387
rect -1285 -407 -1260 -387
rect -1260 -407 -1259 -387
rect -1286 -415 -1259 -407
rect -1226 -387 -1199 -380
rect -1226 -407 -1225 -387
rect -1225 -407 -1200 -387
rect -1200 -407 -1199 -387
rect -1226 -415 -1199 -407
rect -1100 -1080 -1070 -1075
rect -1100 -1100 -1095 -1080
rect -1095 -1100 -1075 -1080
rect -1075 -1100 -1070 -1080
rect -1100 -1105 -1070 -1100
rect -900 -1105 -870 -1075
rect -700 -1105 -670 -1075
rect -500 -1080 -470 -1075
rect -500 -1100 -495 -1080
rect -495 -1100 -475 -1080
rect -475 -1100 -470 -1080
rect -500 -1105 -470 -1100
rect -230 -275 -200 -245
rect -230 -410 -200 -380
rect -45 870 -15 900
rect 65 870 95 900
rect 175 870 205 900
rect 285 870 315 900
rect 395 870 425 900
rect 505 870 535 900
rect 1540 925 1545 945
rect 1545 925 1565 945
rect 1565 925 1570 945
rect 1540 920 1570 925
rect 10 655 40 685
rect 120 655 150 685
rect 230 655 260 685
rect -45 610 -15 640
rect 65 610 95 640
rect 175 610 205 640
rect -100 575 -70 605
rect 145 545 175 550
rect 145 525 150 545
rect 150 525 170 545
rect 170 525 175 545
rect 145 520 175 525
rect 340 655 370 685
rect 450 655 480 685
rect 285 610 315 640
rect 395 610 425 640
rect 505 610 535 640
rect 1155 870 1185 900
rect 1265 870 1295 900
rect 1375 870 1405 900
rect 1485 870 1515 900
rect 1595 870 1625 900
rect 1705 870 1735 900
rect 1210 655 1240 685
rect 1320 655 1350 685
rect 1430 655 1460 685
rect 1155 610 1185 640
rect 1265 610 1295 640
rect 1375 610 1405 640
rect 560 575 590 605
rect 720 600 750 605
rect 720 580 725 600
rect 725 580 745 600
rect 745 580 750 600
rect 720 575 750 580
rect 830 575 860 605
rect 940 600 970 605
rect 940 580 945 600
rect 945 580 965 600
rect 965 580 970 600
rect 940 575 970 580
rect 1100 575 1130 605
rect 795 545 825 550
rect 795 525 800 545
rect 800 525 820 545
rect 820 525 825 545
rect 795 520 825 525
rect 865 545 895 550
rect 865 525 870 545
rect 870 525 890 545
rect 890 525 895 545
rect 865 520 895 525
rect -45 435 -15 465
rect 65 435 95 465
rect 175 435 205 465
rect 230 445 260 475
rect 285 435 315 465
rect 395 435 425 465
rect 505 435 535 465
rect 1540 655 1570 685
rect 1650 655 1680 685
rect 1485 610 1515 640
rect 1595 610 1625 640
rect 1705 610 1735 640
rect 1760 575 1790 605
rect 1515 545 1545 550
rect 1515 525 1520 545
rect 1520 525 1540 545
rect 1540 525 1545 545
rect 1515 520 1545 525
rect 10 245 40 275
rect 120 245 150 275
rect 230 245 260 275
rect 340 245 370 275
rect 450 245 480 275
rect -45 200 -15 230
rect 65 200 95 230
rect 175 200 205 230
rect 285 200 315 230
rect 395 200 425 230
rect 505 200 535 230
rect 445 -40 475 -10
rect -100 -365 -70 -335
rect 775 175 805 205
rect 1155 435 1185 465
rect 1265 435 1295 465
rect 1375 435 1405 465
rect 1430 445 1460 475
rect 1485 435 1515 465
rect 1595 435 1625 465
rect 1705 435 1735 465
rect 1210 245 1240 275
rect 1320 245 1350 275
rect 1430 245 1460 275
rect 1540 245 1570 275
rect 1650 245 1680 275
rect 885 175 915 205
rect 830 120 860 150
rect 885 120 915 150
rect 775 65 805 95
rect 830 65 860 95
rect 775 10 805 40
rect 885 10 915 40
rect 830 -15 860 -10
rect 830 -35 835 -15
rect 835 -35 855 -15
rect 855 -35 860 -15
rect 830 -40 860 -35
rect 1155 200 1185 230
rect 1265 200 1295 230
rect 1375 200 1405 230
rect 1485 200 1515 230
rect 1595 200 1625 230
rect 1705 200 1735 230
rect 560 -365 590 -335
rect 720 -340 750 -335
rect 720 -360 725 -340
rect 725 -360 745 -340
rect 745 -360 750 -340
rect 720 -365 750 -360
rect 830 -365 860 -335
rect 940 -340 970 -335
rect 940 -360 945 -340
rect 945 -360 965 -340
rect 965 -360 970 -340
rect 940 -365 970 -360
rect 1100 -365 1130 -335
rect 1760 -365 1790 -335
rect 1980 1075 2010 1105
rect 1935 730 1965 760
rect 1890 640 1920 670
rect 1935 575 1965 605
rect 1890 -120 1920 -90
rect 1935 -175 1965 -145
rect 1890 -275 1920 -245
rect 2370 1620 2400 1625
rect 2370 1600 2375 1620
rect 2375 1600 2395 1620
rect 2395 1600 2400 1620
rect 2370 1595 2400 1600
rect 2130 1480 2160 1485
rect 2130 1460 2135 1480
rect 2135 1460 2155 1480
rect 2155 1460 2160 1480
rect 2130 1455 2160 1460
rect 2240 1455 2270 1485
rect 2350 1455 2380 1485
rect 2460 1455 2490 1485
rect 2570 1455 2600 1485
rect 2680 1455 2710 1485
rect 2790 1480 2820 1485
rect 2790 1460 2795 1480
rect 2795 1460 2815 1480
rect 2815 1460 2820 1480
rect 2790 1455 2820 1460
rect 3105 1460 3135 1490
rect 2025 870 2055 900
rect 2185 785 2215 815
rect 2295 785 2325 815
rect 2405 785 2435 815
rect 2515 785 2545 815
rect 2625 785 2655 815
rect 2735 785 2765 815
rect 2185 730 2215 760
rect 2625 730 2655 760
rect 2025 685 2055 715
rect 3195 730 3225 760
rect 2460 710 2490 715
rect 2460 690 2465 710
rect 2465 690 2485 710
rect 2485 690 2490 710
rect 2460 685 2490 690
rect 3105 685 3135 715
rect 2130 665 2160 670
rect 2130 645 2135 665
rect 2135 645 2155 665
rect 2155 645 2160 665
rect 2130 640 2160 645
rect 2185 640 2215 670
rect 2295 640 2325 670
rect 2405 640 2435 670
rect 2515 640 2545 670
rect 2625 640 2655 670
rect 2735 640 2765 670
rect 2790 665 2820 670
rect 2790 645 2795 665
rect 2795 645 2815 665
rect 2815 645 2820 665
rect 2790 640 2820 645
rect 2240 385 2270 415
rect 2350 385 2380 415
rect 2460 385 2490 415
rect 2570 385 2600 415
rect 2680 385 2710 415
rect 2925 385 2955 415
rect 2025 310 2055 340
rect 2405 335 2435 340
rect 2405 315 2410 335
rect 2410 315 2430 335
rect 2430 315 2435 335
rect 2405 310 2435 315
rect 2240 235 2270 265
rect 2350 235 2380 265
rect 2460 235 2490 265
rect 2570 235 2600 265
rect 2680 235 2710 265
rect 2880 235 2910 265
rect 2185 -120 2215 -90
rect 2295 -120 2325 -90
rect 2405 -120 2435 -90
rect 2515 -120 2545 -90
rect 2625 -120 2655 -90
rect 2735 -120 2765 -90
rect 2790 -95 2820 -90
rect 2790 -115 2795 -95
rect 2795 -115 2815 -95
rect 2815 -115 2820 -95
rect 2790 -120 2820 -115
rect 2130 -175 2160 -145
rect 2880 -120 2910 -90
rect 3195 320 3225 350
rect 2969 -93 2996 -85
rect 2969 -113 2970 -93
rect 2970 -113 2995 -93
rect 2995 -113 2996 -93
rect 2969 -120 2996 -113
rect 3029 -93 3056 -85
rect 3029 -113 3030 -93
rect 3030 -113 3055 -93
rect 3055 -113 3056 -93
rect 3029 -120 3056 -113
rect 3089 -93 3116 -85
rect 3089 -113 3090 -93
rect 3090 -113 3115 -93
rect 3115 -113 3116 -93
rect 3089 -120 3116 -113
rect 3149 -93 3176 -85
rect 3149 -113 3150 -93
rect 3150 -113 3175 -93
rect 3175 -113 3176 -93
rect 3149 -120 3176 -113
rect 2790 -175 2820 -145
rect 2925 -175 2955 -145
rect 3025 -175 3060 -145
rect 1980 -220 2010 -190
rect 3145 -220 3180 -190
rect 2460 -250 2490 -245
rect 2460 -270 2465 -250
rect 2465 -270 2485 -250
rect 2485 -270 2490 -250
rect 2460 -275 2490 -270
rect 2945 -275 2980 -245
rect 1935 -340 1965 -310
rect 2260 -335 2290 -305
rect 2460 -335 2490 -305
rect 2660 -335 2690 -305
rect 2885 -335 2920 -305
rect 1890 -410 1920 -380
rect 1355 -440 1385 -435
rect 1355 -460 1360 -440
rect 1360 -460 1380 -440
rect 1380 -460 1385 -440
rect 1355 -465 1385 -460
rect 1845 -465 1875 -435
rect 390 -520 420 -490
rect 500 -520 530 -490
rect 610 -520 640 -490
rect 720 -520 750 -490
rect 830 -520 860 -490
rect 940 -520 970 -490
rect 1050 -520 1080 -490
rect 1160 -520 1190 -490
rect 1270 -520 1300 -490
rect 1380 -520 1410 -490
rect 280 -810 310 -805
rect 280 -830 285 -810
rect 285 -830 305 -810
rect 305 -830 310 -810
rect 280 -835 310 -830
rect 335 -835 365 -805
rect 445 -835 475 -805
rect 555 -835 585 -805
rect 665 -835 695 -805
rect 775 -835 805 -805
rect 885 -835 915 -805
rect 995 -835 1025 -805
rect 1105 -835 1135 -805
rect 1215 -835 1245 -805
rect 1325 -835 1355 -805
rect 1435 -810 1465 -805
rect 1435 -830 1440 -810
rect 1440 -830 1460 -810
rect 1460 -830 1465 -810
rect 1435 -835 1465 -830
rect 1935 -835 1965 -805
rect 390 -880 420 -850
rect 500 -880 530 -850
rect 610 -880 640 -850
rect 720 -880 750 -850
rect 830 -880 860 -850
rect 940 -880 970 -850
rect 1050 -880 1080 -850
rect 1160 -880 1190 -850
rect 1270 -880 1300 -850
rect 1380 -880 1410 -850
rect 600 -945 630 -915
rect 710 -945 740 -915
rect 930 -945 960 -915
rect -185 -990 -155 -960
rect 545 -990 575 -960
rect 655 -965 685 -960
rect 655 -985 660 -965
rect 660 -985 680 -965
rect 680 -985 685 -965
rect 655 -990 685 -985
rect 600 -1195 630 -1165
rect 765 -990 795 -960
rect 710 -1195 740 -1165
rect 1100 -965 1130 -960
rect 1100 -985 1105 -965
rect 1105 -985 1125 -965
rect 1125 -985 1130 -965
rect 1100 -990 1130 -985
rect 1270 -990 1300 -960
rect 930 -1195 960 -1165
rect 545 -1240 575 -1210
rect 655 -1240 685 -1210
rect 765 -1240 795 -1210
rect 3195 -335 3225 -305
rect 2889 -387 2916 -380
rect 2889 -407 2890 -387
rect 2890 -407 2915 -387
rect 2915 -407 2916 -387
rect 2889 -415 2916 -407
rect 2949 -387 2976 -380
rect 2949 -407 2950 -387
rect 2950 -407 2975 -387
rect 2975 -407 2976 -387
rect 2949 -415 2976 -407
rect 2160 -1080 2190 -1075
rect 2160 -1100 2165 -1080
rect 2165 -1100 2185 -1080
rect 2185 -1100 2190 -1080
rect 2160 -1105 2190 -1100
rect 2360 -1105 2390 -1075
rect 2560 -1105 2590 -1075
rect 2760 -1080 2790 -1075
rect 2760 -1100 2765 -1080
rect 2765 -1100 2785 -1080
rect 2785 -1100 2790 -1080
rect 2760 -1105 2790 -1100
rect -700 -1285 -670 -1255
rect -275 -1285 -245 -1255
rect 490 -1285 520 -1255
rect 820 -1285 850 -1255
rect 1935 -1285 1965 -1255
rect 2360 -1285 2390 -1255
rect 830 -2455 860 -2425
<< metal2 >>
rect 825 4275 865 4280
rect 825 4245 830 4275
rect 860 4245 865 4275
rect 825 4240 865 4245
rect 210 2780 250 2785
rect 210 2750 215 2780
rect 245 2775 250 2780
rect 620 2780 660 2785
rect 620 2775 625 2780
rect 245 2755 625 2775
rect 245 2750 250 2755
rect 210 2745 250 2750
rect 620 2750 625 2755
rect 655 2750 660 2780
rect 620 2745 660 2750
rect 1030 2780 1070 2785
rect 1030 2750 1035 2780
rect 1065 2775 1070 2780
rect 1440 2780 1480 2785
rect 1440 2775 1445 2780
rect 1065 2755 1445 2775
rect 1065 2750 1070 2755
rect 1030 2745 1070 2750
rect 1440 2750 1445 2755
rect 1475 2750 1480 2780
rect 1440 2745 1480 2750
rect 30 2725 70 2730
rect 30 2695 35 2725
rect 65 2720 70 2725
rect 150 2725 190 2730
rect 150 2720 155 2725
rect 65 2700 155 2720
rect 65 2695 70 2700
rect 30 2690 70 2695
rect 150 2695 155 2700
rect 185 2720 190 2725
rect 210 2725 250 2730
rect 210 2720 215 2725
rect 185 2700 215 2720
rect 185 2695 190 2700
rect 150 2690 190 2695
rect 210 2695 215 2700
rect 245 2695 250 2725
rect 210 2690 250 2695
rect 825 2725 865 2730
rect 825 2695 830 2725
rect 860 2720 865 2725
rect 970 2725 1010 2730
rect 970 2720 975 2725
rect 860 2700 975 2720
rect 860 2695 865 2700
rect 825 2690 865 2695
rect 970 2695 975 2700
rect 1005 2720 1010 2725
rect 1090 2725 1130 2730
rect 1090 2720 1095 2725
rect 1005 2700 1095 2720
rect 1005 2695 1010 2700
rect 970 2690 1010 2695
rect 1090 2695 1095 2700
rect 1125 2720 1130 2725
rect 1150 2725 1190 2730
rect 1150 2720 1155 2725
rect 1125 2700 1155 2720
rect 1125 2695 1130 2700
rect 1090 2690 1130 2695
rect 1150 2695 1155 2700
rect 1185 2695 1190 2725
rect 1150 2690 1190 2695
rect 1440 2725 1480 2730
rect 1440 2695 1445 2725
rect 1475 2720 1480 2725
rect 1500 2725 1540 2730
rect 1500 2720 1505 2725
rect 1475 2700 1505 2720
rect 1475 2695 1480 2700
rect 1440 2690 1480 2695
rect 1500 2695 1505 2700
rect 1535 2720 1540 2725
rect 1620 2725 1660 2730
rect 1620 2720 1625 2725
rect 1535 2700 1625 2720
rect 1535 2695 1540 2700
rect 1500 2690 1540 2695
rect 1620 2695 1625 2700
rect 1655 2695 1660 2725
rect 1620 2690 1660 2695
rect 500 2555 540 2560
rect 500 2525 505 2555
rect 535 2550 540 2555
rect 560 2555 600 2560
rect 560 2550 565 2555
rect 535 2530 565 2550
rect 535 2525 540 2530
rect 500 2520 540 2525
rect 560 2525 565 2530
rect 595 2550 600 2555
rect 680 2555 720 2560
rect 680 2550 685 2555
rect 595 2530 685 2550
rect 595 2525 600 2530
rect 560 2520 600 2525
rect 680 2525 685 2530
rect 715 2550 720 2555
rect 825 2555 865 2560
rect 825 2550 830 2555
rect 715 2530 830 2550
rect 715 2525 720 2530
rect 680 2520 720 2525
rect 825 2525 830 2530
rect 860 2525 865 2555
rect 825 2520 865 2525
rect 75 2305 115 2310
rect 75 2275 80 2305
rect 110 2300 115 2305
rect 139 2305 169 2310
rect 110 2280 139 2300
rect 110 2275 115 2280
rect 75 2270 115 2275
rect 609 2305 639 2310
rect 169 2280 609 2300
rect 139 2270 169 2275
rect 770 2305 810 2310
rect 770 2300 775 2305
rect 639 2280 775 2300
rect 609 2270 639 2275
rect 770 2275 775 2280
rect 805 2300 810 2305
rect 1521 2305 1551 2310
rect 805 2280 1521 2300
rect 805 2275 810 2280
rect 770 2270 810 2275
rect 1521 2270 1551 2275
rect 880 2260 920 2265
rect 880 2230 885 2260
rect 915 2245 920 2260
rect 1045 2250 1085 2255
rect 1045 2245 1050 2250
rect 915 2230 1050 2245
rect 880 2225 1050 2230
rect 1045 2220 1050 2225
rect 1080 2245 1085 2250
rect 1560 2250 1600 2255
rect 1560 2245 1565 2250
rect 1080 2225 1565 2245
rect 1080 2220 1085 2225
rect 1045 2215 1085 2220
rect 1560 2220 1565 2225
rect 1595 2220 1600 2250
rect 1560 2215 1600 2220
rect -805 2205 -765 2210
rect -805 2175 -800 2205
rect -770 2200 -765 2205
rect -235 2205 -195 2210
rect -235 2200 -230 2205
rect -770 2180 -230 2200
rect -770 2175 -765 2180
rect -805 2170 -765 2175
rect -235 2175 -230 2180
rect -200 2200 -195 2205
rect 825 2205 865 2210
rect 825 2200 830 2205
rect -200 2180 830 2200
rect -200 2175 -195 2180
rect -235 2170 -195 2175
rect 825 2175 830 2180
rect 860 2200 865 2205
rect 1885 2205 1925 2210
rect 1885 2200 1890 2205
rect 860 2180 1890 2200
rect 860 2175 865 2180
rect 825 2170 865 2175
rect 1885 2175 1890 2180
rect 1920 2200 1925 2205
rect 2455 2205 2495 2210
rect 2455 2200 2460 2205
rect 1920 2180 2460 2200
rect 1920 2175 1925 2180
rect 1885 2170 1925 2175
rect 2455 2175 2460 2180
rect 2490 2175 2495 2205
rect 2455 2170 2495 2175
rect -1165 2150 -1125 2155
rect -1165 2120 -1160 2150
rect -1130 2145 -1125 2150
rect -1045 2150 -1005 2155
rect -1045 2145 -1040 2150
rect -1130 2125 -1040 2145
rect -1130 2120 -1125 2125
rect -1165 2115 -1125 2120
rect -1045 2120 -1040 2125
rect -1010 2145 -1005 2150
rect -925 2150 -885 2155
rect -925 2145 -920 2150
rect -1010 2125 -920 2145
rect -1010 2120 -1005 2125
rect -1045 2115 -1005 2120
rect -925 2120 -920 2125
rect -890 2145 -885 2150
rect -805 2150 -765 2155
rect -805 2145 -800 2150
rect -890 2125 -800 2145
rect -890 2120 -885 2125
rect -925 2115 -885 2120
rect -805 2120 -800 2125
rect -770 2145 -765 2150
rect -685 2150 -645 2155
rect -685 2145 -680 2150
rect -770 2125 -680 2145
rect -770 2120 -765 2125
rect -805 2115 -765 2120
rect -685 2120 -680 2125
rect -650 2145 -645 2150
rect -565 2150 -525 2155
rect -565 2145 -560 2150
rect -650 2125 -560 2145
rect -650 2120 -645 2125
rect -685 2115 -645 2120
rect -565 2120 -560 2125
rect -530 2145 -525 2150
rect -445 2150 -405 2155
rect -445 2145 -440 2150
rect -530 2125 -440 2145
rect -530 2120 -525 2125
rect -565 2115 -525 2120
rect -445 2120 -440 2125
rect -410 2120 -405 2150
rect -445 2115 -405 2120
rect -280 2150 -240 2155
rect -280 2120 -275 2150
rect -245 2145 -240 2150
rect -40 2150 0 2155
rect -40 2145 -35 2150
rect -245 2125 -35 2145
rect -245 2120 -240 2125
rect -280 2115 -240 2120
rect -40 2120 -35 2125
rect -5 2145 0 2150
rect 80 2150 120 2155
rect 80 2145 85 2150
rect -5 2125 85 2145
rect -5 2120 0 2125
rect -40 2115 0 2120
rect 80 2120 85 2125
rect 115 2145 120 2150
rect 200 2150 240 2155
rect 200 2145 205 2150
rect 115 2125 205 2145
rect 115 2120 120 2125
rect 80 2115 120 2120
rect 200 2120 205 2125
rect 235 2145 240 2150
rect 320 2150 360 2155
rect 320 2145 325 2150
rect 235 2125 325 2145
rect 235 2120 240 2125
rect 200 2115 240 2120
rect 320 2120 325 2125
rect 355 2145 360 2150
rect 440 2150 480 2155
rect 440 2145 445 2150
rect 355 2125 445 2145
rect 355 2120 360 2125
rect 320 2115 360 2120
rect 440 2120 445 2125
rect 475 2145 480 2150
rect 560 2150 600 2155
rect 560 2145 565 2150
rect 475 2125 565 2145
rect 475 2120 480 2125
rect 440 2115 480 2120
rect 560 2120 565 2125
rect 595 2145 600 2150
rect 680 2150 720 2155
rect 680 2145 685 2150
rect 595 2125 685 2145
rect 595 2120 600 2125
rect 560 2115 600 2120
rect 680 2120 685 2125
rect 715 2120 720 2150
rect 680 2115 720 2120
rect 970 2150 1010 2155
rect 970 2120 975 2150
rect 1005 2145 1010 2150
rect 1090 2150 1130 2155
rect 1090 2145 1095 2150
rect 1005 2125 1095 2145
rect 1005 2120 1010 2125
rect 970 2115 1010 2120
rect 1090 2120 1095 2125
rect 1125 2145 1130 2150
rect 1210 2150 1250 2155
rect 1210 2145 1215 2150
rect 1125 2125 1215 2145
rect 1125 2120 1130 2125
rect 1090 2115 1130 2120
rect 1210 2120 1215 2125
rect 1245 2145 1250 2150
rect 1330 2150 1370 2155
rect 1330 2145 1335 2150
rect 1245 2125 1335 2145
rect 1245 2120 1250 2125
rect 1210 2115 1250 2120
rect 1330 2120 1335 2125
rect 1365 2145 1370 2150
rect 1450 2150 1490 2155
rect 1450 2145 1455 2150
rect 1365 2125 1455 2145
rect 1365 2120 1370 2125
rect 1330 2115 1370 2120
rect 1450 2120 1455 2125
rect 1485 2145 1490 2150
rect 1570 2150 1610 2155
rect 1570 2145 1575 2150
rect 1485 2125 1575 2145
rect 1485 2120 1490 2125
rect 1450 2115 1490 2120
rect 1570 2120 1575 2125
rect 1605 2145 1610 2150
rect 1690 2150 1730 2155
rect 1690 2145 1695 2150
rect 1605 2125 1695 2145
rect 1605 2120 1610 2125
rect 1570 2115 1610 2120
rect 1690 2120 1695 2125
rect 1725 2145 1730 2150
rect 1930 2150 1970 2155
rect 1930 2145 1935 2150
rect 1725 2125 1935 2145
rect 1725 2120 1730 2125
rect 1690 2115 1730 2120
rect 1930 2120 1935 2125
rect 1965 2120 1970 2150
rect 1930 2115 1970 2120
rect 2095 2150 2135 2155
rect 2095 2120 2100 2150
rect 2130 2145 2135 2150
rect 2215 2150 2255 2155
rect 2215 2145 2220 2150
rect 2130 2125 2220 2145
rect 2130 2120 2135 2125
rect 2095 2115 2135 2120
rect 2215 2120 2220 2125
rect 2250 2145 2255 2150
rect 2335 2150 2375 2155
rect 2335 2145 2340 2150
rect 2250 2125 2340 2145
rect 2250 2120 2255 2125
rect 2215 2115 2255 2120
rect 2335 2120 2340 2125
rect 2370 2145 2375 2150
rect 2455 2150 2495 2155
rect 2455 2145 2460 2150
rect 2370 2125 2460 2145
rect 2370 2120 2375 2125
rect 2335 2115 2375 2120
rect 2455 2120 2460 2125
rect 2490 2145 2495 2150
rect 2575 2150 2615 2155
rect 2575 2145 2580 2150
rect 2490 2125 2580 2145
rect 2490 2120 2495 2125
rect 2455 2115 2495 2120
rect 2575 2120 2580 2125
rect 2610 2145 2615 2150
rect 2695 2150 2735 2155
rect 2695 2145 2700 2150
rect 2610 2125 2700 2145
rect 2610 2120 2615 2125
rect 2575 2115 2615 2120
rect 2695 2120 2700 2125
rect 2730 2145 2735 2150
rect 2815 2150 2855 2155
rect 2815 2145 2820 2150
rect 2730 2125 2820 2145
rect 2730 2120 2735 2125
rect 2695 2115 2735 2120
rect 2815 2120 2820 2125
rect 2850 2120 2855 2150
rect 2815 2115 2855 2120
rect -1105 1730 -1065 1735
rect -1105 1700 -1100 1730
rect -1070 1725 -1065 1730
rect -985 1730 -945 1735
rect -985 1725 -980 1730
rect -1070 1705 -980 1725
rect -1070 1700 -1065 1705
rect -1105 1695 -1065 1700
rect -985 1700 -980 1705
rect -950 1725 -945 1730
rect -865 1730 -825 1735
rect -865 1725 -860 1730
rect -950 1705 -860 1725
rect -950 1700 -945 1705
rect -985 1695 -945 1700
rect -865 1700 -860 1705
rect -830 1725 -825 1730
rect -745 1730 -705 1735
rect -745 1725 -740 1730
rect -830 1705 -740 1725
rect -830 1700 -825 1705
rect -865 1695 -825 1700
rect -745 1700 -740 1705
rect -710 1725 -705 1730
rect -625 1730 -585 1735
rect -625 1725 -620 1730
rect -710 1705 -620 1725
rect -710 1700 -705 1705
rect -745 1695 -705 1700
rect -625 1700 -620 1705
rect -590 1725 -585 1730
rect -505 1730 -465 1735
rect -505 1725 -500 1730
rect -590 1705 -500 1725
rect -590 1700 -585 1705
rect -625 1695 -585 1700
rect -505 1700 -500 1705
rect -470 1725 -465 1730
rect -280 1730 -240 1735
rect -280 1725 -275 1730
rect -470 1705 -275 1725
rect -470 1700 -465 1705
rect -505 1695 -465 1700
rect -280 1700 -275 1705
rect -245 1700 -240 1730
rect -280 1695 -240 1700
rect 20 1730 60 1735
rect 20 1700 25 1730
rect 55 1725 60 1730
rect 140 1730 180 1735
rect 140 1725 145 1730
rect 55 1705 145 1725
rect 55 1700 60 1705
rect 20 1695 60 1700
rect 140 1700 145 1705
rect 175 1725 180 1730
rect 260 1730 300 1735
rect 260 1725 265 1730
rect 175 1705 265 1725
rect 175 1700 180 1705
rect 140 1695 180 1700
rect 260 1700 265 1705
rect 295 1725 300 1730
rect 380 1730 420 1735
rect 380 1725 385 1730
rect 295 1705 385 1725
rect 295 1700 300 1705
rect 260 1695 300 1700
rect 380 1700 385 1705
rect 415 1725 420 1730
rect 500 1730 540 1735
rect 500 1725 505 1730
rect 415 1705 505 1725
rect 415 1700 420 1705
rect 380 1695 420 1700
rect 500 1700 505 1705
rect 535 1725 540 1730
rect 620 1730 660 1735
rect 620 1725 625 1730
rect 535 1705 625 1725
rect 535 1700 540 1705
rect 500 1695 540 1700
rect 620 1700 625 1705
rect 655 1700 660 1730
rect 620 1695 660 1700
rect 1030 1730 1070 1735
rect 1030 1700 1035 1730
rect 1065 1725 1070 1730
rect 1150 1730 1190 1735
rect 1150 1725 1155 1730
rect 1065 1705 1155 1725
rect 1065 1700 1070 1705
rect 1030 1695 1070 1700
rect 1150 1700 1155 1705
rect 1185 1725 1190 1730
rect 1270 1730 1310 1735
rect 1270 1725 1275 1730
rect 1185 1705 1275 1725
rect 1185 1700 1190 1705
rect 1150 1695 1190 1700
rect 1270 1700 1275 1705
rect 1305 1725 1310 1730
rect 1390 1730 1430 1735
rect 1390 1725 1395 1730
rect 1305 1705 1395 1725
rect 1305 1700 1310 1705
rect 1270 1695 1310 1700
rect 1390 1700 1395 1705
rect 1425 1725 1430 1730
rect 1510 1730 1550 1735
rect 1510 1725 1515 1730
rect 1425 1705 1515 1725
rect 1425 1700 1430 1705
rect 1390 1695 1430 1700
rect 1510 1700 1515 1705
rect 1545 1725 1550 1730
rect 1630 1730 1670 1735
rect 1630 1725 1635 1730
rect 1545 1705 1635 1725
rect 1545 1700 1550 1705
rect 1510 1695 1550 1700
rect 1630 1700 1635 1705
rect 1665 1700 1670 1730
rect 1630 1695 1670 1700
rect 1930 1730 1970 1735
rect 1930 1700 1935 1730
rect 1965 1725 1970 1730
rect 2155 1730 2195 1735
rect 2155 1725 2160 1730
rect 1965 1705 2160 1725
rect 1965 1700 1970 1705
rect 1930 1695 1970 1700
rect 2155 1700 2160 1705
rect 2190 1725 2195 1730
rect 2275 1730 2315 1735
rect 2275 1725 2280 1730
rect 2190 1705 2280 1725
rect 2190 1700 2195 1705
rect 2155 1695 2195 1700
rect 2275 1700 2280 1705
rect 2310 1725 2315 1730
rect 2395 1730 2435 1735
rect 2395 1725 2400 1730
rect 2310 1705 2400 1725
rect 2310 1700 2315 1705
rect 2275 1695 2315 1700
rect 2395 1700 2400 1705
rect 2430 1725 2435 1730
rect 2515 1730 2555 1735
rect 2515 1725 2520 1730
rect 2430 1705 2520 1725
rect 2430 1700 2435 1705
rect 2395 1695 2435 1700
rect 2515 1700 2520 1705
rect 2550 1725 2555 1730
rect 2635 1730 2675 1735
rect 2635 1725 2640 1730
rect 2550 1705 2640 1725
rect 2550 1700 2555 1705
rect 2515 1695 2555 1700
rect 2635 1700 2640 1705
rect 2670 1725 2675 1730
rect 2755 1730 2795 1735
rect 2755 1725 2760 1730
rect 2670 1705 2760 1725
rect 2670 1700 2675 1705
rect 2635 1695 2675 1700
rect 2755 1700 2760 1705
rect 2790 1700 2795 1730
rect 2755 1695 2795 1700
rect -370 1670 -330 1675
rect -370 1640 -365 1670
rect -335 1665 -330 1670
rect 260 1670 300 1675
rect 260 1665 265 1670
rect -335 1645 265 1665
rect -335 1640 -330 1645
rect -370 1635 -330 1640
rect 260 1640 265 1645
rect 295 1640 300 1670
rect 260 1635 300 1640
rect 410 1670 450 1675
rect 410 1640 415 1670
rect 445 1665 450 1670
rect 780 1670 820 1675
rect 780 1665 785 1670
rect 445 1645 785 1665
rect 445 1640 450 1645
rect 410 1635 450 1640
rect 780 1640 785 1645
rect 815 1665 820 1670
rect 1240 1670 1280 1675
rect 1240 1665 1245 1670
rect 815 1645 1245 1665
rect 815 1640 820 1645
rect 780 1635 820 1640
rect 1240 1640 1245 1645
rect 1275 1640 1280 1670
rect 1240 1635 1280 1640
rect 1390 1670 1430 1675
rect 1390 1640 1395 1670
rect 1425 1665 1430 1670
rect 2020 1670 2060 1675
rect 2020 1665 2025 1670
rect 1425 1645 2025 1665
rect 1425 1640 1430 1645
rect 1390 1635 1430 1640
rect 2020 1640 2025 1645
rect 2055 1640 2060 1670
rect 2020 1635 2060 1640
rect -715 1625 -675 1630
rect -715 1595 -710 1625
rect -680 1620 -675 1625
rect 870 1620 875 1630
rect -680 1600 875 1620
rect 905 1620 910 1630
rect 2365 1625 2405 1630
rect 2365 1620 2370 1625
rect 905 1600 2370 1620
rect -680 1595 -675 1600
rect -715 1590 -675 1595
rect 2365 1595 2370 1600
rect 2400 1595 2405 1625
rect 2365 1590 2405 1595
rect 455 1565 495 1570
rect -1450 1540 -1410 1545
rect -1450 1510 -1445 1540
rect -1415 1510 -1410 1540
rect 455 1535 460 1565
rect 490 1560 495 1565
rect 620 1565 660 1570
rect 620 1560 625 1565
rect 490 1540 625 1560
rect 490 1535 495 1540
rect 455 1530 495 1535
rect 620 1535 625 1540
rect 655 1560 660 1565
rect 785 1565 825 1570
rect 785 1560 790 1565
rect 655 1540 790 1560
rect 655 1535 660 1540
rect 620 1530 660 1535
rect 785 1535 790 1540
rect 820 1560 825 1565
rect 865 1565 905 1570
rect 865 1560 870 1565
rect 820 1540 870 1560
rect 820 1535 825 1540
rect 785 1530 825 1535
rect 865 1535 870 1540
rect 900 1560 905 1565
rect 1030 1565 1070 1570
rect 1030 1560 1035 1565
rect 900 1540 1035 1560
rect 900 1535 905 1540
rect 865 1530 905 1535
rect 1030 1535 1035 1540
rect 1065 1560 1070 1565
rect 1195 1565 1235 1570
rect 1195 1560 1200 1565
rect 1065 1540 1200 1560
rect 1065 1535 1070 1540
rect 1030 1530 1070 1535
rect 1195 1535 1200 1540
rect 1230 1560 1235 1565
rect 1885 1565 1925 1570
rect 1885 1560 1890 1565
rect 1230 1540 1890 1560
rect 1230 1535 1235 1540
rect 1195 1530 1235 1535
rect 1885 1535 1890 1540
rect 1920 1535 1925 1565
rect 1885 1530 1925 1535
rect -1450 1505 -1410 1510
rect 565 1520 605 1525
rect 565 1490 570 1520
rect 600 1515 605 1520
rect 675 1520 715 1525
rect 675 1515 680 1520
rect 600 1495 680 1515
rect 600 1490 605 1495
rect -1135 1485 -1095 1490
rect -1135 1455 -1130 1485
rect -1100 1480 -1095 1485
rect -1025 1485 -985 1490
rect -1025 1480 -1020 1485
rect -1100 1460 -1020 1480
rect -1100 1455 -1095 1460
rect -1135 1450 -1095 1455
rect -1025 1455 -1020 1460
rect -990 1480 -985 1485
rect -915 1485 -875 1490
rect -915 1480 -910 1485
rect -990 1460 -910 1480
rect -990 1455 -985 1460
rect -1025 1450 -985 1455
rect -915 1455 -910 1460
rect -880 1480 -875 1485
rect -805 1485 -765 1490
rect -805 1480 -800 1485
rect -880 1460 -800 1480
rect -880 1455 -875 1460
rect -915 1450 -875 1455
rect -805 1455 -800 1460
rect -770 1480 -765 1485
rect -695 1485 -655 1490
rect -695 1480 -690 1485
rect -770 1460 -690 1480
rect -770 1455 -765 1460
rect -805 1450 -765 1455
rect -695 1455 -690 1460
rect -660 1480 -655 1485
rect -585 1485 -545 1490
rect -585 1480 -580 1485
rect -660 1460 -580 1480
rect -660 1455 -655 1460
rect -695 1450 -655 1455
rect -585 1455 -580 1460
rect -550 1480 -545 1485
rect -475 1485 -435 1490
rect -475 1480 -470 1485
rect -550 1460 -470 1480
rect -550 1455 -545 1460
rect -585 1450 -545 1455
rect -475 1455 -470 1460
rect -440 1480 -435 1485
rect -235 1485 -195 1490
rect 565 1485 605 1490
rect 675 1490 680 1495
rect 710 1490 715 1520
rect 675 1485 715 1490
rect 975 1520 1015 1525
rect 975 1490 980 1520
rect 1010 1515 1015 1520
rect 1085 1520 1125 1525
rect 1085 1515 1090 1520
rect 1010 1495 1090 1515
rect 1010 1490 1015 1495
rect 975 1485 1015 1490
rect 1085 1490 1090 1495
rect 1120 1490 1125 1520
rect 3100 1490 3140 1495
rect 1085 1485 1125 1490
rect 1885 1485 1925 1490
rect -235 1480 -230 1485
rect -440 1460 -230 1480
rect -440 1455 -435 1460
rect -475 1450 -435 1455
rect -235 1455 -230 1460
rect -200 1455 -195 1485
rect -235 1450 -195 1455
rect 1885 1455 1890 1485
rect 1920 1480 1925 1485
rect 2125 1485 2165 1490
rect 2125 1480 2130 1485
rect 1920 1460 2130 1480
rect 1920 1455 1925 1460
rect 1885 1450 1925 1455
rect 2125 1455 2130 1460
rect 2160 1480 2165 1485
rect 2235 1485 2275 1490
rect 2235 1480 2240 1485
rect 2160 1460 2240 1480
rect 2160 1455 2165 1460
rect 2125 1450 2165 1455
rect 2235 1455 2240 1460
rect 2270 1480 2275 1485
rect 2345 1485 2385 1490
rect 2345 1480 2350 1485
rect 2270 1460 2350 1480
rect 2270 1455 2275 1460
rect 2235 1450 2275 1455
rect 2345 1455 2350 1460
rect 2380 1480 2385 1485
rect 2455 1485 2495 1490
rect 2455 1480 2460 1485
rect 2380 1460 2460 1480
rect 2380 1455 2385 1460
rect 2345 1450 2385 1455
rect 2455 1455 2460 1460
rect 2490 1480 2495 1485
rect 2565 1485 2605 1490
rect 2565 1480 2570 1485
rect 2490 1460 2570 1480
rect 2490 1455 2495 1460
rect 2455 1450 2495 1455
rect 2565 1455 2570 1460
rect 2600 1480 2605 1485
rect 2675 1485 2715 1490
rect 2675 1480 2680 1485
rect 2600 1460 2680 1480
rect 2600 1455 2605 1460
rect 2565 1450 2605 1455
rect 2675 1455 2680 1460
rect 2710 1480 2715 1485
rect 2785 1485 2825 1490
rect 2785 1480 2790 1485
rect 2710 1460 2790 1480
rect 2710 1455 2715 1460
rect 2675 1450 2715 1455
rect 2785 1455 2790 1460
rect 2820 1455 2825 1485
rect 3100 1460 3105 1490
rect 3135 1460 3140 1490
rect 3100 1455 3140 1460
rect 2785 1450 2825 1455
rect 620 1215 660 1220
rect 620 1210 625 1215
rect 495 1205 625 1210
rect 495 1175 500 1205
rect 530 1190 625 1205
rect 530 1175 535 1190
rect 620 1185 625 1190
rect 655 1210 660 1215
rect 1030 1215 1070 1220
rect 1030 1210 1035 1215
rect 655 1205 1035 1210
rect 655 1190 750 1205
rect 655 1185 660 1190
rect 620 1180 660 1185
rect 495 1170 535 1175
rect 745 1175 750 1190
rect 780 1190 1035 1205
rect 780 1175 785 1190
rect 1030 1185 1035 1190
rect 1065 1210 1070 1215
rect 1065 1190 1075 1210
rect 1065 1185 1070 1190
rect 1030 1180 1070 1185
rect 745 1170 785 1175
rect 545 1155 585 1160
rect 545 1150 550 1155
rect 310 1130 550 1150
rect 545 1125 550 1130
rect 580 1150 585 1155
rect 1095 1155 1135 1160
rect 1095 1150 1100 1155
rect 580 1130 1100 1150
rect 580 1125 585 1130
rect 545 1120 585 1125
rect 1095 1125 1100 1130
rect 1130 1125 1135 1155
rect 1095 1120 1135 1125
rect -325 1105 -285 1110
rect -325 1075 -320 1105
rect -290 1100 -285 1105
rect 690 1105 730 1110
rect 690 1100 695 1105
rect -290 1080 695 1100
rect -290 1075 -285 1080
rect -325 1070 -285 1075
rect 690 1075 695 1080
rect 725 1100 730 1105
rect 965 1105 1005 1110
rect 965 1100 970 1105
rect 725 1080 970 1100
rect 725 1075 730 1080
rect 690 1070 730 1075
rect 965 1075 970 1080
rect 1000 1100 1005 1105
rect 1975 1105 2015 1110
rect 1975 1100 1980 1105
rect 1000 1080 1980 1100
rect 1000 1075 1005 1080
rect 965 1070 1005 1075
rect 1975 1075 1980 1080
rect 2010 1075 2015 1105
rect 1975 1070 2015 1075
rect 795 1060 835 1065
rect 795 1030 800 1060
rect 830 1055 835 1060
rect 905 1060 945 1065
rect 905 1055 910 1060
rect 830 1035 910 1055
rect 830 1030 835 1035
rect 795 1025 835 1030
rect 905 1030 910 1035
rect 940 1030 945 1060
rect 905 1025 945 1030
rect 1155 1010 1195 1015
rect 795 1005 835 1010
rect 795 975 800 1005
rect 830 975 835 1005
rect 795 970 835 975
rect 880 1005 920 1010
rect 880 975 885 1005
rect 915 1000 920 1005
rect 1155 1000 1160 1010
rect 915 980 1160 1000
rect 1190 1005 1195 1010
rect 1840 1010 1880 1015
rect 1840 1005 1845 1010
rect 1190 985 1845 1005
rect 1190 980 1195 985
rect 915 975 920 980
rect 1155 975 1195 980
rect 1840 980 1845 985
rect 1875 980 1880 1010
rect 1840 975 1880 980
rect 880 970 920 975
rect -190 950 -150 955
rect -190 920 -185 950
rect -155 945 -150 950
rect 120 950 150 955
rect -155 925 120 945
rect -155 920 -150 925
rect -190 915 -150 920
rect 1540 950 1570 955
rect 150 925 1540 945
rect 120 915 150 920
rect 1540 915 1570 920
rect -370 900 -330 905
rect -370 870 -365 900
rect -335 895 -330 900
rect -50 900 -10 905
rect -50 895 -45 900
rect -335 875 -45 895
rect -335 870 -330 875
rect -370 865 -330 870
rect -50 870 -45 875
rect -15 895 -10 900
rect 60 900 100 905
rect 60 895 65 900
rect -15 875 65 895
rect -15 870 -10 875
rect -50 865 -10 870
rect 60 870 65 875
rect 95 895 100 900
rect 170 900 210 905
rect 170 895 175 900
rect 95 875 175 895
rect 95 870 100 875
rect 60 865 100 870
rect 170 870 175 875
rect 205 895 210 900
rect 280 900 320 905
rect 280 895 285 900
rect 205 875 285 895
rect 205 870 210 875
rect 170 865 210 870
rect 280 870 285 875
rect 315 895 320 900
rect 390 900 430 905
rect 390 895 395 900
rect 315 875 395 895
rect 315 870 320 875
rect 280 865 320 870
rect 390 870 395 875
rect 425 895 430 900
rect 500 900 540 905
rect 500 895 505 900
rect 425 875 505 895
rect 425 870 430 875
rect 390 865 430 870
rect 500 870 505 875
rect 535 870 540 900
rect 500 865 540 870
rect 1150 900 1190 905
rect 1150 870 1155 900
rect 1185 895 1190 900
rect 1260 900 1300 905
rect 1260 895 1265 900
rect 1185 875 1265 895
rect 1185 870 1190 875
rect 1150 865 1190 870
rect 1260 870 1265 875
rect 1295 895 1300 900
rect 1370 900 1410 905
rect 1370 895 1375 900
rect 1295 875 1375 895
rect 1295 870 1300 875
rect 1260 865 1300 870
rect 1370 870 1375 875
rect 1405 895 1410 900
rect 1480 900 1520 905
rect 1480 895 1485 900
rect 1405 875 1485 895
rect 1405 870 1410 875
rect 1370 865 1410 870
rect 1480 870 1485 875
rect 1515 895 1520 900
rect 1590 900 1630 905
rect 1590 895 1595 900
rect 1515 875 1595 895
rect 1515 870 1520 875
rect 1480 865 1520 870
rect 1590 870 1595 875
rect 1625 895 1630 900
rect 1700 900 1740 905
rect 1700 895 1705 900
rect 1625 875 1705 895
rect 1625 870 1630 875
rect 1590 865 1630 870
rect 1700 870 1705 875
rect 1735 895 1740 900
rect 2020 900 2060 905
rect 2020 895 2025 900
rect 1735 875 2025 895
rect 1735 870 1740 875
rect 1700 865 1740 870
rect 2020 870 2025 875
rect 2055 870 2060 900
rect 2020 865 2060 870
rect -1080 815 -1040 820
rect -1080 785 -1075 815
rect -1045 810 -1040 815
rect -970 815 -930 820
rect -970 810 -965 815
rect -1045 790 -965 810
rect -1045 785 -1040 790
rect -1080 780 -1040 785
rect -970 785 -965 790
rect -935 810 -930 815
rect -860 815 -820 820
rect -860 810 -855 815
rect -935 790 -855 810
rect -935 785 -930 790
rect -970 780 -930 785
rect -860 785 -855 790
rect -825 810 -820 815
rect -750 815 -710 820
rect -750 810 -745 815
rect -825 790 -745 810
rect -825 785 -820 790
rect -860 780 -820 785
rect -750 785 -745 790
rect -715 810 -710 815
rect -640 815 -600 820
rect -640 810 -635 815
rect -715 790 -635 810
rect -715 785 -710 790
rect -750 780 -710 785
rect -640 785 -635 790
rect -605 810 -600 815
rect -530 815 -490 820
rect -530 810 -525 815
rect -605 790 -525 810
rect -605 785 -600 790
rect -640 780 -600 785
rect -530 785 -525 790
rect -495 785 -490 815
rect -530 780 -490 785
rect 2180 815 2220 820
rect 2180 785 2185 815
rect 2215 810 2220 815
rect 2290 815 2330 820
rect 2290 810 2295 815
rect 2215 790 2295 810
rect 2215 785 2220 790
rect 2180 780 2220 785
rect 2290 785 2295 790
rect 2325 810 2330 815
rect 2400 815 2440 820
rect 2400 810 2405 815
rect 2325 790 2405 810
rect 2325 785 2330 790
rect 2290 780 2330 785
rect 2400 785 2405 790
rect 2435 810 2440 815
rect 2510 815 2550 820
rect 2510 810 2515 815
rect 2435 790 2515 810
rect 2435 785 2440 790
rect 2400 780 2440 785
rect 2510 785 2515 790
rect 2545 810 2550 815
rect 2620 815 2660 820
rect 2620 810 2625 815
rect 2545 790 2625 810
rect 2545 785 2550 790
rect 2510 780 2550 785
rect 2620 785 2625 790
rect 2655 810 2660 815
rect 2730 815 2770 820
rect 2730 810 2735 815
rect 2655 790 2735 810
rect 2655 785 2660 790
rect 2620 780 2660 785
rect 2730 785 2735 790
rect 2765 785 2770 815
rect 2730 780 2770 785
rect -280 770 -240 775
rect -1540 760 -1500 765
rect -1540 730 -1535 760
rect -1505 755 -1500 760
rect -970 760 -930 765
rect -970 755 -965 760
rect -1505 735 -965 755
rect -1505 730 -1500 735
rect -1540 725 -1500 730
rect -970 730 -965 735
rect -935 730 -930 760
rect -970 725 -930 730
rect -530 760 -490 765
rect -530 730 -525 760
rect -495 755 -490 760
rect -280 755 -275 770
rect -495 740 -275 755
rect -245 740 -240 770
rect -495 735 -240 740
rect 1930 760 1970 765
rect -495 730 -490 735
rect -530 725 -490 730
rect 1930 730 1935 760
rect 1965 755 1970 760
rect 2180 760 2220 765
rect 2180 755 2185 760
rect 1965 735 2185 755
rect 1965 730 1970 735
rect 1930 725 1970 730
rect 2180 730 2185 735
rect 2215 730 2220 760
rect 2180 725 2220 730
rect 2620 760 2660 765
rect 2620 730 2625 760
rect 2655 755 2660 760
rect 3190 760 3230 765
rect 3190 755 3195 760
rect 2655 735 3195 755
rect 2655 730 2660 735
rect 2620 725 2660 730
rect 3190 730 3195 735
rect 3225 730 3230 760
rect 3190 725 3230 730
rect -1450 715 -1410 720
rect -1450 685 -1445 715
rect -1415 710 -1410 715
rect -805 715 -765 720
rect -805 710 -800 715
rect -1415 690 -800 710
rect -1415 685 -1410 690
rect -1450 680 -1410 685
rect -805 685 -800 690
rect -770 710 -765 715
rect -370 715 -330 720
rect -370 710 -365 715
rect -770 690 -365 710
rect -770 685 -765 690
rect -805 680 -765 685
rect -370 685 -365 690
rect -335 685 -330 715
rect 2020 715 2060 720
rect 2020 685 2025 715
rect 2055 710 2060 715
rect 2455 715 2495 720
rect 2455 710 2460 715
rect 2055 690 2460 710
rect 2055 685 2060 690
rect -370 680 -330 685
rect -1135 670 -1095 675
rect -1135 640 -1130 670
rect -1100 640 -1095 670
rect -1135 635 -1095 640
rect -1080 670 -1040 675
rect -1080 640 -1075 670
rect -1045 665 -1040 670
rect -970 670 -930 675
rect -970 665 -965 670
rect -1045 645 -965 665
rect -1045 640 -1040 645
rect -1080 635 -1040 640
rect -970 640 -965 645
rect -935 665 -930 670
rect -860 670 -820 675
rect -860 665 -855 670
rect -935 645 -855 665
rect -935 640 -930 645
rect -970 635 -930 640
rect -860 640 -855 645
rect -825 665 -820 670
rect -750 670 -710 675
rect -750 665 -745 670
rect -825 645 -745 665
rect -825 640 -820 645
rect -860 635 -820 640
rect -750 640 -745 645
rect -715 665 -710 670
rect -640 670 -600 675
rect -640 665 -635 670
rect -715 645 -635 665
rect -715 640 -710 645
rect -750 635 -710 640
rect -640 640 -635 645
rect -605 665 -600 670
rect -530 670 -490 675
rect -530 665 -525 670
rect -605 645 -525 665
rect -605 640 -600 645
rect -640 635 -600 640
rect -530 640 -525 645
rect -495 640 -490 670
rect -530 635 -490 640
rect -475 670 -435 675
rect -475 640 -470 670
rect -440 665 -435 670
rect -235 670 -195 675
rect -235 665 -230 670
rect -440 645 -230 665
rect -440 640 -435 645
rect -475 635 -435 640
rect -235 640 -230 645
rect -200 640 -195 670
rect 5 655 10 685
rect 40 680 45 685
rect 115 680 120 685
rect 40 660 120 680
rect 40 655 45 660
rect 115 655 120 660
rect 150 680 155 685
rect 225 680 230 685
rect 150 660 230 680
rect 150 655 155 660
rect 225 655 230 660
rect 260 680 265 685
rect 335 680 340 685
rect 260 660 340 680
rect 260 655 265 660
rect 335 655 340 660
rect 370 680 375 685
rect 445 680 450 685
rect 370 660 450 680
rect 370 655 375 660
rect 395 655 425 660
rect 445 655 450 660
rect 480 655 485 685
rect 1205 655 1210 685
rect 1240 680 1245 685
rect 1315 680 1320 685
rect 1240 660 1320 680
rect 1240 655 1245 660
rect 1315 655 1320 660
rect 1350 680 1355 685
rect 1425 680 1430 685
rect 1350 660 1430 680
rect 1350 655 1355 660
rect 1425 655 1430 660
rect 1460 680 1465 685
rect 1535 680 1540 685
rect 1460 660 1540 680
rect 1460 655 1465 660
rect 1535 655 1540 660
rect 1570 680 1575 685
rect 1645 680 1650 685
rect 1570 660 1650 680
rect 1570 655 1575 660
rect 1645 655 1650 660
rect 1680 655 1685 685
rect 2020 680 2060 685
rect 2455 685 2460 690
rect 2490 710 2495 715
rect 3100 715 3140 720
rect 3100 710 3105 715
rect 2490 690 3105 710
rect 2490 685 2495 690
rect 2455 680 2495 685
rect 3100 685 3105 690
rect 3135 685 3140 715
rect 3100 680 3140 685
rect 1885 670 1925 675
rect 1885 640 1890 670
rect 1920 665 1925 670
rect 2125 670 2165 675
rect 2125 665 2130 670
rect 1920 645 2130 665
rect 1920 640 1925 645
rect -235 635 -195 640
rect -50 610 -45 640
rect -15 635 -10 640
rect 60 635 65 640
rect -15 615 65 635
rect -15 610 -10 615
rect 60 610 65 615
rect 95 635 100 640
rect 170 635 175 640
rect 95 615 175 635
rect 95 610 100 615
rect 170 610 175 615
rect 205 635 210 640
rect 280 635 285 640
rect 205 615 285 635
rect 205 610 210 615
rect 280 610 285 615
rect 315 635 320 640
rect 390 635 395 640
rect 315 615 395 635
rect 315 610 320 615
rect 390 610 395 615
rect 425 635 430 640
rect 500 635 505 640
rect 425 615 505 635
rect 425 610 430 615
rect 500 610 505 615
rect 535 610 540 640
rect 1150 610 1155 640
rect 1185 635 1190 640
rect 1260 635 1265 640
rect 1185 615 1265 635
rect 1185 610 1190 615
rect 1260 610 1265 615
rect 1295 635 1300 640
rect 1370 635 1375 640
rect 1295 615 1375 635
rect 1295 610 1300 615
rect 1370 610 1375 615
rect 1405 635 1410 640
rect 1480 635 1485 640
rect 1405 615 1485 635
rect 1405 610 1410 615
rect 1480 610 1485 615
rect 1515 635 1520 640
rect 1590 635 1595 640
rect 1515 615 1595 635
rect 1515 610 1520 615
rect 1590 610 1595 615
rect 1625 635 1630 640
rect 1700 635 1705 640
rect 1625 615 1705 635
rect 1625 610 1630 615
rect 1700 610 1705 615
rect 1735 610 1740 640
rect 1885 635 1925 640
rect 2125 640 2130 645
rect 2160 640 2165 670
rect 2125 635 2165 640
rect 2180 670 2220 675
rect 2180 640 2185 670
rect 2215 665 2220 670
rect 2290 670 2330 675
rect 2290 665 2295 670
rect 2215 645 2295 665
rect 2215 640 2220 645
rect 2180 635 2220 640
rect 2290 640 2295 645
rect 2325 665 2330 670
rect 2400 670 2440 675
rect 2400 665 2405 670
rect 2325 645 2405 665
rect 2325 640 2330 645
rect 2290 635 2330 640
rect 2400 640 2405 645
rect 2435 665 2440 670
rect 2510 670 2550 675
rect 2510 665 2515 670
rect 2435 645 2515 665
rect 2435 640 2440 645
rect 2400 635 2440 640
rect 2510 640 2515 645
rect 2545 665 2550 670
rect 2620 670 2660 675
rect 2620 665 2625 670
rect 2545 645 2625 665
rect 2545 640 2550 645
rect 2510 635 2550 640
rect 2620 640 2625 645
rect 2655 665 2660 670
rect 2730 670 2770 675
rect 2730 665 2735 670
rect 2655 645 2735 665
rect 2655 640 2660 645
rect 2620 635 2660 640
rect 2730 640 2735 645
rect 2765 640 2770 670
rect 2730 635 2770 640
rect 2785 670 2825 675
rect 2785 640 2790 670
rect 2820 640 2825 670
rect 2785 635 2825 640
rect -105 605 -65 610
rect -105 575 -100 605
rect -70 590 -65 605
rect 555 605 595 610
rect 555 590 560 605
rect -70 575 560 590
rect 590 600 595 605
rect 715 605 755 610
rect 715 600 720 605
rect 590 580 720 600
rect 590 575 595 580
rect -105 570 595 575
rect 715 575 720 580
rect 750 600 755 605
rect 825 605 865 610
rect 825 600 830 605
rect 750 580 830 600
rect 750 575 755 580
rect 715 570 755 575
rect 825 575 830 580
rect 860 600 865 605
rect 935 605 975 610
rect 935 600 940 605
rect 860 580 940 600
rect 860 575 865 580
rect 825 570 865 575
rect 935 575 940 580
rect 970 600 975 605
rect 1095 605 1135 610
rect 1095 600 1100 605
rect 970 580 1100 600
rect 970 575 975 580
rect 935 570 975 575
rect 1095 575 1100 580
rect 1130 590 1135 605
rect 1755 605 1795 610
rect 1755 590 1760 605
rect 1130 575 1760 590
rect 1790 600 1795 605
rect 1930 605 1970 610
rect 1930 600 1935 605
rect 1790 580 1935 600
rect 1790 575 1795 580
rect 1095 570 1795 575
rect 1930 575 1935 580
rect 1965 575 1970 605
rect 1930 570 1970 575
rect 145 550 175 555
rect -105 525 145 545
rect 795 550 825 555
rect 175 525 795 545
rect 145 515 175 520
rect 795 515 825 520
rect 865 550 895 555
rect 1515 550 1545 555
rect 895 525 1515 545
rect 865 515 895 520
rect 1545 525 1795 545
rect 1515 515 1545 520
rect 230 475 260 480
rect -50 465 -10 470
rect -50 435 -45 465
rect -15 460 -10 465
rect 60 465 100 470
rect 60 460 65 465
rect -15 440 65 460
rect -15 435 -10 440
rect -50 430 -10 435
rect 60 435 65 440
rect 95 460 100 465
rect 170 465 210 470
rect 170 460 175 465
rect 95 440 175 460
rect 95 435 100 440
rect 60 430 100 435
rect 170 435 175 440
rect 205 460 210 465
rect 205 445 230 460
rect 1430 475 1460 480
rect 280 465 320 470
rect 280 460 285 465
rect 260 445 285 460
rect 205 440 285 445
rect 205 435 210 440
rect 170 430 210 435
rect 280 435 285 440
rect 315 460 320 465
rect 390 465 430 470
rect 390 460 395 465
rect 315 440 395 460
rect 315 435 320 440
rect 280 430 320 435
rect 390 435 395 440
rect 425 460 430 465
rect 500 465 540 470
rect 500 460 505 465
rect 425 440 505 460
rect 425 435 430 440
rect 390 430 430 435
rect 500 435 505 440
rect 535 435 540 465
rect 500 430 540 435
rect 1150 465 1190 470
rect 1150 435 1155 465
rect 1185 460 1190 465
rect 1260 465 1300 470
rect 1260 460 1265 465
rect 1185 440 1265 460
rect 1185 435 1190 440
rect 1150 430 1190 435
rect 1260 435 1265 440
rect 1295 460 1300 465
rect 1370 465 1410 470
rect 1370 460 1375 465
rect 1295 440 1375 460
rect 1295 435 1300 440
rect 1260 430 1300 435
rect 1370 435 1375 440
rect 1405 460 1410 465
rect 1405 445 1430 460
rect 1480 465 1520 470
rect 1480 460 1485 465
rect 1460 445 1485 460
rect 1405 440 1485 445
rect 1405 435 1410 440
rect 1370 430 1410 435
rect 1480 435 1485 440
rect 1515 460 1520 465
rect 1590 465 1630 470
rect 1590 460 1595 465
rect 1515 440 1595 460
rect 1515 435 1520 440
rect 1480 430 1520 435
rect 1590 435 1595 440
rect 1625 460 1630 465
rect 1700 465 1740 470
rect 1700 460 1705 465
rect 1625 440 1705 460
rect 1625 435 1630 440
rect 1590 430 1630 435
rect 1700 435 1705 440
rect 1735 435 1740 465
rect 1700 430 1740 435
rect -1270 415 -1230 420
rect -1270 385 -1265 415
rect -1235 410 -1230 415
rect -1025 415 -985 420
rect -1025 410 -1020 415
rect -1235 390 -1020 410
rect -1235 385 -1230 390
rect -1270 380 -1230 385
rect -1025 385 -1020 390
rect -990 410 -985 415
rect -915 415 -875 420
rect -915 410 -910 415
rect -990 390 -910 410
rect -990 385 -985 390
rect -1025 380 -985 385
rect -915 385 -910 390
rect -880 410 -875 415
rect -805 415 -765 420
rect -805 410 -800 415
rect -880 390 -800 410
rect -880 385 -875 390
rect -915 380 -875 385
rect -805 385 -800 390
rect -770 410 -765 415
rect -695 415 -655 420
rect -695 410 -690 415
rect -770 390 -690 410
rect -770 385 -765 390
rect -805 380 -765 385
rect -695 385 -690 390
rect -660 410 -655 415
rect -585 415 -545 420
rect -585 410 -580 415
rect -660 390 -580 410
rect -660 385 -655 390
rect -695 380 -655 385
rect -585 385 -580 390
rect -550 385 -545 415
rect -585 380 -545 385
rect 2235 415 2275 420
rect 2235 385 2240 415
rect 2270 410 2275 415
rect 2345 415 2385 420
rect 2345 410 2350 415
rect 2270 390 2350 410
rect 2270 385 2275 390
rect 2235 380 2275 385
rect 2345 385 2350 390
rect 2380 410 2385 415
rect 2455 415 2495 420
rect 2455 410 2460 415
rect 2380 390 2460 410
rect 2380 385 2385 390
rect 2345 380 2385 385
rect 2455 385 2460 390
rect 2490 410 2495 415
rect 2565 415 2605 420
rect 2565 410 2570 415
rect 2490 390 2570 410
rect 2490 385 2495 390
rect 2455 380 2495 385
rect 2565 385 2570 390
rect 2600 410 2605 415
rect 2675 415 2715 420
rect 2675 410 2680 415
rect 2600 390 2680 410
rect 2600 385 2605 390
rect 2565 380 2605 385
rect 2675 385 2680 390
rect 2710 410 2715 415
rect 2920 415 2960 420
rect 2920 410 2925 415
rect 2710 390 2925 410
rect 2710 385 2715 390
rect 2675 380 2715 385
rect 2920 385 2925 390
rect 2955 385 2960 415
rect 2920 380 2960 385
rect -1545 350 -1495 360
rect -1545 320 -1535 350
rect -1505 320 -1495 350
rect 3185 350 3235 360
rect -1545 310 -1495 320
rect -750 340 -710 345
rect -750 310 -745 340
rect -715 335 -710 340
rect -370 340 -330 345
rect -370 335 -365 340
rect -715 315 -365 335
rect -715 310 -710 315
rect -750 305 -710 310
rect -370 310 -365 315
rect -335 310 -330 340
rect -370 305 -330 310
rect 2020 340 2060 345
rect 2020 310 2025 340
rect 2055 335 2060 340
rect 2400 340 2440 345
rect 2400 335 2405 340
rect 2055 315 2405 335
rect 2055 310 2060 315
rect 2020 305 2060 310
rect 2400 310 2405 315
rect 2435 310 2440 340
rect 3185 320 3195 350
rect 3225 320 3235 350
rect 3185 310 3235 320
rect 2400 305 2440 310
rect 5 275 45 280
rect -1225 265 -1185 270
rect -1225 235 -1220 265
rect -1190 260 -1185 265
rect -1025 265 -985 270
rect -1025 260 -1020 265
rect -1190 240 -1020 260
rect -1190 235 -1185 240
rect -1225 230 -1185 235
rect -1025 235 -1020 240
rect -990 260 -985 265
rect -915 265 -875 270
rect -915 260 -910 265
rect -990 240 -910 260
rect -990 235 -985 240
rect -1025 230 -985 235
rect -915 235 -910 240
rect -880 260 -875 265
rect -805 265 -765 270
rect -805 260 -800 265
rect -880 240 -800 260
rect -880 235 -875 240
rect -915 230 -875 235
rect -805 235 -800 240
rect -770 260 -765 265
rect -695 265 -655 270
rect -695 260 -690 265
rect -770 240 -690 260
rect -770 235 -765 240
rect -805 230 -765 235
rect -695 235 -690 240
rect -660 260 -655 265
rect -585 265 -545 270
rect -585 260 -580 265
rect -660 240 -580 260
rect -660 235 -655 240
rect -695 230 -655 235
rect -585 235 -580 240
rect -550 235 -545 265
rect 5 245 10 275
rect 40 270 45 275
rect 115 275 155 280
rect 115 270 120 275
rect 40 250 120 270
rect 40 245 45 250
rect 5 240 45 245
rect 115 245 120 250
rect 150 270 155 275
rect 225 275 265 280
rect 225 270 230 275
rect 150 250 230 270
rect 150 245 155 250
rect 115 240 155 245
rect 225 245 230 250
rect 260 270 265 275
rect 335 275 375 280
rect 335 270 340 275
rect 260 250 340 270
rect 260 245 265 250
rect 225 240 265 245
rect 335 245 340 250
rect 370 270 375 275
rect 445 275 485 280
rect 445 270 450 275
rect 370 250 450 270
rect 370 245 375 250
rect 335 240 375 245
rect 445 245 450 250
rect 480 245 485 275
rect 445 240 485 245
rect 1205 275 1245 280
rect 1205 245 1210 275
rect 1240 270 1245 275
rect 1315 275 1355 280
rect 1315 270 1320 275
rect 1240 250 1320 270
rect 1240 245 1245 250
rect 1205 240 1245 245
rect 1315 245 1320 250
rect 1350 270 1355 275
rect 1425 275 1465 280
rect 1425 270 1430 275
rect 1350 250 1430 270
rect 1350 245 1355 250
rect 1315 240 1355 245
rect 1425 245 1430 250
rect 1460 270 1465 275
rect 1535 275 1575 280
rect 1535 270 1540 275
rect 1460 250 1540 270
rect 1460 245 1465 250
rect 1425 240 1465 245
rect 1535 245 1540 250
rect 1570 270 1575 275
rect 1645 275 1685 280
rect 1645 270 1650 275
rect 1570 250 1650 270
rect 1570 245 1575 250
rect 1535 240 1575 245
rect 1645 245 1650 250
rect 1680 245 1685 275
rect 1645 240 1685 245
rect 2235 265 2275 270
rect 2235 235 2240 265
rect 2270 260 2275 265
rect 2345 265 2385 270
rect 2345 260 2350 265
rect 2270 240 2350 260
rect 2270 235 2275 240
rect -585 230 -545 235
rect -50 230 -10 235
rect -50 200 -45 230
rect -15 225 -10 230
rect 60 230 100 235
rect 60 225 65 230
rect -15 205 65 225
rect -15 200 -10 205
rect -50 195 -10 200
rect 60 200 65 205
rect 95 225 100 230
rect 170 230 210 235
rect 170 225 175 230
rect 95 205 175 225
rect 95 200 100 205
rect 60 195 100 200
rect 170 200 175 205
rect 205 225 210 230
rect 280 230 320 235
rect 280 225 285 230
rect 205 205 285 225
rect 205 200 210 205
rect 170 195 210 200
rect 280 200 285 205
rect 315 225 320 230
rect 390 230 430 235
rect 390 225 395 230
rect 315 205 395 225
rect 315 200 320 205
rect 280 195 320 200
rect 390 200 395 205
rect 425 225 430 230
rect 500 230 540 235
rect 500 225 505 230
rect 425 205 505 225
rect 425 200 430 205
rect 390 195 430 200
rect 500 200 505 205
rect 535 225 540 230
rect 1150 230 1190 235
rect 1150 225 1155 230
rect 535 205 1155 225
rect 535 200 540 205
rect 500 195 540 200
rect 770 175 775 205
rect 805 200 810 205
rect 880 200 885 205
rect 805 180 885 200
rect 805 175 810 180
rect 770 170 810 175
rect 880 175 885 180
rect 915 175 920 205
rect 1150 200 1155 205
rect 1185 225 1190 230
rect 1260 230 1300 235
rect 1260 225 1265 230
rect 1185 205 1265 225
rect 1185 200 1190 205
rect 1150 195 1190 200
rect 1260 200 1265 205
rect 1295 225 1300 230
rect 1370 230 1410 235
rect 1370 225 1375 230
rect 1295 205 1375 225
rect 1295 200 1300 205
rect 1260 195 1300 200
rect 1370 200 1375 205
rect 1405 225 1410 230
rect 1480 230 1520 235
rect 1480 225 1485 230
rect 1405 205 1485 225
rect 1405 200 1410 205
rect 1370 195 1410 200
rect 1480 200 1485 205
rect 1515 225 1520 230
rect 1590 230 1630 235
rect 1590 225 1595 230
rect 1515 205 1595 225
rect 1515 200 1520 205
rect 1480 195 1520 200
rect 1590 200 1595 205
rect 1625 225 1630 230
rect 1700 230 1740 235
rect 2235 230 2275 235
rect 2345 235 2350 240
rect 2380 260 2385 265
rect 2455 265 2495 270
rect 2455 260 2460 265
rect 2380 240 2460 260
rect 2380 235 2385 240
rect 2345 230 2385 235
rect 2455 235 2460 240
rect 2490 260 2495 265
rect 2565 265 2605 270
rect 2565 260 2570 265
rect 2490 240 2570 260
rect 2490 235 2495 240
rect 2455 230 2495 235
rect 2565 235 2570 240
rect 2600 260 2605 265
rect 2675 265 2715 270
rect 2675 260 2680 265
rect 2600 240 2680 260
rect 2600 235 2605 240
rect 2565 230 2605 235
rect 2675 235 2680 240
rect 2710 260 2715 265
rect 2875 265 2915 270
rect 2875 260 2880 265
rect 2710 240 2880 260
rect 2710 235 2715 240
rect 2675 230 2715 235
rect 2875 235 2880 240
rect 2910 235 2915 265
rect 2875 230 2915 235
rect 1700 225 1705 230
rect 1625 205 1705 225
rect 1625 200 1630 205
rect 1590 195 1630 200
rect 1700 200 1705 205
rect 1735 200 1740 230
rect 1700 195 1740 200
rect 880 170 920 175
rect 830 150 860 155
rect 880 150 920 155
rect 880 145 885 150
rect 860 125 885 145
rect 830 115 860 120
rect 880 120 885 125
rect 915 120 920 150
rect 880 115 920 120
rect 770 95 810 100
rect 770 65 775 95
rect 805 90 810 95
rect 830 95 860 100
rect 805 70 830 90
rect 805 65 810 70
rect 770 60 810 65
rect 830 60 860 65
rect 770 40 810 45
rect 770 10 775 40
rect 805 35 810 40
rect 880 40 920 45
rect 880 35 885 40
rect 805 15 885 35
rect 805 10 810 15
rect 770 5 810 10
rect 880 10 885 15
rect 915 10 920 40
rect 880 5 920 10
rect 440 -10 480 -5
rect 440 -40 445 -10
rect 475 -15 480 -10
rect 830 -10 860 -5
rect 475 -35 830 -15
rect 475 -40 480 -35
rect 440 -45 480 -40
rect 830 -45 860 -40
rect -1490 -120 -1486 -85
rect -1459 -120 -1426 -85
rect -1399 -120 -1395 -85
rect -1370 -120 -1366 -85
rect -1339 -120 -1335 -85
rect -1310 -120 -1306 -85
rect -1279 -95 -1275 -85
rect -1225 -90 -1185 -85
rect -1225 -95 -1220 -90
rect -1279 -115 -1220 -95
rect -1279 -120 -1275 -115
rect -1225 -120 -1220 -115
rect -1190 -120 -1185 -90
rect -1225 -125 -1185 -120
rect -1135 -90 -1095 -85
rect -1135 -120 -1130 -90
rect -1100 -120 -1095 -90
rect -1135 -125 -1095 -120
rect -1080 -90 -1040 -85
rect -1080 -120 -1075 -90
rect -1045 -95 -1040 -90
rect -970 -90 -930 -85
rect -970 -95 -965 -90
rect -1045 -115 -965 -95
rect -1045 -120 -1040 -115
rect -1080 -125 -1040 -120
rect -970 -120 -965 -115
rect -935 -95 -930 -90
rect -860 -90 -820 -85
rect -860 -95 -855 -90
rect -935 -115 -855 -95
rect -935 -120 -930 -115
rect -970 -125 -930 -120
rect -860 -120 -855 -115
rect -825 -95 -820 -90
rect -750 -90 -710 -85
rect -750 -95 -745 -90
rect -825 -115 -745 -95
rect -825 -120 -820 -115
rect -860 -125 -820 -120
rect -750 -120 -745 -115
rect -715 -95 -710 -90
rect -640 -90 -600 -85
rect -640 -95 -635 -90
rect -715 -115 -635 -95
rect -715 -120 -710 -115
rect -750 -125 -710 -120
rect -640 -120 -635 -115
rect -605 -95 -600 -90
rect -530 -90 -490 -85
rect -530 -95 -525 -90
rect -605 -115 -525 -95
rect -605 -120 -600 -115
rect -640 -125 -600 -120
rect -530 -120 -525 -115
rect -495 -95 -490 -90
rect -235 -90 -195 -85
rect -235 -95 -230 -90
rect -495 -115 -230 -95
rect -495 -120 -490 -115
rect -530 -125 -490 -120
rect -235 -120 -230 -115
rect -200 -120 -195 -90
rect -235 -125 -195 -120
rect 1885 -90 1925 -85
rect 1885 -120 1890 -90
rect 1920 -95 1925 -90
rect 2180 -90 2220 -85
rect 2180 -95 2185 -90
rect 1920 -115 2185 -95
rect 1920 -120 1925 -115
rect 1885 -125 1925 -120
rect 2180 -120 2185 -115
rect 2215 -95 2220 -90
rect 2290 -90 2330 -85
rect 2290 -95 2295 -90
rect 2215 -115 2295 -95
rect 2215 -120 2220 -115
rect 2180 -125 2220 -120
rect 2290 -120 2295 -115
rect 2325 -95 2330 -90
rect 2400 -90 2440 -85
rect 2400 -95 2405 -90
rect 2325 -115 2405 -95
rect 2325 -120 2330 -115
rect 2290 -125 2330 -120
rect 2400 -120 2405 -115
rect 2435 -95 2440 -90
rect 2510 -90 2550 -85
rect 2510 -95 2515 -90
rect 2435 -115 2515 -95
rect 2435 -120 2440 -115
rect 2400 -125 2440 -120
rect 2510 -120 2515 -115
rect 2545 -95 2550 -90
rect 2620 -90 2660 -85
rect 2620 -95 2625 -90
rect 2545 -115 2625 -95
rect 2545 -120 2550 -115
rect 2510 -125 2550 -120
rect 2620 -120 2625 -115
rect 2655 -95 2660 -90
rect 2730 -90 2770 -85
rect 2730 -95 2735 -90
rect 2655 -115 2735 -95
rect 2655 -120 2660 -115
rect 2620 -125 2660 -120
rect 2730 -120 2735 -115
rect 2765 -120 2770 -90
rect 2730 -125 2770 -120
rect 2785 -90 2825 -85
rect 2785 -120 2790 -90
rect 2820 -120 2825 -90
rect 2785 -125 2825 -120
rect 2875 -90 2915 -85
rect 2875 -120 2880 -90
rect 2910 -95 2915 -90
rect 2965 -95 2969 -85
rect 2910 -115 2969 -95
rect 2910 -120 2915 -115
rect 2965 -120 2969 -115
rect 2996 -120 3000 -85
rect 3025 -120 3029 -85
rect 3056 -120 3060 -85
rect 3085 -120 3089 -85
rect 3116 -120 3149 -85
rect 3176 -120 3180 -85
rect 2875 -125 2915 -120
rect -1370 -145 -1335 -140
rect -1270 -145 -1230 -140
rect -1270 -150 -1265 -145
rect -1335 -170 -1265 -150
rect -1370 -180 -1335 -175
rect -1270 -175 -1265 -170
rect -1235 -175 -1230 -145
rect -1270 -180 -1230 -175
rect -1135 -145 -1095 -140
rect -1135 -175 -1130 -145
rect -1100 -150 -1095 -145
rect -475 -145 -435 -140
rect -475 -150 -470 -145
rect -1100 -170 -470 -150
rect -1100 -175 -1095 -170
rect -1135 -180 -1095 -175
rect -475 -175 -470 -170
rect -440 -150 -435 -145
rect -280 -145 -240 -140
rect -280 -150 -275 -145
rect -440 -170 -275 -150
rect -440 -175 -435 -170
rect -280 -175 -275 -170
rect -245 -175 -240 -145
rect 1930 -145 1970 -140
rect 1930 -175 1935 -145
rect 1965 -150 1970 -145
rect 2125 -145 2165 -140
rect 2125 -150 2130 -145
rect 1965 -170 2130 -150
rect 1965 -175 1970 -170
rect 2125 -175 2130 -170
rect 2160 -150 2165 -145
rect 2785 -145 2825 -140
rect 2785 -150 2790 -145
rect 2160 -170 2790 -150
rect 2160 -175 2165 -170
rect -475 -180 -435 -175
rect 2125 -180 2165 -175
rect 2785 -175 2790 -170
rect 2820 -175 2825 -145
rect 2785 -180 2825 -175
rect 2920 -145 2960 -140
rect 2920 -175 2925 -145
rect 2955 -150 2960 -145
rect 3025 -145 3060 -140
rect 2955 -170 3025 -150
rect 2955 -175 2960 -170
rect 2920 -180 2960 -175
rect 3025 -180 3060 -175
rect -1490 -190 -1455 -185
rect 3145 -190 3180 -185
rect -325 -195 -320 -190
rect -1455 -215 -320 -195
rect -1490 -225 -1455 -220
rect -325 -220 -320 -215
rect -290 -220 -285 -190
rect -325 -225 -285 -220
rect 1975 -220 1980 -190
rect 2010 -195 2015 -190
rect 2010 -215 3145 -195
rect 2010 -220 2015 -215
rect 1975 -225 2015 -220
rect 3145 -225 3180 -220
rect -1290 -245 -1255 -240
rect -805 -245 -765 -240
rect -805 -250 -800 -245
rect -1255 -270 -800 -250
rect -1290 -280 -1255 -275
rect -805 -275 -800 -270
rect -770 -250 -765 -245
rect -235 -245 -195 -240
rect -235 -250 -230 -245
rect -770 -270 -230 -250
rect -770 -275 -765 -270
rect -805 -280 -765 -275
rect -235 -275 -230 -270
rect -200 -275 -195 -245
rect -235 -280 -195 -275
rect 1885 -245 1925 -240
rect 1885 -275 1890 -245
rect 1920 -250 1925 -245
rect 2455 -245 2495 -240
rect 2455 -250 2460 -245
rect 1920 -270 2460 -250
rect 1920 -275 1925 -270
rect 1885 -280 1925 -275
rect 2455 -275 2460 -270
rect 2490 -250 2495 -245
rect 2945 -245 2980 -240
rect 2490 -270 2945 -250
rect 2490 -275 2495 -270
rect 2455 -280 2495 -275
rect 2945 -280 2980 -275
rect -1540 -305 -1500 -300
rect -1540 -335 -1535 -305
rect -1505 -310 -1500 -305
rect -1230 -305 -1195 -300
rect -1505 -330 -1230 -310
rect -1505 -335 -1500 -330
rect -1540 -340 -1500 -335
rect -1005 -305 -965 -300
rect -1005 -310 -1000 -305
rect -1195 -330 -1000 -310
rect -1230 -340 -1195 -335
rect -1005 -335 -1000 -330
rect -970 -310 -965 -305
rect -805 -305 -765 -300
rect -805 -310 -800 -305
rect -970 -330 -800 -310
rect -970 -335 -965 -330
rect -1005 -340 -965 -335
rect -805 -335 -800 -330
rect -770 -310 -765 -305
rect -605 -305 -565 -300
rect 2255 -305 2295 -300
rect -605 -310 -600 -305
rect -770 -330 -600 -310
rect -770 -335 -765 -330
rect -805 -340 -765 -335
rect -605 -335 -600 -330
rect -570 -335 -565 -305
rect 1930 -310 1970 -305
rect 1930 -315 1935 -310
rect -605 -340 -565 -335
rect -105 -335 -65 -330
rect -105 -365 -100 -335
rect -70 -340 -65 -335
rect 555 -335 595 -330
rect 555 -340 560 -335
rect -70 -360 560 -340
rect -70 -365 -65 -360
rect -105 -370 -65 -365
rect 555 -365 560 -360
rect 590 -340 595 -335
rect 715 -335 755 -330
rect 715 -340 720 -335
rect 590 -360 720 -340
rect 590 -365 595 -360
rect 555 -370 595 -365
rect 715 -365 720 -360
rect 750 -340 755 -335
rect 825 -335 865 -330
rect 825 -340 830 -335
rect 750 -360 830 -340
rect 750 -365 755 -360
rect 715 -370 755 -365
rect 825 -365 830 -360
rect 860 -340 865 -335
rect 935 -335 975 -330
rect 935 -340 940 -335
rect 860 -360 940 -340
rect 860 -365 865 -360
rect 825 -370 865 -365
rect 935 -365 940 -360
rect 970 -340 975 -335
rect 1095 -335 1135 -330
rect 1095 -340 1100 -335
rect 970 -360 1100 -340
rect 970 -365 975 -360
rect 935 -370 975 -365
rect 1095 -365 1100 -360
rect 1130 -340 1135 -335
rect 1755 -335 1795 -330
rect 1845 -335 1935 -315
rect 1755 -340 1760 -335
rect 1130 -360 1760 -340
rect 1130 -365 1135 -360
rect 1095 -370 1135 -365
rect 1755 -365 1760 -360
rect 1790 -340 1795 -335
rect 1930 -340 1935 -335
rect 1965 -340 1970 -310
rect 2255 -335 2260 -305
rect 2290 -310 2295 -305
rect 2455 -305 2495 -300
rect 2455 -310 2460 -305
rect 2290 -330 2460 -310
rect 2290 -335 2295 -330
rect 2255 -340 2295 -335
rect 2455 -335 2460 -330
rect 2490 -310 2495 -305
rect 2655 -305 2695 -300
rect 2655 -310 2660 -305
rect 2490 -330 2660 -310
rect 2490 -335 2495 -330
rect 2455 -340 2495 -335
rect 2655 -335 2660 -330
rect 2690 -310 2695 -305
rect 2885 -305 2920 -300
rect 2690 -330 2885 -310
rect 2690 -335 2695 -330
rect 2655 -340 2695 -335
rect 3190 -305 3230 -300
rect 3190 -310 3195 -305
rect 2920 -330 3195 -310
rect 2885 -340 2920 -335
rect 3190 -335 3195 -330
rect 3225 -335 3230 -305
rect 3190 -340 3230 -335
rect 1790 -360 1845 -340
rect 1930 -345 1970 -340
rect 1790 -365 1795 -360
rect 1755 -370 1795 -365
rect -235 -380 -195 -375
rect -1290 -415 -1286 -380
rect -1259 -415 -1255 -380
rect -1230 -415 -1226 -380
rect -1199 -415 -1195 -380
rect -235 -410 -230 -380
rect -200 -385 -195 -380
rect 1885 -380 1925 -375
rect 1885 -385 1890 -380
rect -200 -405 1890 -385
rect -200 -410 -195 -405
rect -235 -415 -195 -410
rect 1885 -410 1890 -405
rect 1920 -410 1925 -380
rect 1885 -415 1925 -410
rect 2885 -415 2889 -380
rect 2916 -415 2920 -380
rect 2945 -415 2949 -380
rect 2976 -415 2980 -380
rect 1350 -435 1390 -430
rect 1350 -465 1355 -435
rect 1385 -440 1390 -435
rect 1840 -435 1880 -430
rect 1840 -440 1845 -435
rect 1385 -460 1845 -440
rect 1385 -465 1390 -460
rect 1350 -470 1390 -465
rect 1840 -465 1845 -460
rect 1875 -465 1880 -435
rect 1840 -470 1880 -465
rect 385 -490 425 -485
rect 385 -520 390 -490
rect 420 -495 425 -490
rect 495 -490 535 -485
rect 495 -495 500 -490
rect 420 -515 500 -495
rect 420 -520 425 -515
rect 385 -525 425 -520
rect 495 -520 500 -515
rect 530 -495 535 -490
rect 605 -490 645 -485
rect 605 -495 610 -490
rect 530 -515 610 -495
rect 530 -520 535 -515
rect 495 -525 535 -520
rect 605 -520 610 -515
rect 640 -495 645 -490
rect 715 -490 755 -485
rect 715 -495 720 -490
rect 640 -515 720 -495
rect 640 -520 645 -515
rect 605 -525 645 -520
rect 715 -520 720 -515
rect 750 -495 755 -490
rect 825 -490 865 -485
rect 825 -495 830 -490
rect 750 -515 830 -495
rect 750 -520 755 -515
rect 715 -525 755 -520
rect 825 -520 830 -515
rect 860 -495 865 -490
rect 935 -490 975 -485
rect 935 -495 940 -490
rect 860 -515 940 -495
rect 860 -520 865 -515
rect 825 -525 865 -520
rect 935 -520 940 -515
rect 970 -495 975 -490
rect 1045 -490 1085 -485
rect 1045 -495 1050 -490
rect 970 -515 1050 -495
rect 970 -520 975 -515
rect 935 -525 975 -520
rect 1045 -520 1050 -515
rect 1080 -495 1085 -490
rect 1155 -490 1195 -485
rect 1155 -495 1160 -490
rect 1080 -515 1160 -495
rect 1080 -520 1085 -515
rect 1045 -525 1085 -520
rect 1155 -520 1160 -515
rect 1190 -495 1195 -490
rect 1265 -490 1305 -485
rect 1265 -495 1270 -490
rect 1190 -515 1270 -495
rect 1190 -520 1195 -515
rect 1155 -525 1195 -520
rect 1265 -520 1270 -515
rect 1300 -495 1305 -490
rect 1375 -490 1415 -485
rect 1375 -495 1380 -490
rect 1300 -515 1380 -495
rect 1300 -520 1305 -515
rect 1265 -525 1305 -520
rect 1375 -520 1380 -515
rect 1410 -520 1415 -490
rect 1375 -525 1415 -520
rect 275 -805 315 -800
rect 275 -835 280 -805
rect 310 -810 315 -805
rect 330 -805 370 -800
rect 330 -810 335 -805
rect 310 -830 335 -810
rect 310 -835 315 -830
rect 275 -840 315 -835
rect 330 -835 335 -830
rect 365 -810 370 -805
rect 440 -805 480 -800
rect 440 -810 445 -805
rect 365 -830 445 -810
rect 365 -835 370 -830
rect 330 -840 370 -835
rect 440 -835 445 -830
rect 475 -810 480 -805
rect 550 -805 590 -800
rect 550 -810 555 -805
rect 475 -830 555 -810
rect 475 -835 480 -830
rect 440 -840 480 -835
rect 550 -835 555 -830
rect 585 -810 590 -805
rect 660 -805 700 -800
rect 660 -810 665 -805
rect 585 -830 665 -810
rect 585 -835 590 -830
rect 550 -840 590 -835
rect 660 -835 665 -830
rect 695 -810 700 -805
rect 770 -805 810 -800
rect 770 -810 775 -805
rect 695 -830 775 -810
rect 695 -835 700 -830
rect 660 -840 700 -835
rect 770 -835 775 -830
rect 805 -810 810 -805
rect 880 -805 920 -800
rect 880 -810 885 -805
rect 805 -830 885 -810
rect 805 -835 810 -830
rect 770 -840 810 -835
rect 880 -835 885 -830
rect 915 -810 920 -805
rect 990 -805 1030 -800
rect 990 -810 995 -805
rect 915 -830 995 -810
rect 915 -835 920 -830
rect 880 -840 920 -835
rect 990 -835 995 -830
rect 1025 -810 1030 -805
rect 1100 -805 1140 -800
rect 1100 -810 1105 -805
rect 1025 -830 1105 -810
rect 1025 -835 1030 -830
rect 990 -840 1030 -835
rect 1100 -835 1105 -830
rect 1135 -810 1140 -805
rect 1210 -805 1250 -800
rect 1210 -810 1215 -805
rect 1135 -830 1215 -810
rect 1135 -835 1140 -830
rect 1100 -840 1140 -835
rect 1210 -835 1215 -830
rect 1245 -810 1250 -805
rect 1320 -805 1360 -800
rect 1320 -810 1325 -805
rect 1245 -830 1325 -810
rect 1245 -835 1250 -830
rect 1210 -840 1250 -835
rect 1320 -835 1325 -830
rect 1355 -810 1360 -805
rect 1430 -805 1470 -800
rect 1430 -810 1435 -805
rect 1355 -830 1435 -810
rect 1355 -835 1360 -830
rect 1320 -840 1360 -835
rect 1430 -835 1435 -830
rect 1465 -810 1470 -805
rect 1930 -805 1970 -800
rect 1930 -810 1935 -805
rect 1465 -830 1935 -810
rect 1465 -835 1470 -830
rect 1430 -840 1470 -835
rect 1930 -835 1935 -830
rect 1965 -835 1970 -805
rect 1930 -840 1970 -835
rect 385 -850 425 -845
rect 385 -880 390 -850
rect 420 -855 425 -850
rect 495 -850 535 -845
rect 495 -855 500 -850
rect 420 -875 500 -855
rect 420 -880 425 -875
rect 385 -885 425 -880
rect 495 -880 500 -875
rect 530 -855 535 -850
rect 605 -850 645 -845
rect 605 -855 610 -850
rect 530 -875 610 -855
rect 530 -880 535 -875
rect 495 -885 535 -880
rect 605 -880 610 -875
rect 640 -855 645 -850
rect 715 -850 755 -845
rect 715 -855 720 -850
rect 640 -875 720 -855
rect 640 -880 645 -875
rect 605 -885 645 -880
rect 715 -880 720 -875
rect 750 -855 755 -850
rect 825 -850 865 -845
rect 825 -855 830 -850
rect 750 -875 830 -855
rect 750 -880 755 -875
rect 715 -885 755 -880
rect 825 -880 830 -875
rect 860 -855 865 -850
rect 935 -850 975 -845
rect 935 -855 940 -850
rect 860 -875 940 -855
rect 860 -880 865 -875
rect 825 -885 865 -880
rect 935 -880 940 -875
rect 970 -855 975 -850
rect 1045 -850 1085 -845
rect 1045 -855 1050 -850
rect 970 -875 1050 -855
rect 970 -880 975 -875
rect 935 -885 975 -880
rect 1045 -880 1050 -875
rect 1080 -855 1085 -850
rect 1155 -850 1195 -845
rect 1155 -855 1160 -850
rect 1080 -875 1160 -855
rect 1080 -880 1085 -875
rect 1045 -885 1085 -880
rect 1155 -880 1160 -875
rect 1190 -855 1195 -850
rect 1265 -850 1305 -845
rect 1265 -855 1270 -850
rect 1190 -875 1270 -855
rect 1190 -880 1195 -875
rect 1155 -885 1195 -880
rect 1265 -880 1270 -875
rect 1300 -855 1305 -850
rect 1375 -850 1415 -845
rect 1375 -855 1380 -850
rect 1300 -875 1380 -855
rect 1300 -880 1305 -875
rect 1265 -885 1305 -880
rect 1375 -880 1380 -875
rect 1410 -880 1415 -850
rect 1375 -885 1415 -880
rect 595 -915 635 -910
rect 595 -945 600 -915
rect 630 -920 635 -915
rect 705 -915 745 -910
rect 705 -920 710 -915
rect 630 -940 710 -920
rect 630 -945 635 -940
rect 595 -950 635 -945
rect 705 -945 710 -940
rect 740 -920 745 -915
rect 925 -915 965 -910
rect 925 -920 930 -915
rect 740 -940 930 -920
rect 740 -945 745 -940
rect 705 -950 745 -945
rect 925 -945 930 -940
rect 960 -945 965 -915
rect 925 -950 965 -945
rect -190 -960 -150 -955
rect -190 -990 -185 -960
rect -155 -965 -150 -960
rect 540 -960 580 -955
rect 540 -965 545 -960
rect -155 -985 545 -965
rect -155 -990 -150 -985
rect -190 -995 -150 -990
rect 540 -990 545 -985
rect 575 -965 580 -960
rect 650 -960 690 -955
rect 650 -965 655 -960
rect 575 -985 655 -965
rect 575 -990 580 -985
rect 540 -995 580 -990
rect 650 -990 655 -985
rect 685 -965 690 -960
rect 760 -960 800 -955
rect 760 -965 765 -960
rect 685 -985 765 -965
rect 685 -990 690 -985
rect 650 -995 690 -990
rect 760 -990 765 -985
rect 795 -965 800 -960
rect 1095 -960 1135 -955
rect 1095 -965 1100 -960
rect 795 -985 1100 -965
rect 795 -990 800 -985
rect 760 -995 800 -990
rect 1095 -990 1100 -985
rect 1130 -990 1135 -960
rect 1095 -995 1135 -990
rect 1265 -960 1305 -955
rect 1265 -990 1270 -960
rect 1300 -990 1305 -960
rect 1265 -995 1305 -990
rect -1105 -1075 -1065 -1070
rect -1105 -1105 -1100 -1075
rect -1070 -1080 -1065 -1075
rect -905 -1075 -865 -1070
rect -905 -1080 -900 -1075
rect -1070 -1100 -900 -1080
rect -1070 -1105 -1065 -1100
rect -1105 -1110 -1065 -1105
rect -905 -1105 -900 -1100
rect -870 -1080 -865 -1075
rect -705 -1075 -665 -1070
rect -705 -1080 -700 -1075
rect -870 -1100 -700 -1080
rect -870 -1105 -865 -1100
rect -905 -1110 -865 -1105
rect -705 -1105 -700 -1100
rect -670 -1080 -665 -1075
rect -505 -1075 -465 -1070
rect -505 -1080 -500 -1075
rect -670 -1100 -500 -1080
rect -670 -1105 -665 -1100
rect -705 -1110 -665 -1105
rect -505 -1105 -500 -1100
rect -470 -1105 -465 -1075
rect -505 -1110 -465 -1105
rect 2155 -1075 2195 -1070
rect 2155 -1105 2160 -1075
rect 2190 -1080 2195 -1075
rect 2355 -1075 2395 -1070
rect 2355 -1080 2360 -1075
rect 2190 -1100 2360 -1080
rect 2190 -1105 2195 -1100
rect 2155 -1110 2195 -1105
rect 2355 -1105 2360 -1100
rect 2390 -1080 2395 -1075
rect 2555 -1075 2595 -1070
rect 2555 -1080 2560 -1075
rect 2390 -1100 2560 -1080
rect 2390 -1105 2395 -1100
rect 2355 -1110 2395 -1105
rect 2555 -1105 2560 -1100
rect 2590 -1080 2595 -1075
rect 2755 -1075 2795 -1070
rect 2755 -1080 2760 -1075
rect 2590 -1100 2760 -1080
rect 2590 -1105 2595 -1100
rect 2555 -1110 2595 -1105
rect 2755 -1105 2760 -1100
rect 2790 -1105 2795 -1075
rect 2755 -1110 2795 -1105
rect 595 -1165 635 -1160
rect 595 -1195 600 -1165
rect 630 -1170 635 -1165
rect 705 -1165 745 -1160
rect 705 -1170 710 -1165
rect 630 -1190 710 -1170
rect 630 -1195 635 -1190
rect 595 -1200 635 -1195
rect 705 -1195 710 -1190
rect 740 -1170 745 -1165
rect 925 -1165 965 -1160
rect 925 -1170 930 -1165
rect 740 -1190 930 -1170
rect 740 -1195 745 -1190
rect 705 -1200 745 -1195
rect 925 -1195 930 -1190
rect 960 -1195 965 -1165
rect 925 -1200 965 -1195
rect 540 -1210 580 -1205
rect 540 -1240 545 -1210
rect 575 -1215 580 -1210
rect 650 -1210 690 -1205
rect 650 -1215 655 -1210
rect 575 -1235 655 -1215
rect 575 -1240 580 -1235
rect 540 -1245 580 -1240
rect 650 -1240 655 -1235
rect 685 -1215 690 -1210
rect 760 -1210 800 -1205
rect 760 -1215 765 -1210
rect 685 -1235 765 -1215
rect 685 -1240 690 -1235
rect 650 -1245 690 -1240
rect 760 -1240 765 -1235
rect 795 -1240 800 -1210
rect 760 -1245 800 -1240
rect -705 -1255 -665 -1250
rect -705 -1285 -700 -1255
rect -670 -1260 -665 -1255
rect -280 -1255 -240 -1250
rect -280 -1260 -275 -1255
rect -670 -1280 -275 -1260
rect -670 -1285 -665 -1280
rect -705 -1290 -665 -1285
rect -280 -1285 -275 -1280
rect -245 -1260 -240 -1255
rect 485 -1255 525 -1250
rect 485 -1260 490 -1255
rect -245 -1280 490 -1260
rect -245 -1285 -240 -1280
rect -280 -1290 -240 -1285
rect 485 -1285 490 -1280
rect 520 -1260 525 -1255
rect 815 -1255 855 -1250
rect 815 -1260 820 -1255
rect 520 -1280 820 -1260
rect 520 -1285 525 -1280
rect 485 -1290 525 -1285
rect 815 -1285 820 -1280
rect 850 -1260 855 -1255
rect 1930 -1255 1970 -1250
rect 1930 -1260 1935 -1255
rect 850 -1280 1935 -1260
rect 850 -1285 855 -1280
rect 815 -1290 855 -1285
rect 1930 -1285 1935 -1280
rect 1965 -1260 1970 -1255
rect 2355 -1255 2395 -1250
rect 2355 -1260 2360 -1255
rect 1965 -1280 2360 -1260
rect 1965 -1285 1970 -1280
rect 1930 -1290 1970 -1285
rect 2355 -1285 2360 -1280
rect 2390 -1285 2395 -1255
rect 2355 -1290 2395 -1285
rect 825 -2425 865 -2420
rect 825 -2455 830 -2425
rect 860 -2455 865 -2425
rect 825 -2460 865 -2455
<< via2 >>
rect 830 4245 860 4275
rect -1445 1510 -1415 1540
rect 3105 1460 3135 1490
rect -1535 320 -1505 350
rect 3195 320 3225 350
rect 830 -2455 860 -2425
<< metal3 >>
rect 820 4280 870 4285
rect 820 4240 825 4280
rect 865 4240 870 4280
rect 820 4235 870 4240
rect -3295 3860 -3065 3945
rect -2945 3860 -2715 3945
rect -2595 3860 -2365 3945
rect -3295 3810 -2365 3860
rect -3295 3715 -3065 3810
rect -2945 3715 -2715 3810
rect -2595 3715 -2365 3810
rect -2245 3715 -2015 3945
rect -1895 3715 -1665 3945
rect -1545 3715 -1315 3945
rect -1195 3715 -965 3945
rect -845 3715 -615 3945
rect -495 3715 -265 3945
rect -145 3715 85 3945
rect 205 3715 435 3945
rect 555 3715 785 3945
rect 905 3715 1135 3945
rect 1255 3715 1485 3945
rect 1605 3715 1835 3945
rect 1955 3715 2185 3945
rect 2305 3715 2535 3945
rect 2655 3715 2885 3945
rect 3005 3715 3235 3945
rect 3355 3715 3585 3945
rect 3705 3715 3935 3945
rect 4055 3860 4285 3945
rect 4405 3860 4635 3945
rect 4755 3860 4985 3945
rect 4055 3810 4985 3860
rect 4055 3715 4285 3810
rect 4405 3715 4635 3810
rect 4755 3715 4985 3810
rect -2505 3595 -2455 3715
rect -2155 3595 -2105 3715
rect -1805 3595 -1755 3715
rect -1455 3595 -1405 3715
rect -1105 3595 -1055 3715
rect -755 3595 -705 3715
rect -405 3595 -355 3715
rect -55 3595 -5 3715
rect 295 3595 345 3715
rect 645 3595 695 3715
rect 995 3595 1045 3715
rect 1345 3595 1395 3715
rect 1695 3595 1745 3715
rect 2045 3595 2095 3715
rect 2395 3595 2445 3715
rect 2745 3595 2795 3715
rect 3095 3595 3145 3715
rect 3445 3595 3495 3715
rect 3795 3595 3845 3715
rect 4145 3595 4195 3715
rect -3295 3510 -3065 3595
rect -2945 3510 -2715 3595
rect -2595 3510 -2365 3595
rect -2245 3510 -2015 3595
rect -1895 3510 -1665 3595
rect -1545 3510 -1315 3595
rect -1195 3510 -965 3595
rect -845 3510 -615 3595
rect -495 3510 -265 3595
rect -145 3510 85 3595
rect 205 3510 435 3595
rect 555 3510 785 3595
rect -3295 3460 785 3510
rect -3295 3365 -3065 3460
rect -2945 3365 -2715 3460
rect -2595 3365 -2365 3460
rect -2245 3365 -2015 3460
rect -1895 3365 -1665 3460
rect -1545 3365 -1315 3460
rect -1195 3365 -965 3460
rect -845 3365 -615 3460
rect -495 3365 -265 3460
rect -145 3365 85 3460
rect 205 3365 435 3460
rect 555 3365 785 3460
rect 905 3510 1135 3595
rect 1255 3510 1485 3595
rect 1605 3510 1835 3595
rect 1955 3510 2185 3595
rect 2305 3510 2535 3595
rect 2655 3510 2885 3595
rect 3005 3510 3235 3595
rect 3355 3510 3585 3595
rect 3705 3510 3935 3595
rect 4055 3510 4285 3595
rect 4405 3510 4635 3595
rect 4755 3510 4985 3595
rect 905 3460 4985 3510
rect 905 3365 1135 3460
rect 1255 3365 1485 3460
rect 1605 3365 1835 3460
rect 1955 3365 2185 3460
rect 2305 3365 2535 3460
rect 2655 3365 2885 3460
rect 3005 3365 3235 3460
rect 3355 3365 3585 3460
rect 3705 3365 3935 3460
rect 4055 3365 4285 3460
rect 4405 3365 4635 3460
rect 4755 3365 4985 3460
rect -2505 3245 -2455 3365
rect -1805 3245 -1755 3365
rect -1455 3245 -1405 3365
rect -1105 3245 -1055 3365
rect -755 3245 -705 3365
rect -405 3245 -355 3365
rect -55 3245 -5 3365
rect 295 3245 345 3365
rect 645 3245 695 3365
rect 995 3245 1045 3365
rect 1345 3245 1395 3365
rect 1695 3245 1745 3365
rect 2045 3245 2095 3365
rect 2395 3245 2445 3365
rect 2745 3245 2795 3365
rect 3095 3245 3145 3365
rect 3445 3245 3495 3365
rect 4145 3245 4195 3365
rect -3295 3160 -3065 3245
rect -2945 3160 -2715 3245
rect -2595 3160 -2365 3245
rect -2245 3160 -2015 3245
rect -3295 3110 -2015 3160
rect -3295 3015 -3065 3110
rect -2945 3015 -2715 3110
rect -2595 3015 -2365 3110
rect -2245 3015 -2015 3110
rect -1895 3015 -1665 3245
rect -1545 3015 -1315 3245
rect -1195 3015 -965 3245
rect -845 3015 -615 3245
rect -495 3015 -265 3245
rect -145 3015 85 3245
rect 205 3015 435 3245
rect 555 3015 785 3245
rect 905 3015 1135 3245
rect 1255 3015 1485 3245
rect 1605 3015 1835 3245
rect 1955 3015 2185 3245
rect 2305 3015 2535 3245
rect 2655 3015 2885 3245
rect 3005 3015 3235 3245
rect 3355 3015 3585 3245
rect 3705 3160 3935 3245
rect 4055 3160 4285 3245
rect 4405 3160 4635 3245
rect 4755 3160 4985 3245
rect 3705 3110 4985 3160
rect 3705 3015 3935 3110
rect 4055 3015 4285 3110
rect 4405 3015 4635 3110
rect 4755 3015 4985 3110
rect -2505 2895 -2455 3015
rect -1805 2895 -1755 3015
rect -1455 2895 -1405 3015
rect -1105 2895 -1055 3015
rect -755 2895 -705 3015
rect 2395 2895 2445 3015
rect 2745 2895 2795 3015
rect 3095 2895 3145 3015
rect 3445 2895 3495 3015
rect 4145 2895 4195 3015
rect -3295 2810 -3065 2895
rect -2945 2810 -2715 2895
rect -2595 2810 -2365 2895
rect -2245 2810 -2015 2895
rect -3295 2760 -2015 2810
rect -3295 2665 -3065 2760
rect -2945 2665 -2715 2760
rect -2595 2665 -2365 2760
rect -2245 2665 -2015 2760
rect -1895 2665 -1665 2895
rect -1545 2665 -1315 2895
rect -1195 2665 -965 2895
rect -845 2665 -615 2895
rect 2305 2665 2535 2895
rect 2655 2665 2885 2895
rect 3005 2665 3235 2895
rect 3355 2665 3585 2895
rect 3705 2810 3935 2895
rect 4055 2810 4285 2895
rect 4405 2810 4635 2895
rect 4755 2810 4985 2895
rect 3705 2760 4985 2810
rect 3705 2665 3935 2760
rect 4055 2665 4285 2760
rect 4405 2665 4635 2760
rect 4755 2665 4985 2760
rect -2505 2545 -2455 2665
rect -1455 2545 -1405 2665
rect -1105 2545 -1055 2665
rect -755 2545 -705 2665
rect 2395 2545 2445 2665
rect 2745 2545 2795 2665
rect 3095 2545 3145 2665
rect 4145 2545 4195 2665
rect -3295 2460 -3065 2545
rect -2945 2460 -2715 2545
rect -2595 2460 -2365 2545
rect -2245 2460 -2015 2545
rect -1895 2460 -1665 2545
rect -3295 2410 -1665 2460
rect -3295 2315 -3065 2410
rect -2945 2315 -2715 2410
rect -2595 2315 -2365 2410
rect -2245 2315 -2015 2410
rect -1895 2315 -1665 2410
rect -1545 2315 -1315 2545
rect -1195 2315 -965 2545
rect -845 2315 -615 2545
rect 2305 2315 2535 2545
rect 2655 2315 2885 2545
rect 3005 2315 3235 2545
rect 3355 2460 3585 2545
rect 3705 2460 3935 2545
rect 4055 2460 4285 2545
rect 4405 2460 4635 2545
rect 4755 2460 4985 2545
rect 3355 2410 4985 2460
rect 3355 2315 3585 2410
rect 3705 2315 3935 2410
rect 4055 2315 4285 2410
rect 4405 2315 4635 2410
rect 4755 2315 4985 2410
rect -2505 2195 -2455 2315
rect -3295 2110 -3065 2195
rect -2945 2110 -2715 2195
rect -2595 2110 -2365 2195
rect -2245 2110 -2015 2195
rect -1895 2110 -1665 2195
rect -3295 2060 -1665 2110
rect -3295 1965 -3065 2060
rect -2945 1965 -2715 2060
rect -2595 1965 -2365 2060
rect -2245 1965 -2015 2060
rect -1895 1965 -1665 2060
rect -2505 1845 -2455 1965
rect -3295 1760 -3065 1845
rect -2945 1760 -2715 1845
rect -2595 1760 -2365 1845
rect -2245 1760 -2015 1845
rect -1895 1760 -1665 1845
rect -3295 1710 -1665 1760
rect -3295 1615 -3065 1710
rect -2945 1615 -2715 1710
rect -2595 1615 -2365 1710
rect -2245 1615 -2015 1710
rect -1895 1615 -1665 1710
rect -2505 1495 -2455 1615
rect -1450 1540 -1410 2315
rect -1450 1510 -1445 1540
rect -1415 1510 -1410 1540
rect -1450 1505 -1410 1510
rect -3295 1410 -3065 1495
rect -2945 1410 -2715 1495
rect -2595 1410 -2365 1495
rect -2245 1410 -2015 1495
rect -1895 1410 -1665 1495
rect 3100 1490 3140 2315
rect 4145 2195 4195 2315
rect 3355 2110 3585 2195
rect 3705 2110 3935 2195
rect 4055 2110 4285 2195
rect 4405 2110 4635 2195
rect 4755 2110 4985 2195
rect 3355 2060 4985 2110
rect 3355 1965 3585 2060
rect 3705 1965 3935 2060
rect 4055 1965 4285 2060
rect 4405 1965 4635 2060
rect 4755 1965 4985 2060
rect 4145 1845 4195 1965
rect 3355 1760 3585 1845
rect 3705 1760 3935 1845
rect 4055 1760 4285 1845
rect 4405 1760 4635 1845
rect 4755 1760 4985 1845
rect 3355 1710 4985 1760
rect 3355 1615 3585 1710
rect 3705 1615 3935 1710
rect 4055 1615 4285 1710
rect 4405 1615 4635 1710
rect 4755 1615 4985 1710
rect 4145 1495 4195 1615
rect 3100 1460 3105 1490
rect 3135 1460 3140 1490
rect 3100 1455 3140 1460
rect -3295 1360 -1665 1410
rect -3295 1265 -3065 1360
rect -2945 1265 -2715 1360
rect -2595 1265 -2365 1360
rect -2245 1265 -2015 1360
rect -1895 1265 -1665 1360
rect 3355 1410 3585 1495
rect 3705 1410 3935 1495
rect 4055 1410 4285 1495
rect 4405 1410 4635 1495
rect 4755 1410 4985 1495
rect 3355 1360 4985 1410
rect 3355 1265 3585 1360
rect 3705 1265 3935 1360
rect 4055 1265 4285 1360
rect 4405 1265 4635 1360
rect 4755 1265 4985 1360
rect -2505 1145 -2455 1265
rect 4145 1145 4195 1265
rect -3295 1060 -3065 1145
rect -2945 1060 -2715 1145
rect -2595 1060 -2365 1145
rect -2245 1060 -2015 1145
rect -1895 1060 -1665 1145
rect -3295 1010 -1665 1060
rect -3295 915 -3065 1010
rect -2945 915 -2715 1010
rect -2595 915 -2365 1010
rect -2245 915 -2015 1010
rect -1895 915 -1665 1010
rect 3355 1060 3585 1145
rect 3705 1060 3935 1145
rect 4055 1060 4285 1145
rect 4405 1060 4635 1145
rect 4755 1060 4985 1145
rect 3355 1010 4985 1060
rect 3355 915 3585 1010
rect 3705 915 3935 1010
rect 4055 915 4285 1010
rect 4405 915 4635 1010
rect 4755 915 4985 1010
rect -2505 795 -2455 915
rect 4145 795 4195 915
rect -3295 710 -3065 795
rect -2945 710 -2715 795
rect -2595 710 -2365 795
rect -2245 710 -2015 795
rect -1895 710 -1665 795
rect -3295 660 -1665 710
rect -3295 565 -3065 660
rect -2945 565 -2715 660
rect -2595 565 -2365 660
rect -2245 565 -2015 660
rect -1895 565 -1665 660
rect 3355 710 3585 795
rect 3705 710 3935 795
rect 4055 710 4285 795
rect 4405 710 4635 795
rect 4755 710 4985 795
rect 3355 660 4985 710
rect 3355 565 3585 660
rect 3705 565 3935 660
rect 4055 565 4285 660
rect 4405 565 4635 660
rect 4755 565 4985 660
rect -2505 445 -2455 565
rect 4145 445 4195 565
rect -3295 360 -3065 445
rect -2945 360 -2715 445
rect -2595 360 -2365 445
rect -2245 360 -2015 445
rect -1895 360 -1665 445
rect 3355 360 3585 445
rect 3705 360 3935 445
rect 4055 360 4285 445
rect 4405 360 4635 445
rect 4755 360 4985 445
rect -3295 310 -1665 360
rect -1545 355 -1495 360
rect -1545 315 -1540 355
rect -1500 315 -1495 355
rect -1545 310 -1495 315
rect 3185 355 3235 360
rect 3185 315 3190 355
rect 3230 315 3235 355
rect 3185 310 3235 315
rect 3355 310 4985 360
rect -3295 215 -3065 310
rect -2945 215 -2715 310
rect -2595 215 -2365 310
rect -2245 215 -2015 310
rect -1895 215 -1665 310
rect 3355 215 3585 310
rect 3705 215 3935 310
rect 4055 215 4285 310
rect 4405 215 4635 310
rect 4755 215 4985 310
rect -2505 95 -2455 215
rect 4145 95 4195 215
rect -3295 10 -3065 95
rect -2945 10 -2715 95
rect -2595 10 -2365 95
rect -2245 10 -2015 95
rect -1895 10 -1665 95
rect -3295 -40 -1665 10
rect -3295 -135 -3065 -40
rect -2945 -135 -2715 -40
rect -2595 -135 -2365 -40
rect -2245 -135 -2015 -40
rect -1895 -135 -1665 -40
rect 3355 10 3585 95
rect 3705 10 3935 95
rect 4055 10 4285 95
rect 4405 10 4635 95
rect 4755 10 4985 95
rect 3355 -40 4985 10
rect 3355 -135 3585 -40
rect 3705 -135 3935 -40
rect 4055 -135 4285 -40
rect 4405 -135 4635 -40
rect 4755 -135 4985 -40
rect -2505 -255 -2455 -135
rect 4145 -255 4195 -135
rect -3295 -340 -3065 -255
rect -2945 -340 -2715 -255
rect -2595 -340 -2365 -255
rect -2245 -340 -2015 -255
rect -1895 -340 -1665 -255
rect -3295 -390 -1665 -340
rect -3295 -485 -3065 -390
rect -2945 -485 -2715 -390
rect -2595 -485 -2365 -390
rect -2245 -485 -2015 -390
rect -1895 -485 -1665 -390
rect 3355 -340 3585 -255
rect 3705 -340 3935 -255
rect 4055 -340 4285 -255
rect 4405 -340 4635 -255
rect 4755 -340 4985 -255
rect 3355 -390 4985 -340
rect 3355 -485 3585 -390
rect 3705 -485 3935 -390
rect 4055 -485 4285 -390
rect 4405 -485 4635 -390
rect 4755 -485 4985 -390
rect -2505 -605 -2455 -485
rect 4145 -605 4195 -485
rect -3295 -690 -3065 -605
rect -2945 -690 -2715 -605
rect -2595 -690 -2365 -605
rect -2245 -690 -2015 -605
rect -1895 -690 -1665 -605
rect -3295 -740 -1665 -690
rect -3295 -835 -3065 -740
rect -2945 -835 -2715 -740
rect -2595 -835 -2365 -740
rect -2245 -835 -2015 -740
rect -1895 -835 -1665 -740
rect 3355 -690 3585 -605
rect 3705 -690 3935 -605
rect 4055 -690 4285 -605
rect 4405 -690 4635 -605
rect 4755 -690 4985 -605
rect 3355 -740 4985 -690
rect 3355 -835 3585 -740
rect 3705 -835 3935 -740
rect 4055 -835 4285 -740
rect 4405 -835 4635 -740
rect 4755 -835 4985 -740
rect -2505 -955 -2455 -835
rect 4145 -955 4195 -835
rect -3295 -1040 -3065 -955
rect -2945 -1040 -2715 -955
rect -2595 -1040 -2365 -955
rect -2245 -1040 -2015 -955
rect -1895 -1040 -1665 -955
rect -3295 -1090 -1665 -1040
rect -3295 -1185 -3065 -1090
rect -2945 -1185 -2715 -1090
rect -2595 -1185 -2365 -1090
rect -2245 -1185 -2015 -1090
rect -1895 -1185 -1665 -1090
rect 3355 -1040 3585 -955
rect 3705 -1040 3935 -955
rect 4055 -1040 4285 -955
rect 4405 -1040 4635 -955
rect 4755 -1040 4985 -955
rect 3355 -1090 4985 -1040
rect 3355 -1185 3585 -1090
rect 3705 -1185 3935 -1090
rect 4055 -1185 4285 -1090
rect 4405 -1185 4635 -1090
rect 4755 -1185 4985 -1090
rect -2505 -1305 -2455 -1185
rect 4145 -1305 4195 -1185
rect -3295 -1390 -3065 -1305
rect -2945 -1390 -2715 -1305
rect -2595 -1390 -2365 -1305
rect -2245 -1390 -2015 -1305
rect -1895 -1390 -1665 -1305
rect -3295 -1440 -1665 -1390
rect -3295 -1535 -3065 -1440
rect -2945 -1535 -2715 -1440
rect -2595 -1535 -2365 -1440
rect -2245 -1535 -2015 -1440
rect -1895 -1535 -1665 -1440
rect -1545 -1535 -1315 -1305
rect -1195 -1535 -965 -1305
rect -845 -1535 -615 -1305
rect -495 -1535 -265 -1305
rect -145 -1535 85 -1305
rect 205 -1535 435 -1305
rect 555 -1535 785 -1305
rect 905 -1535 1135 -1305
rect 1255 -1535 1485 -1305
rect 1605 -1535 1835 -1305
rect 1955 -1535 2185 -1305
rect 2305 -1535 2535 -1305
rect 2655 -1535 2885 -1305
rect 3005 -1535 3235 -1305
rect 3355 -1390 3585 -1305
rect 3705 -1390 3935 -1305
rect 4055 -1390 4285 -1305
rect 4405 -1390 4635 -1305
rect 4755 -1390 4985 -1305
rect 3355 -1440 4985 -1390
rect 3355 -1535 3585 -1440
rect 3705 -1535 3935 -1440
rect 4055 -1535 4285 -1440
rect 4405 -1535 4635 -1440
rect 4755 -1535 4985 -1440
rect -2505 -1655 -2455 -1535
rect -1455 -1655 -1405 -1535
rect -1105 -1655 -1055 -1535
rect -755 -1655 -705 -1535
rect -405 -1655 -355 -1535
rect -55 -1655 -5 -1535
rect 295 -1655 345 -1535
rect 645 -1655 695 -1535
rect 995 -1655 1045 -1535
rect 1345 -1655 1395 -1535
rect 1695 -1655 1745 -1535
rect 2045 -1655 2095 -1535
rect 2395 -1655 2445 -1535
rect 2745 -1655 2795 -1535
rect 3095 -1655 3145 -1535
rect 4145 -1655 4195 -1535
rect -3295 -1740 -3065 -1655
rect -2945 -1740 -2715 -1655
rect -2595 -1740 -2365 -1655
rect -2245 -1740 -2015 -1655
rect -1895 -1740 -1665 -1655
rect -1545 -1740 -1315 -1655
rect -1195 -1740 -965 -1655
rect -845 -1740 -615 -1655
rect -495 -1740 -265 -1655
rect -145 -1740 85 -1655
rect 205 -1740 435 -1655
rect 555 -1740 785 -1655
rect -3295 -1790 785 -1740
rect -3295 -1885 -3065 -1790
rect -2945 -1885 -2715 -1790
rect -2595 -1885 -2365 -1790
rect -2245 -1885 -2015 -1790
rect -1895 -1885 -1665 -1790
rect -1545 -1885 -1315 -1790
rect -1195 -1885 -965 -1790
rect -845 -1885 -615 -1790
rect -495 -1885 -265 -1790
rect -145 -1885 85 -1790
rect 205 -1885 435 -1790
rect 555 -1885 785 -1790
rect 905 -1740 1135 -1655
rect 1255 -1740 1485 -1655
rect 1605 -1740 1835 -1655
rect 1955 -1740 2185 -1655
rect 2305 -1740 2535 -1655
rect 2655 -1740 2885 -1655
rect 3005 -1740 3235 -1655
rect 3355 -1740 3585 -1655
rect 3705 -1740 3935 -1655
rect 4055 -1740 4285 -1655
rect 4405 -1740 4635 -1655
rect 4755 -1740 4985 -1655
rect 905 -1790 4985 -1740
rect 905 -1885 1135 -1790
rect 1255 -1885 1485 -1790
rect 1605 -1885 1835 -1790
rect 1955 -1885 2185 -1790
rect 2305 -1885 2535 -1790
rect 2655 -1885 2885 -1790
rect 3005 -1885 3235 -1790
rect 3355 -1885 3585 -1790
rect 3705 -1885 3935 -1790
rect 4055 -1885 4285 -1790
rect 4405 -1885 4635 -1790
rect 4755 -1885 4985 -1790
rect -2505 -2005 -2455 -1885
rect -2155 -2005 -2105 -1885
rect -1805 -2005 -1755 -1885
rect -1455 -2005 -1405 -1885
rect -1105 -2005 -1055 -1885
rect -755 -2005 -705 -1885
rect -405 -2005 -355 -1885
rect -55 -2005 -5 -1885
rect 295 -2005 345 -1885
rect 645 -2005 695 -1885
rect 995 -2005 1045 -1885
rect 1345 -2005 1395 -1885
rect 1695 -2005 1745 -1885
rect 2045 -2005 2095 -1885
rect 2395 -2005 2445 -1885
rect 2745 -2005 2795 -1885
rect 3095 -2005 3145 -1885
rect 3445 -2005 3495 -1885
rect 3795 -2005 3845 -1885
rect 4145 -2005 4195 -1885
rect -3295 -2090 -3065 -2005
rect -2945 -2090 -2715 -2005
rect -2595 -2090 -2365 -2005
rect -3295 -2140 -2365 -2090
rect -3295 -2235 -3065 -2140
rect -2945 -2235 -2715 -2140
rect -2595 -2235 -2365 -2140
rect -2245 -2235 -2015 -2005
rect -1895 -2235 -1665 -2005
rect -1545 -2235 -1315 -2005
rect -1195 -2235 -965 -2005
rect -845 -2235 -615 -2005
rect -495 -2235 -265 -2005
rect -145 -2235 85 -2005
rect 205 -2235 435 -2005
rect 555 -2235 785 -2005
rect 905 -2235 1135 -2005
rect 1255 -2235 1485 -2005
rect 1605 -2235 1835 -2005
rect 1955 -2235 2185 -2005
rect 2305 -2235 2535 -2005
rect 2655 -2235 2885 -2005
rect 3005 -2235 3235 -2005
rect 3355 -2235 3585 -2005
rect 3705 -2235 3935 -2005
rect 4055 -2090 4285 -2005
rect 4405 -2090 4635 -2005
rect 4755 -2090 4985 -2005
rect 4055 -2140 4985 -2090
rect 4055 -2235 4285 -2140
rect 4405 -2235 4635 -2140
rect 4755 -2235 4985 -2140
rect 820 -2420 870 -2415
rect 820 -2460 825 -2420
rect 865 -2460 870 -2420
rect 820 -2465 870 -2460
<< via3 >>
rect 825 4275 865 4280
rect 825 4245 830 4275
rect 830 4245 860 4275
rect 860 4245 865 4275
rect 825 4240 865 4245
rect -1540 350 -1500 355
rect -1540 320 -1535 350
rect -1535 320 -1505 350
rect -1505 320 -1500 350
rect -1540 315 -1500 320
rect 3190 350 3230 355
rect 3190 320 3195 350
rect 3195 320 3225 350
rect 3225 320 3230 350
rect 3190 315 3230 320
rect 825 -2425 865 -2420
rect 825 -2455 830 -2425
rect 830 -2455 860 -2425
rect 860 -2455 865 -2425
rect 825 -2460 865 -2455
<< mimcap >>
rect -3280 3855 -3080 3930
rect -3280 3815 -3200 3855
rect -3160 3815 -3080 3855
rect -3280 3730 -3080 3815
rect -2930 3855 -2730 3930
rect -2930 3815 -2850 3855
rect -2810 3815 -2730 3855
rect -2930 3730 -2730 3815
rect -2580 3855 -2380 3930
rect -2580 3815 -2500 3855
rect -2460 3815 -2380 3855
rect -2580 3730 -2380 3815
rect -2230 3855 -2030 3930
rect -2230 3815 -2150 3855
rect -2110 3815 -2030 3855
rect -2230 3730 -2030 3815
rect -1880 3855 -1680 3930
rect -1880 3815 -1800 3855
rect -1760 3815 -1680 3855
rect -1880 3730 -1680 3815
rect -1530 3855 -1330 3930
rect -1530 3815 -1450 3855
rect -1410 3815 -1330 3855
rect -1530 3730 -1330 3815
rect -1180 3855 -980 3930
rect -1180 3815 -1100 3855
rect -1060 3815 -980 3855
rect -1180 3730 -980 3815
rect -830 3855 -630 3930
rect -830 3815 -750 3855
rect -710 3815 -630 3855
rect -830 3730 -630 3815
rect -480 3855 -280 3930
rect -480 3815 -400 3855
rect -360 3815 -280 3855
rect -480 3730 -280 3815
rect -130 3855 70 3930
rect -130 3815 -50 3855
rect -10 3815 70 3855
rect -130 3730 70 3815
rect 220 3855 420 3930
rect 220 3815 300 3855
rect 340 3815 420 3855
rect 220 3730 420 3815
rect 570 3855 770 3930
rect 570 3815 650 3855
rect 690 3815 770 3855
rect 570 3730 770 3815
rect 920 3855 1120 3930
rect 920 3815 1000 3855
rect 1040 3815 1120 3855
rect 920 3730 1120 3815
rect 1270 3855 1470 3930
rect 1270 3815 1350 3855
rect 1390 3815 1470 3855
rect 1270 3730 1470 3815
rect 1620 3855 1820 3930
rect 1620 3815 1700 3855
rect 1740 3815 1820 3855
rect 1620 3730 1820 3815
rect 1970 3855 2170 3930
rect 1970 3815 2050 3855
rect 2090 3815 2170 3855
rect 1970 3730 2170 3815
rect 2320 3855 2520 3930
rect 2320 3815 2400 3855
rect 2440 3815 2520 3855
rect 2320 3730 2520 3815
rect 2670 3855 2870 3930
rect 2670 3815 2750 3855
rect 2790 3815 2870 3855
rect 2670 3730 2870 3815
rect 3020 3855 3220 3930
rect 3020 3815 3100 3855
rect 3140 3815 3220 3855
rect 3020 3730 3220 3815
rect 3370 3855 3570 3930
rect 3370 3815 3450 3855
rect 3490 3815 3570 3855
rect 3370 3730 3570 3815
rect 3720 3855 3920 3930
rect 3720 3815 3800 3855
rect 3840 3815 3920 3855
rect 3720 3730 3920 3815
rect 4070 3855 4270 3930
rect 4070 3815 4150 3855
rect 4190 3815 4270 3855
rect 4070 3730 4270 3815
rect 4420 3855 4620 3930
rect 4420 3815 4500 3855
rect 4540 3815 4620 3855
rect 4420 3730 4620 3815
rect 4770 3855 4970 3930
rect 4770 3815 4850 3855
rect 4890 3815 4970 3855
rect 4770 3730 4970 3815
rect -3280 3505 -3080 3580
rect -3280 3465 -3200 3505
rect -3160 3465 -3080 3505
rect -3280 3380 -3080 3465
rect -2930 3505 -2730 3580
rect -2930 3465 -2850 3505
rect -2810 3465 -2730 3505
rect -2930 3380 -2730 3465
rect -2580 3505 -2380 3580
rect -2580 3465 -2500 3505
rect -2460 3465 -2380 3505
rect -2580 3380 -2380 3465
rect -2230 3505 -2030 3580
rect -2230 3465 -2150 3505
rect -2110 3465 -2030 3505
rect -2230 3380 -2030 3465
rect -1880 3505 -1680 3580
rect -1880 3465 -1800 3505
rect -1760 3465 -1680 3505
rect -1880 3380 -1680 3465
rect -1530 3505 -1330 3580
rect -1530 3465 -1450 3505
rect -1410 3465 -1330 3505
rect -1530 3380 -1330 3465
rect -1180 3505 -980 3580
rect -1180 3465 -1100 3505
rect -1060 3465 -980 3505
rect -1180 3380 -980 3465
rect -830 3505 -630 3580
rect -830 3465 -750 3505
rect -710 3465 -630 3505
rect -830 3380 -630 3465
rect -480 3505 -280 3580
rect -480 3465 -400 3505
rect -360 3465 -280 3505
rect -480 3380 -280 3465
rect -130 3505 70 3580
rect -130 3465 -50 3505
rect -10 3465 70 3505
rect -130 3380 70 3465
rect 220 3505 420 3580
rect 220 3465 300 3505
rect 340 3465 420 3505
rect 220 3380 420 3465
rect 570 3505 770 3580
rect 570 3465 650 3505
rect 690 3465 770 3505
rect 570 3380 770 3465
rect 920 3505 1120 3580
rect 920 3465 1000 3505
rect 1040 3465 1120 3505
rect 920 3380 1120 3465
rect 1270 3505 1470 3580
rect 1270 3465 1350 3505
rect 1390 3465 1470 3505
rect 1270 3380 1470 3465
rect 1620 3505 1820 3580
rect 1620 3465 1700 3505
rect 1740 3465 1820 3505
rect 1620 3380 1820 3465
rect 1970 3505 2170 3580
rect 1970 3465 2050 3505
rect 2090 3465 2170 3505
rect 1970 3380 2170 3465
rect 2320 3505 2520 3580
rect 2320 3465 2400 3505
rect 2440 3465 2520 3505
rect 2320 3380 2520 3465
rect 2670 3505 2870 3580
rect 2670 3465 2750 3505
rect 2790 3465 2870 3505
rect 2670 3380 2870 3465
rect 3020 3505 3220 3580
rect 3020 3465 3100 3505
rect 3140 3465 3220 3505
rect 3020 3380 3220 3465
rect 3370 3505 3570 3580
rect 3370 3465 3450 3505
rect 3490 3465 3570 3505
rect 3370 3380 3570 3465
rect 3720 3505 3920 3580
rect 3720 3465 3800 3505
rect 3840 3465 3920 3505
rect 3720 3380 3920 3465
rect 4070 3505 4270 3580
rect 4070 3465 4150 3505
rect 4190 3465 4270 3505
rect 4070 3380 4270 3465
rect 4420 3505 4620 3580
rect 4420 3465 4500 3505
rect 4540 3465 4620 3505
rect 4420 3380 4620 3465
rect 4770 3505 4970 3580
rect 4770 3465 4850 3505
rect 4890 3465 4970 3505
rect 4770 3380 4970 3465
rect -3280 3155 -3080 3230
rect -3280 3115 -3200 3155
rect -3160 3115 -3080 3155
rect -3280 3030 -3080 3115
rect -2930 3155 -2730 3230
rect -2930 3115 -2850 3155
rect -2810 3115 -2730 3155
rect -2930 3030 -2730 3115
rect -2580 3155 -2380 3230
rect -2580 3115 -2500 3155
rect -2460 3115 -2380 3155
rect -2580 3030 -2380 3115
rect -2230 3155 -2030 3230
rect -2230 3115 -2150 3155
rect -2110 3115 -2030 3155
rect -2230 3030 -2030 3115
rect -1880 3155 -1680 3230
rect -1880 3115 -1800 3155
rect -1760 3115 -1680 3155
rect -1880 3030 -1680 3115
rect -1530 3155 -1330 3230
rect -1530 3115 -1450 3155
rect -1410 3115 -1330 3155
rect -1530 3030 -1330 3115
rect -1180 3155 -980 3230
rect -1180 3115 -1100 3155
rect -1060 3115 -980 3155
rect -1180 3030 -980 3115
rect -830 3155 -630 3230
rect -830 3115 -750 3155
rect -710 3115 -630 3155
rect -830 3030 -630 3115
rect -480 3155 -280 3230
rect -480 3115 -400 3155
rect -360 3115 -280 3155
rect -480 3030 -280 3115
rect -130 3145 70 3230
rect -130 3105 -50 3145
rect -10 3105 70 3145
rect -130 3030 70 3105
rect 220 3145 420 3230
rect 220 3105 300 3145
rect 340 3105 420 3145
rect 220 3030 420 3105
rect 570 3145 770 3230
rect 570 3105 650 3145
rect 690 3105 770 3145
rect 570 3030 770 3105
rect 920 3145 1120 3230
rect 920 3105 1000 3145
rect 1040 3105 1120 3145
rect 920 3030 1120 3105
rect 1270 3145 1470 3230
rect 1270 3105 1350 3145
rect 1390 3105 1470 3145
rect 1270 3030 1470 3105
rect 1620 3145 1820 3230
rect 1620 3105 1700 3145
rect 1740 3105 1820 3145
rect 1620 3030 1820 3105
rect 1970 3155 2170 3230
rect 1970 3115 2050 3155
rect 2090 3115 2170 3155
rect 1970 3030 2170 3115
rect 2320 3155 2520 3230
rect 2320 3115 2400 3155
rect 2440 3115 2520 3155
rect 2320 3030 2520 3115
rect 2670 3155 2870 3230
rect 2670 3115 2750 3155
rect 2790 3115 2870 3155
rect 2670 3030 2870 3115
rect 3020 3155 3220 3230
rect 3020 3115 3100 3155
rect 3140 3115 3220 3155
rect 3020 3030 3220 3115
rect 3370 3155 3570 3230
rect 3370 3115 3450 3155
rect 3490 3115 3570 3155
rect 3370 3030 3570 3115
rect 3720 3155 3920 3230
rect 3720 3115 3800 3155
rect 3840 3115 3920 3155
rect 3720 3030 3920 3115
rect 4070 3155 4270 3230
rect 4070 3115 4150 3155
rect 4190 3115 4270 3155
rect 4070 3030 4270 3115
rect 4420 3155 4620 3230
rect 4420 3115 4500 3155
rect 4540 3115 4620 3155
rect 4420 3030 4620 3115
rect 4770 3155 4970 3230
rect 4770 3115 4850 3155
rect 4890 3115 4970 3155
rect 4770 3030 4970 3115
rect -3280 2805 -3080 2880
rect -3280 2765 -3200 2805
rect -3160 2765 -3080 2805
rect -3280 2680 -3080 2765
rect -2930 2805 -2730 2880
rect -2930 2765 -2850 2805
rect -2810 2765 -2730 2805
rect -2930 2680 -2730 2765
rect -2580 2805 -2380 2880
rect -2580 2765 -2500 2805
rect -2460 2765 -2380 2805
rect -2580 2680 -2380 2765
rect -2230 2805 -2030 2880
rect -2230 2765 -2150 2805
rect -2110 2765 -2030 2805
rect -2230 2680 -2030 2765
rect -1880 2805 -1680 2880
rect -1880 2765 -1800 2805
rect -1760 2765 -1680 2805
rect -1880 2680 -1680 2765
rect -1530 2805 -1330 2880
rect -1530 2765 -1450 2805
rect -1410 2765 -1330 2805
rect -1530 2680 -1330 2765
rect -1180 2805 -980 2880
rect -1180 2765 -1100 2805
rect -1060 2765 -980 2805
rect -1180 2680 -980 2765
rect -830 2805 -630 2880
rect -830 2765 -750 2805
rect -710 2765 -630 2805
rect -830 2680 -630 2765
rect 2320 2805 2520 2880
rect 2320 2765 2400 2805
rect 2440 2765 2520 2805
rect 2320 2680 2520 2765
rect 2670 2805 2870 2880
rect 2670 2765 2750 2805
rect 2790 2765 2870 2805
rect 2670 2680 2870 2765
rect 3020 2805 3220 2880
rect 3020 2765 3100 2805
rect 3140 2765 3220 2805
rect 3020 2680 3220 2765
rect 3370 2805 3570 2880
rect 3370 2765 3450 2805
rect 3490 2765 3570 2805
rect 3370 2680 3570 2765
rect 3720 2805 3920 2880
rect 3720 2765 3800 2805
rect 3840 2765 3920 2805
rect 3720 2680 3920 2765
rect 4070 2805 4270 2880
rect 4070 2765 4150 2805
rect 4190 2765 4270 2805
rect 4070 2680 4270 2765
rect 4420 2805 4620 2880
rect 4420 2765 4500 2805
rect 4540 2765 4620 2805
rect 4420 2680 4620 2765
rect 4770 2805 4970 2880
rect 4770 2765 4850 2805
rect 4890 2765 4970 2805
rect 4770 2680 4970 2765
rect -3280 2455 -3080 2530
rect -3280 2415 -3200 2455
rect -3160 2415 -3080 2455
rect -3280 2330 -3080 2415
rect -2930 2455 -2730 2530
rect -2930 2415 -2850 2455
rect -2810 2415 -2730 2455
rect -2930 2330 -2730 2415
rect -2580 2455 -2380 2530
rect -2580 2415 -2500 2455
rect -2460 2415 -2380 2455
rect -2580 2330 -2380 2415
rect -2230 2455 -2030 2530
rect -2230 2415 -2150 2455
rect -2110 2415 -2030 2455
rect -2230 2330 -2030 2415
rect -1880 2455 -1680 2530
rect -1880 2415 -1800 2455
rect -1760 2415 -1680 2455
rect -1880 2330 -1680 2415
rect -1530 2455 -1330 2530
rect -1530 2415 -1450 2455
rect -1410 2415 -1330 2455
rect -1530 2330 -1330 2415
rect -1180 2455 -980 2530
rect -1180 2415 -1100 2455
rect -1060 2415 -980 2455
rect -1180 2330 -980 2415
rect -830 2455 -630 2530
rect -830 2415 -750 2455
rect -710 2415 -630 2455
rect -830 2330 -630 2415
rect 2320 2455 2520 2530
rect 2320 2415 2400 2455
rect 2440 2415 2520 2455
rect 2320 2330 2520 2415
rect 2670 2455 2870 2530
rect 2670 2415 2750 2455
rect 2790 2415 2870 2455
rect 2670 2330 2870 2415
rect 3020 2455 3220 2530
rect 3020 2415 3100 2455
rect 3140 2415 3220 2455
rect 3020 2330 3220 2415
rect 3370 2455 3570 2530
rect 3370 2415 3450 2455
rect 3490 2415 3570 2455
rect 3370 2330 3570 2415
rect 3720 2455 3920 2530
rect 3720 2415 3800 2455
rect 3840 2415 3920 2455
rect 3720 2330 3920 2415
rect 4070 2455 4270 2530
rect 4070 2415 4150 2455
rect 4190 2415 4270 2455
rect 4070 2330 4270 2415
rect 4420 2455 4620 2530
rect 4420 2415 4500 2455
rect 4540 2415 4620 2455
rect 4420 2330 4620 2415
rect 4770 2455 4970 2530
rect 4770 2415 4850 2455
rect 4890 2415 4970 2455
rect 4770 2330 4970 2415
rect -3280 2105 -3080 2180
rect -3280 2065 -3200 2105
rect -3160 2065 -3080 2105
rect -3280 1980 -3080 2065
rect -2930 2105 -2730 2180
rect -2930 2065 -2850 2105
rect -2810 2065 -2730 2105
rect -2930 1980 -2730 2065
rect -2580 2105 -2380 2180
rect -2580 2065 -2500 2105
rect -2460 2065 -2380 2105
rect -2580 1980 -2380 2065
rect -2230 2105 -2030 2180
rect -2230 2065 -2150 2105
rect -2110 2065 -2030 2105
rect -2230 1980 -2030 2065
rect -1880 2105 -1680 2180
rect -1880 2065 -1800 2105
rect -1760 2065 -1680 2105
rect -1880 1980 -1680 2065
rect 3370 2105 3570 2180
rect 3370 2065 3450 2105
rect 3490 2065 3570 2105
rect 3370 1980 3570 2065
rect 3720 2105 3920 2180
rect 3720 2065 3800 2105
rect 3840 2065 3920 2105
rect 3720 1980 3920 2065
rect 4070 2105 4270 2180
rect 4070 2065 4150 2105
rect 4190 2065 4270 2105
rect 4070 1980 4270 2065
rect 4420 2105 4620 2180
rect 4420 2065 4500 2105
rect 4540 2065 4620 2105
rect 4420 1980 4620 2065
rect 4770 2105 4970 2180
rect 4770 2065 4850 2105
rect 4890 2065 4970 2105
rect 4770 1980 4970 2065
rect -3280 1755 -3080 1830
rect -3280 1715 -3200 1755
rect -3160 1715 -3080 1755
rect -3280 1630 -3080 1715
rect -2930 1755 -2730 1830
rect -2930 1715 -2850 1755
rect -2810 1715 -2730 1755
rect -2930 1630 -2730 1715
rect -2580 1755 -2380 1830
rect -2580 1715 -2500 1755
rect -2460 1715 -2380 1755
rect -2580 1630 -2380 1715
rect -2230 1755 -2030 1830
rect -2230 1715 -2150 1755
rect -2110 1715 -2030 1755
rect -2230 1630 -2030 1715
rect -1880 1755 -1680 1830
rect -1880 1715 -1800 1755
rect -1760 1715 -1680 1755
rect -1880 1630 -1680 1715
rect 3370 1755 3570 1830
rect 3370 1715 3450 1755
rect 3490 1715 3570 1755
rect 3370 1630 3570 1715
rect 3720 1755 3920 1830
rect 3720 1715 3800 1755
rect 3840 1715 3920 1755
rect 3720 1630 3920 1715
rect 4070 1755 4270 1830
rect 4070 1715 4150 1755
rect 4190 1715 4270 1755
rect 4070 1630 4270 1715
rect 4420 1755 4620 1830
rect 4420 1715 4500 1755
rect 4540 1715 4620 1755
rect 4420 1630 4620 1715
rect 4770 1755 4970 1830
rect 4770 1715 4850 1755
rect 4890 1715 4970 1755
rect 4770 1630 4970 1715
rect -3280 1405 -3080 1480
rect -3280 1365 -3200 1405
rect -3160 1365 -3080 1405
rect -3280 1280 -3080 1365
rect -2930 1405 -2730 1480
rect -2930 1365 -2850 1405
rect -2810 1365 -2730 1405
rect -2930 1280 -2730 1365
rect -2580 1405 -2380 1480
rect -2580 1365 -2500 1405
rect -2460 1365 -2380 1405
rect -2580 1280 -2380 1365
rect -2230 1405 -2030 1480
rect -2230 1365 -2150 1405
rect -2110 1365 -2030 1405
rect -2230 1280 -2030 1365
rect -1880 1405 -1680 1480
rect -1880 1365 -1800 1405
rect -1760 1365 -1680 1405
rect -1880 1280 -1680 1365
rect 3370 1405 3570 1480
rect 3370 1365 3450 1405
rect 3490 1365 3570 1405
rect 3370 1280 3570 1365
rect 3720 1405 3920 1480
rect 3720 1365 3800 1405
rect 3840 1365 3920 1405
rect 3720 1280 3920 1365
rect 4070 1405 4270 1480
rect 4070 1365 4150 1405
rect 4190 1365 4270 1405
rect 4070 1280 4270 1365
rect 4420 1405 4620 1480
rect 4420 1365 4500 1405
rect 4540 1365 4620 1405
rect 4420 1280 4620 1365
rect 4770 1405 4970 1480
rect 4770 1365 4850 1405
rect 4890 1365 4970 1405
rect 4770 1280 4970 1365
rect -3280 1055 -3080 1130
rect -3280 1015 -3200 1055
rect -3160 1015 -3080 1055
rect -3280 930 -3080 1015
rect -2930 1055 -2730 1130
rect -2930 1015 -2850 1055
rect -2810 1015 -2730 1055
rect -2930 930 -2730 1015
rect -2580 1055 -2380 1130
rect -2580 1015 -2500 1055
rect -2460 1015 -2380 1055
rect -2580 930 -2380 1015
rect -2230 1055 -2030 1130
rect -2230 1015 -2150 1055
rect -2110 1015 -2030 1055
rect -2230 930 -2030 1015
rect -1880 1055 -1680 1130
rect -1880 1015 -1800 1055
rect -1760 1015 -1680 1055
rect -1880 930 -1680 1015
rect 3370 1055 3570 1130
rect 3370 1015 3450 1055
rect 3490 1015 3570 1055
rect 3370 930 3570 1015
rect 3720 1055 3920 1130
rect 3720 1015 3800 1055
rect 3840 1015 3920 1055
rect 3720 930 3920 1015
rect 4070 1055 4270 1130
rect 4070 1015 4150 1055
rect 4190 1015 4270 1055
rect 4070 930 4270 1015
rect 4420 1055 4620 1130
rect 4420 1015 4500 1055
rect 4540 1015 4620 1055
rect 4420 930 4620 1015
rect 4770 1055 4970 1130
rect 4770 1015 4850 1055
rect 4890 1015 4970 1055
rect 4770 930 4970 1015
rect -3280 705 -3080 780
rect -3280 665 -3200 705
rect -3160 665 -3080 705
rect -3280 580 -3080 665
rect -2930 705 -2730 780
rect -2930 665 -2850 705
rect -2810 665 -2730 705
rect -2930 580 -2730 665
rect -2580 705 -2380 780
rect -2580 665 -2500 705
rect -2460 665 -2380 705
rect -2580 580 -2380 665
rect -2230 705 -2030 780
rect -2230 665 -2150 705
rect -2110 665 -2030 705
rect -2230 580 -2030 665
rect -1880 705 -1680 780
rect -1880 665 -1800 705
rect -1760 665 -1680 705
rect -1880 580 -1680 665
rect 3370 705 3570 780
rect 3370 665 3450 705
rect 3490 665 3570 705
rect 3370 580 3570 665
rect 3720 705 3920 780
rect 3720 665 3800 705
rect 3840 665 3920 705
rect 3720 580 3920 665
rect 4070 705 4270 780
rect 4070 665 4150 705
rect 4190 665 4270 705
rect 4070 580 4270 665
rect 4420 705 4620 780
rect 4420 665 4500 705
rect 4540 665 4620 705
rect 4420 580 4620 665
rect 4770 705 4970 780
rect 4770 665 4850 705
rect 4890 665 4970 705
rect 4770 580 4970 665
rect -3280 355 -3080 430
rect -3280 315 -3200 355
rect -3160 315 -3080 355
rect -3280 230 -3080 315
rect -2930 355 -2730 430
rect -2930 315 -2850 355
rect -2810 315 -2730 355
rect -2930 230 -2730 315
rect -2580 355 -2380 430
rect -2580 315 -2500 355
rect -2460 315 -2380 355
rect -2580 230 -2380 315
rect -2230 355 -2030 430
rect -2230 315 -2150 355
rect -2110 315 -2030 355
rect -2230 230 -2030 315
rect -1880 355 -1680 430
rect -1880 315 -1800 355
rect -1760 315 -1680 355
rect -1880 230 -1680 315
rect 3370 355 3570 430
rect 3370 315 3450 355
rect 3490 315 3570 355
rect 3370 230 3570 315
rect 3720 355 3920 430
rect 3720 315 3800 355
rect 3840 315 3920 355
rect 3720 230 3920 315
rect 4070 355 4270 430
rect 4070 315 4150 355
rect 4190 315 4270 355
rect 4070 230 4270 315
rect 4420 355 4620 430
rect 4420 315 4500 355
rect 4540 315 4620 355
rect 4420 230 4620 315
rect 4770 355 4970 430
rect 4770 315 4850 355
rect 4890 315 4970 355
rect 4770 230 4970 315
rect -3280 5 -3080 80
rect -3280 -35 -3200 5
rect -3160 -35 -3080 5
rect -3280 -120 -3080 -35
rect -2930 5 -2730 80
rect -2930 -35 -2850 5
rect -2810 -35 -2730 5
rect -2930 -120 -2730 -35
rect -2580 5 -2380 80
rect -2580 -35 -2500 5
rect -2460 -35 -2380 5
rect -2580 -120 -2380 -35
rect -2230 5 -2030 80
rect -2230 -35 -2150 5
rect -2110 -35 -2030 5
rect -2230 -120 -2030 -35
rect -1880 5 -1680 80
rect -1880 -35 -1800 5
rect -1760 -35 -1680 5
rect -1880 -120 -1680 -35
rect 3370 5 3570 80
rect 3370 -35 3450 5
rect 3490 -35 3570 5
rect 3370 -120 3570 -35
rect 3720 5 3920 80
rect 3720 -35 3800 5
rect 3840 -35 3920 5
rect 3720 -120 3920 -35
rect 4070 5 4270 80
rect 4070 -35 4150 5
rect 4190 -35 4270 5
rect 4070 -120 4270 -35
rect 4420 5 4620 80
rect 4420 -35 4500 5
rect 4540 -35 4620 5
rect 4420 -120 4620 -35
rect 4770 5 4970 80
rect 4770 -35 4850 5
rect 4890 -35 4970 5
rect 4770 -120 4970 -35
rect -3280 -345 -3080 -270
rect -3280 -385 -3200 -345
rect -3160 -385 -3080 -345
rect -3280 -470 -3080 -385
rect -2930 -345 -2730 -270
rect -2930 -385 -2850 -345
rect -2810 -385 -2730 -345
rect -2930 -470 -2730 -385
rect -2580 -345 -2380 -270
rect -2580 -385 -2500 -345
rect -2460 -385 -2380 -345
rect -2580 -470 -2380 -385
rect -2230 -345 -2030 -270
rect -2230 -385 -2150 -345
rect -2110 -385 -2030 -345
rect -2230 -470 -2030 -385
rect -1880 -345 -1680 -270
rect -1880 -385 -1800 -345
rect -1760 -385 -1680 -345
rect -1880 -470 -1680 -385
rect 3370 -345 3570 -270
rect 3370 -385 3450 -345
rect 3490 -385 3570 -345
rect 3370 -470 3570 -385
rect 3720 -345 3920 -270
rect 3720 -385 3800 -345
rect 3840 -385 3920 -345
rect 3720 -470 3920 -385
rect 4070 -345 4270 -270
rect 4070 -385 4150 -345
rect 4190 -385 4270 -345
rect 4070 -470 4270 -385
rect 4420 -345 4620 -270
rect 4420 -385 4500 -345
rect 4540 -385 4620 -345
rect 4420 -470 4620 -385
rect 4770 -345 4970 -270
rect 4770 -385 4850 -345
rect 4890 -385 4970 -345
rect 4770 -470 4970 -385
rect -3280 -695 -3080 -620
rect -3280 -735 -3200 -695
rect -3160 -735 -3080 -695
rect -3280 -820 -3080 -735
rect -2930 -695 -2730 -620
rect -2930 -735 -2850 -695
rect -2810 -735 -2730 -695
rect -2930 -820 -2730 -735
rect -2580 -695 -2380 -620
rect -2580 -735 -2500 -695
rect -2460 -735 -2380 -695
rect -2580 -820 -2380 -735
rect -2230 -695 -2030 -620
rect -2230 -735 -2150 -695
rect -2110 -735 -2030 -695
rect -2230 -820 -2030 -735
rect -1880 -695 -1680 -620
rect -1880 -735 -1800 -695
rect -1760 -735 -1680 -695
rect -1880 -820 -1680 -735
rect 3370 -695 3570 -620
rect 3370 -735 3450 -695
rect 3490 -735 3570 -695
rect 3370 -820 3570 -735
rect 3720 -695 3920 -620
rect 3720 -735 3800 -695
rect 3840 -735 3920 -695
rect 3720 -820 3920 -735
rect 4070 -695 4270 -620
rect 4070 -735 4150 -695
rect 4190 -735 4270 -695
rect 4070 -820 4270 -735
rect 4420 -695 4620 -620
rect 4420 -735 4500 -695
rect 4540 -735 4620 -695
rect 4420 -820 4620 -735
rect 4770 -695 4970 -620
rect 4770 -735 4850 -695
rect 4890 -735 4970 -695
rect 4770 -820 4970 -735
rect -3280 -1045 -3080 -970
rect -3280 -1085 -3200 -1045
rect -3160 -1085 -3080 -1045
rect -3280 -1170 -3080 -1085
rect -2930 -1045 -2730 -970
rect -2930 -1085 -2850 -1045
rect -2810 -1085 -2730 -1045
rect -2930 -1170 -2730 -1085
rect -2580 -1045 -2380 -970
rect -2580 -1085 -2500 -1045
rect -2460 -1085 -2380 -1045
rect -2580 -1170 -2380 -1085
rect -2230 -1045 -2030 -970
rect -2230 -1085 -2150 -1045
rect -2110 -1085 -2030 -1045
rect -2230 -1170 -2030 -1085
rect -1880 -1045 -1680 -970
rect -1880 -1085 -1800 -1045
rect -1760 -1085 -1680 -1045
rect -1880 -1170 -1680 -1085
rect 3370 -1045 3570 -970
rect 3370 -1085 3450 -1045
rect 3490 -1085 3570 -1045
rect 3370 -1170 3570 -1085
rect 3720 -1045 3920 -970
rect 3720 -1085 3800 -1045
rect 3840 -1085 3920 -1045
rect 3720 -1170 3920 -1085
rect 4070 -1045 4270 -970
rect 4070 -1085 4150 -1045
rect 4190 -1085 4270 -1045
rect 4070 -1170 4270 -1085
rect 4420 -1045 4620 -970
rect 4420 -1085 4500 -1045
rect 4540 -1085 4620 -1045
rect 4420 -1170 4620 -1085
rect 4770 -1045 4970 -970
rect 4770 -1085 4850 -1045
rect 4890 -1085 4970 -1045
rect 4770 -1170 4970 -1085
rect -3280 -1395 -3080 -1320
rect -3280 -1435 -3200 -1395
rect -3160 -1435 -3080 -1395
rect -3280 -1520 -3080 -1435
rect -2930 -1395 -2730 -1320
rect -2930 -1435 -2850 -1395
rect -2810 -1435 -2730 -1395
rect -2930 -1520 -2730 -1435
rect -2580 -1395 -2380 -1320
rect -2580 -1435 -2500 -1395
rect -2460 -1435 -2380 -1395
rect -2580 -1520 -2380 -1435
rect -2230 -1395 -2030 -1320
rect -2230 -1435 -2150 -1395
rect -2110 -1435 -2030 -1395
rect -2230 -1520 -2030 -1435
rect -1880 -1395 -1680 -1320
rect -1880 -1435 -1800 -1395
rect -1760 -1435 -1680 -1395
rect -1880 -1520 -1680 -1435
rect -1530 -1395 -1330 -1320
rect -1530 -1435 -1450 -1395
rect -1410 -1435 -1330 -1395
rect -1530 -1520 -1330 -1435
rect -1180 -1395 -980 -1320
rect -1180 -1435 -1100 -1395
rect -1060 -1435 -980 -1395
rect -1180 -1520 -980 -1435
rect -830 -1395 -630 -1320
rect -830 -1435 -750 -1395
rect -710 -1435 -630 -1395
rect -830 -1520 -630 -1435
rect -480 -1395 -280 -1320
rect -480 -1435 -400 -1395
rect -360 -1435 -280 -1395
rect -480 -1520 -280 -1435
rect -130 -1395 70 -1320
rect -130 -1435 -50 -1395
rect -10 -1435 70 -1395
rect -130 -1520 70 -1435
rect 220 -1395 420 -1320
rect 220 -1435 300 -1395
rect 340 -1435 420 -1395
rect 220 -1520 420 -1435
rect 570 -1395 770 -1320
rect 570 -1435 650 -1395
rect 690 -1435 770 -1395
rect 570 -1520 770 -1435
rect 920 -1395 1120 -1320
rect 920 -1435 1000 -1395
rect 1040 -1435 1120 -1395
rect 920 -1520 1120 -1435
rect 1270 -1395 1470 -1320
rect 1270 -1435 1350 -1395
rect 1390 -1435 1470 -1395
rect 1270 -1520 1470 -1435
rect 1620 -1395 1820 -1320
rect 1620 -1435 1700 -1395
rect 1740 -1435 1820 -1395
rect 1620 -1520 1820 -1435
rect 1970 -1395 2170 -1320
rect 1970 -1435 2050 -1395
rect 2090 -1435 2170 -1395
rect 1970 -1520 2170 -1435
rect 2320 -1395 2520 -1320
rect 2320 -1435 2400 -1395
rect 2440 -1435 2520 -1395
rect 2320 -1520 2520 -1435
rect 2670 -1395 2870 -1320
rect 2670 -1435 2750 -1395
rect 2790 -1435 2870 -1395
rect 2670 -1520 2870 -1435
rect 3020 -1395 3220 -1320
rect 3020 -1435 3100 -1395
rect 3140 -1435 3220 -1395
rect 3020 -1520 3220 -1435
rect 3370 -1395 3570 -1320
rect 3370 -1435 3450 -1395
rect 3490 -1435 3570 -1395
rect 3370 -1520 3570 -1435
rect 3720 -1395 3920 -1320
rect 3720 -1435 3800 -1395
rect 3840 -1435 3920 -1395
rect 3720 -1520 3920 -1435
rect 4070 -1395 4270 -1320
rect 4070 -1435 4150 -1395
rect 4190 -1435 4270 -1395
rect 4070 -1520 4270 -1435
rect 4420 -1395 4620 -1320
rect 4420 -1435 4500 -1395
rect 4540 -1435 4620 -1395
rect 4420 -1520 4620 -1435
rect 4770 -1395 4970 -1320
rect 4770 -1435 4850 -1395
rect 4890 -1435 4970 -1395
rect 4770 -1520 4970 -1435
rect -3280 -1745 -3080 -1670
rect -3280 -1785 -3200 -1745
rect -3160 -1785 -3080 -1745
rect -3280 -1870 -3080 -1785
rect -2930 -1745 -2730 -1670
rect -2930 -1785 -2850 -1745
rect -2810 -1785 -2730 -1745
rect -2930 -1870 -2730 -1785
rect -2580 -1745 -2380 -1670
rect -2580 -1785 -2500 -1745
rect -2460 -1785 -2380 -1745
rect -2580 -1870 -2380 -1785
rect -2230 -1745 -2030 -1670
rect -2230 -1785 -2150 -1745
rect -2110 -1785 -2030 -1745
rect -2230 -1870 -2030 -1785
rect -1880 -1745 -1680 -1670
rect -1880 -1785 -1800 -1745
rect -1760 -1785 -1680 -1745
rect -1880 -1870 -1680 -1785
rect -1530 -1745 -1330 -1670
rect -1530 -1785 -1450 -1745
rect -1410 -1785 -1330 -1745
rect -1530 -1870 -1330 -1785
rect -1180 -1745 -980 -1670
rect -1180 -1785 -1100 -1745
rect -1060 -1785 -980 -1745
rect -1180 -1870 -980 -1785
rect -830 -1745 -630 -1670
rect -830 -1785 -750 -1745
rect -710 -1785 -630 -1745
rect -830 -1870 -630 -1785
rect -480 -1745 -280 -1670
rect -480 -1785 -400 -1745
rect -360 -1785 -280 -1745
rect -480 -1870 -280 -1785
rect -130 -1745 70 -1670
rect -130 -1785 -50 -1745
rect -10 -1785 70 -1745
rect -130 -1870 70 -1785
rect 220 -1745 420 -1670
rect 220 -1785 300 -1745
rect 340 -1785 420 -1745
rect 220 -1870 420 -1785
rect 570 -1745 770 -1670
rect 570 -1785 650 -1745
rect 690 -1785 770 -1745
rect 570 -1870 770 -1785
rect 920 -1745 1120 -1670
rect 920 -1785 1000 -1745
rect 1040 -1785 1120 -1745
rect 920 -1870 1120 -1785
rect 1270 -1745 1470 -1670
rect 1270 -1785 1350 -1745
rect 1390 -1785 1470 -1745
rect 1270 -1870 1470 -1785
rect 1620 -1745 1820 -1670
rect 1620 -1785 1700 -1745
rect 1740 -1785 1820 -1745
rect 1620 -1870 1820 -1785
rect 1970 -1745 2170 -1670
rect 1970 -1785 2050 -1745
rect 2090 -1785 2170 -1745
rect 1970 -1870 2170 -1785
rect 2320 -1745 2520 -1670
rect 2320 -1785 2400 -1745
rect 2440 -1785 2520 -1745
rect 2320 -1870 2520 -1785
rect 2670 -1745 2870 -1670
rect 2670 -1785 2750 -1745
rect 2790 -1785 2870 -1745
rect 2670 -1870 2870 -1785
rect 3020 -1745 3220 -1670
rect 3020 -1785 3100 -1745
rect 3140 -1785 3220 -1745
rect 3020 -1870 3220 -1785
rect 3370 -1745 3570 -1670
rect 3370 -1785 3450 -1745
rect 3490 -1785 3570 -1745
rect 3370 -1870 3570 -1785
rect 3720 -1745 3920 -1670
rect 3720 -1785 3800 -1745
rect 3840 -1785 3920 -1745
rect 3720 -1870 3920 -1785
rect 4070 -1745 4270 -1670
rect 4070 -1785 4150 -1745
rect 4190 -1785 4270 -1745
rect 4070 -1870 4270 -1785
rect 4420 -1745 4620 -1670
rect 4420 -1785 4500 -1745
rect 4540 -1785 4620 -1745
rect 4420 -1870 4620 -1785
rect 4770 -1745 4970 -1670
rect 4770 -1785 4850 -1745
rect 4890 -1785 4970 -1745
rect 4770 -1870 4970 -1785
rect -3280 -2095 -3080 -2020
rect -3280 -2135 -3200 -2095
rect -3160 -2135 -3080 -2095
rect -3280 -2220 -3080 -2135
rect -2930 -2095 -2730 -2020
rect -2930 -2135 -2850 -2095
rect -2810 -2135 -2730 -2095
rect -2930 -2220 -2730 -2135
rect -2580 -2095 -2380 -2020
rect -2580 -2135 -2500 -2095
rect -2460 -2135 -2380 -2095
rect -2580 -2220 -2380 -2135
rect -2230 -2095 -2030 -2020
rect -2230 -2135 -2150 -2095
rect -2110 -2135 -2030 -2095
rect -2230 -2220 -2030 -2135
rect -1880 -2095 -1680 -2020
rect -1880 -2135 -1800 -2095
rect -1760 -2135 -1680 -2095
rect -1880 -2220 -1680 -2135
rect -1530 -2095 -1330 -2020
rect -1530 -2135 -1450 -2095
rect -1410 -2135 -1330 -2095
rect -1530 -2220 -1330 -2135
rect -1180 -2095 -980 -2020
rect -1180 -2135 -1100 -2095
rect -1060 -2135 -980 -2095
rect -1180 -2220 -980 -2135
rect -830 -2095 -630 -2020
rect -830 -2135 -750 -2095
rect -710 -2135 -630 -2095
rect -830 -2220 -630 -2135
rect -480 -2095 -280 -2020
rect -480 -2135 -400 -2095
rect -360 -2135 -280 -2095
rect -480 -2220 -280 -2135
rect -130 -2095 70 -2020
rect -130 -2135 -50 -2095
rect -10 -2135 70 -2095
rect -130 -2220 70 -2135
rect 220 -2095 420 -2020
rect 220 -2135 300 -2095
rect 340 -2135 420 -2095
rect 220 -2220 420 -2135
rect 570 -2095 770 -2020
rect 570 -2135 650 -2095
rect 690 -2135 770 -2095
rect 570 -2220 770 -2135
rect 920 -2095 1120 -2020
rect 920 -2135 1000 -2095
rect 1040 -2135 1120 -2095
rect 920 -2220 1120 -2135
rect 1270 -2095 1470 -2020
rect 1270 -2135 1350 -2095
rect 1390 -2135 1470 -2095
rect 1270 -2220 1470 -2135
rect 1620 -2095 1820 -2020
rect 1620 -2135 1700 -2095
rect 1740 -2135 1820 -2095
rect 1620 -2220 1820 -2135
rect 1970 -2095 2170 -2020
rect 1970 -2135 2050 -2095
rect 2090 -2135 2170 -2095
rect 1970 -2220 2170 -2135
rect 2320 -2095 2520 -2020
rect 2320 -2135 2400 -2095
rect 2440 -2135 2520 -2095
rect 2320 -2220 2520 -2135
rect 2670 -2095 2870 -2020
rect 2670 -2135 2750 -2095
rect 2790 -2135 2870 -2095
rect 2670 -2220 2870 -2135
rect 3020 -2095 3220 -2020
rect 3020 -2135 3100 -2095
rect 3140 -2135 3220 -2095
rect 3020 -2220 3220 -2135
rect 3370 -2095 3570 -2020
rect 3370 -2135 3450 -2095
rect 3490 -2135 3570 -2095
rect 3370 -2220 3570 -2135
rect 3720 -2095 3920 -2020
rect 3720 -2135 3800 -2095
rect 3840 -2135 3920 -2095
rect 3720 -2220 3920 -2135
rect 4070 -2095 4270 -2020
rect 4070 -2135 4150 -2095
rect 4190 -2135 4270 -2095
rect 4070 -2220 4270 -2135
rect 4420 -2095 4620 -2020
rect 4420 -2135 4500 -2095
rect 4540 -2135 4620 -2095
rect 4420 -2220 4620 -2135
rect 4770 -2095 4970 -2020
rect 4770 -2135 4850 -2095
rect 4890 -2135 4970 -2095
rect 4770 -2220 4970 -2135
<< mimcapcontact >>
rect -3200 3815 -3160 3855
rect -2850 3815 -2810 3855
rect -2500 3815 -2460 3855
rect -2150 3815 -2110 3855
rect -1800 3815 -1760 3855
rect -1450 3815 -1410 3855
rect -1100 3815 -1060 3855
rect -750 3815 -710 3855
rect -400 3815 -360 3855
rect -50 3815 -10 3855
rect 300 3815 340 3855
rect 650 3815 690 3855
rect 1000 3815 1040 3855
rect 1350 3815 1390 3855
rect 1700 3815 1740 3855
rect 2050 3815 2090 3855
rect 2400 3815 2440 3855
rect 2750 3815 2790 3855
rect 3100 3815 3140 3855
rect 3450 3815 3490 3855
rect 3800 3815 3840 3855
rect 4150 3815 4190 3855
rect 4500 3815 4540 3855
rect 4850 3815 4890 3855
rect -3200 3465 -3160 3505
rect -2850 3465 -2810 3505
rect -2500 3465 -2460 3505
rect -2150 3465 -2110 3505
rect -1800 3465 -1760 3505
rect -1450 3465 -1410 3505
rect -1100 3465 -1060 3505
rect -750 3465 -710 3505
rect -400 3465 -360 3505
rect -50 3465 -10 3505
rect 300 3465 340 3505
rect 650 3465 690 3505
rect 1000 3465 1040 3505
rect 1350 3465 1390 3505
rect 1700 3465 1740 3505
rect 2050 3465 2090 3505
rect 2400 3465 2440 3505
rect 2750 3465 2790 3505
rect 3100 3465 3140 3505
rect 3450 3465 3490 3505
rect 3800 3465 3840 3505
rect 4150 3465 4190 3505
rect 4500 3465 4540 3505
rect 4850 3465 4890 3505
rect -3200 3115 -3160 3155
rect -2850 3115 -2810 3155
rect -2500 3115 -2460 3155
rect -2150 3115 -2110 3155
rect -1800 3115 -1760 3155
rect -1450 3115 -1410 3155
rect -1100 3115 -1060 3155
rect -750 3115 -710 3155
rect -400 3115 -360 3155
rect -50 3105 -10 3145
rect 300 3105 340 3145
rect 650 3105 690 3145
rect 1000 3105 1040 3145
rect 1350 3105 1390 3145
rect 1700 3105 1740 3145
rect 2050 3115 2090 3155
rect 2400 3115 2440 3155
rect 2750 3115 2790 3155
rect 3100 3115 3140 3155
rect 3450 3115 3490 3155
rect 3800 3115 3840 3155
rect 4150 3115 4190 3155
rect 4500 3115 4540 3155
rect 4850 3115 4890 3155
rect -3200 2765 -3160 2805
rect -2850 2765 -2810 2805
rect -2500 2765 -2460 2805
rect -2150 2765 -2110 2805
rect -1800 2765 -1760 2805
rect -1450 2765 -1410 2805
rect -1100 2765 -1060 2805
rect -750 2765 -710 2805
rect 2400 2765 2440 2805
rect 2750 2765 2790 2805
rect 3100 2765 3140 2805
rect 3450 2765 3490 2805
rect 3800 2765 3840 2805
rect 4150 2765 4190 2805
rect 4500 2765 4540 2805
rect 4850 2765 4890 2805
rect -3200 2415 -3160 2455
rect -2850 2415 -2810 2455
rect -2500 2415 -2460 2455
rect -2150 2415 -2110 2455
rect -1800 2415 -1760 2455
rect -1450 2415 -1410 2455
rect -1100 2415 -1060 2455
rect -750 2415 -710 2455
rect 2400 2415 2440 2455
rect 2750 2415 2790 2455
rect 3100 2415 3140 2455
rect 3450 2415 3490 2455
rect 3800 2415 3840 2455
rect 4150 2415 4190 2455
rect 4500 2415 4540 2455
rect 4850 2415 4890 2455
rect -3200 2065 -3160 2105
rect -2850 2065 -2810 2105
rect -2500 2065 -2460 2105
rect -2150 2065 -2110 2105
rect -1800 2065 -1760 2105
rect 3450 2065 3490 2105
rect 3800 2065 3840 2105
rect 4150 2065 4190 2105
rect 4500 2065 4540 2105
rect 4850 2065 4890 2105
rect -3200 1715 -3160 1755
rect -2850 1715 -2810 1755
rect -2500 1715 -2460 1755
rect -2150 1715 -2110 1755
rect -1800 1715 -1760 1755
rect 3450 1715 3490 1755
rect 3800 1715 3840 1755
rect 4150 1715 4190 1755
rect 4500 1715 4540 1755
rect 4850 1715 4890 1755
rect -3200 1365 -3160 1405
rect -2850 1365 -2810 1405
rect -2500 1365 -2460 1405
rect -2150 1365 -2110 1405
rect -1800 1365 -1760 1405
rect 3450 1365 3490 1405
rect 3800 1365 3840 1405
rect 4150 1365 4190 1405
rect 4500 1365 4540 1405
rect 4850 1365 4890 1405
rect -3200 1015 -3160 1055
rect -2850 1015 -2810 1055
rect -2500 1015 -2460 1055
rect -2150 1015 -2110 1055
rect -1800 1015 -1760 1055
rect 3450 1015 3490 1055
rect 3800 1015 3840 1055
rect 4150 1015 4190 1055
rect 4500 1015 4540 1055
rect 4850 1015 4890 1055
rect -3200 665 -3160 705
rect -2850 665 -2810 705
rect -2500 665 -2460 705
rect -2150 665 -2110 705
rect -1800 665 -1760 705
rect 3450 665 3490 705
rect 3800 665 3840 705
rect 4150 665 4190 705
rect 4500 665 4540 705
rect 4850 665 4890 705
rect -3200 315 -3160 355
rect -2850 315 -2810 355
rect -2500 315 -2460 355
rect -2150 315 -2110 355
rect -1800 315 -1760 355
rect 3450 315 3490 355
rect 3800 315 3840 355
rect 4150 315 4190 355
rect 4500 315 4540 355
rect 4850 315 4890 355
rect -3200 -35 -3160 5
rect -2850 -35 -2810 5
rect -2500 -35 -2460 5
rect -2150 -35 -2110 5
rect -1800 -35 -1760 5
rect 3450 -35 3490 5
rect 3800 -35 3840 5
rect 4150 -35 4190 5
rect 4500 -35 4540 5
rect 4850 -35 4890 5
rect -3200 -385 -3160 -345
rect -2850 -385 -2810 -345
rect -2500 -385 -2460 -345
rect -2150 -385 -2110 -345
rect -1800 -385 -1760 -345
rect 3450 -385 3490 -345
rect 3800 -385 3840 -345
rect 4150 -385 4190 -345
rect 4500 -385 4540 -345
rect 4850 -385 4890 -345
rect -3200 -735 -3160 -695
rect -2850 -735 -2810 -695
rect -2500 -735 -2460 -695
rect -2150 -735 -2110 -695
rect -1800 -735 -1760 -695
rect 3450 -735 3490 -695
rect 3800 -735 3840 -695
rect 4150 -735 4190 -695
rect 4500 -735 4540 -695
rect 4850 -735 4890 -695
rect -3200 -1085 -3160 -1045
rect -2850 -1085 -2810 -1045
rect -2500 -1085 -2460 -1045
rect -2150 -1085 -2110 -1045
rect -1800 -1085 -1760 -1045
rect 3450 -1085 3490 -1045
rect 3800 -1085 3840 -1045
rect 4150 -1085 4190 -1045
rect 4500 -1085 4540 -1045
rect 4850 -1085 4890 -1045
rect -3200 -1435 -3160 -1395
rect -2850 -1435 -2810 -1395
rect -2500 -1435 -2460 -1395
rect -2150 -1435 -2110 -1395
rect -1800 -1435 -1760 -1395
rect -1450 -1435 -1410 -1395
rect -1100 -1435 -1060 -1395
rect -750 -1435 -710 -1395
rect -400 -1435 -360 -1395
rect -50 -1435 -10 -1395
rect 300 -1435 340 -1395
rect 650 -1435 690 -1395
rect 1000 -1435 1040 -1395
rect 1350 -1435 1390 -1395
rect 1700 -1435 1740 -1395
rect 2050 -1435 2090 -1395
rect 2400 -1435 2440 -1395
rect 2750 -1435 2790 -1395
rect 3100 -1435 3140 -1395
rect 3450 -1435 3490 -1395
rect 3800 -1435 3840 -1395
rect 4150 -1435 4190 -1395
rect 4500 -1435 4540 -1395
rect 4850 -1435 4890 -1395
rect -3200 -1785 -3160 -1745
rect -2850 -1785 -2810 -1745
rect -2500 -1785 -2460 -1745
rect -2150 -1785 -2110 -1745
rect -1800 -1785 -1760 -1745
rect -1450 -1785 -1410 -1745
rect -1100 -1785 -1060 -1745
rect -750 -1785 -710 -1745
rect -400 -1785 -360 -1745
rect -50 -1785 -10 -1745
rect 300 -1785 340 -1745
rect 650 -1785 690 -1745
rect 1000 -1785 1040 -1745
rect 1350 -1785 1390 -1745
rect 1700 -1785 1740 -1745
rect 2050 -1785 2090 -1745
rect 2400 -1785 2440 -1745
rect 2750 -1785 2790 -1745
rect 3100 -1785 3140 -1745
rect 3450 -1785 3490 -1745
rect 3800 -1785 3840 -1745
rect 4150 -1785 4190 -1745
rect 4500 -1785 4540 -1745
rect 4850 -1785 4890 -1745
rect -3200 -2135 -3160 -2095
rect -2850 -2135 -2810 -2095
rect -2500 -2135 -2460 -2095
rect -2150 -2135 -2110 -2095
rect -1800 -2135 -1760 -2095
rect -1450 -2135 -1410 -2095
rect -1100 -2135 -1060 -2095
rect -750 -2135 -710 -2095
rect -400 -2135 -360 -2095
rect -50 -2135 -10 -2095
rect 300 -2135 340 -2095
rect 650 -2135 690 -2095
rect 1000 -2135 1040 -2095
rect 1350 -2135 1390 -2095
rect 1700 -2135 1740 -2095
rect 2050 -2135 2090 -2095
rect 2400 -2135 2440 -2095
rect 2750 -2135 2790 -2095
rect 3100 -2135 3140 -2095
rect 3450 -2135 3490 -2095
rect 3800 -2135 3840 -2095
rect 4150 -2135 4190 -2095
rect 4500 -2135 4540 -2095
rect 4850 -2135 4890 -2095
<< metal4 >>
rect -3850 4280 5140 4285
rect -3850 4240 825 4280
rect 865 4240 5140 4280
rect -3850 4235 5140 4240
rect -3205 3855 -2455 3860
rect -3205 3815 -3200 3855
rect -3160 3815 -2850 3855
rect -2810 3815 -2500 3855
rect -2460 3815 -2455 3855
rect -3205 3810 -2455 3815
rect -2505 3510 -2455 3810
rect -2155 3855 -2105 3860
rect -2155 3815 -2150 3855
rect -2110 3815 -2105 3855
rect -2155 3510 -2105 3815
rect -1805 3855 -1755 3860
rect -1805 3815 -1800 3855
rect -1760 3815 -1755 3855
rect -1805 3510 -1755 3815
rect -1455 3855 -1405 3860
rect -1455 3815 -1450 3855
rect -1410 3815 -1405 3855
rect -1455 3510 -1405 3815
rect -1105 3855 -1055 3860
rect -1105 3815 -1100 3855
rect -1060 3815 -1055 3855
rect -1105 3510 -1055 3815
rect -755 3855 -705 3860
rect -755 3815 -750 3855
rect -710 3815 -705 3855
rect -755 3510 -705 3815
rect -405 3855 -355 3860
rect -405 3815 -400 3855
rect -360 3815 -355 3855
rect -405 3510 -355 3815
rect -55 3855 -5 3860
rect -55 3815 -50 3855
rect -10 3815 -5 3855
rect -55 3510 -5 3815
rect 295 3855 345 3860
rect 295 3815 300 3855
rect 340 3815 345 3855
rect 295 3510 345 3815
rect 645 3855 695 3860
rect 645 3815 650 3855
rect 690 3815 695 3855
rect 645 3510 695 3815
rect -3205 3505 695 3510
rect -3205 3465 -3200 3505
rect -3160 3465 -2850 3505
rect -2810 3465 -2500 3505
rect -2460 3465 -2150 3505
rect -2110 3465 -1800 3505
rect -1760 3465 -1450 3505
rect -1410 3465 -1100 3505
rect -1060 3465 -750 3505
rect -710 3465 -400 3505
rect -360 3465 -50 3505
rect -10 3465 300 3505
rect 340 3465 650 3505
rect 690 3465 695 3505
rect -3205 3460 695 3465
rect -2505 3160 -2455 3460
rect -3205 3155 -2105 3160
rect -3205 3115 -3200 3155
rect -3160 3115 -2850 3155
rect -2810 3115 -2500 3155
rect -2460 3115 -2150 3155
rect -2110 3115 -2105 3155
rect -3205 3110 -2105 3115
rect -1805 3155 -1755 3460
rect -1805 3115 -1800 3155
rect -1760 3115 -1755 3155
rect -2505 2810 -2455 3110
rect -3205 2805 -2105 2810
rect -3205 2765 -3200 2805
rect -3160 2765 -2850 2805
rect -2810 2765 -2500 2805
rect -2460 2765 -2150 2805
rect -2110 2765 -2105 2805
rect -3205 2760 -2105 2765
rect -1805 2805 -1755 3115
rect -1805 2765 -1800 2805
rect -1760 2765 -1755 2805
rect -1805 2760 -1755 2765
rect -1455 3155 -1405 3460
rect -1455 3115 -1450 3155
rect -1410 3115 -1405 3155
rect -1455 2805 -1405 3115
rect -1455 2765 -1450 2805
rect -1410 2765 -1405 2805
rect -2505 2460 -2455 2760
rect -3205 2455 -1755 2460
rect -3205 2415 -3200 2455
rect -3160 2415 -2850 2455
rect -2810 2415 -2500 2455
rect -2460 2415 -2150 2455
rect -2110 2415 -1800 2455
rect -1760 2415 -1755 2455
rect -3205 2410 -1755 2415
rect -1455 2455 -1405 2765
rect -1455 2415 -1450 2455
rect -1410 2415 -1405 2455
rect -1455 2410 -1405 2415
rect -1105 3155 -1055 3460
rect -1105 3115 -1100 3155
rect -1060 3115 -1055 3155
rect -1105 2805 -1055 3115
rect -1105 2765 -1100 2805
rect -1060 2765 -1055 2805
rect -1105 2455 -1055 2765
rect -1105 2415 -1100 2455
rect -1060 2415 -1055 2455
rect -1105 2410 -1055 2415
rect -755 3155 -705 3460
rect -755 3115 -750 3155
rect -710 3115 -705 3155
rect -755 2805 -705 3115
rect -405 3155 -355 3460
rect -405 3115 -400 3155
rect -360 3115 -355 3155
rect -405 3110 -355 3115
rect -55 3145 -5 3460
rect -55 3105 -50 3145
rect -10 3105 -5 3145
rect -55 3100 -5 3105
rect 295 3145 345 3460
rect 295 3105 300 3145
rect 340 3105 345 3145
rect 295 3100 345 3105
rect 645 3145 695 3460
rect 645 3105 650 3145
rect 690 3105 695 3145
rect 645 3100 695 3105
rect 995 3855 1045 3860
rect 995 3815 1000 3855
rect 1040 3815 1045 3855
rect 995 3510 1045 3815
rect 1345 3855 1395 3860
rect 1345 3815 1350 3855
rect 1390 3815 1395 3855
rect 1345 3510 1395 3815
rect 1695 3855 1745 3860
rect 1695 3815 1700 3855
rect 1740 3815 1745 3855
rect 1695 3510 1745 3815
rect 2045 3855 2095 3860
rect 2045 3815 2050 3855
rect 2090 3815 2095 3855
rect 2045 3510 2095 3815
rect 2395 3855 2445 3860
rect 2395 3815 2400 3855
rect 2440 3815 2445 3855
rect 2395 3510 2445 3815
rect 2745 3855 2795 3860
rect 2745 3815 2750 3855
rect 2790 3815 2795 3855
rect 2745 3510 2795 3815
rect 3095 3855 3145 3860
rect 3095 3815 3100 3855
rect 3140 3815 3145 3855
rect 3095 3510 3145 3815
rect 3445 3855 3495 3860
rect 3445 3815 3450 3855
rect 3490 3815 3495 3855
rect 3445 3510 3495 3815
rect 3795 3855 3845 3860
rect 3795 3815 3800 3855
rect 3840 3815 3845 3855
rect 3795 3510 3845 3815
rect 4145 3855 4895 3860
rect 4145 3815 4150 3855
rect 4190 3815 4500 3855
rect 4540 3815 4850 3855
rect 4890 3815 4895 3855
rect 4145 3810 4895 3815
rect 4145 3510 4195 3810
rect 995 3505 4895 3510
rect 995 3465 1000 3505
rect 1040 3465 1350 3505
rect 1390 3465 1700 3505
rect 1740 3465 2050 3505
rect 2090 3465 2400 3505
rect 2440 3465 2750 3505
rect 2790 3465 3100 3505
rect 3140 3465 3450 3505
rect 3490 3465 3800 3505
rect 3840 3465 4150 3505
rect 4190 3465 4500 3505
rect 4540 3465 4850 3505
rect 4890 3465 4895 3505
rect 995 3460 4895 3465
rect 995 3145 1045 3460
rect 995 3105 1000 3145
rect 1040 3105 1045 3145
rect 995 3100 1045 3105
rect 1345 3145 1395 3460
rect 1345 3105 1350 3145
rect 1390 3105 1395 3145
rect 1345 3100 1395 3105
rect 1695 3145 1745 3460
rect 1695 3105 1700 3145
rect 1740 3105 1745 3145
rect 2045 3155 2095 3460
rect 2045 3115 2050 3155
rect 2090 3115 2095 3155
rect 2045 3110 2095 3115
rect 2395 3155 2445 3460
rect 2395 3115 2400 3155
rect 2440 3115 2445 3155
rect 1695 3100 1745 3105
rect -755 2765 -750 2805
rect -710 2765 -705 2805
rect -755 2455 -705 2765
rect -755 2415 -750 2455
rect -710 2415 -705 2455
rect -755 2410 -705 2415
rect 2395 2805 2445 3115
rect 2395 2765 2400 2805
rect 2440 2765 2445 2805
rect 2395 2455 2445 2765
rect 2395 2415 2400 2455
rect 2440 2415 2445 2455
rect 2395 2410 2445 2415
rect 2745 3155 2795 3460
rect 2745 3115 2750 3155
rect 2790 3115 2795 3155
rect 2745 2805 2795 3115
rect 2745 2765 2750 2805
rect 2790 2765 2795 2805
rect 2745 2455 2795 2765
rect 2745 2415 2750 2455
rect 2790 2415 2795 2455
rect 2745 2410 2795 2415
rect 3095 3155 3145 3460
rect 3095 3115 3100 3155
rect 3140 3115 3145 3155
rect 3095 2805 3145 3115
rect 3095 2765 3100 2805
rect 3140 2765 3145 2805
rect 3095 2455 3145 2765
rect 3445 3155 3495 3460
rect 4145 3160 4195 3460
rect 3445 3115 3450 3155
rect 3490 3115 3495 3155
rect 3445 2805 3495 3115
rect 3795 3155 4895 3160
rect 3795 3115 3800 3155
rect 3840 3115 4150 3155
rect 4190 3115 4500 3155
rect 4540 3115 4850 3155
rect 4890 3115 4895 3155
rect 3795 3110 4895 3115
rect 4145 2810 4195 3110
rect 3445 2765 3450 2805
rect 3490 2765 3495 2805
rect 3445 2760 3495 2765
rect 3795 2805 4895 2810
rect 3795 2765 3800 2805
rect 3840 2765 4150 2805
rect 4190 2765 4500 2805
rect 4540 2765 4850 2805
rect 4890 2765 4895 2805
rect 3795 2760 4895 2765
rect 4145 2460 4195 2760
rect 3095 2415 3100 2455
rect 3140 2415 3145 2455
rect 3095 2410 3145 2415
rect 3445 2455 4895 2460
rect 3445 2415 3450 2455
rect 3490 2415 3800 2455
rect 3840 2415 4150 2455
rect 4190 2415 4500 2455
rect 4540 2415 4850 2455
rect 4890 2415 4895 2455
rect 3445 2410 4895 2415
rect -2505 2110 -2455 2410
rect 4145 2110 4195 2410
rect -3205 2105 -1755 2110
rect -3205 2065 -3200 2105
rect -3160 2065 -2850 2105
rect -2810 2065 -2500 2105
rect -2460 2065 -2150 2105
rect -2110 2065 -1800 2105
rect -1760 2065 -1755 2105
rect -3205 2060 -1755 2065
rect 3445 2105 4895 2110
rect 3445 2065 3450 2105
rect 3490 2065 3800 2105
rect 3840 2065 4150 2105
rect 4190 2065 4500 2105
rect 4540 2065 4850 2105
rect 4890 2065 4895 2105
rect 3445 2060 4895 2065
rect -2505 1760 -2455 2060
rect 4145 1760 4195 2060
rect -3205 1755 -1755 1760
rect -3205 1715 -3200 1755
rect -3160 1715 -2850 1755
rect -2810 1715 -2500 1755
rect -2460 1715 -2150 1755
rect -2110 1715 -1800 1755
rect -1760 1715 -1755 1755
rect -3205 1710 -1755 1715
rect 3445 1755 4895 1760
rect 3445 1715 3450 1755
rect 3490 1715 3800 1755
rect 3840 1715 4150 1755
rect 4190 1715 4500 1755
rect 4540 1715 4850 1755
rect 4890 1715 4895 1755
rect 3445 1710 4895 1715
rect -2505 1410 -2455 1710
rect 4145 1410 4195 1710
rect -3205 1405 -1755 1410
rect -3205 1365 -3200 1405
rect -3160 1365 -2850 1405
rect -2810 1365 -2500 1405
rect -2460 1365 -2150 1405
rect -2110 1365 -1800 1405
rect -1760 1365 -1755 1405
rect -3205 1360 -1755 1365
rect 3445 1405 4895 1410
rect 3445 1365 3450 1405
rect 3490 1365 3800 1405
rect 3840 1365 4150 1405
rect 4190 1365 4500 1405
rect 4540 1365 4850 1405
rect 4890 1365 4895 1405
rect 3445 1360 4895 1365
rect -2505 1060 -2455 1360
rect 4145 1060 4195 1360
rect -3205 1055 -1755 1060
rect -3205 1015 -3200 1055
rect -3160 1015 -2850 1055
rect -2810 1015 -2500 1055
rect -2460 1015 -2150 1055
rect -2110 1015 -1800 1055
rect -1760 1015 -1755 1055
rect -3205 1010 -1755 1015
rect 3445 1055 4895 1060
rect 3445 1015 3450 1055
rect 3490 1015 3800 1055
rect 3840 1015 4150 1055
rect 4190 1015 4500 1055
rect 4540 1015 4850 1055
rect 4890 1015 4895 1055
rect 3445 1010 4895 1015
rect -2505 710 -2455 1010
rect 4145 710 4195 1010
rect -3205 705 -1755 710
rect -3205 665 -3200 705
rect -3160 665 -2850 705
rect -2810 665 -2500 705
rect -2460 665 -2150 705
rect -2110 665 -1800 705
rect -1760 665 -1755 705
rect -3205 660 -1755 665
rect 3445 705 4895 710
rect 3445 665 3450 705
rect 3490 665 3800 705
rect 3840 665 4150 705
rect 4190 665 4500 705
rect 4540 665 4850 705
rect 4890 665 4895 705
rect 3445 660 4895 665
rect -2505 360 -2455 660
rect 4145 360 4195 660
rect -3205 355 -1495 360
rect -3205 315 -3200 355
rect -3160 315 -2850 355
rect -2810 315 -2500 355
rect -2460 315 -2150 355
rect -2110 315 -1800 355
rect -1760 315 -1540 355
rect -1500 315 -1495 355
rect -3205 310 -1495 315
rect 3185 355 4895 360
rect 3185 315 3190 355
rect 3230 315 3450 355
rect 3490 315 3800 355
rect 3840 315 4150 355
rect 4190 315 4500 355
rect 4540 315 4850 355
rect 4890 315 4895 355
rect 3185 310 4895 315
rect -2505 10 -2455 310
rect 4145 10 4195 310
rect -3205 5 -1755 10
rect -3205 -35 -3200 5
rect -3160 -35 -2850 5
rect -2810 -35 -2500 5
rect -2460 -35 -2150 5
rect -2110 -35 -1800 5
rect -1760 -35 -1755 5
rect -3205 -40 -1755 -35
rect 3445 5 4895 10
rect 3445 -35 3450 5
rect 3490 -35 3800 5
rect 3840 -35 4150 5
rect 4190 -35 4500 5
rect 4540 -35 4850 5
rect 4890 -35 4895 5
rect 3445 -40 4895 -35
rect -2505 -340 -2455 -40
rect 4145 -340 4195 -40
rect -3205 -345 -1755 -340
rect -3205 -385 -3200 -345
rect -3160 -385 -2850 -345
rect -2810 -385 -2500 -345
rect -2460 -385 -2150 -345
rect -2110 -385 -1800 -345
rect -1760 -385 -1755 -345
rect -3205 -390 -1755 -385
rect 3445 -345 4895 -340
rect 3445 -385 3450 -345
rect 3490 -385 3800 -345
rect 3840 -385 4150 -345
rect 4190 -385 4500 -345
rect 4540 -385 4850 -345
rect 4890 -385 4895 -345
rect 3445 -390 4895 -385
rect -2505 -690 -2455 -390
rect 4145 -690 4195 -390
rect -3205 -695 -1755 -690
rect -3205 -735 -3200 -695
rect -3160 -735 -2850 -695
rect -2810 -735 -2500 -695
rect -2460 -735 -2150 -695
rect -2110 -735 -1800 -695
rect -1760 -735 -1755 -695
rect -3205 -740 -1755 -735
rect 3445 -695 4895 -690
rect 3445 -735 3450 -695
rect 3490 -735 3800 -695
rect 3840 -735 4150 -695
rect 4190 -735 4500 -695
rect 4540 -735 4850 -695
rect 4890 -735 4895 -695
rect 3445 -740 4895 -735
rect -2505 -1040 -2455 -740
rect 4145 -1040 4195 -740
rect -3205 -1045 -1755 -1040
rect -3205 -1085 -3200 -1045
rect -3160 -1085 -2850 -1045
rect -2810 -1085 -2500 -1045
rect -2460 -1085 -2150 -1045
rect -2110 -1085 -1800 -1045
rect -1760 -1085 -1755 -1045
rect -3205 -1090 -1755 -1085
rect 3445 -1045 4895 -1040
rect 3445 -1085 3450 -1045
rect 3490 -1085 3800 -1045
rect 3840 -1085 4150 -1045
rect 4190 -1085 4500 -1045
rect 4540 -1085 4850 -1045
rect 4890 -1085 4895 -1045
rect 3445 -1090 4895 -1085
rect -2505 -1390 -2455 -1090
rect 4145 -1390 4195 -1090
rect -3205 -1395 -1755 -1390
rect -3205 -1435 -3200 -1395
rect -3160 -1435 -2850 -1395
rect -2810 -1435 -2500 -1395
rect -2460 -1435 -2150 -1395
rect -2110 -1435 -1800 -1395
rect -1760 -1435 -1755 -1395
rect -3205 -1440 -1755 -1435
rect -1455 -1395 -1405 -1390
rect -1455 -1435 -1450 -1395
rect -1410 -1435 -1405 -1395
rect -2505 -1740 -2455 -1440
rect -1455 -1740 -1405 -1435
rect -1105 -1395 -1055 -1390
rect -1105 -1435 -1100 -1395
rect -1060 -1435 -1055 -1395
rect -1105 -1740 -1055 -1435
rect -755 -1395 -705 -1390
rect -755 -1435 -750 -1395
rect -710 -1435 -705 -1395
rect -755 -1740 -705 -1435
rect -405 -1395 -355 -1390
rect -405 -1435 -400 -1395
rect -360 -1435 -355 -1395
rect -405 -1740 -355 -1435
rect -55 -1395 -5 -1390
rect -55 -1435 -50 -1395
rect -10 -1435 -5 -1395
rect -55 -1740 -5 -1435
rect 295 -1395 345 -1390
rect 295 -1435 300 -1395
rect 340 -1435 345 -1395
rect 295 -1740 345 -1435
rect 645 -1395 695 -1390
rect 645 -1435 650 -1395
rect 690 -1435 695 -1395
rect 645 -1740 695 -1435
rect -3205 -1745 695 -1740
rect -3205 -1785 -3200 -1745
rect -3160 -1785 -2850 -1745
rect -2810 -1785 -2500 -1745
rect -2460 -1785 -2150 -1745
rect -2110 -1785 -1800 -1745
rect -1760 -1785 -1450 -1745
rect -1410 -1785 -1100 -1745
rect -1060 -1785 -750 -1745
rect -710 -1785 -400 -1745
rect -360 -1785 -50 -1745
rect -10 -1785 300 -1745
rect 340 -1785 650 -1745
rect 690 -1785 695 -1745
rect -3205 -1790 695 -1785
rect -2505 -2090 -2455 -1790
rect -3205 -2095 -2455 -2090
rect -3205 -2135 -3200 -2095
rect -3160 -2135 -2850 -2095
rect -2810 -2135 -2500 -2095
rect -2460 -2135 -2455 -2095
rect -3205 -2140 -2455 -2135
rect -2155 -2095 -2105 -1790
rect -2155 -2135 -2150 -2095
rect -2110 -2135 -2105 -2095
rect -2155 -2140 -2105 -2135
rect -1805 -2095 -1755 -1790
rect -1805 -2135 -1800 -2095
rect -1760 -2135 -1755 -2095
rect -1805 -2140 -1755 -2135
rect -1455 -2095 -1405 -1790
rect -1455 -2135 -1450 -2095
rect -1410 -2135 -1405 -2095
rect -1455 -2140 -1405 -2135
rect -1105 -2095 -1055 -1790
rect -1105 -2135 -1100 -2095
rect -1060 -2135 -1055 -2095
rect -1105 -2140 -1055 -2135
rect -755 -2095 -705 -1790
rect -755 -2135 -750 -2095
rect -710 -2135 -705 -2095
rect -755 -2140 -705 -2135
rect -405 -2095 -355 -1790
rect -405 -2135 -400 -2095
rect -360 -2135 -355 -2095
rect -405 -2140 -355 -2135
rect -55 -2095 -5 -1790
rect -55 -2135 -50 -2095
rect -10 -2135 -5 -2095
rect -55 -2140 -5 -2135
rect 295 -2095 345 -1790
rect 295 -2135 300 -2095
rect 340 -2135 345 -2095
rect 295 -2140 345 -2135
rect 645 -2095 695 -1790
rect 645 -2135 650 -2095
rect 690 -2135 695 -2095
rect 645 -2140 695 -2135
rect 995 -1395 1045 -1390
rect 995 -1435 1000 -1395
rect 1040 -1435 1045 -1395
rect 995 -1740 1045 -1435
rect 1345 -1395 1395 -1390
rect 1345 -1435 1350 -1395
rect 1390 -1435 1395 -1395
rect 1345 -1740 1395 -1435
rect 1695 -1395 1745 -1390
rect 1695 -1435 1700 -1395
rect 1740 -1435 1745 -1395
rect 1695 -1740 1745 -1435
rect 2045 -1395 2095 -1390
rect 2045 -1435 2050 -1395
rect 2090 -1435 2095 -1395
rect 2045 -1740 2095 -1435
rect 2395 -1395 2445 -1390
rect 2395 -1435 2400 -1395
rect 2440 -1435 2445 -1395
rect 2395 -1740 2445 -1435
rect 2745 -1395 2795 -1390
rect 2745 -1435 2750 -1395
rect 2790 -1435 2795 -1395
rect 2745 -1740 2795 -1435
rect 3095 -1395 3145 -1390
rect 3095 -1435 3100 -1395
rect 3140 -1435 3145 -1395
rect 3095 -1740 3145 -1435
rect 3445 -1395 4895 -1390
rect 3445 -1435 3450 -1395
rect 3490 -1435 3800 -1395
rect 3840 -1435 4150 -1395
rect 4190 -1435 4500 -1395
rect 4540 -1435 4850 -1395
rect 4890 -1435 4895 -1395
rect 3445 -1440 4895 -1435
rect 4145 -1740 4195 -1440
rect 995 -1745 4895 -1740
rect 995 -1785 1000 -1745
rect 1040 -1785 1350 -1745
rect 1390 -1785 1700 -1745
rect 1740 -1785 2050 -1745
rect 2090 -1785 2400 -1745
rect 2440 -1785 2750 -1745
rect 2790 -1785 3100 -1745
rect 3140 -1785 3450 -1745
rect 3490 -1785 3800 -1745
rect 3840 -1785 4150 -1745
rect 4190 -1785 4500 -1745
rect 4540 -1785 4850 -1745
rect 4890 -1785 4895 -1745
rect 995 -1790 4895 -1785
rect 995 -2095 1045 -1790
rect 995 -2135 1000 -2095
rect 1040 -2135 1045 -2095
rect 995 -2140 1045 -2135
rect 1345 -2095 1395 -1790
rect 1345 -2135 1350 -2095
rect 1390 -2135 1395 -2095
rect 1345 -2140 1395 -2135
rect 1695 -2095 1745 -1790
rect 1695 -2135 1700 -2095
rect 1740 -2135 1745 -2095
rect 1695 -2140 1745 -2135
rect 2045 -2095 2095 -1790
rect 2045 -2135 2050 -2095
rect 2090 -2135 2095 -2095
rect 2045 -2140 2095 -2135
rect 2395 -2095 2445 -1790
rect 2395 -2135 2400 -2095
rect 2440 -2135 2445 -2095
rect 2395 -2140 2445 -2135
rect 2745 -2095 2795 -1790
rect 2745 -2135 2750 -2095
rect 2790 -2135 2795 -2095
rect 2745 -2140 2795 -2135
rect 3095 -2095 3145 -1790
rect 3095 -2135 3100 -2095
rect 3140 -2135 3145 -2095
rect 3095 -2140 3145 -2135
rect 3445 -2095 3495 -1790
rect 3445 -2135 3450 -2095
rect 3490 -2135 3495 -2095
rect 3445 -2140 3495 -2135
rect 3795 -2095 3845 -1790
rect 3795 -2135 3800 -2095
rect 3840 -2135 3845 -2095
rect 3795 -2140 3845 -2135
rect 4145 -2090 4195 -1790
rect 4145 -2095 4895 -2090
rect 4145 -2135 4150 -2095
rect 4190 -2135 4500 -2095
rect 4540 -2135 4850 -2095
rect 4890 -2135 4895 -2095
rect 4145 -2140 4895 -2135
rect -3850 -2420 5140 -2415
rect -3850 -2460 825 -2420
rect 865 -2460 5140 -2420
rect -3850 -2465 5140 -2460
<< labels >>
flabel metal3 3100 1595 3100 1595 7 FreeSans 240 0 -80 0 cap_res_X
flabel metal3 -1410 1610 -1410 1610 3 FreeSans 240 0 80 0 cap_res_Y
flabel metal4 -3850 -2440 -3850 -2440 7 FreeSans 240 0 -80 0 GNDA
port 16 w
flabel metal2 1310 2775 1310 2775 1 FreeSans 240 0 0 80 Vb2_Vb3
flabel metal2 400 2775 400 2775 1 FreeSans 240 0 0 80 Vb2_2
flabel metal2 310 1140 310 1140 7 FreeSans 240 0 -80 0 V_err_amp_ref
port 12 w
flabel metal2 1525 1100 1525 1100 1 FreeSans 240 0 0 160 V_tot
flabel metal2 1070 1200 1070 1200 3 FreeSans 240 0 80 0 V_err_gate
port 13 e
flabel metal2 945 1045 945 1045 3 FreeSans 240 0 80 0 err_amp_mir
flabel metal1 -350 305 -350 305 5 FreeSans 240 0 0 -80 Y
flabel metal1 1970 2135 1970 2135 3 FreeSans 240 0 80 0 VD3
flabel metal2 1470 1005 1470 1005 1 FreeSans 240 0 0 80 err_amp_out
flabel metal2 -105 535 -105 535 7 FreeSans 240 0 -80 0 VIN+
port 14 w
flabel metal2 1795 535 1795 535 3 FreeSans 240 0 80 0 VIN-
port 15 e
flabel metal1 2040 305 2040 305 5 FreeSans 240 0 0 -80 X
flabel metal1 3210 -340 3210 -340 5 FreeSans 240 0 0 -80 VOUT-
port 9 s
flabel metal1 -1520 -340 -1520 -340 5 FreeSans 240 0 0 -80 VOUT+
port 10 s
flabel metal2 845 945 845 945 1 FreeSans 240 0 0 80 Vb1
port 6 n
flabel metal4 -3850 4260 -3850 4260 7 FreeSans 240 0 -80 0 VDDA
port 1 w
flabel metal2 2260 1600 2260 1600 5 FreeSans 240 0 0 -80 Vb3
port 4 s
flabel metal2 1070 1665 1070 1665 1 FreeSans 240 0 0 80 Vb2
port 5 n
flabel metal1 2895 270 2895 270 1 FreeSans 240 0 0 80 V_CMFB_S2
port 7 n
flabel metal1 2940 420 2940 420 1 FreeSans 240 0 0 80 V_CMFB_S1
port 2 n
flabel metal2 1125 1505 1125 1505 3 FreeSans 240 0 80 0 V_err_p
flabel metal1 565 1505 565 1505 7 FreeSans 240 0 -80 0 V_err_mir_p
flabel metal1 -280 2135 -280 2135 7 FreeSans 240 0 -80 0 VD4
flabel metal1 -1250 420 -1250 420 1 FreeSans 240 0 0 80 V_CMFB_S3
port 3 n
flabel metal1 -1205 270 -1205 270 1 FreeSans 240 0 0 80 V_CMFB_S4
port 8 n
flabel metal1 235 560 235 560 7 FreeSans 240 0 -80 0 VD2
flabel metal1 1455 560 1455 560 3 FreeSans 240 0 80 0 VD1
flabel metal2 965 -1180 965 -1180 3 FreeSans 240 0 80 0 Vb1_2
flabel metal2 1570 -405 1570 -405 5 FreeSans 240 0 0 -80 V_b_2nd_stage
flabel metal2 460 -5 460 -5 1 FreeSans 240 0 0 80 V_tail_gate
port 11 n
flabel metal1 920 25 920 25 3 FreeSans 240 0 80 0 V_p_mir
flabel metal1 1265 -165 1265 -165 3 FreeSans 240 0 80 0 V_source
<< end >>
