* PEX produced on Sun Jul 13 02:46:43 PM CEST 2025 using /foss/tools/osic-multitool/iic-pex.sh with m=3 and s=1
* NGSPICE file created from bgr_opamp_dummy_magic_10.ext - technology: sky130A

.subckt bgr_opamp_dummy_magic_10 VDDA GNDA VOUT+ VOUT- VIN+ VIN-
X0 GNDA.t201 bgr_0.NFET_GATE_10uA.t5 two_stage_opamp_dummy_magic_14_0.Vb3.t2 GNDA.t200 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X1 bgr_0.V_TOP.t9 VDDA.t372 VDDA.t374 VDDA.t373 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.45 ps=2.9 w=1 l=0.15
X2 VOUT-.t19 two_stage_opamp_dummy_magic_14_0.cap_res_X.t138 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3 VOUT+.t19 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t138 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.t9 two_stage_opamp_dummy_magic_14_0.X.t25 VDDA.t75 GNDA.t60 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X5 VOUT+.t20 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t137 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6 GNDA.t312 two_stage_opamp_dummy_magic_14_0.V_b_2nd_stage.t2 VOUT-.t18 GNDA.t311 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X7 VDDA.t29 bgr_0.V_TOP.t14 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.t3 VDDA.t28 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X8 VDDA.t371 VDDA.t369 two_stage_opamp_dummy_magic_14_0.err_amp_out.t3 VDDA.t370 sky130_fd_pr__pfet_01v8 ad=1 pd=5.8 as=0.5 ps=2.9 w=2.5 l=0.15
X9 VOUT+.t21 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t136 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X10 two_stage_opamp_dummy_magic_14_0.V_source.t29 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t12 GNDA.t305 GNDA.t304 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X11 bgr_0.Vin+.t3 bgr_0.V_TOP.t15 VDDA.t97 VDDA.t96 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X12 VDDA.t261 two_stage_opamp_dummy_magic_14_0.Vb3.t8 two_stage_opamp_dummy_magic_14_0.VD3.t29 VDDA.t260 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X13 GNDA.t21 VDDA.t366 VDDA.t368 VDDA.t367 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X14 VDDA.t18 bgr_0.V_mir1.t17 bgr_0.1st_Vout_1.t5 VDDA.t17 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X15 VOUT+.t22 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t135 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X16 bgr_0.1st_Vout_2.t11 bgr_0.cap_res2.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X17 two_stage_opamp_dummy_magic_14_0.X.t23 two_stage_opamp_dummy_magic_14_0.Vb2.t11 two_stage_opamp_dummy_magic_14_0.VD3.t35 two_stage_opamp_dummy_magic_14_0.VD3.t34 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X18 VOUT+.t23 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t134 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X19 bgr_0.1st_Vout_2.t3 bgr_0.V_CUR_REF_REG.t3 bgr_0.V_p_2.t9 GNDA.t96 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X20 VOUT+.t24 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t133 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X21 VOUT+.t25 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t132 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X22 a_7460_23988.t1 bgr_0.Vin+.t4 GNDA.t2 sky130_fd_pr__res_xhigh_po_0p35 l=6
X23 VDDA.t163 two_stage_opamp_dummy_magic_14_0.V_err_gate.t6 two_stage_opamp_dummy_magic_14_0.V_err_mir_p.t1 VDDA.t162 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X24 two_stage_opamp_dummy_magic_14_0.VD2.t12 two_stage_opamp_dummy_magic_14_0.Vb1.t6 two_stage_opamp_dummy_magic_14_0.Y.t16 GNDA.t160 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X25 VOUT+.t26 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t131 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X26 two_stage_opamp_dummy_magic_14_0.VD2.t11 two_stage_opamp_dummy_magic_14_0.Vb1.t7 two_stage_opamp_dummy_magic_14_0.Y.t15 GNDA.t131 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X27 bgr_0.1st_Vout_2.t12 bgr_0.cap_res2.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X28 VDDA.t365 VDDA.t363 bgr_0.NFET_GATE_10uA.t0 VDDA.t364 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X29 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t7 bgr_0.PFET_GATE_10uA.t10 VDDA.t200 VDDA.t199 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X30 VDDA.t47 bgr_0.PFET_GATE_10uA.t11 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t2 VDDA.t46 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X31 VOUT-.t20 two_stage_opamp_dummy_magic_14_0.cap_res_X.t137 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X32 VOUT-.t21 two_stage_opamp_dummy_magic_14_0.cap_res_X.t136 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X33 VOUT-.t22 two_stage_opamp_dummy_magic_14_0.cap_res_X.t135 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X34 two_stage_opamp_dummy_magic_14_0.V_source.t2 VIN-.t0 two_stage_opamp_dummy_magic_14_0.VD1.t9 GNDA.t3 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X35 VOUT+.t27 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t130 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X36 bgr_0.1st_Vout_1.t11 bgr_0.cap_res1.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X37 bgr_0.1st_Vout_2.t9 bgr_0.V_mir2.t17 VDDA.t395 VDDA.t394 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X38 VDDA.t99 bgr_0.V_TOP.t16 bgr_0.Vin-.t3 VDDA.t98 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X39 bgr_0.1st_Vout_1.t7 bgr_0.Vin+.t6 bgr_0.V_p_1.t9 GNDA.t123 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X40 GNDA.t86 VDDA.t415 bgr_0.V_p_2.t10 GNDA.t85 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=1 ps=5.8 w=2.5 l=5
X41 VDDA.t259 two_stage_opamp_dummy_magic_14_0.Vb3.t9 two_stage_opamp_dummy_magic_14_0.VD3.t28 VDDA.t258 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X42 VOUT+.t28 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t129 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X43 bgr_0.cap_res2.t20 bgr_0.PFET_GATE_10uA.t6 GNDA.t10 sky130_fd_pr__res_high_po_0p35 l=2.05
X44 bgr_0.1st_Vout_1.t12 bgr_0.cap_res1.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X45 GNDA.t293 GNDA.t291 two_stage_opamp_dummy_magic_14_0.err_amp_out.t2 GNDA.t292 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=0.5 ps=2.9 w=2.5 l=0.15
X46 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.t9 two_stage_opamp_dummy_magic_14_0.Y.t25 VDDA.t198 GNDA.t136 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X47 two_stage_opamp_dummy_magic_14_0.V_source.t36 VIN+.t0 two_stage_opamp_dummy_magic_14_0.VD2.t20 GNDA.t93 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X48 VOUT+.t29 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t128 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X49 VOUT-.t23 two_stage_opamp_dummy_magic_14_0.cap_res_X.t134 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X50 VOUT-.t24 two_stage_opamp_dummy_magic_14_0.cap_res_X.t133 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X51 VOUT-.t25 two_stage_opamp_dummy_magic_14_0.cap_res_X.t132 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X52 VDDA.t399 bgr_0.1st_Vout_1.t13 bgr_0.V_TOP.t11 VDDA.t398 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X53 GNDA.t135 two_stage_opamp_dummy_magic_14_0.Y.t26 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.t9 VDDA.t197 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X54 bgr_0.V_TOP.t17 VDDA.t100 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X55 VOUT-.t26 two_stage_opamp_dummy_magic_14_0.cap_res_X.t131 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X56 two_stage_opamp_dummy_magic_14_0.VD4.t37 VDDA.t360 VDDA.t362 VDDA.t361 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X57 GNDA.t290 GNDA.t288 bgr_0.NFET_GATE_10uA.t1 GNDA.t289 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X58 bgr_0.START_UP.t3 bgr_0.V_TOP.t18 VDDA.t102 VDDA.t101 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X59 VOUT-.t27 two_stage_opamp_dummy_magic_14_0.cap_res_X.t130 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X60 two_stage_opamp_dummy_magic_14_0.V_err_gate.t2 bgr_0.NFET_GATE_10uA.t6 GNDA.t199 GNDA.t198 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X61 bgr_0.1st_Vout_1.t9 bgr_0.Vin+.t7 bgr_0.V_p_1.t8 GNDA.t124 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.2
X62 VOUT-.t28 two_stage_opamp_dummy_magic_14_0.cap_res_X.t129 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X63 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.t8 two_stage_opamp_dummy_magic_14_0.X.t26 VDDA.t39 GNDA.t30 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X64 VOUT+.t30 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t127 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X65 bgr_0.1st_Vout_1.t14 bgr_0.cap_res1.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X66 two_stage_opamp_dummy_magic_14_0.V_err_p.t1 two_stage_opamp_dummy_magic_14_0.V_err_gate.t7 VDDA.t191 VDDA.t190 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X67 bgr_0.V_TOP.t19 VDDA.t103 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X68 bgr_0.V_mir2.t11 bgr_0.V_mir2.t10 VDDA.t87 VDDA.t86 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X69 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.t16 VDDA.t357 VDDA.t359 VDDA.t358 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X70 VOUT-.t29 two_stage_opamp_dummy_magic_14_0.cap_res_X.t128 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X71 VOUT-.t2 two_stage_opamp_dummy_magic_14_0.X.t27 VDDA.t41 VDDA.t40 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X72 two_stage_opamp_dummy_magic_14_0.VD1.t19 two_stage_opamp_dummy_magic_14_0.Vb1.t8 two_stage_opamp_dummy_magic_14_0.X.t6 GNDA.t17 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X73 VOUT+.t0 a_5980_2720.t0 GNDA.t16 sky130_fd_pr__res_xhigh_po_0p35 l=2.63
X74 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.t14 bgr_0.PFET_GATE_10uA.t12 VDDA.t9 VDDA.t8 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X75 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.t10 VDDA.t354 VDDA.t356 VDDA.t355 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X76 VDDA.t14 bgr_0.PFET_GATE_10uA.t13 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.t13 VDDA.t13 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X77 VOUT+.t31 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t126 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X78 bgr_0.V_TOP.t20 VDDA.t104 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X79 bgr_0.1st_Vout_2.t7 bgr_0.V_CUR_REF_REG.t4 bgr_0.V_p_2.t8 GNDA.t159 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X80 two_stage_opamp_dummy_magic_14_0.VD4.t19 two_stage_opamp_dummy_magic_14_0.Vb2.t12 two_stage_opamp_dummy_magic_14_0.Y.t7 two_stage_opamp_dummy_magic_14_0.VD4.t18 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X81 VOUT+.t2 two_stage_opamp_dummy_magic_14_0.V_b_2nd_stage.t3 GNDA.t19 GNDA.t18 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X82 VDDA.t120 two_stage_opamp_dummy_magic_14_0.Y.t27 VOUT+.t10 VDDA.t119 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X83 two_stage_opamp_dummy_magic_14_0.VD2.t10 two_stage_opamp_dummy_magic_14_0.Vb1.t9 two_stage_opamp_dummy_magic_14_0.Y.t18 GNDA.t0 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X84 VOUT-.t30 two_stage_opamp_dummy_magic_14_0.cap_res_X.t127 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X85 two_stage_opamp_dummy_magic_14_0.VD4.t35 two_stage_opamp_dummy_magic_14_0.Vb3.t10 VDDA.t257 VDDA.t256 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X86 VOUT-.t31 two_stage_opamp_dummy_magic_14_0.cap_res_X.t126 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X87 VOUT-.t32 two_stage_opamp_dummy_magic_14_0.cap_res_X.t125 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X88 VOUT-.t3 a_14010_2720.t0 GNDA.t38 sky130_fd_pr__res_xhigh_po_0p35 l=2.63
X89 bgr_0.PFET_GATE_10uA.t5 bgr_0.1st_Vout_2.t13 VDDA.t405 VDDA.t404 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X90 VOUT-.t33 two_stage_opamp_dummy_magic_14_0.cap_res_X.t124 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X91 bgr_0.V_TOP.t21 VDDA.t121 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X92 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.t9 two_stage_opamp_dummy_magic_14_0.X.t28 GNDA.t8 VDDA.t10 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X93 GNDA.t287 GNDA.t285 two_stage_opamp_dummy_magic_14_0.V_source.t30 GNDA.t286 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=0.5 ps=2.9 w=2.5 l=0.15
X94 bgr_0.START_UP_NFET1.t0 bgr_0.START_UP_NFET1 GNDA.t128 GNDA.t127 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X95 VDDA.t353 VDDA.t351 GNDA.t84 VDDA.t352 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X96 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.t8 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.t6 two_stage_opamp_dummy_magic_14_0.Vb3.t1 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.t7 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X97 two_stage_opamp_dummy_magic_14_0.VD3.t17 two_stage_opamp_dummy_magic_14_0.Vb2.t13 two_stage_opamp_dummy_magic_14_0.X.t14 two_stage_opamp_dummy_magic_14_0.VD3.t16 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X98 VOUT+.t32 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t125 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X99 GNDA.t37 two_stage_opamp_dummy_magic_14_0.err_amp_mir.t0 two_stage_opamp_dummy_magic_14_0.err_amp_mir.t1 GNDA.t36 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X100 two_stage_opamp_dummy_magic_14_0.V_source.t34 VIN+.t1 two_stage_opamp_dummy_magic_14_0.VD2.t18 GNDA.t160 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X101 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.t8 two_stage_opamp_dummy_magic_14_0.Y.t28 VDDA.t71 GNDA.t54 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X102 two_stage_opamp_dummy_magic_14_0.V_source.t10 VIN+.t2 two_stage_opamp_dummy_magic_14_0.VD2.t1 GNDA.t131 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X103 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t10 GNDA.t282 GNDA.t284 GNDA.t283 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X104 VOUT+.t33 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t124 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X105 bgr_0.V_TOP.t22 VDDA.t122 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X106 GNDA.t197 bgr_0.NFET_GATE_10uA.t7 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.t12 GNDA.t196 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X107 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.t11 bgr_0.NFET_GATE_10uA.t8 GNDA.t195 GNDA.t194 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X108 two_stage_opamp_dummy_magic_14_0.VD4.t17 two_stage_opamp_dummy_magic_14_0.Vb2.t14 two_stage_opamp_dummy_magic_14_0.Y.t5 two_stage_opamp_dummy_magic_14_0.VD4.t16 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X109 GNDA.t53 two_stage_opamp_dummy_magic_14_0.Y.t29 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.t8 VDDA.t70 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X110 VOUT-.t34 two_stage_opamp_dummy_magic_14_0.cap_res_X.t123 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X111 VOUT-.t35 two_stage_opamp_dummy_magic_14_0.cap_res_X.t122 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X112 VOUT-.t36 two_stage_opamp_dummy_magic_14_0.cap_res_X.t121 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X113 VOUT-.t37 two_stage_opamp_dummy_magic_14_0.cap_res_X.t120 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X114 bgr_0.1st_Vout_2.t14 bgr_0.cap_res2.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X115 VOUT+.t34 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t123 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X116 VOUT+.t35 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t122 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X117 VOUT+.t36 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t121 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X118 VOUT+.t37 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t120 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X119 VOUT+.t38 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t119 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X120 a_12530_23988.t1 bgr_0.Vin-.t6 GNDA.t126 sky130_fd_pr__res_xhigh_po_0p35 l=6
X121 two_stage_opamp_dummy_magic_14_0.VD3.t27 two_stage_opamp_dummy_magic_14_0.Vb3.t11 VDDA.t255 VDDA.t254 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X122 two_stage_opamp_dummy_magic_14_0.VD3.t5 two_stage_opamp_dummy_magic_14_0.Vb2.t15 two_stage_opamp_dummy_magic_14_0.X.t3 two_stage_opamp_dummy_magic_14_0.VD3.t4 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X123 VOUT-.t38 two_stage_opamp_dummy_magic_14_0.cap_res_X.t119 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X124 VOUT-.t39 two_stage_opamp_dummy_magic_14_0.cap_res_X.t118 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X125 bgr_0.1st_Vout_2.t2 bgr_0.V_mir2.t18 VDDA.t45 VDDA.t44 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X126 two_stage_opamp_dummy_magic_14_0.V_err_p.t3 two_stage_opamp_dummy_magic_14_0.V_tot.t4 two_stage_opamp_dummy_magic_14_0.err_amp_mir.t4 VDDA.t376 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X127 VOUT-.t0 two_stage_opamp_dummy_magic_14_0.X.t29 VDDA.t12 VDDA.t11 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X128 two_stage_opamp_dummy_magic_14_0.VD1.t18 two_stage_opamp_dummy_magic_14_0.Vb1.t10 two_stage_opamp_dummy_magic_14_0.X.t1 GNDA.t6 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X129 VOUT-.t40 two_stage_opamp_dummy_magic_14_0.cap_res_X.t117 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X130 VOUT-.t41 two_stage_opamp_dummy_magic_14_0.cap_res_X.t116 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X131 bgr_0.1st_Vout_2.t15 bgr_0.cap_res2.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X132 VOUT-.t42 two_stage_opamp_dummy_magic_14_0.cap_res_X.t115 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X133 VOUT+.t39 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t118 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X134 two_stage_opamp_dummy_magic_14_0.V_p_mir.t3 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t13 GNDA.t307 GNDA.t306 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X135 two_stage_opamp_dummy_magic_14_0.V_source.t28 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t14 GNDA.t74 GNDA.t73 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X136 two_stage_opamp_dummy_magic_14_0.VD2.t9 two_stage_opamp_dummy_magic_14_0.Vb1.t11 two_stage_opamp_dummy_magic_14_0.Y.t17 GNDA.t130 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X137 VOUT-.t43 two_stage_opamp_dummy_magic_14_0.cap_res_X.t114 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X138 VOUT+.t40 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t117 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X139 VOUT+.t41 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t116 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X140 bgr_0.1st_Vout_1.t15 bgr_0.cap_res1.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X141 VOUT+.t42 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t115 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X142 bgr_0.V_mir1.t1 bgr_0.Vin-.t8 bgr_0.V_p_1.t4 GNDA.t69 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X143 bgr_0.V_mir1.t14 bgr_0.V_mir1.t13 VDDA.t43 VDDA.t42 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X144 two_stage_opamp_dummy_magic_14_0.VD3.t26 two_stage_opamp_dummy_magic_14_0.Vb3.t12 VDDA.t253 VDDA.t252 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X145 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t1 VIN-.t1 two_stage_opamp_dummy_magic_14_0.V_p_mir.t1 GNDA.t35 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X146 two_stage_opamp_dummy_magic_14_0.V_source.t4 VIN-.t2 two_stage_opamp_dummy_magic_14_0.VD1.t8 GNDA.t17 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X147 GNDA.t97 a_7580_22380.t1 GNDA.t2 sky130_fd_pr__res_xhigh_po_0p35 l=6
X148 VOUT-.t44 two_stage_opamp_dummy_magic_14_0.cap_res_X.t113 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X149 VOUT-.t45 two_stage_opamp_dummy_magic_14_0.cap_res_X.t112 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X150 VOUT+.t43 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t114 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X151 GNDA.t72 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t15 two_stage_opamp_dummy_magic_14_0.V_source.t27 GNDA.t71 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X152 VOUT-.t46 two_stage_opamp_dummy_magic_14_0.cap_res_X.t111 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X153 VOUT-.t47 two_stage_opamp_dummy_magic_14_0.cap_res_X.t110 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X154 GNDA.t122 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t16 two_stage_opamp_dummy_magic_14_0.V_source.t26 GNDA.t121 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X155 VDDA.t219 bgr_0.PFET_GATE_10uA.t14 two_stage_opamp_dummy_magic_14_0.Vb1.t3 VDDA.t218 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X156 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.t8 two_stage_opamp_dummy_magic_14_0.X.t30 GNDA.t61 VDDA.t76 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X157 VOUT-.t48 two_stage_opamp_dummy_magic_14_0.cap_res_X.t109 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X158 bgr_0.V_TOP.t23 VDDA.t123 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X159 two_stage_opamp_dummy_magic_14_0.V_source.t0 VIN+.t3 two_stage_opamp_dummy_magic_14_0.VD2.t0 GNDA.t0 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X160 VDDA.t350 VDDA.t348 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.t15 VDDA.t349 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X161 VOUT-.t49 two_stage_opamp_dummy_magic_14_0.cap_res_X.t108 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X162 VOUT-.t50 two_stage_opamp_dummy_magic_14_0.cap_res_X.t107 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X163 GNDA.t78 two_stage_opamp_dummy_magic_14_0.V_b_2nd_stage.t4 VOUT+.t11 GNDA.t77 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X164 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.t13 bgr_0.PFET_GATE_10uA.t15 VDDA.t215 VDDA.t214 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X165 a_5700_5524.t1 two_stage_opamp_dummy_magic_14_0.V_tot.t3 GNDA.t120 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X166 VOUT+.t44 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t113 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X167 VOUT+.t45 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t112 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X168 VDDA.t251 two_stage_opamp_dummy_magic_14_0.Vb3.t13 two_stage_opamp_dummy_magic_14_0.VD4.t34 VDDA.t250 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X169 VOUT+.t1 two_stage_opamp_dummy_magic_14_0.Y.t30 VDDA.t20 VDDA.t19 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X170 GNDA.t115 VDDA.t345 VDDA.t347 VDDA.t346 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X171 bgr_0.V_mir1.t15 bgr_0.Vin-.t9 bgr_0.V_p_1.t3 GNDA.t301 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X172 VOUT+.t46 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t111 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X173 VOUT+.t47 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t110 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X174 two_stage_opamp_dummy_magic_14_0.VD3.t15 two_stage_opamp_dummy_magic_14_0.Vb2.t16 two_stage_opamp_dummy_magic_14_0.X.t13 two_stage_opamp_dummy_magic_14_0.VD3.t14 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X175 bgr_0.START_UP.t2 bgr_0.V_TOP.t24 VDDA.t407 VDDA.t406 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X176 VOUT-.t51 two_stage_opamp_dummy_magic_14_0.cap_res_X.t106 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X177 bgr_0.PFET_GATE_10uA.t4 bgr_0.1st_Vout_2.t16 VDDA.t157 VDDA.t156 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X178 VDDA.t159 bgr_0.V_mir1.t18 bgr_0.1st_Vout_1.t4 VDDA.t158 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X179 VOUT+.t48 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t109 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X180 VOUT+.t49 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t108 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X181 VOUT-.t52 two_stage_opamp_dummy_magic_14_0.cap_res_X.t105 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X182 VOUT-.t53 two_stage_opamp_dummy_magic_14_0.cap_res_X.t104 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X183 two_stage_opamp_dummy_magic_14_0.Vb2.t8 bgr_0.NFET_GATE_10uA.t9 GNDA.t193 GNDA.t192 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X184 VDDA.t249 two_stage_opamp_dummy_magic_14_0.Vb3.t14 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.t9 VDDA.t248 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X185 GNDA.t191 bgr_0.NFET_GATE_10uA.t10 two_stage_opamp_dummy_magic_14_0.Vb2.t7 GNDA.t190 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X186 VOUT+.t50 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t107 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X187 bgr_0.V_TOP.t25 VDDA.t408 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X188 GNDA.t189 bgr_0.NFET_GATE_10uA.t11 two_stage_opamp_dummy_magic_14_0.Vb2.t6 GNDA.t188 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X189 two_stage_opamp_dummy_magic_14_0.Y.t11 two_stage_opamp_dummy_magic_14_0.Vb2.t17 two_stage_opamp_dummy_magic_14_0.VD4.t15 two_stage_opamp_dummy_magic_14_0.VD4.t14 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X190 VOUT+.t51 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t106 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X191 VOUT-.t54 two_stage_opamp_dummy_magic_14_0.cap_res_X.t103 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X192 VOUT-.t8 two_stage_opamp_dummy_magic_14_0.X.t31 VDDA.t78 VDDA.t77 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X193 two_stage_opamp_dummy_magic_14_0.VD1.t17 two_stage_opamp_dummy_magic_14_0.Vb1.t12 two_stage_opamp_dummy_magic_14_0.X.t17 GNDA.t7 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X194 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.t7 two_stage_opamp_dummy_magic_14_0.Y.t31 GNDA.t297 VDDA.t385 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X195 VDDA.t247 two_stage_opamp_dummy_magic_14_0.Vb3.t15 two_stage_opamp_dummy_magic_14_0.VD4.t33 VDDA.t246 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X196 VOUT+.t52 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t105 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X197 VOUT+.t53 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t104 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X198 VOUT+.t54 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t103 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X199 VOUT+.t55 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t102 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X200 two_stage_opamp_dummy_magic_14_0.VD3.t25 two_stage_opamp_dummy_magic_14_0.Vb3.t16 VDDA.t245 VDDA.t244 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X201 VDDA.t410 bgr_0.V_TOP.t26 bgr_0.Vin+.t2 VDDA.t409 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X202 two_stage_opamp_dummy_magic_14_0.V_source.t25 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t17 GNDA.t303 GNDA.t302 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X203 bgr_0.1st_Vout_2.t1 bgr_0.V_mir2.t19 VDDA.t37 VDDA.t36 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X204 VOUT-.t55 two_stage_opamp_dummy_magic_14_0.cap_res_X.t102 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X205 two_stage_opamp_dummy_magic_14_0.V_b_2nd_stage.t1 a_14010_2720.t1 GNDA.t119 sky130_fd_pr__res_xhigh_po_0p35 l=2.63
X206 bgr_0.V_TOP.t3 bgr_0.1st_Vout_1.t16 VDDA.t155 VDDA.t154 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X207 bgr_0.V_CUR_REF_REG.t2 VDDA.t342 VDDA.t344 VDDA.t343 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X208 VOUT-.t56 two_stage_opamp_dummy_magic_14_0.cap_res_X.t101 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X209 VOUT-.t57 two_stage_opamp_dummy_magic_14_0.cap_res_X.t100 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X210 VOUT-.t58 two_stage_opamp_dummy_magic_14_0.cap_res_X.t99 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X211 VOUT+.t56 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t101 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X212 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t6 bgr_0.PFET_GATE_10uA.t16 VDDA.t165 VDDA.t164 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X213 VOUT-.t59 two_stage_opamp_dummy_magic_14_0.cap_res_X.t98 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X214 two_stage_opamp_dummy_magic_14_0.V_source.t8 VIN-.t3 two_stage_opamp_dummy_magic_14_0.VD1.t7 GNDA.t6 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X215 VDDA.t149 two_stage_opamp_dummy_magic_14_0.X.t32 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.t7 GNDA.t101 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X216 two_stage_opamp_dummy_magic_14_0.X.t24 two_stage_opamp_dummy_magic_14_0.Vb2.t18 two_stage_opamp_dummy_magic_14_0.VD3.t37 two_stage_opamp_dummy_magic_14_0.VD3.t36 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X217 VOUT+.t57 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t100 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X218 GNDA.t316 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t18 two_stage_opamp_dummy_magic_14_0.V_source.t24 GNDA.t315 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X219 VOUT+.t58 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t99 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X220 bgr_0.1st_Vout_2.t17 bgr_0.cap_res2.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X221 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.t7 two_stage_opamp_dummy_magic_14_0.X.t33 GNDA.t102 VDDA.t150 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X222 two_stage_opamp_dummy_magic_14_0.Y.t9 two_stage_opamp_dummy_magic_14_0.Vb2.t19 two_stage_opamp_dummy_magic_14_0.VD4.t13 two_stage_opamp_dummy_magic_14_0.VD4.t12 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X223 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.t7 two_stage_opamp_dummy_magic_14_0.Y.t32 VDDA.t387 GNDA.t299 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X224 bgr_0.Vin+.t5 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t0 GNDA.t50 sky130_fd_pr__res_xhigh_po_0p35 l=2.3
X225 two_stage_opamp_dummy_magic_14_0.V_source.t32 VIN+.t4 two_stage_opamp_dummy_magic_14_0.VD2.t16 GNDA.t130 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X226 VOUT+.t59 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t98 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X227 VOUT+.t60 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t97 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X228 VOUT-.t60 two_stage_opamp_dummy_magic_14_0.cap_res_X.t97 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X229 VOUT-.t61 two_stage_opamp_dummy_magic_14_0.cap_res_X.t96 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X230 bgr_0.1st_Vout_2.t18 bgr_0.cap_res2.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X231 bgr_0.Vin+.t1 bgr_0.V_TOP.t27 VDDA.t106 VDDA.t105 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X232 VOUT-.t62 two_stage_opamp_dummy_magic_14_0.cap_res_X.t95 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X233 VDDA.t341 VDDA.t339 bgr_0.PFET_GATE_10uA.t9 VDDA.t340 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.2
X234 VOUT+.t61 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t96 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X235 VDDA.t108 bgr_0.V_TOP.t28 bgr_0.Vin+.t0 VDDA.t107 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X236 VOUT+.t6 two_stage_opamp_dummy_magic_14_0.Y.t33 VDDA.t58 VDDA.t57 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X237 VOUT+.t62 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t95 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X238 a_5580_5524.t0 two_stage_opamp_dummy_magic_14_0.V_tot.t2 GNDA.t109 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X239 bgr_0.1st_Vout_1.t17 bgr_0.cap_res1.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X240 GNDA.t34 a_12410_22380.t0 GNDA.t33 sky130_fd_pr__res_xhigh_po_0p35 l=6
X241 GNDA.t187 bgr_0.NFET_GATE_10uA.t12 two_stage_opamp_dummy_magic_14_0.Vb3.t3 GNDA.t186 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X242 VOUT-.t63 two_stage_opamp_dummy_magic_14_0.cap_res_X.t94 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X243 VOUT-.t64 two_stage_opamp_dummy_magic_14_0.cap_res_X.t93 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X244 VDDA.t243 two_stage_opamp_dummy_magic_14_0.Vb3.t17 two_stage_opamp_dummy_magic_14_0.VD3.t24 VDDA.t242 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X245 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t0 two_stage_opamp_dummy_magic_14_0.Y.t12 GNDA.t108 sky130_fd_pr__res_high_po_1p41 l=1.41
X246 VOUT+.t63 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t94 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X247 bgr_0.cap_res1.t20 bgr_0.V_TOP.t12 GNDA.t308 sky130_fd_pr__res_high_po_0p35 l=2.05
X248 two_stage_opamp_dummy_magic_14_0.Vb3.t5 bgr_0.NFET_GATE_10uA.t13 GNDA.t185 GNDA.t184 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X249 bgr_0.V_mir2.t9 bgr_0.V_mir2.t8 VDDA.t85 VDDA.t84 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X250 VDDA.t338 VDDA.t336 bgr_0.V_TOP.t8 VDDA.t337 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X251 two_stage_opamp_dummy_magic_14_0.X.t12 two_stage_opamp_dummy_magic_14_0.Vb2.t20 two_stage_opamp_dummy_magic_14_0.VD3.t13 two_stage_opamp_dummy_magic_14_0.VD3.t12 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X252 VOUT+.t64 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t93 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X253 VOUT+.t65 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t92 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X254 bgr_0.1st_Vout_1.t18 bgr_0.cap_res1.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X255 VOUT-.t65 two_stage_opamp_dummy_magic_14_0.cap_res_X.t92 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X256 VOUT+.t66 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t91 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X257 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.t2 bgr_0.V_TOP.t29 VDDA.t110 VDDA.t109 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X258 bgr_0.1st_Vout_2.t19 bgr_0.cap_res2.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X259 VOUT-.t12 two_stage_opamp_dummy_magic_14_0.X.t34 VDDA.t142 VDDA.t141 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X260 VOUT-.t66 two_stage_opamp_dummy_magic_14_0.cap_res_X.t91 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X261 GNDA.t14 a_13060_22630.t0 GNDA.t13 sky130_fd_pr__res_xhigh_po_0p35 l=4
X262 VOUT-.t13 two_stage_opamp_dummy_magic_14_0.X.t35 VDDA.t144 VDDA.t143 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X263 two_stage_opamp_dummy_magic_14_0.VD1.t16 two_stage_opamp_dummy_magic_14_0.Vb1.t13 two_stage_opamp_dummy_magic_14_0.X.t16 GNDA.t98 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X264 VOUT+.t67 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t90 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X265 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.t6 two_stage_opamp_dummy_magic_14_0.Y.t34 GNDA.t142 VDDA.t211 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X266 VDDA.t335 VDDA.t333 GNDA.t161 VDDA.t334 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X267 bgr_0.1st_Vout_1.t3 bgr_0.V_mir1.t19 VDDA.t161 VDDA.t160 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X268 bgr_0.1st_Vout_1.t19 bgr_0.cap_res1.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X269 two_stage_opamp_dummy_magic_14_0.X.t22 two_stage_opamp_dummy_magic_14_0.Vb2.t21 two_stage_opamp_dummy_magic_14_0.VD3.t33 two_stage_opamp_dummy_magic_14_0.VD3.t32 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X270 VOUT-.t67 two_stage_opamp_dummy_magic_14_0.cap_res_X.t90 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X271 two_stage_opamp_dummy_magic_14_0.V_err_gate.t4 VDDA.t330 VDDA.t332 VDDA.t331 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=1 ps=5.8 w=2.5 l=0.15
X272 two_stage_opamp_dummy_magic_14_0.V_source.t23 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t19 GNDA.t296 GNDA.t295 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X273 VDDA.t241 two_stage_opamp_dummy_magic_14_0.Vb3.t18 two_stage_opamp_dummy_magic_14_0.VD3.t23 VDDA.t240 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X274 bgr_0.NFET_GATE_10uA.t2 bgr_0.PFET_GATE_10uA.t17 VDDA.t91 VDDA.t90 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X275 VDDA.t7 bgr_0.PFET_GATE_10uA.t18 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t0 VDDA.t6 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X276 two_stage_opamp_dummy_magic_14_0.Y.t6 two_stage_opamp_dummy_magic_14_0.Vb2.t22 two_stage_opamp_dummy_magic_14_0.VD4.t11 two_stage_opamp_dummy_magic_14_0.VD4.t10 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X277 VOUT+.t68 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t89 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X278 VOUT+.t69 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t88 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X279 bgr_0.1st_Vout_1.t20 bgr_0.cap_res1.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X280 GNDA.t23 two_stage_opamp_dummy_magic_14_0.V_b_2nd_stage.t5 VOUT-.t1 GNDA.t22 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X281 bgr_0.V_p_2.t4 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.t7 bgr_0.V_mir2.t16 GNDA.t39 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X282 VDDA.t79 two_stage_opamp_dummy_magic_14_0.X.t36 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.t6 GNDA.t62 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X283 two_stage_opamp_dummy_magic_14_0.V_source.t3 VIN-.t4 two_stage_opamp_dummy_magic_14_0.VD1.t6 GNDA.t7 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X284 VDDA.t132 bgr_0.V_TOP.t30 bgr_0.START_UP.t1 VDDA.t131 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X285 VOUT+.t70 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t87 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X286 VOUT-.t68 two_stage_opamp_dummy_magic_14_0.cap_res_X.t89 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X287 GNDA.t107 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t20 two_stage_opamp_dummy_magic_14_0.V_source.t22 GNDA.t106 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X288 VOUT-.t69 two_stage_opamp_dummy_magic_14_0.cap_res_X.t88 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X289 a_5700_5524.t0 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.t10 GNDA.t32 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X290 VOUT+.t71 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t86 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X291 VOUT+.t72 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t85 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X292 bgr_0.V_TOP.t31 VDDA.t133 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X293 bgr_0.V_TOP.t10 bgr_0.1st_Vout_1.t21 VDDA.t397 VDDA.t396 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X294 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.t6 two_stage_opamp_dummy_magic_14_0.X.t37 GNDA.t63 VDDA.t80 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X295 two_stage_opamp_dummy_magic_14_0.X.t10 two_stage_opamp_dummy_magic_14_0.Vb1.t14 two_stage_opamp_dummy_magic_14_0.VD1.t15 GNDA.t87 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X296 VOUT+.t73 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t84 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X297 two_stage_opamp_dummy_magic_14_0.VD4.t32 two_stage_opamp_dummy_magic_14_0.Vb3.t19 VDDA.t239 VDDA.t238 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X298 two_stage_opamp_dummy_magic_14_0.X.t2 two_stage_opamp_dummy_magic_14_0.Vb2.t23 two_stage_opamp_dummy_magic_14_0.VD3.t3 two_stage_opamp_dummy_magic_14_0.VD3.t2 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X299 VDDA.t329 VDDA.t327 two_stage_opamp_dummy_magic_14_0.V_err_gate.t3 VDDA.t328 sky130_fd_pr__pfet_01v8 ad=1 pd=5.8 as=0.5 ps=2.9 w=2.5 l=0.15
X300 GNDA.t281 GNDA.t279 VOUT-.t15 GNDA.t280 sky130_fd_pr__nfet_01v8 ad=2.8 pd=14.8 as=1.4 ps=7.4 w=7 l=0.6
X301 VOUT+.t5 two_stage_opamp_dummy_magic_14_0.Y.t35 VDDA.t56 VDDA.t55 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X302 VOUT-.t70 two_stage_opamp_dummy_magic_14_0.cap_res_X.t87 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X303 GNDA.t41 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t21 two_stage_opamp_dummy_magic_14_0.V_source.t21 GNDA.t40 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X304 two_stage_opamp_dummy_magic_14_0.Y.t21 two_stage_opamp_dummy_magic_14_0.Vb1.t15 two_stage_opamp_dummy_magic_14_0.VD2.t8 GNDA.t105 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X305 VOUT-.t71 two_stage_opamp_dummy_magic_14_0.cap_res_X.t86 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X306 bgr_0.V_TOP.t13 bgr_0.1st_Vout_1.t22 VDDA.t412 VDDA.t411 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X307 VOUT+.t74 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t83 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X308 VOUT+.t75 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t82 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X309 VOUT+.t76 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t81 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X310 bgr_0.NFET_GATE_10uA.t4 bgr_0.NFET_GATE_10uA.t3 GNDA.t183 GNDA.t182 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X311 GNDA.t181 bgr_0.NFET_GATE_10uA.t14 two_stage_opamp_dummy_magic_14_0.Vb3.t4 GNDA.t180 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X312 VOUT+.t77 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t80 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X313 bgr_0.V_TOP.t32 VDDA.t134 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X314 a_6810_23838.t0 a_6930_22664.t0 GNDA.t65 sky130_fd_pr__res_xhigh_po_0p35 l=3.83
X315 VDDA.t326 VDDA.t324 VDDA.t326 VDDA.t325 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0 ps=0 w=3.5 l=0.2
X316 two_stage_opamp_dummy_magic_14_0.VD4.t9 two_stage_opamp_dummy_magic_14_0.Vb2.t24 two_stage_opamp_dummy_magic_14_0.Y.t3 two_stage_opamp_dummy_magic_14_0.VD4.t8 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X317 bgr_0.1st_Vout_2.t20 bgr_0.cap_res2.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X318 VOUT-.t72 two_stage_opamp_dummy_magic_14_0.cap_res_X.t85 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X319 VOUT-.t73 two_stage_opamp_dummy_magic_14_0.cap_res_X.t84 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X320 VDDA.t169 two_stage_opamp_dummy_magic_14_0.Y.t36 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.t6 GNDA.t114 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X321 VOUT-.t74 two_stage_opamp_dummy_magic_14_0.cap_res_X.t83 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X322 VOUT+.t78 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t79 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X323 two_stage_opamp_dummy_magic_14_0.VD4.t31 two_stage_opamp_dummy_magic_14_0.Vb3.t20 VDDA.t237 VDDA.t236 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X324 VOUT-.t17 VDDA.t321 VDDA.t323 VDDA.t322 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=2.4 ps=12.8 w=6 l=0.15
X325 VDDA.t5 bgr_0.PFET_GATE_10uA.t19 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.t12 VDDA.t4 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X326 VDDA.t320 VDDA.t318 two_stage_opamp_dummy_magic_14_0.VD3.t31 VDDA.t319 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X327 VOUT-.t75 two_stage_opamp_dummy_magic_14_0.cap_res_X.t82 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X328 bgr_0.1st_Vout_1.t23 bgr_0.cap_res1.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X329 bgr_0.V_mir1.t12 bgr_0.V_mir1.t11 VDDA.t206 VDDA.t205 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X330 VDDA.t389 bgr_0.V_TOP.t33 bgr_0.START_UP.t0 VDDA.t388 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X331 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.t5 two_stage_opamp_dummy_magic_14_0.Y.t37 GNDA.t141 VDDA.t210 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X332 VOUT-.t76 two_stage_opamp_dummy_magic_14_0.cap_res_X.t81 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X333 bgr_0.1st_Vout_2.t21 bgr_0.cap_res2.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X334 VOUT+.t79 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t78 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X335 VOUT+.t80 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t77 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X336 a_7460_23988.t0 a_7580_22380.t0 GNDA.t2 sky130_fd_pr__res_xhigh_po_0p35 l=6
X337 bgr_0.V_p_2.t7 bgr_0.V_CUR_REF_REG.t5 bgr_0.1st_Vout_2.t5 GNDA.t145 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X338 VOUT-.t77 two_stage_opamp_dummy_magic_14_0.cap_res_X.t80 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X339 two_stage_opamp_dummy_magic_14_0.V_source.t20 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t22 GNDA.t45 GNDA.t44 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X340 VOUT+.t81 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t76 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X341 two_stage_opamp_dummy_magic_14_0.VD3.t19 two_stage_opamp_dummy_magic_14_0.Vb2.t25 two_stage_opamp_dummy_magic_14_0.X.t15 two_stage_opamp_dummy_magic_14_0.VD3.t18 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X342 VDDA.t147 two_stage_opamp_dummy_magic_14_0.X.t38 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.t5 GNDA.t99 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X343 bgr_0.1st_Vout_2.t22 bgr_0.cap_res2.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X344 two_stage_opamp_dummy_magic_14_0.VD4.t7 two_stage_opamp_dummy_magic_14_0.Vb2.t26 two_stage_opamp_dummy_magic_14_0.Y.t10 two_stage_opamp_dummy_magic_14_0.VD4.t6 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X345 two_stage_opamp_dummy_magic_14_0.V_source.t9 VIN-.t5 two_stage_opamp_dummy_magic_14_0.VD1.t5 GNDA.t98 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X346 GNDA.t138 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t23 two_stage_opamp_dummy_magic_14_0.V_source.t19 GNDA.t137 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X347 bgr_0.1st_Vout_1.t6 bgr_0.Vin+.t8 bgr_0.V_p_1.t7 GNDA.t11 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X348 VDDA.t204 bgr_0.V_mir2.t20 bgr_0.1st_Vout_2.t4 VDDA.t203 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X349 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.t5 two_stage_opamp_dummy_magic_14_0.X.t39 GNDA.t100 VDDA.t148 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X350 VOUT-.t78 two_stage_opamp_dummy_magic_14_0.cap_res_X.t79 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X351 VOUT-.t79 two_stage_opamp_dummy_magic_14_0.cap_res_X.t78 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X352 bgr_0.1st_Vout_1.t24 bgr_0.cap_res1.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X353 GNDA.t218 GNDA.t217 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t8 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X354 VOUT-.t80 two_stage_opamp_dummy_magic_14_0.cap_res_X.t77 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X355 bgr_0.1st_Vout_2.t23 bgr_0.cap_res2.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X356 GNDA.t179 bgr_0.NFET_GATE_10uA.t15 two_stage_opamp_dummy_magic_14_0.Vb2.t5 GNDA.t178 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X357 two_stage_opamp_dummy_magic_14_0.Vb2.t4 bgr_0.NFET_GATE_10uA.t16 GNDA.t177 GNDA.t176 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X358 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.t13 GNDA.t214 GNDA.t216 GNDA.t215 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X359 VOUT+.t82 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t75 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X360 GNDA.t209 GNDA.t278 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t7 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X361 GNDA.t277 GNDA.t275 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.t14 GNDA.t276 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X362 GNDA.t274 GNDA.t272 two_stage_opamp_dummy_magic_14_0.Vb2.t10 GNDA.t273 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X363 VOUT-.t81 two_stage_opamp_dummy_magic_14_0.cap_res_X.t76 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X364 two_stage_opamp_dummy_magic_14_0.V_err_mir_p.t0 two_stage_opamp_dummy_magic_14_0.V_err_gate.t8 VDDA.t173 VDDA.t172 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X365 VOUT+.t83 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t74 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X366 bgr_0.PFET_GATE_10uA.t8 VDDA.t315 VDDA.t317 VDDA.t316 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.2
X367 two_stage_opamp_dummy_magic_14_0.VD3.t22 two_stage_opamp_dummy_magic_14_0.Vb3.t21 VDDA.t235 VDDA.t234 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X368 VOUT+.t84 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t73 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X369 bgr_0.1st_Vout_1.t2 bgr_0.V_mir1.t20 VDDA.t185 VDDA.t184 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X370 VOUT+.t4 two_stage_opamp_dummy_magic_14_0.Y.t38 VDDA.t54 VDDA.t53 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X371 two_stage_opamp_dummy_magic_14_0.Y.t14 two_stage_opamp_dummy_magic_14_0.Vb1.t16 two_stage_opamp_dummy_magic_14_0.VD2.t7 GNDA.t83 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X372 two_stage_opamp_dummy_magic_14_0.Vb2_2.t2 two_stage_opamp_dummy_magic_14_0.Vb2.t27 VDDA.t208 VDDA.t207 sky130_fd_pr__pfet_01v8 ad=0.36 pd=2.2 as=0.36 ps=2.2 w=1.8 l=0.2
X373 VOUT-.t82 two_stage_opamp_dummy_magic_14_0.cap_res_X.t75 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X374 VOUT-.t14 GNDA.t269 GNDA.t271 GNDA.t270 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=2.8 ps=14.8 w=7 l=0.6
X375 two_stage_opamp_dummy_magic_14_0.VD4.t30 two_stage_opamp_dummy_magic_14_0.Vb3.t22 VDDA.t233 VDDA.t232 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X376 bgr_0.V_p_2.t6 bgr_0.V_CUR_REF_REG.t6 bgr_0.1st_Vout_2.t10 GNDA.t314 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.2
X377 VOUT-.t83 two_stage_opamp_dummy_magic_14_0.cap_res_X.t74 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X378 two_stage_opamp_dummy_magic_14_0.VD1.t4 VIN-.t6 two_stage_opamp_dummy_magic_14_0.V_source.t40 GNDA.t87 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X379 VOUT+.t85 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t72 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X380 GNDA.t209 GNDA.t268 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t6 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X381 VOUT-.t84 two_stage_opamp_dummy_magic_14_0.cap_res_X.t73 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X382 VOUT+.t86 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t71 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X383 GNDA.t209 GNDA.t208 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t5 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X384 VOUT-.t85 two_stage_opamp_dummy_magic_14_0.cap_res_X.t72 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X385 VDDA.t168 two_stage_opamp_dummy_magic_14_0.Y.t39 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.t5 GNDA.t113 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X386 two_stage_opamp_dummy_magic_14_0.VD2.t15 VIN+.t5 two_stage_opamp_dummy_magic_14_0.V_source.t31 GNDA.t105 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X387 VDDA.t181 bgr_0.V_mir2.t6 bgr_0.V_mir2.t7 VDDA.t180 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X388 VOUT+.t87 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t70 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X389 VOUT+.t88 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t69 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X390 VOUT+.t89 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t68 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X391 VOUT+.t90 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t67 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X392 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.t4 two_stage_opamp_dummy_magic_14_0.Y.t40 GNDA.t140 VDDA.t209 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X393 bgr_0.V_p_2.t5 bgr_0.V_CUR_REF_REG.t7 bgr_0.1st_Vout_2.t6 GNDA.t148 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X394 two_stage_opamp_dummy_magic_14_0.VD4.t25 two_stage_opamp_dummy_magic_14_0.VD4.t23 two_stage_opamp_dummy_magic_14_0.Y.t1 two_stage_opamp_dummy_magic_14_0.VD4.t24 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X395 VOUT+.t91 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t66 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X396 two_stage_opamp_dummy_magic_14_0.err_amp_mir.t2 GNDA.t265 GNDA.t267 GNDA.t266 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=1 ps=5.8 w=2.5 l=0.15
X397 a_13180_23838.t0 bgr_0.V_CUR_REF_REG.t0 GNDA.t64 sky130_fd_pr__res_xhigh_po_0p35 l=4
X398 VOUT-.t86 two_stage_opamp_dummy_magic_14_0.cap_res_X.t71 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X399 bgr_0.V_TOP.t34 VDDA.t390 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X400 VOUT-.t87 two_stage_opamp_dummy_magic_14_0.cap_res_X.t70 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X401 VOUT-.t88 two_stage_opamp_dummy_magic_14_0.cap_res_X.t69 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X402 VOUT-.t89 two_stage_opamp_dummy_magic_14_0.cap_res_X.t68 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X403 VOUT-.t90 two_stage_opamp_dummy_magic_14_0.cap_res_X.t67 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X404 VDDA.t139 two_stage_opamp_dummy_magic_14_0.X.t40 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.t4 GNDA.t94 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X405 VOUT-.t91 two_stage_opamp_dummy_magic_14_0.cap_res_X.t66 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X406 VOUT+.t92 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t65 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X407 bgr_0.V_TOP.t35 VDDA.t391 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X408 a_5580_5524.t1 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.t10 GNDA.t112 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X409 VDDA.t140 two_stage_opamp_dummy_magic_14_0.X.t41 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.t3 GNDA.t95 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X410 VDDA.t231 two_stage_opamp_dummy_magic_14_0.Vb3.t23 two_stage_opamp_dummy_magic_14_0.VD4.t29 VDDA.t230 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X411 VDDA.t130 bgr_0.1st_Vout_2.t24 bgr_0.PFET_GATE_10uA.t3 VDDA.t129 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X412 VDDA.t314 VDDA.t312 two_stage_opamp_dummy_magic_14_0.Vb1.t5 VDDA.t313 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X413 two_stage_opamp_dummy_magic_14_0.err_amp_out.t0 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.t8 two_stage_opamp_dummy_magic_14_0.V_err_p.t2 VDDA.t170 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X414 VOUT+.t93 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t64 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X415 two_stage_opamp_dummy_magic_14_0.Vb1.t4 VDDA.t309 VDDA.t311 VDDA.t310 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X416 VDDA.t136 two_stage_opamp_dummy_magic_14_0.X.t42 VOUT-.t10 VDDA.t135 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X417 two_stage_opamp_dummy_magic_14_0.X.t4 two_stage_opamp_dummy_magic_14_0.Vb1.t17 two_stage_opamp_dummy_magic_14_0.VD1.t14 GNDA.t24 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X418 VOUT-.t92 two_stage_opamp_dummy_magic_14_0.cap_res_X.t65 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X419 VDDA.t308 VDDA.t306 VOUT-.t16 VDDA.t307 sky130_fd_pr__pfet_01v8 ad=2.4 pd=12.8 as=1.2 ps=6.4 w=6 l=0.15
X420 VOUT+.t94 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t63 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X421 VOUT+.t95 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t62 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X422 VOUT+.t96 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t61 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X423 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.t12 bgr_0.PFET_GATE_10uA.t20 VDDA.t22 VDDA.t21 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X424 two_stage_opamp_dummy_magic_14_0.VD3.t11 two_stage_opamp_dummy_magic_14_0.VD3.t9 two_stage_opamp_dummy_magic_14_0.X.t7 two_stage_opamp_dummy_magic_14_0.VD3.t10 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X425 VOUT-.t93 two_stage_opamp_dummy_magic_14_0.cap_res_X.t64 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X426 VOUT-.t94 two_stage_opamp_dummy_magic_14_0.cap_res_X.t63 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X427 VDDA.t49 bgr_0.PFET_GATE_10uA.t21 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.t11 VDDA.t48 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X428 VOUT-.t95 two_stage_opamp_dummy_magic_14_0.cap_res_X.t62 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X429 VOUT+.t9 two_stage_opamp_dummy_magic_14_0.Y.t41 VDDA.t118 VDDA.t117 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X430 VOUT-.t96 two_stage_opamp_dummy_magic_14_0.cap_res_X.t61 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X431 two_stage_opamp_dummy_magic_14_0.V_err_mir_p.t2 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.t9 two_stage_opamp_dummy_magic_14_0.V_err_gate.t0 VDDA.t171 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X432 two_stage_opamp_dummy_magic_14_0.Y.t22 two_stage_opamp_dummy_magic_14_0.Vb1.t18 two_stage_opamp_dummy_magic_14_0.VD2.t6 GNDA.t46 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X433 two_stage_opamp_dummy_magic_14_0.cap_res_X.t0 two_stage_opamp_dummy_magic_14_0.X.t8 GNDA.t67 sky130_fd_pr__res_high_po_1p41 l=1.41
X434 VOUT-.t97 two_stage_opamp_dummy_magic_14_0.cap_res_X.t60 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X435 bgr_0.V_TOP.t36 VDDA.t23 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X436 VOUT-.t98 two_stage_opamp_dummy_magic_14_0.cap_res_X.t59 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X437 bgr_0.Vin-.t2 bgr_0.V_TOP.t37 VDDA.t25 VDDA.t24 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X438 two_stage_opamp_dummy_magic_14_0.Y.t8 two_stage_opamp_dummy_magic_14_0.Vb2.t28 two_stage_opamp_dummy_magic_14_0.VD4.t5 two_stage_opamp_dummy_magic_14_0.VD4.t4 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X439 VOUT-.t99 two_stage_opamp_dummy_magic_14_0.cap_res_X.t58 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X440 VDDA.t305 VDDA.t302 VDDA.t304 VDDA.t303 sky130_fd_pr__pfet_01v8 ad=0.72 pd=4.4 as=0 ps=0 w=1.8 l=0.2
X441 VOUT+.t97 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t60 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X442 a_14170_5524.t1 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.t14 GNDA.t313 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X443 VOUT+.t98 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t59 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X444 VDDA.t229 two_stage_opamp_dummy_magic_14_0.Vb3.t24 two_stage_opamp_dummy_magic_14_0.VD4.t28 VDDA.t228 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X445 VOUT+.t99 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t58 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X446 GNDA.t175 bgr_0.NFET_GATE_10uA.t17 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.t13 GNDA.t174 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X447 bgr_0.1st_Vout_1.t1 bgr_0.V_mir1.t21 VDDA.t187 VDDA.t186 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X448 two_stage_opamp_dummy_magic_14_0.Vb2.t9 GNDA.t262 GNDA.t264 GNDA.t263 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X449 VOUT+.t100 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t57 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X450 VOUT+.t101 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t56 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X451 VOUT+.t102 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t55 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X452 bgr_0.1st_Vout_1.t25 bgr_0.cap_res1.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X453 GNDA.t318 two_stage_opamp_dummy_magic_14_0.V_b_2nd_stage.t6 VOUT+.t18 GNDA.t317 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X454 VOUT-.t100 two_stage_opamp_dummy_magic_14_0.cap_res_X.t57 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X455 bgr_0.1st_Vout_2.t25 bgr_0.cap_res2.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X456 two_stage_opamp_dummy_magic_14_0.err_amp_out.t1 two_stage_opamp_dummy_magic_14_0.err_amp_mir.t5 GNDA.t117 GNDA.t116 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X457 VDDA.t196 two_stage_opamp_dummy_magic_14_0.Y.t42 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.t4 GNDA.t134 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X458 VOUT+.t103 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t54 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X459 two_stage_opamp_dummy_magic_14_0.VD2.t17 VIN+.t6 two_stage_opamp_dummy_magic_14_0.V_source.t33 GNDA.t83 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X460 VOUT-.t101 two_stage_opamp_dummy_magic_14_0.cap_res_X.t56 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X461 bgr_0.1st_Vout_1.t26 bgr_0.cap_res1.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X462 VOUT-.t102 two_stage_opamp_dummy_magic_14_0.cap_res_X.t55 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X463 VOUT-.t103 two_stage_opamp_dummy_magic_14_0.cap_res_X.t54 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X464 VOUT-.t104 two_stage_opamp_dummy_magic_14_0.cap_res_X.t53 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X465 VDDA.t227 two_stage_opamp_dummy_magic_14_0.Vb3.t25 two_stage_opamp_dummy_magic_14_0.VD4.t27 VDDA.t226 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X466 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t8 bgr_0.PFET_GATE_10uA.t22 VDDA.t213 VDDA.t212 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X467 VOUT-.t105 two_stage_opamp_dummy_magic_14_0.cap_res_X.t52 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X468 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.t1 bgr_0.V_TOP.t38 VDDA.t27 VDDA.t26 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X469 VOUT+.t104 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t53 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X470 GNDA.t261 GNDA.t259 VOUT+.t14 GNDA.t260 sky130_fd_pr__nfet_01v8 ad=2.8 pd=14.8 as=1.4 ps=7.4 w=7 l=0.6
X471 VDDA.t183 bgr_0.V_mir2.t4 bgr_0.V_mir2.t5 VDDA.t182 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X472 VOUT+.t105 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t52 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X473 VDDA.t167 bgr_0.V_mir1.t9 bgr_0.V_mir1.t10 VDDA.t166 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X474 VDDA.t112 bgr_0.PFET_GATE_10uA.t23 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t5 VDDA.t111 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X475 bgr_0.V_p_1.t2 bgr_0.Vin-.t10 bgr_0.V_mir1.t16 GNDA.t310 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X476 VDDA.t265 GNDA.t256 GNDA.t258 GNDA.t257 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=1.2 ps=6.8 w=3 l=0.15
X477 two_stage_opamp_dummy_magic_14_0.Vb2.t2 two_stage_opamp_dummy_magic_14_0.Vb2_2.t7 two_stage_opamp_dummy_magic_14_0.Vb2_2.t9 two_stage_opamp_dummy_magic_14_0.Vb2_2.t8 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X478 VOUT+.t106 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t51 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X479 bgr_0.1st_Vout_1.t27 bgr_0.cap_res1.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X480 bgr_0.1st_Vout_2.t26 bgr_0.cap_res2.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X481 VDDA.t189 two_stage_opamp_dummy_magic_14_0.V_err_gate.t9 two_stage_opamp_dummy_magic_14_0.V_err_p.t0 VDDA.t188 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X482 VOUT+.t107 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t50 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X483 two_stage_opamp_dummy_magic_14_0.X.t9 two_stage_opamp_dummy_magic_14_0.Vb1.t19 two_stage_opamp_dummy_magic_14_0.VD1.t13 GNDA.t25 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X484 VOUT+.t108 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t49 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X485 VDDA.t138 two_stage_opamp_dummy_magic_14_0.X.t43 VOUT-.t11 VDDA.t137 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X486 bgr_0.V_TOP.t7 VDDA.t299 VDDA.t301 VDDA.t300 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.2
X487 VOUT+.t109 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t48 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X488 bgr_0.1st_Vout_1.t28 bgr_0.cap_res1.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X489 VOUT-.t106 two_stage_opamp_dummy_magic_14_0.cap_res_X.t51 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X490 VDDA.t298 VDDA.t296 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.t6 VDDA.t297 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.8 as=0.6 ps=3.4 w=3 l=0.5
X491 VDDA.t295 VDDA.t293 two_stage_opamp_dummy_magic_14_0.Vb2_2.t3 VDDA.t294 sky130_fd_pr__pfet_01v8 ad=0.72 pd=4.4 as=0.36 ps=2.2 w=1.8 l=0.2
X492 a_14290_5524.t0 two_stage_opamp_dummy_magic_14_0.V_tot.t1 GNDA.t92 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X493 VOUT+.t16 VDDA.t290 VDDA.t292 VDDA.t291 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=2.4 ps=12.8 w=6 l=0.15
X494 VDDA.t289 VDDA.t287 two_stage_opamp_dummy_magic_14_0.VD4.t36 VDDA.t288 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X495 two_stage_opamp_dummy_magic_14_0.Y.t19 two_stage_opamp_dummy_magic_14_0.Vb1.t20 two_stage_opamp_dummy_magic_14_0.VD2.t5 GNDA.t149 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X496 bgr_0.V_p_1.t1 bgr_0.Vin-.t11 bgr_0.V_mir1.t0 GNDA.t9 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X497 VOUT+.t110 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t47 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X498 VOUT-.t107 two_stage_opamp_dummy_magic_14_0.cap_res_X.t50 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X499 VOUT+.t111 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t46 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X500 VOUT+.t112 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t45 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X501 VOUT+.t113 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t44 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X502 bgr_0.1st_Vout_1.t29 bgr_0.cap_res1.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X503 two_stage_opamp_dummy_magic_14_0.Vb3.t7 GNDA.t253 GNDA.t255 GNDA.t254 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X504 VOUT+.t114 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t43 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X505 bgr_0.Vin-.t4 bgr_0.START_UP.t6 bgr_0.V_TOP.t0 VDDA.t32 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X506 GNDA.t252 GNDA.t250 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t9 GNDA.t251 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X507 two_stage_opamp_dummy_magic_14_0.VD1.t3 VIN-.t7 two_stage_opamp_dummy_magic_14_0.V_source.t39 GNDA.t24 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X508 bgr_0.V_TOP.t2 bgr_0.START_UP.t7 bgr_0.Vin-.t5 VDDA.t153 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X509 VOUT-.t108 two_stage_opamp_dummy_magic_14_0.cap_res_X.t49 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X510 VOUT+.t115 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t42 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X511 VOUT+.t116 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t41 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X512 two_stage_opamp_dummy_magic_14_0.V_source.t18 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t24 GNDA.t158 GNDA.t157 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X513 VDDA.t403 bgr_0.1st_Vout_2.t27 bgr_0.PFET_GATE_10uA.t2 VDDA.t402 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X514 bgr_0.V_mir1.t8 bgr_0.V_mir1.t7 VDDA.t384 VDDA.t383 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X515 VOUT-.t109 two_stage_opamp_dummy_magic_14_0.cap_res_X.t48 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X516 VOUT-.t110 two_stage_opamp_dummy_magic_14_0.cap_res_X.t47 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X517 two_stage_opamp_dummy_magic_14_0.V_source.t1 two_stage_opamp_dummy_magic_14_0.err_amp_out.t4 GNDA.t147 GNDA.t146 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X518 GNDA.t59 two_stage_opamp_dummy_magic_14_0.X.t44 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.t4 VDDA.t72 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X519 VOUT-.t111 two_stage_opamp_dummy_magic_14_0.cap_res_X.t46 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X520 GNDA.t209 GNDA.t249 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t4 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X521 bgr_0.START_UP.t5 bgr_0.START_UP.t4 bgr_0.START_UP_NFET1.t0 GNDA.t139 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X522 bgr_0.V_p_2.t0 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.t10 bgr_0.V_mir2.t15 GNDA.t118 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X523 two_stage_opamp_dummy_magic_14_0.VD2.t2 VIN+.t7 two_stage_opamp_dummy_magic_14_0.V_source.t11 GNDA.t46 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X524 VDDA.t116 two_stage_opamp_dummy_magic_14_0.Y.t43 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.t3 GNDA.t76 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X525 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.t3 two_stage_opamp_dummy_magic_14_0.Y.t44 GNDA.t52 VDDA.t69 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X526 VDDA.t195 two_stage_opamp_dummy_magic_14_0.Y.t45 VOUT+.t12 VDDA.t194 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X527 VOUT+.t117 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t40 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X528 VOUT+.t118 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t39 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X529 VOUT-.t112 two_stage_opamp_dummy_magic_14_0.cap_res_X.t45 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X530 bgr_0.1st_Vout_2.t28 bgr_0.cap_res2.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X531 VOUT-.t113 two_stage_opamp_dummy_magic_14_0.cap_res_X.t44 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X532 VOUT+.t119 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t38 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X533 VDDA.t378 bgr_0.PFET_GATE_10uA.t24 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t11 VDDA.t377 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X534 VDDA.t34 bgr_0.V_mir2.t21 bgr_0.1st_Vout_2.t0 VDDA.t33 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X535 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t3 bgr_0.PFET_GATE_10uA.t25 VDDA.t89 VDDA.t88 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X536 VOUT-.t114 two_stage_opamp_dummy_magic_14_0.cap_res_X.t43 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X537 bgr_0.V_p_1.t0 bgr_0.Vin-.t12 bgr_0.V_mir1.t2 GNDA.t129 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.2
X538 two_stage_opamp_dummy_magic_14_0.VD4.t26 two_stage_opamp_dummy_magic_14_0.Vb3.t26 VDDA.t225 VDDA.t224 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X539 GNDA.t209 GNDA.t245 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t3 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X540 bgr_0.1st_Vout_2.t29 bgr_0.cap_res2.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X541 VOUT-.t115 two_stage_opamp_dummy_magic_14_0.cap_res_X.t42 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X542 VOUT-.t116 two_stage_opamp_dummy_magic_14_0.cap_res_X.t41 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X543 VOUT+.t120 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t37 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X544 VOUT+.t13 GNDA.t246 GNDA.t248 GNDA.t247 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=2.8 ps=14.8 w=7 l=0.6
X545 two_stage_opamp_dummy_magic_14_0.err_amp_mir.t3 VDDA.t284 VDDA.t286 VDDA.t285 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=1 ps=5.8 w=2.5 l=0.15
X546 VOUT-.t117 two_stage_opamp_dummy_magic_14_0.cap_res_X.t40 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X547 VOUT+.t121 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t36 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X548 bgr_0.1st_Vout_1.t30 bgr_0.cap_res1.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X549 GNDA.t218 GNDA.t244 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t2 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X550 two_stage_opamp_dummy_magic_14_0.X.t20 GNDA.t242 GNDA.t243 GNDA.t230 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X551 VDDA.t74 two_stage_opamp_dummy_magic_14_0.X.t45 VOUT-.t7 VDDA.t73 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X552 two_stage_opamp_dummy_magic_14_0.X.t18 two_stage_opamp_dummy_magic_14_0.Vb1.t21 two_stage_opamp_dummy_magic_14_0.VD1.t12 GNDA.t68 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X553 GNDA.t103 a_6930_22664.t1 GNDA.t65 sky130_fd_pr__res_xhigh_po_0p35 l=3.83
X554 VOUT+.t122 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t35 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X555 GNDA.t209 GNDA.t241 bgr_0.Vin-.t7 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X556 VOUT+.t123 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t34 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X557 bgr_0.1st_Vout_2.t30 bgr_0.cap_res2.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X558 VDDA.t223 two_stage_opamp_dummy_magic_14_0.Vb3.t27 two_stage_opamp_dummy_magic_14_0.VD3.t21 VDDA.t222 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X559 GNDA.t82 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t25 two_stage_opamp_dummy_magic_14_0.V_source.t17 GNDA.t81 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X560 GNDA.t240 GNDA.t237 GNDA.t239 GNDA.t238 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=0 ps=0 w=2.5 l=0.15
X561 two_stage_opamp_dummy_magic_14_0.Y.t24 GNDA.t235 GNDA.t236 GNDA.t222 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X562 VOUT+.t3 two_stage_opamp_dummy_magic_14_0.V_b_2nd_stage.t7 GNDA.t28 GNDA.t27 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X563 VOUT+.t124 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t33 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X564 GNDA.t173 bgr_0.NFET_GATE_10uA.t18 two_stage_opamp_dummy_magic_14_0.V_err_gate.t1 GNDA.t172 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X565 bgr_0.Vin-.t1 bgr_0.V_TOP.t39 VDDA.t1 VDDA.t0 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X566 a_14290_5524.t1 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.t16 GNDA.t300 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X567 a_12530_23988.t0 a_12410_22380.t1 GNDA.t66 sky130_fd_pr__res_xhigh_po_0p35 l=6
X568 two_stage_opamp_dummy_magic_14_0.Vb3.t6 bgr_0.NFET_GATE_10uA.t19 GNDA.t171 GNDA.t170 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X569 bgr_0.1st_Vout_2.t31 bgr_0.cap_res2.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X570 two_stage_opamp_dummy_magic_14_0.V_p_mir.t0 VIN+.t8 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t4 GNDA.t70 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X571 two_stage_opamp_dummy_magic_14_0.VD1.t2 VIN-.t8 two_stage_opamp_dummy_magic_14_0.V_source.t6 GNDA.t25 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X572 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.t2 two_stage_opamp_dummy_magic_14_0.X.t46 VDDA.t62 GNDA.t48 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X573 GNDA.t234 GNDA.t232 VDDA.t264 GNDA.t233 sky130_fd_pr__nfet_01v8 ad=1.2 pd=6.8 as=0.6 ps=3.4 w=3 l=0.15
X574 VOUT-.t118 two_stage_opamp_dummy_magic_14_0.cap_res_X.t39 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X575 VDDA.t380 bgr_0.V_mir2.t2 bgr_0.V_mir2.t3 VDDA.t379 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X576 two_stage_opamp_dummy_magic_14_0.V_source.t16 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t26 GNDA.t144 GNDA.t143 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X577 VOUT+.t125 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t32 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X578 bgr_0.1st_Vout_1.t31 bgr_0.cap_res1.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X579 bgr_0.1st_Vout_2.t32 bgr_0.cap_res2.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X580 two_stage_opamp_dummy_magic_14_0.V_source.t5 two_stage_opamp_dummy_magic_14_0.Vb1.t1 two_stage_opamp_dummy_magic_14_0.Vb1.t2 GNDA.t20 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=2.9
X581 bgr_0.V_p_1.t10 VDDA.t416 GNDA.t152 GNDA.t151 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=1.01 ps=6.15 w=2.5 l=5
X582 GNDA.t49 two_stage_opamp_dummy_magic_14_0.X.t47 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.t3 VDDA.t63 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X583 VDDA.t386 two_stage_opamp_dummy_magic_14_0.Y.t46 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.t2 GNDA.t298 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X584 VDDA.t283 VDDA.t281 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.t15 VDDA.t282 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X585 two_stage_opamp_dummy_magic_14_0.VD2.t21 VIN+.t9 two_stage_opamp_dummy_magic_14_0.V_source.t38 GNDA.t149 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X586 VOUT+.t126 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t31 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X587 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.t11 bgr_0.PFET_GATE_10uA.t26 VDDA.t152 VDDA.t151 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X588 VOUT-.t119 two_stage_opamp_dummy_magic_14_0.cap_res_X.t38 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X589 VOUT-.t120 two_stage_opamp_dummy_magic_14_0.cap_res_X.t37 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X590 a_13180_23838.t1 a_13060_22630.t1 GNDA.t150 sky130_fd_pr__res_xhigh_po_0p35 l=4
X591 VOUT+.t127 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t30 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X592 VOUT+.t128 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t29 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X593 VOUT+.t129 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t28 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X594 VDDA.t393 two_stage_opamp_dummy_magic_14_0.Y.t47 VOUT+.t17 VDDA.t392 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X595 VDDA.t280 VDDA.t278 VOUT+.t15 VDDA.t279 sky130_fd_pr__pfet_01v8 ad=2.4 pd=12.8 as=1.2 ps=6.4 w=6 l=0.15
X596 bgr_0.V_p_1.t6 bgr_0.Vin+.t9 bgr_0.1st_Vout_1.t8 GNDA.t12 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X597 VDDA.t179 bgr_0.V_mir1.t22 bgr_0.1st_Vout_1.t0 VDDA.t178 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X598 bgr_0.V_TOP.t40 VDDA.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X599 two_stage_opamp_dummy_magic_14_0.Vb2_2.t1 two_stage_opamp_dummy_magic_14_0.Vb2.t0 two_stage_opamp_dummy_magic_14_0.Vb2.t1 two_stage_opamp_dummy_magic_14_0.Vb2_2.t0 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X600 VOUT-.t121 two_stage_opamp_dummy_magic_14_0.cap_res_X.t36 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X601 VOUT-.t122 two_stage_opamp_dummy_magic_14_0.cap_res_X.t35 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X602 VOUT-.t123 two_stage_opamp_dummy_magic_14_0.cap_res_X.t34 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X603 VOUT-.t124 two_stage_opamp_dummy_magic_14_0.cap_res_X.t33 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X604 VOUT+.t130 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t27 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X605 VOUT+.t131 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t26 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X606 VDDA.t60 two_stage_opamp_dummy_magic_14_0.X.t48 VOUT-.t4 VDDA.t59 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X607 two_stage_opamp_dummy_magic_14_0.X.t21 two_stage_opamp_dummy_magic_14_0.Vb1.t22 two_stage_opamp_dummy_magic_14_0.VD1.t11 GNDA.t294 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X608 bgr_0.V_TOP.t41 VDDA.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X609 a_14170_5524.t0 two_stage_opamp_dummy_magic_14_0.V_tot.t0 GNDA.t31 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X610 bgr_0.V_p_1.t5 bgr_0.Vin+.t10 bgr_0.1st_Vout_1.t10 GNDA.t125 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X611 VDDA.t277 VDDA.t275 bgr_0.V_TOP.t6 VDDA.t276 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.2
X612 VOUT-.t125 two_stage_opamp_dummy_magic_14_0.cap_res_X.t32 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X613 two_stage_opamp_dummy_magic_14_0.Vb2.t3 bgr_0.NFET_GATE_10uA.t20 GNDA.t169 GNDA.t168 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X614 GNDA.t167 bgr_0.NFET_GATE_10uA.t21 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.t10 GNDA.t166 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X615 GNDA.t26 two_stage_opamp_dummy_magic_14_0.Y.t48 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.t2 VDDA.t35 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X616 VOUT-.t126 two_stage_opamp_dummy_magic_14_0.cap_res_X.t31 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X617 VOUT-.t127 two_stage_opamp_dummy_magic_14_0.cap_res_X.t30 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X618 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.t12 bgr_0.NFET_GATE_10uA.t22 GNDA.t165 GNDA.t164 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X619 bgr_0.V_TOP.t42 VDDA.t50 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X620 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.t5 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.t2 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.t4 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.t3 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0 ps=0 w=3.5 l=0.2
X621 bgr_0.V_TOP.t43 VDDA.t51 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X622 GNDA.t156 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t27 two_stage_opamp_dummy_magic_14_0.V_source.t15 GNDA.t155 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X623 two_stage_opamp_dummy_magic_14_0.Y.t20 two_stage_opamp_dummy_magic_14_0.Vb1.t23 two_stage_opamp_dummy_magic_14_0.VD2.t4 GNDA.t104 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X624 VOUT-.t128 two_stage_opamp_dummy_magic_14_0.cap_res_X.t29 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X625 VOUT-.t129 two_stage_opamp_dummy_magic_14_0.cap_res_X.t28 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X626 VDDA.t382 bgr_0.V_mir2.t22 bgr_0.1st_Vout_2.t8 VDDA.t381 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X627 two_stage_opamp_dummy_magic_14_0.VD4.t3 two_stage_opamp_dummy_magic_14_0.Vb2.t29 two_stage_opamp_dummy_magic_14_0.Y.t4 two_stage_opamp_dummy_magic_14_0.VD4.t2 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X628 VOUT-.t130 two_stage_opamp_dummy_magic_14_0.cap_res_X.t27 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X629 VDDA.t65 bgr_0.1st_Vout_1.t32 bgr_0.V_TOP.t1 VDDA.t64 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X630 VOUT+.t132 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t25 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X631 VOUT-.t131 two_stage_opamp_dummy_magic_14_0.cap_res_X.t26 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X632 VOUT-.t132 two_stage_opamp_dummy_magic_14_0.cap_res_X.t25 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X633 two_stage_opamp_dummy_magic_14_0.VD1.t21 GNDA.t229 GNDA.t231 GNDA.t230 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X634 two_stage_opamp_dummy_magic_14_0.VD1.t1 VIN-.t9 two_stage_opamp_dummy_magic_14_0.V_source.t7 GNDA.t68 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X635 VOUT+.t133 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t24 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X636 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.t1 two_stage_opamp_dummy_magic_14_0.X.t49 VDDA.t61 GNDA.t47 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X637 two_stage_opamp_dummy_magic_14_0.V_source.t14 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t28 GNDA.t43 GNDA.t42 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X638 VOUT+.t134 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t23 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X639 GNDA.t88 two_stage_opamp_dummy_magic_14_0.X.t50 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.t2 VDDA.t124 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X640 bgr_0.V_TOP.t44 VDDA.t52 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X641 VDDA.t263 GNDA.t226 GNDA.t228 GNDA.t227 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=1.2 ps=6.8 w=3 l=0.15
X642 GNDA.t225 GNDA.t224 two_stage_opamp_dummy_magic_14_0.X.t19 GNDA.t211 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X643 two_stage_opamp_dummy_magic_14_0.VD2.t14 GNDA.t221 GNDA.t223 GNDA.t222 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X644 two_stage_opamp_dummy_magic_14_0.VD3.t30 VDDA.t272 VDDA.t274 VDDA.t273 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X645 two_stage_opamp_dummy_magic_14_0.V_b_2nd_stage.t0 a_5980_2720.t1 GNDA.t91 sky130_fd_pr__res_xhigh_po_0p35 l=2.63
X646 VOUT-.t133 two_stage_opamp_dummy_magic_14_0.cap_res_X.t24 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X647 VOUT-.t5 two_stage_opamp_dummy_magic_14_0.V_b_2nd_stage.t8 GNDA.t56 GNDA.t55 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X648 two_stage_opamp_dummy_magic_14_0.VD3.t1 two_stage_opamp_dummy_magic_14_0.Vb2.t30 two_stage_opamp_dummy_magic_14_0.X.t0 two_stage_opamp_dummy_magic_14_0.VD3.t0 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X649 bgr_0.V_TOP.t45 VDDA.t92 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X650 bgr_0.V_mir2.t1 bgr_0.V_mir2.t0 VDDA.t202 VDDA.t201 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X651 VDDA.t401 bgr_0.V_mir1.t5 bgr_0.V_mir1.t6 VDDA.t400 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X652 VDDA.t68 two_stage_opamp_dummy_magic_14_0.Y.t49 VOUT+.t7 VDDA.t67 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X653 VOUT-.t134 two_stage_opamp_dummy_magic_14_0.cap_res_X.t23 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X654 GNDA.t220 GNDA.t219 two_stage_opamp_dummy_magic_14_0.Y.t23 GNDA.t203 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X655 VOUT-.t135 two_stage_opamp_dummy_magic_14_0.cap_res_X.t22 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X656 VOUT-.t136 two_stage_opamp_dummy_magic_14_0.cap_res_X.t21 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X657 bgr_0.V_mir2.t14 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.t11 bgr_0.V_p_2.t3 GNDA.t1 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.2
X658 VOUT+.t135 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t22 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X659 VOUT+.t136 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t21 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X660 bgr_0.PFET_GATE_10uA.t7 VDDA.t417 GNDA.t153 GNDA.t1 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=1 ps=5.8 w=2.5 l=5
X661 VOUT+.t137 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t20 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X662 bgr_0.1st_Vout_1.t33 bgr_0.cap_res1.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X663 VOUT-.t137 two_stage_opamp_dummy_magic_14_0.cap_res_X.t20 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X664 two_stage_opamp_dummy_magic_14_0.Vb1.t0 bgr_0.PFET_GATE_10uA.t27 VDDA.t31 VDDA.t30 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X665 VDDA.t94 bgr_0.V_TOP.t46 bgr_0.Vin-.t0 VDDA.t93 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X666 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.t1 two_stage_opamp_dummy_magic_14_0.Y.t50 VDDA.t193 GNDA.t133 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X667 VOUT+.t138 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X668 VOUT-.t6 two_stage_opamp_dummy_magic_14_0.V_b_2nd_stage.t9 GNDA.t58 GNDA.t57 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X669 VDDA.t126 two_stage_opamp_dummy_magic_14_0.X.t51 VOUT-.t9 VDDA.t125 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X670 VOUT-.t138 two_stage_opamp_dummy_magic_14_0.cap_res_X.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X671 bgr_0.PFET_GATE_10uA.t1 bgr_0.1st_Vout_2.t33 VDDA.t16 VDDA.t15 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X672 two_stage_opamp_dummy_magic_14_0.VD3.t20 two_stage_opamp_dummy_magic_14_0.Vb3.t28 VDDA.t221 VDDA.t220 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X673 VOUT+.t139 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X674 VDDA.t146 bgr_0.PFET_GATE_10uA.t28 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.t10 VDDA.t145 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X675 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.t14 VDDA.t269 VDDA.t271 VDDA.t270 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X676 VOUT-.t139 two_stage_opamp_dummy_magic_14_0.cap_res_X.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X677 GNDA.t132 two_stage_opamp_dummy_magic_14_0.Y.t51 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.t1 VDDA.t192 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X678 VOUT-.t140 two_stage_opamp_dummy_magic_14_0.cap_res_X.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X679 VOUT+.t140 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X680 GNDA.t80 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t29 two_stage_opamp_dummy_magic_14_0.V_source.t13 GNDA.t79 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X681 VDDA.t177 bgr_0.1st_Vout_2.t34 bgr_0.PFET_GATE_10uA.t0 VDDA.t176 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X682 VOUT+.t141 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X683 VOUT+.t142 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X684 VOUT+.t143 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X685 VOUT+.t144 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X686 bgr_0.1st_Vout_1.t34 bgr_0.cap_res1.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X687 bgr_0.1st_Vout_2.t35 bgr_0.cap_res2.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X688 VOUT-.t141 two_stage_opamp_dummy_magic_14_0.cap_res_X.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X689 bgr_0.V_mir2.t13 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.t12 bgr_0.V_p_2.t2 GNDA.t15 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X690 two_stage_opamp_dummy_magic_14_0.VD1.t0 VIN-.t10 two_stage_opamp_dummy_magic_14_0.V_source.t37 GNDA.t294 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X691 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.t0 two_stage_opamp_dummy_magic_14_0.X.t52 VDDA.t127 GNDA.t89 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X692 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.t11 bgr_0.NFET_GATE_10uA.t23 GNDA.t163 GNDA.t162 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X693 GNDA.t90 two_stage_opamp_dummy_magic_14_0.X.t53 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.t1 VDDA.t128 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X694 VOUT-.t142 two_stage_opamp_dummy_magic_14_0.cap_res_X.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X695 VOUT-.t143 two_stage_opamp_dummy_magic_14_0.cap_res_X.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X696 two_stage_opamp_dummy_magic_14_0.V_source.t12 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t30 GNDA.t111 GNDA.t110 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X697 GNDA.t209 GNDA.t213 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t1 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X698 VOUT-.t144 two_stage_opamp_dummy_magic_14_0.cap_res_X.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X699 GNDA.t29 two_stage_opamp_dummy_magic_14_0.X.t54 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.t0 VDDA.t38 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X700 VOUT+.t145 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X701 bgr_0.1st_Vout_1.t35 bgr_0.cap_res1.t0 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X702 two_stage_opamp_dummy_magic_14_0.VD1.t10 two_stage_opamp_dummy_magic_14_0.Vb1.t24 two_stage_opamp_dummy_magic_14_0.X.t11 GNDA.t3 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X703 VOUT-.t145 two_stage_opamp_dummy_magic_14_0.cap_res_X.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X704 VDDA.t175 bgr_0.1st_Vout_1.t36 bgr_0.V_TOP.t4 VDDA.t174 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X705 two_stage_opamp_dummy_magic_14_0.VD2.t19 VIN+.t10 two_stage_opamp_dummy_magic_14_0.V_source.t35 GNDA.t104 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X706 GNDA.t154 VDDA.t418 bgr_0.V_TOP.t5 GNDA.t129 sky130_fd_pr__nfet_01v8 ad=1.01 pd=6.15 as=1 ps=5.8 w=2.5 l=5
X707 bgr_0.V_TOP.t47 VDDA.t95 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X708 VOUT-.t146 two_stage_opamp_dummy_magic_14_0.cap_res_X.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X709 VDDA.t82 bgr_0.V_TOP.t48 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.t0 VDDA.t81 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X710 two_stage_opamp_dummy_magic_14_0.V_err_gate.t5 two_stage_opamp_dummy_magic_14_0.V_tot.t5 two_stage_opamp_dummy_magic_14_0.V_err_mir_p.t3 VDDA.t375 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X711 VOUT+.t146 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X712 VOUT+.t147 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X713 VDDA.t115 two_stage_opamp_dummy_magic_14_0.Y.t52 VOUT+.t8 VDDA.t114 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X714 VOUT+.t148 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X715 VOUT-.t147 two_stage_opamp_dummy_magic_14_0.cap_res_X.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X716 two_stage_opamp_dummy_magic_14_0.Vb2_2.t6 two_stage_opamp_dummy_magic_14_0.Vb2_2.t4 two_stage_opamp_dummy_magic_14_0.Vb2_2.t6 two_stage_opamp_dummy_magic_14_0.Vb2_2.t5 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0 ps=0 w=3.5 l=0.2
X717 two_stage_opamp_dummy_magic_14_0.Y.t0 two_stage_opamp_dummy_magic_14_0.VD4.t20 two_stage_opamp_dummy_magic_14_0.VD4.t22 two_stage_opamp_dummy_magic_14_0.VD4.t21 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X718 two_stage_opamp_dummy_magic_14_0.VD2.t3 two_stage_opamp_dummy_magic_14_0.Vb1.t25 two_stage_opamp_dummy_magic_14_0.Y.t13 GNDA.t93 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X719 VOUT-.t148 two_stage_opamp_dummy_magic_14_0.cap_res_X.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X720 bgr_0.V_mir2.t12 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.t13 bgr_0.V_p_2.t1 GNDA.t309 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X721 VOUT+.t149 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X722 VDDA.t217 bgr_0.PFET_GATE_10uA.t29 bgr_0.V_CUR_REF_REG.t1 VDDA.t216 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X723 VOUT+.t150 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X724 VOUT-.t149 two_stage_opamp_dummy_magic_14_0.cap_res_X.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X725 VOUT+.t151 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X726 GNDA.t212 GNDA.t210 two_stage_opamp_dummy_magic_14_0.VD1.t20 GNDA.t211 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X727 VOUT-.t150 two_stage_opamp_dummy_magic_14_0.cap_res_X.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X728 VOUT-.t151 two_stage_opamp_dummy_magic_14_0.cap_res_X.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X729 VOUT+.t152 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X730 VOUT-.t152 two_stage_opamp_dummy_magic_14_0.cap_res_X.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X731 VOUT-.t153 two_stage_opamp_dummy_magic_14_0.cap_res_X.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X732 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.t0 two_stage_opamp_dummy_magic_14_0.Y.t53 VDDA.t66 GNDA.t51 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X733 GNDA.t207 GNDA.t205 VDDA.t262 GNDA.t206 sky130_fd_pr__nfet_01v8 ad=1.2 pd=6.8 as=0.6 ps=3.4 w=3 l=0.15
X734 GNDA.t204 GNDA.t202 two_stage_opamp_dummy_magic_14_0.VD2.t13 GNDA.t203 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X735 bgr_0.V_TOP.t49 VDDA.t83 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X736 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.t5 VDDA.t266 VDDA.t268 VDDA.t267 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=1.2 ps=6.8 w=3 l=0.5
X737 two_stage_opamp_dummy_magic_14_0.Vb3.t0 two_stage_opamp_dummy_magic_14_0.Vb2.t31 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.t1 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.t0 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X738 two_stage_opamp_dummy_magic_14_0.X.t5 two_stage_opamp_dummy_magic_14_0.VD3.t6 two_stage_opamp_dummy_magic_14_0.VD3.t8 two_stage_opamp_dummy_magic_14_0.VD3.t7 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X739 VOUT+.t153 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X740 VOUT-.t154 two_stage_opamp_dummy_magic_14_0.cap_res_X.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X741 VOUT+.t154 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X742 VOUT-.t155 two_stage_opamp_dummy_magic_14_0.cap_res_X.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X743 bgr_0.1st_Vout_2.t36 bgr_0.cap_res2.t0 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X744 GNDA.t75 two_stage_opamp_dummy_magic_14_0.Y.t54 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.t0 VDDA.t113 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X745 VDDA.t414 bgr_0.V_mir1.t3 bgr_0.V_mir1.t4 VDDA.t413 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X746 VOUT+.t155 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X747 two_stage_opamp_dummy_magic_14_0.Y.t2 two_stage_opamp_dummy_magic_14_0.Vb2.t32 two_stage_opamp_dummy_magic_14_0.VD4.t1 two_stage_opamp_dummy_magic_14_0.VD4.t0 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X748 VOUT+.t156 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X749 GNDA.t5 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t31 two_stage_opamp_dummy_magic_14_0.V_p_mir.t2 GNDA.t4 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X750 a_6810_23838.t1 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.t4 GNDA.t65 sky130_fd_pr__res_xhigh_po_0p35 l=3.83
X751 VOUT-.t156 two_stage_opamp_dummy_magic_14_0.cap_res_X.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
R0 bgr_0.NFET_GATE_10uA.n19 bgr_0.NFET_GATE_10uA.t3 384.967
R1 bgr_0.NFET_GATE_10uA.n10 bgr_0.NFET_GATE_10uA.t10 369.534
R2 bgr_0.NFET_GATE_10uA.n9 bgr_0.NFET_GATE_10uA.t22 369.534
R3 bgr_0.NFET_GATE_10uA.n7 bgr_0.NFET_GATE_10uA.t7 369.534
R4 bgr_0.NFET_GATE_10uA.n4 bgr_0.NFET_GATE_10uA.t16 369.534
R5 bgr_0.NFET_GATE_10uA.n1 bgr_0.NFET_GATE_10uA.t12 369.534
R6 bgr_0.NFET_GATE_10uA.t3 bgr_0.NFET_GATE_10uA.n18 369.534
R7 bgr_0.NFET_GATE_10uA bgr_0.NFET_GATE_10uA.n20 366.553
R8 bgr_0.NFET_GATE_10uA.n12 bgr_0.NFET_GATE_10uA.t9 192.8
R9 bgr_0.NFET_GATE_10uA.n11 bgr_0.NFET_GATE_10uA.t17 192.8
R10 bgr_0.NFET_GATE_10uA.n10 bgr_0.NFET_GATE_10uA.t23 192.8
R11 bgr_0.NFET_GATE_10uA.n9 bgr_0.NFET_GATE_10uA.t11 192.8
R12 bgr_0.NFET_GATE_10uA.n7 bgr_0.NFET_GATE_10uA.t20 192.8
R13 bgr_0.NFET_GATE_10uA.n4 bgr_0.NFET_GATE_10uA.t21 192.8
R14 bgr_0.NFET_GATE_10uA.n5 bgr_0.NFET_GATE_10uA.t8 192.8
R15 bgr_0.NFET_GATE_10uA.n6 bgr_0.NFET_GATE_10uA.t15 192.8
R16 bgr_0.NFET_GATE_10uA.n3 bgr_0.NFET_GATE_10uA.t19 192.8
R17 bgr_0.NFET_GATE_10uA.n2 bgr_0.NFET_GATE_10uA.t5 192.8
R18 bgr_0.NFET_GATE_10uA.n1 bgr_0.NFET_GATE_10uA.t13 192.8
R19 bgr_0.NFET_GATE_10uA.n18 bgr_0.NFET_GATE_10uA.t18 192.8
R20 bgr_0.NFET_GATE_10uA.n17 bgr_0.NFET_GATE_10uA.t6 192.8
R21 bgr_0.NFET_GATE_10uA.n16 bgr_0.NFET_GATE_10uA.t14 192.8
R22 bgr_0.NFET_GATE_10uA.n12 bgr_0.NFET_GATE_10uA.n11 176.733
R23 bgr_0.NFET_GATE_10uA.n11 bgr_0.NFET_GATE_10uA.n10 176.733
R24 bgr_0.NFET_GATE_10uA.n5 bgr_0.NFET_GATE_10uA.n4 176.733
R25 bgr_0.NFET_GATE_10uA.n6 bgr_0.NFET_GATE_10uA.n5 176.733
R26 bgr_0.NFET_GATE_10uA.n3 bgr_0.NFET_GATE_10uA.n2 176.733
R27 bgr_0.NFET_GATE_10uA.n2 bgr_0.NFET_GATE_10uA.n1 176.733
R28 bgr_0.NFET_GATE_10uA.n18 bgr_0.NFET_GATE_10uA.n17 176.733
R29 bgr_0.NFET_GATE_10uA.n17 bgr_0.NFET_GATE_10uA.n16 176.733
R30 bgr_0.NFET_GATE_10uA.n14 bgr_0.NFET_GATE_10uA.n13 169.852
R31 bgr_0.NFET_GATE_10uA.n14 bgr_0.NFET_GATE_10uA.n8 169.852
R32 bgr_0.NFET_GATE_10uA.n15 bgr_0.NFET_GATE_10uA.n14 166.133
R33 bgr_0.NFET_GATE_10uA.n19 bgr_0.NFET_GATE_10uA.n0 126.877
R34 bgr_0.NFET_GATE_10uA.n13 bgr_0.NFET_GATE_10uA.n12 56.2338
R35 bgr_0.NFET_GATE_10uA.n13 bgr_0.NFET_GATE_10uA.n9 56.2338
R36 bgr_0.NFET_GATE_10uA.n8 bgr_0.NFET_GATE_10uA.n7 56.2338
R37 bgr_0.NFET_GATE_10uA.n8 bgr_0.NFET_GATE_10uA.n6 56.2338
R38 bgr_0.NFET_GATE_10uA.n15 bgr_0.NFET_GATE_10uA.n3 56.2338
R39 bgr_0.NFET_GATE_10uA.n16 bgr_0.NFET_GATE_10uA.n15 56.2338
R40 bgr_0.NFET_GATE_10uA.n20 bgr_0.NFET_GATE_10uA.t0 39.4005
R41 bgr_0.NFET_GATE_10uA.n20 bgr_0.NFET_GATE_10uA.t2 39.4005
R42 bgr_0.NFET_GATE_10uA bgr_0.NFET_GATE_10uA.n19 30.6442
R43 bgr_0.NFET_GATE_10uA.n0 bgr_0.NFET_GATE_10uA.t1 24.0005
R44 bgr_0.NFET_GATE_10uA.n0 bgr_0.NFET_GATE_10uA.t4 24.0005
R45 two_stage_opamp_dummy_magic_14_0.Vb3.n25 two_stage_opamp_dummy_magic_14_0.Vb3.t14 650.511
R46 two_stage_opamp_dummy_magic_14_0.Vb3.n19 two_stage_opamp_dummy_magic_14_0.Vb3.t13 611.739
R47 two_stage_opamp_dummy_magic_14_0.Vb3.n15 two_stage_opamp_dummy_magic_14_0.Vb3.t22 611.739
R48 two_stage_opamp_dummy_magic_14_0.Vb3.n10 two_stage_opamp_dummy_magic_14_0.Vb3.t8 611.739
R49 two_stage_opamp_dummy_magic_14_0.Vb3.n6 two_stage_opamp_dummy_magic_14_0.Vb3.t16 611.739
R50 two_stage_opamp_dummy_magic_14_0.Vb3.n19 two_stage_opamp_dummy_magic_14_0.Vb3.t19 421.75
R51 two_stage_opamp_dummy_magic_14_0.Vb3.n20 two_stage_opamp_dummy_magic_14_0.Vb3.t23 421.75
R52 two_stage_opamp_dummy_magic_14_0.Vb3.n21 two_stage_opamp_dummy_magic_14_0.Vb3.t26 421.75
R53 two_stage_opamp_dummy_magic_14_0.Vb3.n22 two_stage_opamp_dummy_magic_14_0.Vb3.t25 421.75
R54 two_stage_opamp_dummy_magic_14_0.Vb3.n15 two_stage_opamp_dummy_magic_14_0.Vb3.t24 421.75
R55 two_stage_opamp_dummy_magic_14_0.Vb3.n16 two_stage_opamp_dummy_magic_14_0.Vb3.t20 421.75
R56 two_stage_opamp_dummy_magic_14_0.Vb3.n17 two_stage_opamp_dummy_magic_14_0.Vb3.t15 421.75
R57 two_stage_opamp_dummy_magic_14_0.Vb3.n18 two_stage_opamp_dummy_magic_14_0.Vb3.t10 421.75
R58 two_stage_opamp_dummy_magic_14_0.Vb3.n10 two_stage_opamp_dummy_magic_14_0.Vb3.t11 421.75
R59 two_stage_opamp_dummy_magic_14_0.Vb3.n11 two_stage_opamp_dummy_magic_14_0.Vb3.t17 421.75
R60 two_stage_opamp_dummy_magic_14_0.Vb3.n12 two_stage_opamp_dummy_magic_14_0.Vb3.t21 421.75
R61 two_stage_opamp_dummy_magic_14_0.Vb3.n13 two_stage_opamp_dummy_magic_14_0.Vb3.t27 421.75
R62 two_stage_opamp_dummy_magic_14_0.Vb3.n6 two_stage_opamp_dummy_magic_14_0.Vb3.t18 421.75
R63 two_stage_opamp_dummy_magic_14_0.Vb3.n7 two_stage_opamp_dummy_magic_14_0.Vb3.t12 421.75
R64 two_stage_opamp_dummy_magic_14_0.Vb3.n8 two_stage_opamp_dummy_magic_14_0.Vb3.t9 421.75
R65 two_stage_opamp_dummy_magic_14_0.Vb3.n9 two_stage_opamp_dummy_magic_14_0.Vb3.t28 421.75
R66 two_stage_opamp_dummy_magic_14_0.Vb3.n24 two_stage_opamp_dummy_magic_14_0.Vb3.n23 176.185
R67 two_stage_opamp_dummy_magic_14_0.Vb3.n24 two_stage_opamp_dummy_magic_14_0.Vb3.n14 175.624
R68 two_stage_opamp_dummy_magic_14_0.Vb3.n20 two_stage_opamp_dummy_magic_14_0.Vb3.n19 167.094
R69 two_stage_opamp_dummy_magic_14_0.Vb3.n21 two_stage_opamp_dummy_magic_14_0.Vb3.n20 167.094
R70 two_stage_opamp_dummy_magic_14_0.Vb3.n22 two_stage_opamp_dummy_magic_14_0.Vb3.n21 167.094
R71 two_stage_opamp_dummy_magic_14_0.Vb3.n16 two_stage_opamp_dummy_magic_14_0.Vb3.n15 167.094
R72 two_stage_opamp_dummy_magic_14_0.Vb3.n17 two_stage_opamp_dummy_magic_14_0.Vb3.n16 167.094
R73 two_stage_opamp_dummy_magic_14_0.Vb3.n18 two_stage_opamp_dummy_magic_14_0.Vb3.n17 167.094
R74 two_stage_opamp_dummy_magic_14_0.Vb3.n11 two_stage_opamp_dummy_magic_14_0.Vb3.n10 167.094
R75 two_stage_opamp_dummy_magic_14_0.Vb3.n12 two_stage_opamp_dummy_magic_14_0.Vb3.n11 167.094
R76 two_stage_opamp_dummy_magic_14_0.Vb3.n13 two_stage_opamp_dummy_magic_14_0.Vb3.n12 167.094
R77 two_stage_opamp_dummy_magic_14_0.Vb3.n7 two_stage_opamp_dummy_magic_14_0.Vb3.n6 167.094
R78 two_stage_opamp_dummy_magic_14_0.Vb3.n8 two_stage_opamp_dummy_magic_14_0.Vb3.n7 167.094
R79 two_stage_opamp_dummy_magic_14_0.Vb3.n9 two_stage_opamp_dummy_magic_14_0.Vb3.n8 167.094
R80 two_stage_opamp_dummy_magic_14_0.Vb3.n26 two_stage_opamp_dummy_magic_14_0.Vb3.n5 161.631
R81 two_stage_opamp_dummy_magic_14_0.Vb3.n2 two_stage_opamp_dummy_magic_14_0.Vb3.n0 139.639
R82 two_stage_opamp_dummy_magic_14_0.Vb3.n2 two_stage_opamp_dummy_magic_14_0.Vb3.n1 139.638
R83 two_stage_opamp_dummy_magic_14_0.Vb3.n4 two_stage_opamp_dummy_magic_14_0.Vb3.n3 134.577
R84 two_stage_opamp_dummy_magic_14_0.Vb3.n23 two_stage_opamp_dummy_magic_14_0.Vb3.n22 49.8072
R85 two_stage_opamp_dummy_magic_14_0.Vb3.n23 two_stage_opamp_dummy_magic_14_0.Vb3.n18 49.8072
R86 two_stage_opamp_dummy_magic_14_0.Vb3.n14 two_stage_opamp_dummy_magic_14_0.Vb3.n13 49.8072
R87 two_stage_opamp_dummy_magic_14_0.Vb3.n14 two_stage_opamp_dummy_magic_14_0.Vb3.n9 49.8072
R88 bgr_0.VB3_CUR_BIAS two_stage_opamp_dummy_magic_14_0.Vb3.n26 48.0943
R89 bgr_0.VB3_CUR_BIAS two_stage_opamp_dummy_magic_14_0.Vb3.n4 41.063
R90 two_stage_opamp_dummy_magic_14_0.Vb3.n3 two_stage_opamp_dummy_magic_14_0.Vb3.t2 24.0005
R91 two_stage_opamp_dummy_magic_14_0.Vb3.n3 two_stage_opamp_dummy_magic_14_0.Vb3.t5 24.0005
R92 two_stage_opamp_dummy_magic_14_0.Vb3.n1 two_stage_opamp_dummy_magic_14_0.Vb3.t3 24.0005
R93 two_stage_opamp_dummy_magic_14_0.Vb3.n1 two_stage_opamp_dummy_magic_14_0.Vb3.t7 24.0005
R94 two_stage_opamp_dummy_magic_14_0.Vb3.n0 two_stage_opamp_dummy_magic_14_0.Vb3.t4 24.0005
R95 two_stage_opamp_dummy_magic_14_0.Vb3.n0 two_stage_opamp_dummy_magic_14_0.Vb3.t6 24.0005
R96 two_stage_opamp_dummy_magic_14_0.Vb3.n25 two_stage_opamp_dummy_magic_14_0.Vb3.n24 13.7349
R97 two_stage_opamp_dummy_magic_14_0.Vb3.n5 two_stage_opamp_dummy_magic_14_0.Vb3.t1 11.2576
R98 two_stage_opamp_dummy_magic_14_0.Vb3.n5 two_stage_opamp_dummy_magic_14_0.Vb3.t0 11.2576
R99 two_stage_opamp_dummy_magic_14_0.Vb3.n4 two_stage_opamp_dummy_magic_14_0.Vb3.n2 4.5005
R100 two_stage_opamp_dummy_magic_14_0.Vb3.n26 two_stage_opamp_dummy_magic_14_0.Vb3.n25 1.438
R101 GNDA.n82 GNDA.n37 22479.7
R102 GNDA.n784 GNDA.n783 15367.3
R103 GNDA.n80 GNDA.n36 13534.7
R104 GNDA.n368 GNDA.n35 13528.5
R105 GNDA.n367 GNDA.n366 13200
R106 GNDA.n782 GNDA.n781 12810.6
R107 GNDA.n785 GNDA.n784 11953.3
R108 GNDA.n785 GNDA.n371 11890.5
R109 GNDA.n369 GNDA.n33 11872.4
R110 GNDA.n366 GNDA.n37 11747.6
R111 GNDA.n366 GNDA.n365 11747.6
R112 GNDA.n368 GNDA.n367 11178.4
R113 GNDA.n779 GNDA.n371 9950.42
R114 GNDA.n784 GNDA.n781 9950.42
R115 GNDA.n369 GNDA.n368 9632.43
R116 GNDA.n780 GNDA.n779 9384.59
R117 GNDA.n781 GNDA.n780 9384.59
R118 GNDA.n2441 GNDA.n369 9001.83
R119 GNDA.n2442 GNDA.n33 8211.75
R120 GNDA.n81 GNDA.n37 7737.08
R121 GNDA.n370 GNDA.n34 7427.52
R122 GNDA.n36 GNDA.n35 4761.61
R123 GNDA.n2439 GNDA.n371 4448.89
R124 GNDA.n786 GNDA.n785 3974.19
R125 GNDA.n367 GNDA.n36 3961.87
R126 GNDA.n347 GNDA.n37 3482.21
R127 GNDA.n365 GNDA.n364 3482.21
R128 GNDA.t108 GNDA.n2441 3375.81
R129 GNDA.n780 GNDA.n34 3105.87
R130 GNDA.n2441 GNDA.n34 2321.1
R131 GNDA.n35 GNDA.n34 2315.79
R132 GNDA.t31 GNDA.n82 2006.86
R133 GNDA.n2441 GNDA.n2440 2001.83
R134 GNDA.n80 GNDA.n34 1779.93
R135 GNDA.n783 GNDA.n782 1460.18
R136 GNDA.t67 GNDA.n81 1440.97
R137 GNDA.n779 GNDA.n370 1440.71
R138 GNDA.n2440 GNDA.n370 1440.71
R139 GNDA.n1665 GNDA.n1664 1336.64
R140 GNDA.n2439 GNDA.t85 1258.74
R141 GNDA.n1690 GNDA.n1084 1214.72
R142 GNDA.n1696 GNDA.n1084 1214.72
R143 GNDA.n1697 GNDA.n1696 1214.72
R144 GNDA.n1697 GNDA.n1080 1214.72
R145 GNDA.n1703 GNDA.n1080 1214.72
R146 GNDA.n1705 GNDA.n1075 1214.72
R147 GNDA.n1711 GNDA.n1075 1214.72
R148 GNDA.n1712 GNDA.n1711 1214.72
R149 GNDA.n1712 GNDA.n1071 1214.72
R150 GNDA.n1718 GNDA.n1071 1214.72
R151 GNDA.n663 GNDA.n373 1212.88
R152 GNDA.n877 GNDA.n876 1185.07
R153 GNDA.n878 GNDA.n877 1185.07
R154 GNDA.n782 GNDA.n34 1167.58
R155 GNDA.n365 GNDA.n33 1158.42
R156 GNDA.n783 GNDA.t308 1012.83
R157 GNDA.n2440 GNDA.n2439 869.924
R158 GNDA.n1703 GNDA.t209 823.313
R159 GNDA.n198 GNDA.t256 762.534
R160 GNDA.n194 GNDA.t232 762.534
R161 GNDA.n2556 GNDA.t205 762.534
R162 GNDA.n14 GNDA.t226 762.534
R163 GNDA.n82 GNDA.t67 702.521
R164 GNDA.n2456 GNDA.n2455 692.506
R165 GNDA.n2552 GNDA.n2551 692.506
R166 GNDA.n208 GNDA.n207 692.506
R167 GNDA.n190 GNDA.n189 692.506
R168 GNDA.n2500 GNDA.n2499 692.506
R169 GNDA.n2540 GNDA.n2539 692.506
R170 GNDA.n117 GNDA.n114 692.506
R171 GNDA.n178 GNDA.n177 692.506
R172 GNDA.n2427 GNDA.n2426 686.717
R173 GNDA.n363 GNDA.n362 686.717
R174 GNDA.n346 GNDA.n345 686.717
R175 GNDA.n324 GNDA.n323 686.717
R176 GNDA.n335 GNDA.n334 686.717
R177 GNDA.n314 GNDA.n313 686.717
R178 GNDA.n276 GNDA.n275 686.717
R179 GNDA.n286 GNDA.n285 686.717
R180 GNDA.n295 GNDA.n56 686.717
R181 GNDA.n306 GNDA.n64 686.717
R182 GNDA.n213 GNDA.n212 686.717
R183 GNDA.n229 GNDA.n228 686.717
R184 GNDA.n266 GNDA.n265 686.717
R185 GNDA.n2430 GNDA.n373 686.717
R186 GNDA.n2430 GNDA.n372 686.717
R187 GNDA.n258 GNDA.n214 686.717
R188 GNDA.n232 GNDA.n231 686.717
R189 GNDA.n349 GNDA.n348 686.717
R190 GNDA.n355 GNDA.n38 686.717
R191 GNDA.n2418 GNDA.n384 686.717
R192 GNDA.n2225 GNDA.n2214 686.717
R193 GNDA.n233 GNDA.t237 682.201
R194 GNDA.n1300 GNDA.n1296 669.307
R195 GNDA.n257 GNDA.t285 650.067
R196 GNDA.n350 GNDA.t291 650.067
R197 GNDA.n354 GNDA.t265 650.067
R198 GNDA.n2324 GNDA.n2323 585.001
R199 GNDA.n2344 GNDA.n2343 585.001
R200 GNDA.n2338 GNDA.n419 585.001
R201 GNDA.n2376 GNDA.n2375 585.001
R202 GNDA.n2386 GNDA.n2385 585.001
R203 GNDA.n2437 GNDA.n2436 585.001
R204 GNDA.n2174 GNDA.n2173 585
R205 GNDA.n2172 GNDA.n2135 585
R206 GNDA.n2171 GNDA.n2170 585
R207 GNDA.n2169 GNDA.n2168 585
R208 GNDA.n2167 GNDA.n2166 585
R209 GNDA.n2165 GNDA.n2164 585
R210 GNDA.n2163 GNDA.n2162 585
R211 GNDA.n2161 GNDA.n2160 585
R212 GNDA.n2159 GNDA.n2158 585
R213 GNDA.n2157 GNDA.n2156 585
R214 GNDA.n475 GNDA.n474 585
R215 GNDA.n2176 GNDA.n475 585
R216 GNDA.n2179 GNDA.n2178 585
R217 GNDA.n2179 GNDA.n472 585
R218 GNDA.n1366 GNDA.n1365 585
R219 GNDA.n1364 GNDA.n1363 585
R220 GNDA.n1362 GNDA.n1361 585
R221 GNDA.n1360 GNDA.n1359 585
R222 GNDA.n1358 GNDA.n1357 585
R223 GNDA.n1356 GNDA.n1355 585
R224 GNDA.n1354 GNDA.n1353 585
R225 GNDA.n1352 GNDA.n1351 585
R226 GNDA.n1350 GNDA.n1349 585
R227 GNDA.n1348 GNDA.n1347 585
R228 GNDA.n1346 GNDA.n482 585
R229 GNDA.n2176 GNDA.n482 585
R230 GNDA.n1128 GNDA.n1127 585
R231 GNDA.n1128 GNDA.n1126 585
R232 GNDA.n2176 GNDA.n2130 585
R233 GNDA.n963 GNDA.n962 585
R234 GNDA.n961 GNDA.n960 585
R235 GNDA.n959 GNDA.n958 585
R236 GNDA.n957 GNDA.n956 585
R237 GNDA.n955 GNDA.n954 585
R238 GNDA.n953 GNDA.n952 585
R239 GNDA.n951 GNDA.n950 585
R240 GNDA.n949 GNDA.n948 585
R241 GNDA.n947 GNDA.n946 585
R242 GNDA.n945 GNDA.n944 585
R243 GNDA.n943 GNDA.n942 585
R244 GNDA.n1717 GNDA.n1070 585
R245 GNDA.n1718 GNDA.n1717 585
R246 GNDA.n1716 GNDA.n1715 585
R247 GNDA.n1716 GNDA.n1071 585
R248 GNDA.n1714 GNDA.n1072 585
R249 GNDA.n1712 GNDA.n1072 585
R250 GNDA.n1710 GNDA.n1073 585
R251 GNDA.n1711 GNDA.n1710 585
R252 GNDA.n1709 GNDA.n1708 585
R253 GNDA.n1709 GNDA.n1075 585
R254 GNDA.n1077 GNDA.n1076 585
R255 GNDA.n1705 GNDA.n1076 585
R256 GNDA.n1702 GNDA.n1079 585
R257 GNDA.n1703 GNDA.n1702 585
R258 GNDA.n1701 GNDA.n1700 585
R259 GNDA.n1701 GNDA.n1080 585
R260 GNDA.n1699 GNDA.n1081 585
R261 GNDA.n1697 GNDA.n1081 585
R262 GNDA.n1695 GNDA.n1082 585
R263 GNDA.n1696 GNDA.n1695 585
R264 GNDA.n1694 GNDA.n1693 585
R265 GNDA.n1694 GNDA.n1084 585
R266 GNDA.n1086 GNDA.n1085 585
R267 GNDA.n1690 GNDA.n1085 585
R268 GNDA.n1691 GNDA.n1086 585
R269 GNDA.n1691 GNDA.n1690 585
R270 GNDA.n1693 GNDA.n1692 585
R271 GNDA.n1692 GNDA.n1084 585
R272 GNDA.n1083 GNDA.n1082 585
R273 GNDA.n1696 GNDA.n1083 585
R274 GNDA.n1699 GNDA.n1698 585
R275 GNDA.n1698 GNDA.n1697 585
R276 GNDA.n1700 GNDA.n1078 585
R277 GNDA.n1080 GNDA.n1078 585
R278 GNDA.n1704 GNDA.n1079 585
R279 GNDA.n1704 GNDA.n1703 585
R280 GNDA.n1706 GNDA.n1077 585
R281 GNDA.n1706 GNDA.n1705 585
R282 GNDA.n1708 GNDA.n1707 585
R283 GNDA.n1707 GNDA.n1075 585
R284 GNDA.n1074 GNDA.n1073 585
R285 GNDA.n1711 GNDA.n1074 585
R286 GNDA.n1714 GNDA.n1713 585
R287 GNDA.n1713 GNDA.n1712 585
R288 GNDA.n1715 GNDA.n1069 585
R289 GNDA.n1071 GNDA.n1069 585
R290 GNDA.n1719 GNDA.n1070 585
R291 GNDA.n1719 GNDA.n1718 585
R292 GNDA.n2050 GNDA.n911 585
R293 GNDA.n2053 GNDA.n2052 585
R294 GNDA.n915 GNDA.n914 585
R295 GNDA.n1760 GNDA.n1759 585
R296 GNDA.n1761 GNDA.n1758 585
R297 GNDA.n1755 GNDA.n1754 585
R298 GNDA.n1767 GNDA.n1753 585
R299 GNDA.n1768 GNDA.n1752 585
R300 GNDA.n1769 GNDA.n1751 585
R301 GNDA.n1749 GNDA.n1748 585
R302 GNDA.n1774 GNDA.n1747 585
R303 GNDA.n1775 GNDA.n1746 585
R304 GNDA.n1776 GNDA.n1775 585
R305 GNDA.n1774 GNDA.n1773 585
R306 GNDA.n1772 GNDA.n1749 585
R307 GNDA.n1770 GNDA.n1769 585
R308 GNDA.n1768 GNDA.n1750 585
R309 GNDA.n1767 GNDA.n1766 585
R310 GNDA.n1764 GNDA.n1755 585
R311 GNDA.n1762 GNDA.n1761 585
R312 GNDA.n1760 GNDA.n1757 585
R313 GNDA.n914 GNDA.n913 585
R314 GNDA.n2054 GNDA.n2053 585
R315 GNDA.n2056 GNDA.n911 585
R316 GNDA.n2046 GNDA.n2045 585
R317 GNDA.n984 GNDA.n940 585
R318 GNDA.n983 GNDA.n982 585
R319 GNDA.n981 GNDA.n980 585
R320 GNDA.n979 GNDA.n978 585
R321 GNDA.n977 GNDA.n976 585
R322 GNDA.n975 GNDA.n974 585
R323 GNDA.n973 GNDA.n972 585
R324 GNDA.n971 GNDA.n970 585
R325 GNDA.n969 GNDA.n968 585
R326 GNDA.n967 GNDA.n966 585
R327 GNDA.n965 GNDA.n964 585
R328 GNDA.n1745 GNDA.n1744 585
R329 GNDA.n1743 GNDA.n1742 585
R330 GNDA.n1741 GNDA.n1740 585
R331 GNDA.n1739 GNDA.n1738 585
R332 GNDA.n1737 GNDA.n1736 585
R333 GNDA.n1735 GNDA.n1734 585
R334 GNDA.n1733 GNDA.n1732 585
R335 GNDA.n1731 GNDA.n1730 585
R336 GNDA.n1729 GNDA.n1728 585
R337 GNDA.n1727 GNDA.n1726 585
R338 GNDA.n1725 GNDA.n1724 585
R339 GNDA.n988 GNDA.n985 585
R340 GNDA.n1800 GNDA.n1799 585
R341 GNDA.n1798 GNDA.n1797 585
R342 GNDA.n1796 GNDA.n1795 585
R343 GNDA.n1794 GNDA.n1793 585
R344 GNDA.n1792 GNDA.n1791 585
R345 GNDA.n1790 GNDA.n1789 585
R346 GNDA.n1788 GNDA.n1787 585
R347 GNDA.n1786 GNDA.n1785 585
R348 GNDA.n1784 GNDA.n1783 585
R349 GNDA.n1782 GNDA.n1781 585
R350 GNDA.n1780 GNDA.n1779 585
R351 GNDA.n1778 GNDA.n1777 585
R352 GNDA.n1515 GNDA.n1514 585
R353 GNDA.n1512 GNDA.n1125 585
R354 GNDA.n1131 GNDA.n1130 585
R355 GNDA.n1507 GNDA.n1506 585
R356 GNDA.n1505 GNDA.n1504 585
R357 GNDA.n1431 GNDA.n1135 585
R358 GNDA.n1433 GNDA.n1432 585
R359 GNDA.n1438 GNDA.n1437 585
R360 GNDA.n1436 GNDA.n1429 585
R361 GNDA.n1444 GNDA.n1443 585
R362 GNDA.n1446 GNDA.n1445 585
R363 GNDA.n1427 GNDA.n1426 585
R364 GNDA.n1721 GNDA.n1066 585
R365 GNDA.n1067 GNDA.n1066 585
R366 GNDA.n1272 GNDA.n1271 585
R367 GNDA.n1269 GNDA.n1268 585
R368 GNDA.n1267 GNDA.n1266 585
R369 GNDA.n1183 GNDA.n1159 585
R370 GNDA.n1185 GNDA.n1184 585
R371 GNDA.n1189 GNDA.n1188 585
R372 GNDA.n1191 GNDA.n1190 585
R373 GNDA.n1198 GNDA.n1197 585
R374 GNDA.n1196 GNDA.n1181 585
R375 GNDA.n1204 GNDA.n1203 585
R376 GNDA.n1206 GNDA.n1205 585
R377 GNDA.n1179 GNDA.n1178 585
R378 GNDA.n1721 GNDA.n1720 585
R379 GNDA.n1720 GNDA.n1067 585
R380 GNDA.n1594 GNDA.n1068 585
R381 GNDA.n1595 GNDA.n1531 585
R382 GNDA.n1605 GNDA.n1604 585
R383 GNDA.n1607 GNDA.n1529 585
R384 GNDA.n1610 GNDA.n1609 585
R385 GNDA.n1611 GNDA.n1525 585
R386 GNDA.n1620 GNDA.n1619 585
R387 GNDA.n1622 GNDA.n1524 585
R388 GNDA.n1625 GNDA.n1624 585
R389 GNDA.n1626 GNDA.n1518 585
R390 GNDA.n1635 GNDA.n1634 585
R391 GNDA.n1637 GNDA.n1112 585
R392 GNDA.n1667 GNDA.n1666 585
R393 GNDA.n1666 GNDA.n1665 585
R394 GNDA.n1668 GNDA.n1099 585
R395 GNDA.n1099 GNDA.n1098 585
R396 GNDA.n1670 GNDA.n1669 585
R397 GNDA.n1671 GNDA.n1670 585
R398 GNDA.n1096 GNDA.n1095 585
R399 GNDA.n1672 GNDA.n1096 585
R400 GNDA.n1675 GNDA.n1674 585
R401 GNDA.n1674 GNDA.n1673 585
R402 GNDA.n1676 GNDA.n1094 585
R403 GNDA.n1097 GNDA.n1094 585
R404 GNDA.n1678 GNDA.n1677 585
R405 GNDA.n1679 GNDA.n1678 585
R406 GNDA.n1093 GNDA.n1092 585
R407 GNDA.n1680 GNDA.n1093 585
R408 GNDA.n1683 GNDA.n1682 585
R409 GNDA.n1682 GNDA.n1681 585
R410 GNDA.n1684 GNDA.n1090 585
R411 GNDA.n1090 GNDA.n1089 585
R412 GNDA.n1686 GNDA.n1685 585
R413 GNDA.n1687 GNDA.n1686 585
R414 GNDA.n1091 GNDA.n1087 585
R415 GNDA.n1688 GNDA.n1087 585
R416 GNDA.n1301 GNDA.n1297 585
R417 GNDA.n1303 GNDA.n1302 585
R418 GNDA.t209 GNDA.n1303 585
R419 GNDA.n1310 GNDA.n1309 585
R420 GNDA.n1310 GNDA.n1088 585
R421 GNDA.n1311 GNDA.n1307 585
R422 GNDA.n1312 GNDA.n1311 585
R423 GNDA.n1315 GNDA.n1314 585
R424 GNDA.n1314 GNDA.n1313 585
R425 GNDA.n1316 GNDA.n1305 585
R426 GNDA.n1305 GNDA.n1304 585
R427 GNDA.n1318 GNDA.n1317 585
R428 GNDA.n1319 GNDA.n1318 585
R429 GNDA.n1306 GNDA.n1295 585
R430 GNDA.n1320 GNDA.n1295 585
R431 GNDA.n1323 GNDA.n1322 585
R432 GNDA.n1322 GNDA.n1321 585
R433 GNDA.n1324 GNDA.n1293 585
R434 GNDA.n1293 GNDA.n1292 585
R435 GNDA.n1326 GNDA.n1325 585
R436 GNDA.n1327 GNDA.n1326 585
R437 GNDA.n1290 GNDA.n1289 585
R438 GNDA.n1328 GNDA.n1290 585
R439 GNDA.n1331 GNDA.n1330 585
R440 GNDA.n1330 GNDA.n1329 585
R441 GNDA.n1332 GNDA.n1288 585
R442 GNDA.n1291 GNDA.n1288 585
R443 GNDA.n1390 GNDA.n1335 585
R444 GNDA.n1390 GNDA.n1389 585
R445 GNDA.n1384 GNDA.n1334 585
R446 GNDA.n1388 GNDA.n1334 585
R447 GNDA.n1386 GNDA.n1385 585
R448 GNDA.n1387 GNDA.n1386 585
R449 GNDA.n1383 GNDA.n1337 585
R450 GNDA.n1337 GNDA.n1336 585
R451 GNDA.n1382 GNDA.n1381 585
R452 GNDA.n1381 GNDA.n1380 585
R453 GNDA.n1339 GNDA.n1338 585
R454 GNDA.n1379 GNDA.n1339 585
R455 GNDA.n1377 GNDA.n1376 585
R456 GNDA.n1378 GNDA.n1377 585
R457 GNDA.n1375 GNDA.n1341 585
R458 GNDA.n1341 GNDA.n1340 585
R459 GNDA.n1374 GNDA.n1373 585
R460 GNDA.n1373 GNDA.n1372 585
R461 GNDA.n1343 GNDA.n1342 585
R462 GNDA.n1371 GNDA.n1343 585
R463 GNDA.n1369 GNDA.n1368 585
R464 GNDA.n1370 GNDA.n1369 585
R465 GNDA.n1367 GNDA.n1345 585
R466 GNDA.n1345 GNDA.n1344 585
R467 GNDA.n1424 GNDA.n1423 585
R468 GNDA.n1412 GNDA.n1156 585
R469 GNDA.n1413 GNDA.n1275 585
R470 GNDA.n1416 GNDA.n1415 585
R471 GNDA.n1278 GNDA.n1277 585
R472 GNDA.n1409 GNDA.n1408 585
R473 GNDA.n1283 GNDA.n1282 585
R474 GNDA.n1402 GNDA.n1401 585
R475 GNDA.n1400 GNDA.n1399 585
R476 GNDA.n1398 GNDA.n1287 585
R477 GNDA.n1286 GNDA.n1285 585
R478 GNDA.n1392 GNDA.n1391 585
R479 GNDA.n1425 GNDA.n986 585
R480 GNDA.n1425 GNDA.n1067 585
R481 GNDA.n1393 GNDA.n1392 585
R482 GNDA.n1395 GNDA.n1285 585
R483 GNDA.n1398 GNDA.n1397 585
R484 GNDA.n1399 GNDA.n1284 585
R485 GNDA.n1403 GNDA.n1402 585
R486 GNDA.n1405 GNDA.n1283 585
R487 GNDA.n1408 GNDA.n1407 585
R488 GNDA.n1277 GNDA.n1276 585
R489 GNDA.n1417 GNDA.n1416 585
R490 GNDA.n1419 GNDA.n1275 585
R491 GNDA.n1420 GNDA.n1156 585
R492 GNDA.n1423 GNDA.n1422 585
R493 GNDA.n1273 GNDA.n986 585
R494 GNDA.n1273 GNDA.n1067 585
R495 GNDA.n2022 GNDA.n1010 585
R496 GNDA.n2023 GNDA.n1008 585
R497 GNDA.n2024 GNDA.n1007 585
R498 GNDA.n1005 GNDA.n1003 585
R499 GNDA.n2030 GNDA.n1002 585
R500 GNDA.n2031 GNDA.n1000 585
R501 GNDA.n2032 GNDA.n999 585
R502 GNDA.n997 GNDA.n995 585
R503 GNDA.n2037 GNDA.n994 585
R504 GNDA.n2038 GNDA.n992 585
R505 GNDA.n991 GNDA.n987 585
R506 GNDA.n2043 GNDA.n941 585
R507 GNDA.n2043 GNDA.n2042 585
R508 GNDA.n2040 GNDA.n987 585
R509 GNDA.n2039 GNDA.n2038 585
R510 GNDA.n2037 GNDA.n2036 585
R511 GNDA.n2035 GNDA.n995 585
R512 GNDA.n2033 GNDA.n2032 585
R513 GNDA.n2031 GNDA.n996 585
R514 GNDA.n2030 GNDA.n2029 585
R515 GNDA.n2027 GNDA.n1003 585
R516 GNDA.n2025 GNDA.n2024 585
R517 GNDA.n2023 GNDA.n1004 585
R518 GNDA.n2022 GNDA.n2021 585
R519 GNDA.n2348 GNDA.n2347 585
R520 GNDA.n2349 GNDA.n465 585
R521 GNDA.n2350 GNDA.n464 585
R522 GNDA.n462 GNDA.n460 585
R523 GNDA.n2356 GNDA.n459 585
R524 GNDA.n2357 GNDA.n457 585
R525 GNDA.n2358 GNDA.n456 585
R526 GNDA.n454 GNDA.n452 585
R527 GNDA.n2363 GNDA.n451 585
R528 GNDA.n2364 GNDA.n449 585
R529 GNDA.n448 GNDA.n444 585
R530 GNDA.n2369 GNDA.n440 585
R531 GNDA.n2369 GNDA.n2368 585
R532 GNDA.n2366 GNDA.n444 585
R533 GNDA.n2365 GNDA.n2364 585
R534 GNDA.n2363 GNDA.n2362 585
R535 GNDA.n2361 GNDA.n452 585
R536 GNDA.n2359 GNDA.n2358 585
R537 GNDA.n2357 GNDA.n453 585
R538 GNDA.n2356 GNDA.n2355 585
R539 GNDA.n2353 GNDA.n460 585
R540 GNDA.n2351 GNDA.n2350 585
R541 GNDA.n2349 GNDA.n461 585
R542 GNDA.n2348 GNDA.n467 585
R543 GNDA.n886 GNDA.n606 585
R544 GNDA.n887 GNDA.n604 585
R545 GNDA.n888 GNDA.n603 585
R546 GNDA.n601 GNDA.n599 585
R547 GNDA.n894 GNDA.n598 585
R548 GNDA.n895 GNDA.n596 585
R549 GNDA.n896 GNDA.n595 585
R550 GNDA.n593 GNDA.n591 585
R551 GNDA.n901 GNDA.n590 585
R552 GNDA.n902 GNDA.n588 585
R553 GNDA.n587 GNDA.n583 585
R554 GNDA.n907 GNDA.n582 585
R555 GNDA.n907 GNDA.n906 585
R556 GNDA.n904 GNDA.n583 585
R557 GNDA.n903 GNDA.n902 585
R558 GNDA.n901 GNDA.n900 585
R559 GNDA.n899 GNDA.n591 585
R560 GNDA.n897 GNDA.n896 585
R561 GNDA.n895 GNDA.n592 585
R562 GNDA.n894 GNDA.n893 585
R563 GNDA.n891 GNDA.n599 585
R564 GNDA.n889 GNDA.n888 585
R565 GNDA.n887 GNDA.n600 585
R566 GNDA.n886 GNDA.n885 585
R567 GNDA.n2372 GNDA.n2371 585
R568 GNDA.n441 GNDA.n439 585
R569 GNDA.n2138 GNDA.n2137 585
R570 GNDA.n2140 GNDA.n2139 585
R571 GNDA.n2142 GNDA.n2141 585
R572 GNDA.n2144 GNDA.n2143 585
R573 GNDA.n2146 GNDA.n2145 585
R574 GNDA.n2148 GNDA.n2147 585
R575 GNDA.n2150 GNDA.n2149 585
R576 GNDA.n2152 GNDA.n2151 585
R577 GNDA.n2154 GNDA.n2153 585
R578 GNDA.n2155 GNDA.n2136 585
R579 GNDA.n581 GNDA.n580 585
R580 GNDA.n579 GNDA.n578 585
R581 GNDA.n577 GNDA.n576 585
R582 GNDA.n575 GNDA.n574 585
R583 GNDA.n573 GNDA.n572 585
R584 GNDA.n571 GNDA.n570 585
R585 GNDA.n569 GNDA.n568 585
R586 GNDA.n567 GNDA.n566 585
R587 GNDA.n565 GNDA.n564 585
R588 GNDA.n563 GNDA.n562 585
R589 GNDA.n561 GNDA.n560 585
R590 GNDA.n445 GNDA.n442 585
R591 GNDA.n643 GNDA.n642 585
R592 GNDA.n641 GNDA.n640 585
R593 GNDA.n639 GNDA.n638 585
R594 GNDA.n637 GNDA.n636 585
R595 GNDA.n635 GNDA.n634 585
R596 GNDA.n633 GNDA.n632 585
R597 GNDA.n631 GNDA.n630 585
R598 GNDA.n629 GNDA.n628 585
R599 GNDA.n627 GNDA.n626 585
R600 GNDA.n625 GNDA.n624 585
R601 GNDA.n623 GNDA.n622 585
R602 GNDA.n584 GNDA.n559 585
R603 GNDA.n557 GNDA.n443 585
R604 GNDA.n2058 GNDA.n557 585
R605 GNDA.n2129 GNDA.n2128 585
R606 GNDA.n2126 GNDA.n2125 585
R607 GNDA.n2124 GNDA.n2123 585
R608 GNDA.n534 GNDA.n496 585
R609 GNDA.n554 GNDA.n553 585
R610 GNDA.n550 GNDA.n533 585
R611 GNDA.n537 GNDA.n536 585
R612 GNDA.n545 GNDA.n544 585
R613 GNDA.n543 GNDA.n542 585
R614 GNDA.n517 GNDA.n516 585
R615 GNDA.n2063 GNDA.n2062 585
R616 GNDA.n1011 GNDA.n518 585
R617 GNDA.n909 GNDA.n558 585
R618 GNDA.n2058 GNDA.n558 585
R619 GNDA.n556 GNDA.n443 585
R620 GNDA.n2058 GNDA.n556 585
R621 GNDA.n2018 GNDA.n2017 585
R622 GNDA.n2015 GNDA.n2014 585
R623 GNDA.n2013 GNDA.n2012 585
R624 GNDA.n1929 GNDA.n1014 585
R625 GNDA.n1931 GNDA.n1930 585
R626 GNDA.n1935 GNDA.n1934 585
R627 GNDA.n1937 GNDA.n1936 585
R628 GNDA.n1944 GNDA.n1943 585
R629 GNDA.n1942 GNDA.n1927 585
R630 GNDA.n1950 GNDA.n1949 585
R631 GNDA.n1952 GNDA.n1951 585
R632 GNDA.n1925 GNDA.n1924 585
R633 GNDA.n2057 GNDA.n909 585
R634 GNDA.n2058 GNDA.n2057 585
R635 GNDA.n1922 GNDA.n910 585
R636 GNDA.n1920 GNDA.n1919 585
R637 GNDA.n1918 GNDA.n1917 585
R638 GNDA.n1834 GNDA.n1035 585
R639 GNDA.n1836 GNDA.n1835 585
R640 GNDA.n1840 GNDA.n1839 585
R641 GNDA.n1842 GNDA.n1841 585
R642 GNDA.n1849 GNDA.n1848 585
R643 GNDA.n1847 GNDA.n1832 585
R644 GNDA.n1855 GNDA.n1854 585
R645 GNDA.n1857 GNDA.n1856 585
R646 GNDA.n1830 GNDA.n1829 585
R647 GNDA.n664 GNDA.n614 585
R648 GNDA.n667 GNDA.n666 585
R649 GNDA.n666 GNDA.n665 585
R650 GNDA.n613 GNDA.n612 585
R651 GNDA.n662 GNDA.n613 585
R652 GNDA.n660 GNDA.n659 585
R653 GNDA.n661 GNDA.n660 585
R654 GNDA.n658 GNDA.n616 585
R655 GNDA.n616 GNDA.n615 585
R656 GNDA.n657 GNDA.n656 585
R657 GNDA.n656 GNDA.n387 585
R658 GNDA.n655 GNDA.n617 585
R659 GNDA.n655 GNDA.n386 585
R660 GNDA.n654 GNDA.n619 585
R661 GNDA.n654 GNDA.n653 585
R662 GNDA.n648 GNDA.n618 585
R663 GNDA.n652 GNDA.n618 585
R664 GNDA.n650 GNDA.n649 585
R665 GNDA.n651 GNDA.n650 585
R666 GNDA.n647 GNDA.n621 585
R667 GNDA.n621 GNDA.n620 585
R668 GNDA.n646 GNDA.n645 585
R669 GNDA.n645 GNDA.n644 585
R670 GNDA.n663 GNDA.n610 585
R671 GNDA.n1826 GNDA.n1825 585
R672 GNDA.n1824 GNDA.n1823 585
R673 GNDA.n1824 GNDA.n1056 585
R674 GNDA.n1822 GNDA.n1057 585
R675 GNDA.n1818 GNDA.n1057 585
R676 GNDA.n1821 GNDA.n1820 585
R677 GNDA.n1820 GNDA.n1819 585
R678 GNDA.n1059 GNDA.n1058 585
R679 GNDA.n1817 GNDA.n1059 585
R680 GNDA.n1815 GNDA.n1814 585
R681 GNDA.n1816 GNDA.n1815 585
R682 GNDA.n1813 GNDA.n1060 585
R683 GNDA.n1809 GNDA.n1060 585
R684 GNDA.n1812 GNDA.n1811 585
R685 GNDA.n1811 GNDA.n1810 585
R686 GNDA.n1062 GNDA.n1061 585
R687 GNDA.n1808 GNDA.n1062 585
R688 GNDA.n1806 GNDA.n1805 585
R689 GNDA.n1807 GNDA.n1806 585
R690 GNDA.n1804 GNDA.n1064 585
R691 GNDA.n1064 GNDA.n1063 585
R692 GNDA.n1803 GNDA.n1802 585
R693 GNDA.n1802 GNDA.n1801 585
R694 GNDA.n1828 GNDA.n1827 585
R695 GNDA.n1641 GNDA.n1640 585
R696 GNDA.n1644 GNDA.n1111 585
R697 GNDA.n1111 GNDA.n1110 585
R698 GNDA.n1646 GNDA.n1645 585
R699 GNDA.n1647 GNDA.n1646 585
R700 GNDA.n1108 GNDA.n1107 585
R701 GNDA.n1648 GNDA.n1108 585
R702 GNDA.n1651 GNDA.n1650 585
R703 GNDA.n1650 GNDA.n1649 585
R704 GNDA.n1652 GNDA.n1106 585
R705 GNDA.n1109 GNDA.n1106 585
R706 GNDA.n1654 GNDA.n1653 585
R707 GNDA.n1655 GNDA.n1654 585
R708 GNDA.n1105 GNDA.n1104 585
R709 GNDA.n1656 GNDA.n1105 585
R710 GNDA.n1659 GNDA.n1658 585
R711 GNDA.n1658 GNDA.n1657 585
R712 GNDA.n1660 GNDA.n1103 585
R713 GNDA.n1103 GNDA.n1102 585
R714 GNDA.n1662 GNDA.n1661 585
R715 GNDA.n1663 GNDA.n1662 585
R716 GNDA.n1101 GNDA.n1100 585
R717 GNDA.n1664 GNDA.n1101 585
R718 GNDA.n1639 GNDA.n1638 585
R719 GNDA.n92 GNDA.n91 585
R720 GNDA.n175 GNDA.n90 585
R721 GNDA.n179 GNDA.n90 585
R722 GNDA.n174 GNDA.n173 585
R723 GNDA.n172 GNDA.n171 585
R724 GNDA.n170 GNDA.n169 585
R725 GNDA.n168 GNDA.n167 585
R726 GNDA.n166 GNDA.n165 585
R727 GNDA.n164 GNDA.n163 585
R728 GNDA.n162 GNDA.n161 585
R729 GNDA.n160 GNDA.n159 585
R730 GNDA.n158 GNDA.n157 585
R731 GNDA.n156 GNDA.n155 585
R732 GNDA.n153 GNDA.n89 585
R733 GNDA.n179 GNDA.n89 585
R734 GNDA.n264 GNDA.n216 585
R735 GNDA.n262 GNDA.n215 585
R736 GNDA.n267 GNDA.n215 585
R737 GNDA.n261 GNDA.n260 585
R738 GNDA.n227 GNDA.n222 585
R739 GNDA.n225 GNDA.n221 585
R740 GNDA.n230 GNDA.n221 585
R741 GNDA.n224 GNDA.n220 585
R742 GNDA.n116 GNDA.n115 585
R743 GNDA.n113 GNDA.n112 585
R744 GNDA.n112 GNDA.n71 585
R745 GNDA.n121 GNDA.n120 585
R746 GNDA.n123 GNDA.n111 585
R747 GNDA.n126 GNDA.n125 585
R748 GNDA.n109 GNDA.n108 585
R749 GNDA.n131 GNDA.n130 585
R750 GNDA.n133 GNDA.n107 585
R751 GNDA.n136 GNDA.n135 585
R752 GNDA.n105 GNDA.n104 585
R753 GNDA.n141 GNDA.n140 585
R754 GNDA.n143 GNDA.n103 585
R755 GNDA.n145 GNDA.n144 585
R756 GNDA.n144 GNDA.n71 585
R757 GNDA.n2504 GNDA.n2503 585
R758 GNDA.n2537 GNDA.n2502 585
R759 GNDA.n2541 GNDA.n2502 585
R760 GNDA.n2536 GNDA.n2535 585
R761 GNDA.n2534 GNDA.n2533 585
R762 GNDA.n2532 GNDA.n2531 585
R763 GNDA.n2530 GNDA.n2529 585
R764 GNDA.n2528 GNDA.n2527 585
R765 GNDA.n2526 GNDA.n2525 585
R766 GNDA.n2524 GNDA.n2523 585
R767 GNDA.n2522 GNDA.n2521 585
R768 GNDA.n2520 GNDA.n2519 585
R769 GNDA.n2518 GNDA.n2517 585
R770 GNDA.n2515 GNDA.n24 585
R771 GNDA.n2541 GNDA.n24 585
R772 GNDA.n2460 GNDA.n2459 585
R773 GNDA.n2497 GNDA.n2458 585
R774 GNDA.n2501 GNDA.n2458 585
R775 GNDA.n2496 GNDA.n2495 585
R776 GNDA.n2494 GNDA.n2493 585
R777 GNDA.n2492 GNDA.n2491 585
R778 GNDA.n2490 GNDA.n2489 585
R779 GNDA.n2488 GNDA.n2487 585
R780 GNDA.n2486 GNDA.n2485 585
R781 GNDA.n2484 GNDA.n2483 585
R782 GNDA.n2482 GNDA.n2481 585
R783 GNDA.n2480 GNDA.n2479 585
R784 GNDA.n2478 GNDA.n2477 585
R785 GNDA.n2475 GNDA.n30 585
R786 GNDA.n2501 GNDA.n30 585
R787 GNDA.n182 GNDA.n181 585
R788 GNDA.n187 GNDA.n180 585
R789 GNDA.n191 GNDA.n180 585
R790 GNDA.n186 GNDA.n185 585
R791 GNDA.n184 GNDA.n79 585
R792 GNDA.n193 GNDA.n192 585
R793 GNDA.n192 GNDA.n191 585
R794 GNDA.n211 GNDA.n70 585
R795 GNDA.n279 GNDA.n278 585
R796 GNDA.n278 GNDA.n277 585
R797 GNDA.n304 GNDA.n65 585
R798 GNDA.n310 GNDA.n309 585
R799 GNDA.n315 GNDA.n310 585
R800 GNDA.n293 GNDA.n292 585
R801 GNDA.n298 GNDA.n57 585
R802 GNDA.n336 GNDA.n57 585
R803 GNDA.n287 GNDA.n283 585
R804 GNDA.n289 GNDA.n288 585
R805 GNDA.n288 GNDA.n17 585
R806 GNDA.n76 GNDA.n75 585
R807 GNDA.n205 GNDA.n74 585
R808 GNDA.n209 GNDA.n74 585
R809 GNDA.n204 GNDA.n203 585
R810 GNDA.n202 GNDA.n201 585
R811 GNDA.n199 GNDA.n73 585
R812 GNDA.n209 GNDA.n73 585
R813 GNDA.n274 GNDA.n269 585
R814 GNDA.n272 GNDA.n268 585
R815 GNDA.n277 GNDA.n268 585
R816 GNDA.n312 GNDA.n63 585
R817 GNDA.n317 GNDA.n316 585
R818 GNDA.n316 GNDA.n315 585
R819 GNDA.n333 GNDA.n59 585
R820 GNDA.n331 GNDA.n58 585
R821 GNDA.n336 GNDA.n58 585
R822 GNDA.n2544 GNDA.n2543 585
R823 GNDA.n2549 GNDA.n2542 585
R824 GNDA.n2553 GNDA.n2542 585
R825 GNDA.n2548 GNDA.n2547 585
R826 GNDA.n2546 GNDA.n16 585
R827 GNDA.n2555 GNDA.n2554 585
R828 GNDA.n2554 GNDA.n2553 585
R829 GNDA.n2445 GNDA.n2444 585
R830 GNDA.n2453 GNDA.n2443 585
R831 GNDA.n2457 GNDA.n2443 585
R832 GNDA.n2452 GNDA.n2451 585
R833 GNDA.n2450 GNDA.n2449 585
R834 GNDA.n2447 GNDA.n32 585
R835 GNDA.n2457 GNDA.n32 585
R836 GNDA.n325 GNDA.n321 585
R837 GNDA.n327 GNDA.n326 585
R838 GNDA.n326 GNDA.n17 585
R839 GNDA.n344 GNDA.n339 585
R840 GNDA.n342 GNDA.n338 585
R841 GNDA.n347 GNDA.n338 585
R842 GNDA.n341 GNDA.n55 585
R843 GNDA.n361 GNDA.n40 585
R844 GNDA.n359 GNDA.n39 585
R845 GNDA.n364 GNDA.n39 585
R846 GNDA.n358 GNDA.n357 585
R847 GNDA.n2421 GNDA.n383 585
R848 GNDA.n2424 GNDA.n2423 585
R849 GNDA.n2425 GNDA.n2424 585
R850 GNDA.n2416 GNDA.n2415 585
R851 GNDA.n2346 GNDA.n471 585
R852 GNDA.n2346 GNDA.n2345 585
R853 GNDA.n2321 GNDA.n2320 585
R854 GNDA.n2322 GNDA.n2321 585
R855 GNDA.n2318 GNDA.n473 585
R856 GNDA.n2187 GNDA.n473 585
R857 GNDA.n2185 GNDA.n2181 585
R858 GNDA.n2188 GNDA.n2185 585
R859 GNDA.n2313 GNDA.n2312 585
R860 GNDA.n2312 GNDA.n2311 585
R861 GNDA.n2190 GNDA.n2186 585
R862 GNDA.n2310 GNDA.n2186 585
R863 GNDA.n2308 GNDA.n2307 585
R864 GNDA.n2309 GNDA.n2308 585
R865 GNDA.n2233 GNDA.n2189 585
R866 GNDA.n2230 GNDA.n2189 585
R867 GNDA.n2235 GNDA.n2232 585
R868 GNDA.n2232 GNDA.n2231 585
R869 GNDA.n2241 GNDA.n2240 585
R870 GNDA.n2242 GNDA.n2241 585
R871 GNDA.n2212 GNDA.n2211 585
R872 GNDA.n2243 GNDA.n2212 585
R873 GNDA.n2247 GNDA.n2246 585
R874 GNDA.n2246 GNDA.n2245 585
R875 GNDA.n2209 GNDA.n470 585
R876 GNDA.n2244 GNDA.n470 585
R877 GNDA.n882 GNDA.n881 585
R878 GNDA.n881 GNDA.n417 585
R879 GNDA.n743 GNDA.n471 585
R880 GNDA.n744 GNDA.n743 585
R881 GNDA.n748 GNDA.n746 585
R882 GNDA.n746 GNDA.n745 585
R883 GNDA.n874 GNDA.n873 585
R884 GNDA.n875 GNDA.n874 585
R885 GNDA.n750 GNDA.n747 585
R886 GNDA.n755 GNDA.n747 585
R887 GNDA.n868 GNDA.n867 585
R888 GNDA.n867 GNDA.n866 585
R889 GNDA.n757 GNDA.n754 585
R890 GNDA.n865 GNDA.n754 585
R891 GNDA.n863 GNDA.n862 585
R892 GNDA.n864 GNDA.n863 585
R893 GNDA.n788 GNDA.n756 585
R894 GNDA.n787 GNDA.n756 585
R895 GNDA.n795 GNDA.n794 585
R896 GNDA.n796 GNDA.n795 585
R897 GNDA.n790 GNDA.n778 585
R898 GNDA.n797 GNDA.n778 585
R899 GNDA.n800 GNDA.n799 585
R900 GNDA.n799 GNDA.n798 585
R901 GNDA.n801 GNDA.n740 585
R902 GNDA.n742 GNDA.n740 585
R903 GNDA.n880 GNDA.n741 585
R904 GNDA.n880 GNDA.n879 585
R905 GNDA.n883 GNDA.n882 585
R906 GNDA.n883 GNDA.n414 585
R907 GNDA.n738 GNDA.n413 585
R908 GNDA.n2387 GNDA.n413 585
R909 GNDA.n2389 GNDA.n411 585
R910 GNDA.n2389 GNDA.n2388 585
R911 GNDA.n2405 GNDA.n2404 585
R912 GNDA.n2404 GNDA.n2403 585
R913 GNDA.n2392 GNDA.n2390 585
R914 GNDA.n2402 GNDA.n2390 585
R915 GNDA.n2400 GNDA.n2399 585
R916 GNDA.n2401 GNDA.n2400 585
R917 GNDA.n2395 GNDA.n388 585
R918 GNDA.n2391 GNDA.n388 585
R919 GNDA.n2413 GNDA.n2412 585
R920 GNDA.n2414 GNDA.n2413 585
R921 GNDA.n390 GNDA.n389 585
R922 GNDA.n671 GNDA.n389 585
R923 GNDA.n676 GNDA.n675 585
R924 GNDA.n677 GNDA.n676 585
R925 GNDA.n609 GNDA.n608 585
R926 GNDA.n678 GNDA.n609 585
R927 GNDA.n681 GNDA.n680 585
R928 GNDA.n680 GNDA.n679 585
R929 GNDA.n670 GNDA.n669 585
R930 GNDA.n670 GNDA.n374 585
R931 GNDA.n2228 GNDA.n2227 585
R932 GNDA.n2229 GNDA.n2228 585
R933 GNDA.n2217 GNDA.n2215 585
R934 GNDA.n2221 GNDA.n2220 585
R935 GNDA.n2223 GNDA.n2222 585
R936 GNDA.n81 GNDA.n80 519.423
R937 GNDA.n1718 GNDA.t209 512.884
R938 GNDA.n152 GNDA.t279 505.467
R939 GNDA.n146 GNDA.t269 505.467
R940 GNDA.n2514 GNDA.t259 505.467
R941 GNDA.n2474 GNDA.t246 505.467
R942 GNDA.n280 GNDA.t210 499.442
R943 GNDA.n290 GNDA.t221 499.442
R944 GNDA.n271 GNDA.t224 489.401
R945 GNDA.n318 GNDA.t242 489.401
R946 GNDA.n330 GNDA.t219 489.401
R947 GNDA.n328 GNDA.t235 489.401
R948 GNDA.n67 GNDA.t250 475.976
R949 GNDA.n67 GNDA.t229 475.976
R950 GNDA.n299 GNDA.t202 475.976
R951 GNDA.n299 GNDA.t282 475.976
R952 GNDA.n277 GNDA.n209 445.375
R953 GNDA.n2553 GNDA.n17 445.375
R954 GNDA.t85 GNDA.n372 433.382
R955 GNDA.n2325 GNDA.t272 409.067
R956 GNDA.n2342 GNDA.t214 409.067
R957 GNDA.n2339 GNDA.t288 409.067
R958 GNDA.n2377 GNDA.t253 409.067
R959 GNDA.n2384 GNDA.t275 409.067
R960 GNDA.n2435 GNDA.t262 409.067
R961 GNDA.n1705 GNDA.t209 391.411
R962 GNDA.n347 GNDA.t292 364.418
R963 GNDA.n364 GNDA.t266 364.418
R964 GNDA.n921 GNDA.t209 172.876
R965 GNDA.n2049 GNDA.t209 172.876
R966 GNDA.t209 GNDA.n418 172.876
R967 GNDA.t209 GNDA.n421 172.876
R968 GNDA.n922 GNDA.t209 172.615
R969 GNDA.n912 GNDA.t209 172.615
R970 GNDA.t209 GNDA.n420 172.615
R971 GNDA.t209 GNDA.n385 172.615
R972 GNDA.t292 GNDA.t116 296.933
R973 GNDA.t36 GNDA.t266 296.933
R974 GNDA.t139 GNDA.t209 294.625
R975 GNDA.n177 GNDA.n176 267.125
R976 GNDA.n154 GNDA.n101 267.125
R977 GNDA.n118 GNDA.n117 267.125
R978 GNDA.n139 GNDA.n102 267.125
R979 GNDA.n207 GNDA.n206 267.125
R980 GNDA.n200 GNDA.n77 267.125
R981 GNDA.n189 GNDA.n188 267.125
R982 GNDA.n183 GNDA.n78 267.125
R983 GNDA.n2551 GNDA.n2550 267.125
R984 GNDA.n2545 GNDA.n15 267.125
R985 GNDA.n2455 GNDA.n2454 267.125
R986 GNDA.n2448 GNDA.n2446 267.125
R987 GNDA.n2539 GNDA.n2538 267.125
R988 GNDA.n2516 GNDA.n2513 267.125
R989 GNDA.n2499 GNDA.n2498 267.125
R990 GNDA.n2476 GNDA.n2469 267.125
R991 GNDA.n2177 GNDA.n2176 264.301
R992 GNDA.n2176 GNDA.n483 264.301
R993 GNDA.n492 GNDA.n490 264.301
R994 GNDA.n668 GNDA.n611 264.301
R995 GNDA.n1055 GNDA.n1054 264.301
R996 GNDA.n1643 GNDA.n1642 264.301
R997 GNDA.n645 GNDA.n643 259.416
R998 GNDA.n582 GNDA.n581 259.416
R999 GNDA.n1391 GNDA.n1390 259.416
R1000 GNDA.n2372 GNDA.n440 259.416
R1001 GNDA.n2046 GNDA.n941 259.416
R1002 GNDA.n1802 GNDA.n1800 259.416
R1003 GNDA.n1746 GNDA.n1745 259.416
R1004 GNDA.n1666 GNDA.n1101 259.416
R1005 GNDA.n1310 GNDA.n1085 259.416
R1006 GNDA.n1483 GNDA.n1152 258.334
R1007 GNDA.n2284 GNDA.n2207 258.334
R1008 GNDA.n2102 GNDA.n2101 258.334
R1009 GNDA.n1991 GNDA.n1990 258.334
R1010 GNDA.n1896 GNDA.n1895 258.334
R1011 GNDA.n1245 GNDA.n1244 258.334
R1012 GNDA.n1579 GNDA.n1537 258.334
R1013 GNDA.n838 GNDA.n774 258.334
R1014 GNDA.n720 GNDA.n719 258.334
R1015 GNDA.n2176 GNDA.n2175 254.34
R1016 GNDA.n2176 GNDA.n2134 254.34
R1017 GNDA.n2176 GNDA.n2133 254.34
R1018 GNDA.n2176 GNDA.n2132 254.34
R1019 GNDA.n2176 GNDA.n2131 254.34
R1020 GNDA.n2176 GNDA.n477 254.34
R1021 GNDA.n2176 GNDA.n478 254.34
R1022 GNDA.n2176 GNDA.n479 254.34
R1023 GNDA.n2176 GNDA.n480 254.34
R1024 GNDA.n2176 GNDA.n481 254.34
R1025 GNDA.n2176 GNDA.n484 254.34
R1026 GNDA.n2176 GNDA.n485 254.34
R1027 GNDA.n2176 GNDA.n486 254.34
R1028 GNDA.n2176 GNDA.n487 254.34
R1029 GNDA.n2176 GNDA.n488 254.34
R1030 GNDA.n2176 GNDA.n489 254.34
R1031 GNDA.n2051 GNDA.n2049 254.34
R1032 GNDA.n2049 GNDA.n920 254.34
R1033 GNDA.n2049 GNDA.n919 254.34
R1034 GNDA.n2049 GNDA.n918 254.34
R1035 GNDA.n2049 GNDA.n917 254.34
R1036 GNDA.n2049 GNDA.n916 254.34
R1037 GNDA.n1723 GNDA.n912 254.34
R1038 GNDA.n1771 GNDA.n912 254.34
R1039 GNDA.n1765 GNDA.n912 254.34
R1040 GNDA.n1763 GNDA.n912 254.34
R1041 GNDA.n1756 GNDA.n912 254.34
R1042 GNDA.n2055 GNDA.n912 254.34
R1043 GNDA.n2048 GNDA.n2047 254.34
R1044 GNDA.n2048 GNDA.n939 254.34
R1045 GNDA.n2048 GNDA.n938 254.34
R1046 GNDA.n2048 GNDA.n937 254.34
R1047 GNDA.n2048 GNDA.n936 254.34
R1048 GNDA.n2048 GNDA.n935 254.34
R1049 GNDA.n2048 GNDA.n934 254.34
R1050 GNDA.n2048 GNDA.n933 254.34
R1051 GNDA.n2048 GNDA.n932 254.34
R1052 GNDA.n2048 GNDA.n931 254.34
R1053 GNDA.n2048 GNDA.n930 254.34
R1054 GNDA.n2048 GNDA.n929 254.34
R1055 GNDA.n2048 GNDA.n928 254.34
R1056 GNDA.n2048 GNDA.n927 254.34
R1057 GNDA.n2048 GNDA.n926 254.34
R1058 GNDA.n2048 GNDA.n925 254.34
R1059 GNDA.n2048 GNDA.n924 254.34
R1060 GNDA.n2048 GNDA.n923 254.34
R1061 GNDA.n1517 GNDA.n1516 254.34
R1062 GNDA.n1517 GNDA.n1124 254.34
R1063 GNDA.n1517 GNDA.n1123 254.34
R1064 GNDA.n1517 GNDA.n1122 254.34
R1065 GNDA.n1517 GNDA.n1121 254.34
R1066 GNDA.n1517 GNDA.n1120 254.34
R1067 GNDA.n1517 GNDA.n1119 254.34
R1068 GNDA.n1517 GNDA.n1118 254.34
R1069 GNDA.n1517 GNDA.n1117 254.34
R1070 GNDA.n1517 GNDA.n1116 254.34
R1071 GNDA.n1517 GNDA.n1115 254.34
R1072 GNDA.n1517 GNDA.n1114 254.34
R1073 GNDA.n1530 GNDA.n1517 254.34
R1074 GNDA.n1606 GNDA.n1517 254.34
R1075 GNDA.n1608 GNDA.n1517 254.34
R1076 GNDA.n1621 GNDA.n1517 254.34
R1077 GNDA.n1623 GNDA.n1517 254.34
R1078 GNDA.n1636 GNDA.n1517 254.34
R1079 GNDA.n1411 GNDA.n1155 254.34
R1080 GNDA.n1414 GNDA.n1411 254.34
R1081 GNDA.n1411 GNDA.n1410 254.34
R1082 GNDA.n1411 GNDA.n1281 254.34
R1083 GNDA.n1411 GNDA.n1280 254.34
R1084 GNDA.n1411 GNDA.n1279 254.34
R1085 GNDA.n1394 GNDA.n1274 254.34
R1086 GNDA.n1396 GNDA.n1274 254.34
R1087 GNDA.n1404 GNDA.n1274 254.34
R1088 GNDA.n1406 GNDA.n1274 254.34
R1089 GNDA.n1418 GNDA.n1274 254.34
R1090 GNDA.n1421 GNDA.n1274 254.34
R1091 GNDA.n1009 GNDA.n921 254.34
R1092 GNDA.n1006 GNDA.n921 254.34
R1093 GNDA.n1001 GNDA.n921 254.34
R1094 GNDA.n998 GNDA.n921 254.34
R1095 GNDA.n993 GNDA.n921 254.34
R1096 GNDA.n990 GNDA.n921 254.34
R1097 GNDA.n2041 GNDA.n922 254.34
R1098 GNDA.n989 GNDA.n922 254.34
R1099 GNDA.n2034 GNDA.n922 254.34
R1100 GNDA.n2028 GNDA.n922 254.34
R1101 GNDA.n2026 GNDA.n922 254.34
R1102 GNDA.n2020 GNDA.n922 254.34
R1103 GNDA.n469 GNDA.n418 254.34
R1104 GNDA.n463 GNDA.n418 254.34
R1105 GNDA.n458 GNDA.n418 254.34
R1106 GNDA.n455 GNDA.n418 254.34
R1107 GNDA.n450 GNDA.n418 254.34
R1108 GNDA.n447 GNDA.n418 254.34
R1109 GNDA.n2367 GNDA.n420 254.34
R1110 GNDA.n446 GNDA.n420 254.34
R1111 GNDA.n2360 GNDA.n420 254.34
R1112 GNDA.n2354 GNDA.n420 254.34
R1113 GNDA.n2352 GNDA.n420 254.34
R1114 GNDA.n466 GNDA.n420 254.34
R1115 GNDA.n605 GNDA.n421 254.34
R1116 GNDA.n602 GNDA.n421 254.34
R1117 GNDA.n597 GNDA.n421 254.34
R1118 GNDA.n594 GNDA.n421 254.34
R1119 GNDA.n589 GNDA.n421 254.34
R1120 GNDA.n586 GNDA.n421 254.34
R1121 GNDA.n905 GNDA.n385 254.34
R1122 GNDA.n585 GNDA.n385 254.34
R1123 GNDA.n898 GNDA.n385 254.34
R1124 GNDA.n892 GNDA.n385 254.34
R1125 GNDA.n890 GNDA.n385 254.34
R1126 GNDA.n884 GNDA.n385 254.34
R1127 GNDA.n2374 GNDA.n2373 254.34
R1128 GNDA.n2374 GNDA.n438 254.34
R1129 GNDA.n2374 GNDA.n437 254.34
R1130 GNDA.n2374 GNDA.n436 254.34
R1131 GNDA.n2374 GNDA.n435 254.34
R1132 GNDA.n2374 GNDA.n434 254.34
R1133 GNDA.n2374 GNDA.n433 254.34
R1134 GNDA.n2374 GNDA.n432 254.34
R1135 GNDA.n2374 GNDA.n431 254.34
R1136 GNDA.n2374 GNDA.n430 254.34
R1137 GNDA.n2374 GNDA.n429 254.34
R1138 GNDA.n2374 GNDA.n428 254.34
R1139 GNDA.n2374 GNDA.n427 254.34
R1140 GNDA.n2374 GNDA.n426 254.34
R1141 GNDA.n2374 GNDA.n425 254.34
R1142 GNDA.n2374 GNDA.n424 254.34
R1143 GNDA.n2374 GNDA.n423 254.34
R1144 GNDA.n2374 GNDA.n422 254.34
R1145 GNDA.n2060 GNDA.n491 254.34
R1146 GNDA.n2060 GNDA.n495 254.34
R1147 GNDA.n2060 GNDA.n555 254.34
R1148 GNDA.n2060 GNDA.n532 254.34
R1149 GNDA.n2060 GNDA.n531 254.34
R1150 GNDA.n2061 GNDA.n2060 254.34
R1151 GNDA.n2060 GNDA.n530 254.34
R1152 GNDA.n2060 GNDA.n529 254.34
R1153 GNDA.n2060 GNDA.n528 254.34
R1154 GNDA.n2060 GNDA.n527 254.34
R1155 GNDA.n2060 GNDA.n526 254.34
R1156 GNDA.n2060 GNDA.n525 254.34
R1157 GNDA.n2060 GNDA.n524 254.34
R1158 GNDA.n2060 GNDA.n523 254.34
R1159 GNDA.n2060 GNDA.n522 254.34
R1160 GNDA.n2060 GNDA.n521 254.34
R1161 GNDA.n2060 GNDA.n520 254.34
R1162 GNDA.n2060 GNDA.n519 254.34
R1163 GNDA.t209 GNDA.n1296 250.349
R1164 GNDA.n906 GNDA.n584 249.663
R1165 GNDA.n2368 GNDA.n445 249.663
R1166 GNDA.n1365 GNDA.n1345 249.663
R1167 GNDA.n2174 GNDA.n2136 249.663
R1168 GNDA.n964 GNDA.n963 249.663
R1169 GNDA.n1777 GNDA.n1776 249.663
R1170 GNDA.n2042 GNDA.n988 249.663
R1171 GNDA.n1691 GNDA.n1087 249.663
R1172 GNDA.n1393 GNDA.n1288 249.663
R1173 GNDA.n2424 GNDA.n383 246.25
R1174 GNDA.n2424 GNDA.n2415 246.25
R1175 GNDA.n40 GNDA.n39 246.25
R1176 GNDA.n357 GNDA.n39 246.25
R1177 GNDA.n339 GNDA.n338 246.25
R1178 GNDA.n338 GNDA.n55 246.25
R1179 GNDA.n326 GNDA.n325 246.25
R1180 GNDA.n2444 GNDA.n2443 246.25
R1181 GNDA.n2451 GNDA.n2443 246.25
R1182 GNDA.n2449 GNDA.n32 246.25
R1183 GNDA.n2543 GNDA.n2542 246.25
R1184 GNDA.n2547 GNDA.n2542 246.25
R1185 GNDA.n2554 GNDA.n16 246.25
R1186 GNDA.n59 GNDA.n58 246.25
R1187 GNDA.n316 GNDA.n63 246.25
R1188 GNDA.n269 GNDA.n268 246.25
R1189 GNDA.n75 GNDA.n74 246.25
R1190 GNDA.n203 GNDA.n74 246.25
R1191 GNDA.n201 GNDA.n73 246.25
R1192 GNDA.n288 GNDA.n287 246.25
R1193 GNDA.n292 GNDA.n57 246.25
R1194 GNDA.n310 GNDA.n65 246.25
R1195 GNDA.n278 GNDA.n70 246.25
R1196 GNDA.n181 GNDA.n180 246.25
R1197 GNDA.n185 GNDA.n180 246.25
R1198 GNDA.n192 GNDA.n79 246.25
R1199 GNDA.n2459 GNDA.n2458 246.25
R1200 GNDA.n2495 GNDA.n2458 246.25
R1201 GNDA.n2493 GNDA.n2492 246.25
R1202 GNDA.n2489 GNDA.n2488 246.25
R1203 GNDA.n2485 GNDA.n2484 246.25
R1204 GNDA.n2481 GNDA.n2480 246.25
R1205 GNDA.n2477 GNDA.n30 246.25
R1206 GNDA.n2503 GNDA.n2502 246.25
R1207 GNDA.n2535 GNDA.n2502 246.25
R1208 GNDA.n2533 GNDA.n2532 246.25
R1209 GNDA.n2529 GNDA.n2528 246.25
R1210 GNDA.n2525 GNDA.n2524 246.25
R1211 GNDA.n2521 GNDA.n2520 246.25
R1212 GNDA.n2517 GNDA.n24 246.25
R1213 GNDA.n115 GNDA.n112 246.25
R1214 GNDA.n121 GNDA.n112 246.25
R1215 GNDA.n125 GNDA.n123 246.25
R1216 GNDA.n131 GNDA.n108 246.25
R1217 GNDA.n135 GNDA.n133 246.25
R1218 GNDA.n141 GNDA.n104 246.25
R1219 GNDA.n144 GNDA.n143 246.25
R1220 GNDA.n222 GNDA.n221 246.25
R1221 GNDA.n221 GNDA.n220 246.25
R1222 GNDA.n216 GNDA.n215 246.25
R1223 GNDA.n260 GNDA.n215 246.25
R1224 GNDA.n91 GNDA.n90 246.25
R1225 GNDA.n173 GNDA.n90 246.25
R1226 GNDA.n171 GNDA.n170 246.25
R1227 GNDA.n167 GNDA.n166 246.25
R1228 GNDA.n163 GNDA.n162 246.25
R1229 GNDA.n159 GNDA.n158 246.25
R1230 GNDA.n155 GNDA.n89 246.25
R1231 GNDA.n2228 GNDA.n2215 246.25
R1232 GNDA.n2222 GNDA.n2221 246.25
R1233 GNDA.n2431 GNDA.n2430 241.643
R1234 GNDA.n179 GNDA.n178 241.643
R1235 GNDA.n179 GNDA.n84 241.643
R1236 GNDA.n179 GNDA.n85 241.643
R1237 GNDA.n179 GNDA.n86 241.643
R1238 GNDA.n179 GNDA.n87 241.643
R1239 GNDA.n179 GNDA.n88 241.643
R1240 GNDA.n267 GNDA.n266 241.643
R1241 GNDA.n267 GNDA.n214 241.643
R1242 GNDA.n230 GNDA.n229 241.643
R1243 GNDA.n231 GNDA.n230 241.643
R1244 GNDA.n114 GNDA.n71 241.643
R1245 GNDA.n122 GNDA.n71 241.643
R1246 GNDA.n124 GNDA.n71 241.643
R1247 GNDA.n132 GNDA.n71 241.643
R1248 GNDA.n134 GNDA.n71 241.643
R1249 GNDA.n142 GNDA.n71 241.643
R1250 GNDA.n2541 GNDA.n2540 241.643
R1251 GNDA.n2541 GNDA.n19 241.643
R1252 GNDA.n2541 GNDA.n20 241.643
R1253 GNDA.n2541 GNDA.n21 241.643
R1254 GNDA.n2541 GNDA.n22 241.643
R1255 GNDA.n2541 GNDA.n23 241.643
R1256 GNDA.n2501 GNDA.n2500 241.643
R1257 GNDA.n2501 GNDA.n25 241.643
R1258 GNDA.n2501 GNDA.n26 241.643
R1259 GNDA.n2501 GNDA.n27 241.643
R1260 GNDA.n2501 GNDA.n28 241.643
R1261 GNDA.n2501 GNDA.n29 241.643
R1262 GNDA.n191 GNDA.n190 241.643
R1263 GNDA.n191 GNDA.n83 241.643
R1264 GNDA.n277 GNDA.n213 241.643
R1265 GNDA.n315 GNDA.n64 241.643
R1266 GNDA.n336 GNDA.n56 241.643
R1267 GNDA.n286 GNDA.n17 241.643
R1268 GNDA.n209 GNDA.n208 241.643
R1269 GNDA.n209 GNDA.n72 241.643
R1270 GNDA.n277 GNDA.n276 241.643
R1271 GNDA.n315 GNDA.n314 241.643
R1272 GNDA.n336 GNDA.n335 241.643
R1273 GNDA.n2553 GNDA.n2552 241.643
R1274 GNDA.n2553 GNDA.n18 241.643
R1275 GNDA.n2457 GNDA.n2456 241.643
R1276 GNDA.n2457 GNDA.n31 241.643
R1277 GNDA.n324 GNDA.n17 241.643
R1278 GNDA.n347 GNDA.n346 241.643
R1279 GNDA.n348 GNDA.n347 241.643
R1280 GNDA.n364 GNDA.n363 241.643
R1281 GNDA.n364 GNDA.n38 241.643
R1282 GNDA.n2426 GNDA.n2425 241.643
R1283 GNDA.n2425 GNDA.n384 241.643
R1284 GNDA.n2229 GNDA.n2213 241.643
R1285 GNDA.n2229 GNDA.n2214 241.643
R1286 GNDA.n44 GNDA.n42 206.052
R1287 GNDA.n5 GNDA.n3 206.052
R1288 GNDA.n50 GNDA.n49 205.488
R1289 GNDA.n48 GNDA.n47 205.488
R1290 GNDA.n46 GNDA.n45 205.488
R1291 GNDA.n44 GNDA.n43 205.488
R1292 GNDA.n11 GNDA.n10 205.488
R1293 GNDA.n9 GNDA.n8 205.488
R1294 GNDA.n7 GNDA.n6 205.488
R1295 GNDA.n5 GNDA.n4 205.488
R1296 GNDA.n52 GNDA.n51 200.988
R1297 GNDA.n13 GNDA.n12 200.988
R1298 GNDA.n670 GNDA.n610 197
R1299 GNDA.n881 GNDA.n880 197
R1300 GNDA.n1426 GNDA.n1425 197
R1301 GNDA.n2346 GNDA.n470 197
R1302 GNDA.n557 GNDA.n518 197
R1303 GNDA.n1829 GNDA.n1828 197
R1304 GNDA.n1924 GNDA.n558 197
R1305 GNDA.n1638 GNDA.n1637 197
R1306 GNDA.n1178 GNDA.n1066 197
R1307 GNDA.n1303 GNDA.n1297 197
R1308 GNDA.n883 GNDA.n413 187.249
R1309 GNDA.n746 GNDA.n743 187.249
R1310 GNDA.n1515 GNDA.n1126 187.249
R1311 GNDA.n2321 GNDA.n472 187.249
R1312 GNDA.n2130 GNDA.n2129 187.249
R1313 GNDA.n2057 GNDA.n910 187.249
R1314 GNDA.n2017 GNDA.n556 187.249
R1315 GNDA.n1720 GNDA.n1068 187.249
R1316 GNDA.n1273 GNDA.n1272 187.249
R1317 GNDA.n2427 GNDA.n382 185
R1318 GNDA.n2419 GNDA.n2418 185
R1319 GNDA.n118 GNDA.n113 185
R1320 GNDA.n120 GNDA.n119 185
R1321 GNDA.n111 GNDA.n110 185
R1322 GNDA.n127 GNDA.n126 185
R1323 GNDA.n128 GNDA.n109 185
R1324 GNDA.n130 GNDA.n129 185
R1325 GNDA.n107 GNDA.n106 185
R1326 GNDA.n137 GNDA.n136 185
R1327 GNDA.n138 GNDA.n105 185
R1328 GNDA.n140 GNDA.n139 185
R1329 GNDA.n265 GNDA.n217 185
R1330 GNDA.n228 GNDA.n223 185
R1331 GNDA.n212 GNDA.n210 185
R1332 GNDA.n307 GNDA.n306 185
R1333 GNDA.n309 GNDA.n66 185
R1334 GNDA.n296 GNDA.n295 185
R1335 GNDA.n298 GNDA.n291 185
R1336 GNDA.n285 GNDA.n284 185
R1337 GNDA.n206 GNDA.n205 185
R1338 GNDA.n204 GNDA.n77 185
R1339 GNDA.n188 GNDA.n187 185
R1340 GNDA.n186 GNDA.n183 185
R1341 GNDA.n275 GNDA.n270 185
R1342 GNDA.n313 GNDA.n311 185
R1343 GNDA.n334 GNDA.n60 185
R1344 GNDA.n323 GNDA.n322 185
R1345 GNDA.n345 GNDA.n340 185
R1346 GNDA.n362 GNDA.n41 185
R1347 GNDA.n2550 GNDA.n2549 185
R1348 GNDA.n2548 GNDA.n2545 185
R1349 GNDA.n2454 GNDA.n2453 185
R1350 GNDA.n2452 GNDA.n2446 185
R1351 GNDA.n2538 GNDA.n2537 185
R1352 GNDA.n2536 GNDA.n2505 185
R1353 GNDA.n2534 GNDA.n2506 185
R1354 GNDA.n2531 GNDA.n2507 185
R1355 GNDA.n2530 GNDA.n2508 185
R1356 GNDA.n2527 GNDA.n2509 185
R1357 GNDA.n2526 GNDA.n2510 185
R1358 GNDA.n2523 GNDA.n2511 185
R1359 GNDA.n2522 GNDA.n2512 185
R1360 GNDA.n2519 GNDA.n2513 185
R1361 GNDA.n2498 GNDA.n2497 185
R1362 GNDA.n2496 GNDA.n2461 185
R1363 GNDA.n2494 GNDA.n2462 185
R1364 GNDA.n2491 GNDA.n2463 185
R1365 GNDA.n2490 GNDA.n2464 185
R1366 GNDA.n2487 GNDA.n2465 185
R1367 GNDA.n2486 GNDA.n2466 185
R1368 GNDA.n2483 GNDA.n2467 185
R1369 GNDA.n2482 GNDA.n2468 185
R1370 GNDA.n2479 GNDA.n2469 185
R1371 GNDA.n176 GNDA.n175 185
R1372 GNDA.n174 GNDA.n93 185
R1373 GNDA.n172 GNDA.n94 185
R1374 GNDA.n169 GNDA.n95 185
R1375 GNDA.n168 GNDA.n96 185
R1376 GNDA.n165 GNDA.n97 185
R1377 GNDA.n164 GNDA.n98 185
R1378 GNDA.n161 GNDA.n99 185
R1379 GNDA.n160 GNDA.n100 185
R1380 GNDA.n157 GNDA.n101 185
R1381 GNDA.n1485 GNDA.n1152 185
R1382 GNDA.n1499 GNDA.n1498 185
R1383 GNDA.n1497 GNDA.n1153 185
R1384 GNDA.n1496 GNDA.n1495 185
R1385 GNDA.n1494 GNDA.n1493 185
R1386 GNDA.n1492 GNDA.n1491 185
R1387 GNDA.n1490 GNDA.n1489 185
R1388 GNDA.n1488 GNDA.n1487 185
R1389 GNDA.n1486 GNDA.n1129 185
R1390 GNDA.n1468 GNDA.n1467 185
R1391 GNDA.n1470 GNDA.n1469 185
R1392 GNDA.n1472 GNDA.n1471 185
R1393 GNDA.n1474 GNDA.n1473 185
R1394 GNDA.n1476 GNDA.n1475 185
R1395 GNDA.n1478 GNDA.n1477 185
R1396 GNDA.n1480 GNDA.n1479 185
R1397 GNDA.n1482 GNDA.n1481 185
R1398 GNDA.n1484 GNDA.n1483 185
R1399 GNDA.n1450 GNDA.n1449 185
R1400 GNDA.n1452 GNDA.n1451 185
R1401 GNDA.n1454 GNDA.n1453 185
R1402 GNDA.n1456 GNDA.n1455 185
R1403 GNDA.n1458 GNDA.n1457 185
R1404 GNDA.n1460 GNDA.n1459 185
R1405 GNDA.n1462 GNDA.n1461 185
R1406 GNDA.n1464 GNDA.n1463 185
R1407 GNDA.n1466 GNDA.n1465 185
R1408 GNDA.n1448 GNDA.n1447 185
R1409 GNDA.n1442 GNDA.n1441 185
R1410 GNDA.n1440 GNDA.n1439 185
R1411 GNDA.n1435 GNDA.n1434 185
R1412 GNDA.n1430 GNDA.n1137 185
R1413 GNDA.n1503 GNDA.n1502 185
R1414 GNDA.n1136 GNDA.n1134 185
R1415 GNDA.n1509 GNDA.n1508 185
R1416 GNDA.n1511 GNDA.n1510 185
R1417 GNDA.n2286 GNDA.n2207 185
R1418 GNDA.n2300 GNDA.n2299 185
R1419 GNDA.n2298 GNDA.n2208 185
R1420 GNDA.n2297 GNDA.n2296 185
R1421 GNDA.n2295 GNDA.n2294 185
R1422 GNDA.n2293 GNDA.n2292 185
R1423 GNDA.n2291 GNDA.n2290 185
R1424 GNDA.n2289 GNDA.n2288 185
R1425 GNDA.n2287 GNDA.n2180 185
R1426 GNDA.n2269 GNDA.n2268 185
R1427 GNDA.n2271 GNDA.n2270 185
R1428 GNDA.n2273 GNDA.n2272 185
R1429 GNDA.n2275 GNDA.n2274 185
R1430 GNDA.n2277 GNDA.n2276 185
R1431 GNDA.n2279 GNDA.n2278 185
R1432 GNDA.n2281 GNDA.n2280 185
R1433 GNDA.n2283 GNDA.n2282 185
R1434 GNDA.n2285 GNDA.n2284 185
R1435 GNDA.n2251 GNDA.n2250 185
R1436 GNDA.n2253 GNDA.n2252 185
R1437 GNDA.n2255 GNDA.n2254 185
R1438 GNDA.n2257 GNDA.n2256 185
R1439 GNDA.n2259 GNDA.n2258 185
R1440 GNDA.n2261 GNDA.n2260 185
R1441 GNDA.n2263 GNDA.n2262 185
R1442 GNDA.n2265 GNDA.n2264 185
R1443 GNDA.n2267 GNDA.n2266 185
R1444 GNDA.n2249 GNDA.n2248 185
R1445 GNDA.n2239 GNDA.n2238 185
R1446 GNDA.n2237 GNDA.n2236 185
R1447 GNDA.n2234 GNDA.n2192 185
R1448 GNDA.n2306 GNDA.n2305 185
R1449 GNDA.n2303 GNDA.n2191 185
R1450 GNDA.n2302 GNDA.n2184 185
R1451 GNDA.n2315 GNDA.n2314 185
R1452 GNDA.n2317 GNDA.n2316 185
R1453 GNDA.n2103 GNDA.n2102 185
R1454 GNDA.n2105 GNDA.n2104 185
R1455 GNDA.n2107 GNDA.n2106 185
R1456 GNDA.n2109 GNDA.n2108 185
R1457 GNDA.n2111 GNDA.n2110 185
R1458 GNDA.n2113 GNDA.n2112 185
R1459 GNDA.n2115 GNDA.n2114 185
R1460 GNDA.n2117 GNDA.n2116 185
R1461 GNDA.n2118 GNDA.n493 185
R1462 GNDA.n2085 GNDA.n2084 185
R1463 GNDA.n2087 GNDA.n2086 185
R1464 GNDA.n2089 GNDA.n2088 185
R1465 GNDA.n2091 GNDA.n2090 185
R1466 GNDA.n2093 GNDA.n2092 185
R1467 GNDA.n2095 GNDA.n2094 185
R1468 GNDA.n2097 GNDA.n2096 185
R1469 GNDA.n2099 GNDA.n2098 185
R1470 GNDA.n2101 GNDA.n2100 185
R1471 GNDA.n2067 GNDA.n2066 185
R1472 GNDA.n2069 GNDA.n2068 185
R1473 GNDA.n2071 GNDA.n2070 185
R1474 GNDA.n2073 GNDA.n2072 185
R1475 GNDA.n2075 GNDA.n2074 185
R1476 GNDA.n2077 GNDA.n2076 185
R1477 GNDA.n2079 GNDA.n2078 185
R1478 GNDA.n2081 GNDA.n2080 185
R1479 GNDA.n2083 GNDA.n2082 185
R1480 GNDA.n2065 GNDA.n2064 185
R1481 GNDA.n541 GNDA.n540 185
R1482 GNDA.n539 GNDA.n538 185
R1483 GNDA.n547 GNDA.n546 185
R1484 GNDA.n549 GNDA.n548 185
R1485 GNDA.n552 GNDA.n551 185
R1486 GNDA.n535 GNDA.n498 185
R1487 GNDA.n2122 GNDA.n2121 185
R1488 GNDA.n497 GNDA.n494 185
R1489 GNDA.n1992 GNDA.n1991 185
R1490 GNDA.n1994 GNDA.n1993 185
R1491 GNDA.n1996 GNDA.n1995 185
R1492 GNDA.n1998 GNDA.n1997 185
R1493 GNDA.n2000 GNDA.n1999 185
R1494 GNDA.n2002 GNDA.n2001 185
R1495 GNDA.n2004 GNDA.n2003 185
R1496 GNDA.n2006 GNDA.n2005 185
R1497 GNDA.n2007 GNDA.n1012 185
R1498 GNDA.n1974 GNDA.n1973 185
R1499 GNDA.n1976 GNDA.n1975 185
R1500 GNDA.n1978 GNDA.n1977 185
R1501 GNDA.n1980 GNDA.n1979 185
R1502 GNDA.n1982 GNDA.n1981 185
R1503 GNDA.n1984 GNDA.n1983 185
R1504 GNDA.n1986 GNDA.n1985 185
R1505 GNDA.n1988 GNDA.n1987 185
R1506 GNDA.n1990 GNDA.n1989 185
R1507 GNDA.n1956 GNDA.n1955 185
R1508 GNDA.n1958 GNDA.n1957 185
R1509 GNDA.n1960 GNDA.n1959 185
R1510 GNDA.n1962 GNDA.n1961 185
R1511 GNDA.n1964 GNDA.n1963 185
R1512 GNDA.n1966 GNDA.n1965 185
R1513 GNDA.n1968 GNDA.n1967 185
R1514 GNDA.n1970 GNDA.n1969 185
R1515 GNDA.n1972 GNDA.n1971 185
R1516 GNDA.n1954 GNDA.n1953 185
R1517 GNDA.n1948 GNDA.n1947 185
R1518 GNDA.n1946 GNDA.n1945 185
R1519 GNDA.n1941 GNDA.n1940 185
R1520 GNDA.n1939 GNDA.n1938 185
R1521 GNDA.n1933 GNDA.n1932 185
R1522 GNDA.n1928 GNDA.n1016 185
R1523 GNDA.n2011 GNDA.n2010 185
R1524 GNDA.n1015 GNDA.n1013 185
R1525 GNDA.n1897 GNDA.n1896 185
R1526 GNDA.n1899 GNDA.n1898 185
R1527 GNDA.n1901 GNDA.n1900 185
R1528 GNDA.n1903 GNDA.n1902 185
R1529 GNDA.n1905 GNDA.n1904 185
R1530 GNDA.n1907 GNDA.n1906 185
R1531 GNDA.n1909 GNDA.n1908 185
R1532 GNDA.n1911 GNDA.n1910 185
R1533 GNDA.n1912 GNDA.n1033 185
R1534 GNDA.n1879 GNDA.n1878 185
R1535 GNDA.n1881 GNDA.n1880 185
R1536 GNDA.n1883 GNDA.n1882 185
R1537 GNDA.n1885 GNDA.n1884 185
R1538 GNDA.n1887 GNDA.n1886 185
R1539 GNDA.n1889 GNDA.n1888 185
R1540 GNDA.n1891 GNDA.n1890 185
R1541 GNDA.n1893 GNDA.n1892 185
R1542 GNDA.n1895 GNDA.n1894 185
R1543 GNDA.n1861 GNDA.n1860 185
R1544 GNDA.n1863 GNDA.n1862 185
R1545 GNDA.n1865 GNDA.n1864 185
R1546 GNDA.n1867 GNDA.n1866 185
R1547 GNDA.n1869 GNDA.n1868 185
R1548 GNDA.n1871 GNDA.n1870 185
R1549 GNDA.n1873 GNDA.n1872 185
R1550 GNDA.n1875 GNDA.n1874 185
R1551 GNDA.n1877 GNDA.n1876 185
R1552 GNDA.n1859 GNDA.n1858 185
R1553 GNDA.n1853 GNDA.n1852 185
R1554 GNDA.n1851 GNDA.n1850 185
R1555 GNDA.n1846 GNDA.n1845 185
R1556 GNDA.n1844 GNDA.n1843 185
R1557 GNDA.n1838 GNDA.n1837 185
R1558 GNDA.n1833 GNDA.n1037 185
R1559 GNDA.n1916 GNDA.n1915 185
R1560 GNDA.n1036 GNDA.n1034 185
R1561 GNDA.n1246 GNDA.n1245 185
R1562 GNDA.n1248 GNDA.n1247 185
R1563 GNDA.n1250 GNDA.n1249 185
R1564 GNDA.n1252 GNDA.n1251 185
R1565 GNDA.n1254 GNDA.n1253 185
R1566 GNDA.n1256 GNDA.n1255 185
R1567 GNDA.n1258 GNDA.n1257 185
R1568 GNDA.n1260 GNDA.n1259 185
R1569 GNDA.n1261 GNDA.n1157 185
R1570 GNDA.n1228 GNDA.n1227 185
R1571 GNDA.n1230 GNDA.n1229 185
R1572 GNDA.n1232 GNDA.n1231 185
R1573 GNDA.n1234 GNDA.n1233 185
R1574 GNDA.n1236 GNDA.n1235 185
R1575 GNDA.n1238 GNDA.n1237 185
R1576 GNDA.n1240 GNDA.n1239 185
R1577 GNDA.n1242 GNDA.n1241 185
R1578 GNDA.n1244 GNDA.n1243 185
R1579 GNDA.n1210 GNDA.n1209 185
R1580 GNDA.n1212 GNDA.n1211 185
R1581 GNDA.n1214 GNDA.n1213 185
R1582 GNDA.n1216 GNDA.n1215 185
R1583 GNDA.n1218 GNDA.n1217 185
R1584 GNDA.n1220 GNDA.n1219 185
R1585 GNDA.n1222 GNDA.n1221 185
R1586 GNDA.n1224 GNDA.n1223 185
R1587 GNDA.n1226 GNDA.n1225 185
R1588 GNDA.n1579 GNDA.n1578 185
R1589 GNDA.n1581 GNDA.n1536 185
R1590 GNDA.n1584 GNDA.n1583 185
R1591 GNDA.n1585 GNDA.n1535 185
R1592 GNDA.n1587 GNDA.n1586 185
R1593 GNDA.n1589 GNDA.n1534 185
R1594 GNDA.n1592 GNDA.n1591 185
R1595 GNDA.n1593 GNDA.n1533 185
R1596 GNDA.n1598 GNDA.n1597 185
R1597 GNDA.n1561 GNDA.n1541 185
R1598 GNDA.n1563 GNDA.n1562 185
R1599 GNDA.n1565 GNDA.n1540 185
R1600 GNDA.n1568 GNDA.n1567 185
R1601 GNDA.n1569 GNDA.n1539 185
R1602 GNDA.n1571 GNDA.n1570 185
R1603 GNDA.n1573 GNDA.n1538 185
R1604 GNDA.n1576 GNDA.n1575 185
R1605 GNDA.n1577 GNDA.n1537 185
R1606 GNDA.n1632 GNDA.n1631 185
R1607 GNDA.n1546 GNDA.n1520 185
R1608 GNDA.n1548 GNDA.n1547 185
R1609 GNDA.n1550 GNDA.n1544 185
R1610 GNDA.n1552 GNDA.n1551 185
R1611 GNDA.n1553 GNDA.n1543 185
R1612 GNDA.n1555 GNDA.n1554 185
R1613 GNDA.n1557 GNDA.n1542 185
R1614 GNDA.n1560 GNDA.n1559 185
R1615 GNDA.n1630 GNDA.n1519 185
R1616 GNDA.n1628 GNDA.n1627 185
R1617 GNDA.n1523 GNDA.n1522 185
R1618 GNDA.n1618 GNDA.n1617 185
R1619 GNDA.n1615 GNDA.n1526 185
R1620 GNDA.n1613 GNDA.n1612 185
R1621 GNDA.n1528 GNDA.n1527 185
R1622 GNDA.n1603 GNDA.n1602 185
R1623 GNDA.n1600 GNDA.n1532 185
R1624 GNDA.n1208 GNDA.n1207 185
R1625 GNDA.n1202 GNDA.n1201 185
R1626 GNDA.n1200 GNDA.n1199 185
R1627 GNDA.n1195 GNDA.n1194 185
R1628 GNDA.n1193 GNDA.n1192 185
R1629 GNDA.n1187 GNDA.n1186 185
R1630 GNDA.n1182 GNDA.n1161 185
R1631 GNDA.n1265 GNDA.n1264 185
R1632 GNDA.n1160 GNDA.n1158 185
R1633 GNDA.n840 GNDA.n774 185
R1634 GNDA.n855 GNDA.n854 185
R1635 GNDA.n853 GNDA.n775 185
R1636 GNDA.n852 GNDA.n851 185
R1637 GNDA.n850 GNDA.n849 185
R1638 GNDA.n848 GNDA.n847 185
R1639 GNDA.n846 GNDA.n845 185
R1640 GNDA.n844 GNDA.n843 185
R1641 GNDA.n842 GNDA.n841 185
R1642 GNDA.n823 GNDA.n822 185
R1643 GNDA.n825 GNDA.n824 185
R1644 GNDA.n827 GNDA.n826 185
R1645 GNDA.n829 GNDA.n828 185
R1646 GNDA.n831 GNDA.n830 185
R1647 GNDA.n833 GNDA.n832 185
R1648 GNDA.n835 GNDA.n834 185
R1649 GNDA.n837 GNDA.n836 185
R1650 GNDA.n839 GNDA.n838 185
R1651 GNDA.n805 GNDA.n804 185
R1652 GNDA.n807 GNDA.n806 185
R1653 GNDA.n809 GNDA.n808 185
R1654 GNDA.n811 GNDA.n810 185
R1655 GNDA.n813 GNDA.n812 185
R1656 GNDA.n815 GNDA.n814 185
R1657 GNDA.n817 GNDA.n816 185
R1658 GNDA.n819 GNDA.n818 185
R1659 GNDA.n821 GNDA.n820 185
R1660 GNDA.n803 GNDA.n802 185
R1661 GNDA.n791 GNDA.n777 185
R1662 GNDA.n793 GNDA.n792 185
R1663 GNDA.n789 GNDA.n759 185
R1664 GNDA.n861 GNDA.n860 185
R1665 GNDA.n858 GNDA.n758 185
R1666 GNDA.n857 GNDA.n753 185
R1667 GNDA.n870 GNDA.n869 185
R1668 GNDA.n872 GNDA.n871 185
R1669 GNDA.n721 GNDA.n720 185
R1670 GNDA.n723 GNDA.n722 185
R1671 GNDA.n725 GNDA.n724 185
R1672 GNDA.n727 GNDA.n726 185
R1673 GNDA.n729 GNDA.n728 185
R1674 GNDA.n731 GNDA.n730 185
R1675 GNDA.n733 GNDA.n732 185
R1676 GNDA.n735 GNDA.n734 185
R1677 GNDA.n736 GNDA.n409 185
R1678 GNDA.n703 GNDA.n702 185
R1679 GNDA.n705 GNDA.n704 185
R1680 GNDA.n707 GNDA.n706 185
R1681 GNDA.n709 GNDA.n708 185
R1682 GNDA.n711 GNDA.n710 185
R1683 GNDA.n713 GNDA.n712 185
R1684 GNDA.n715 GNDA.n714 185
R1685 GNDA.n717 GNDA.n716 185
R1686 GNDA.n719 GNDA.n718 185
R1687 GNDA.n685 GNDA.n684 185
R1688 GNDA.n687 GNDA.n686 185
R1689 GNDA.n689 GNDA.n688 185
R1690 GNDA.n691 GNDA.n690 185
R1691 GNDA.n693 GNDA.n692 185
R1692 GNDA.n695 GNDA.n694 185
R1693 GNDA.n697 GNDA.n696 185
R1694 GNDA.n699 GNDA.n698 185
R1695 GNDA.n701 GNDA.n700 185
R1696 GNDA.n683 GNDA.n682 185
R1697 GNDA.n674 GNDA.n673 185
R1698 GNDA.n672 GNDA.n392 185
R1699 GNDA.n2411 GNDA.n2410 185
R1700 GNDA.n2394 GNDA.n391 185
R1701 GNDA.n2398 GNDA.n2397 185
R1702 GNDA.n2396 GNDA.n2393 185
R1703 GNDA.n412 GNDA.n410 185
R1704 GNDA.n2407 GNDA.n2406 185
R1705 GNDA.n2227 GNDA.n2216 185
R1706 GNDA.n2220 GNDA.n2216 185
R1707 GNDA.n2227 GNDA.n2226 185
R1708 GNDA.n2226 GNDA.n2225 185
R1709 GNDA.n1389 GNDA.t209 183.948
R1710 GNDA.n1689 GNDA.n1088 183.948
R1711 GNDA.n1291 GNDA.t209 180.013
R1712 GNDA.n1689 GNDA.n1688 180.013
R1713 GNDA.n645 GNDA.n621 175.546
R1714 GNDA.n650 GNDA.n621 175.546
R1715 GNDA.n650 GNDA.n618 175.546
R1716 GNDA.n654 GNDA.n618 175.546
R1717 GNDA.n655 GNDA.n654 175.546
R1718 GNDA.n656 GNDA.n655 175.546
R1719 GNDA.n656 GNDA.n616 175.546
R1720 GNDA.n660 GNDA.n616 175.546
R1721 GNDA.n660 GNDA.n613 175.546
R1722 GNDA.n666 GNDA.n613 175.546
R1723 GNDA.n666 GNDA.n614 175.546
R1724 GNDA.n624 GNDA.n623 175.546
R1725 GNDA.n628 GNDA.n627 175.546
R1726 GNDA.n632 GNDA.n631 175.546
R1727 GNDA.n636 GNDA.n635 175.546
R1728 GNDA.n640 GNDA.n639 175.546
R1729 GNDA.n2389 GNDA.n413 175.546
R1730 GNDA.n2404 GNDA.n2389 175.546
R1731 GNDA.n2404 GNDA.n2390 175.546
R1732 GNDA.n2400 GNDA.n2390 175.546
R1733 GNDA.n2400 GNDA.n388 175.546
R1734 GNDA.n2413 GNDA.n388 175.546
R1735 GNDA.n2413 GNDA.n389 175.546
R1736 GNDA.n676 GNDA.n389 175.546
R1737 GNDA.n676 GNDA.n609 175.546
R1738 GNDA.n680 GNDA.n609 175.546
R1739 GNDA.n680 GNDA.n670 175.546
R1740 GNDA.n904 GNDA.n903 175.546
R1741 GNDA.n900 GNDA.n899 175.546
R1742 GNDA.n897 GNDA.n592 175.546
R1743 GNDA.n893 GNDA.n891 175.546
R1744 GNDA.n889 GNDA.n600 175.546
R1745 GNDA.n588 GNDA.n587 175.546
R1746 GNDA.n593 GNDA.n590 175.546
R1747 GNDA.n596 GNDA.n595 175.546
R1748 GNDA.n601 GNDA.n598 175.546
R1749 GNDA.n604 GNDA.n603 175.546
R1750 GNDA.n562 GNDA.n561 175.546
R1751 GNDA.n566 GNDA.n565 175.546
R1752 GNDA.n570 GNDA.n569 175.546
R1753 GNDA.n574 GNDA.n573 175.546
R1754 GNDA.n578 GNDA.n577 175.546
R1755 GNDA.n874 GNDA.n746 175.546
R1756 GNDA.n874 GNDA.n747 175.546
R1757 GNDA.n867 GNDA.n747 175.546
R1758 GNDA.n867 GNDA.n754 175.546
R1759 GNDA.n863 GNDA.n754 175.546
R1760 GNDA.n863 GNDA.n756 175.546
R1761 GNDA.n795 GNDA.n756 175.546
R1762 GNDA.n795 GNDA.n778 175.546
R1763 GNDA.n799 GNDA.n778 175.546
R1764 GNDA.n799 GNDA.n740 175.546
R1765 GNDA.n880 GNDA.n740 175.546
R1766 GNDA.n2366 GNDA.n2365 175.546
R1767 GNDA.n2362 GNDA.n2361 175.546
R1768 GNDA.n2359 GNDA.n453 175.546
R1769 GNDA.n2355 GNDA.n2353 175.546
R1770 GNDA.n2351 GNDA.n461 175.546
R1771 GNDA.n1287 GNDA.n1286 175.546
R1772 GNDA.n1401 GNDA.n1400 175.546
R1773 GNDA.n1409 GNDA.n1282 175.546
R1774 GNDA.n1415 GNDA.n1278 175.546
R1775 GNDA.n1413 GNDA.n1412 175.546
R1776 GNDA.n1369 GNDA.n1345 175.546
R1777 GNDA.n1369 GNDA.n1343 175.546
R1778 GNDA.n1373 GNDA.n1343 175.546
R1779 GNDA.n1373 GNDA.n1341 175.546
R1780 GNDA.n1377 GNDA.n1341 175.546
R1781 GNDA.n1377 GNDA.n1339 175.546
R1782 GNDA.n1381 GNDA.n1339 175.546
R1783 GNDA.n1381 GNDA.n1337 175.546
R1784 GNDA.n1386 GNDA.n1337 175.546
R1785 GNDA.n1386 GNDA.n1334 175.546
R1786 GNDA.n1390 GNDA.n1334 175.546
R1787 GNDA.n1130 GNDA.n1125 175.546
R1788 GNDA.n1506 GNDA.n1505 175.546
R1789 GNDA.n1432 GNDA.n1431 175.546
R1790 GNDA.n1437 GNDA.n1436 175.546
R1791 GNDA.n1445 GNDA.n1444 175.546
R1792 GNDA.n1363 GNDA.n1362 175.546
R1793 GNDA.n1359 GNDA.n1358 175.546
R1794 GNDA.n1355 GNDA.n1354 175.546
R1795 GNDA.n1351 GNDA.n1350 175.546
R1796 GNDA.n1347 GNDA.n482 175.546
R1797 GNDA.n1127 GNDA.n482 175.546
R1798 GNDA.n449 GNDA.n448 175.546
R1799 GNDA.n454 GNDA.n451 175.546
R1800 GNDA.n457 GNDA.n456 175.546
R1801 GNDA.n462 GNDA.n459 175.546
R1802 GNDA.n465 GNDA.n464 175.546
R1803 GNDA.n2153 GNDA.n2152 175.546
R1804 GNDA.n2149 GNDA.n2148 175.546
R1805 GNDA.n2145 GNDA.n2144 175.546
R1806 GNDA.n2141 GNDA.n2140 175.546
R1807 GNDA.n2137 GNDA.n439 175.546
R1808 GNDA.n2321 GNDA.n473 175.546
R1809 GNDA.n2185 GNDA.n473 175.546
R1810 GNDA.n2312 GNDA.n2185 175.546
R1811 GNDA.n2312 GNDA.n2186 175.546
R1812 GNDA.n2308 GNDA.n2186 175.546
R1813 GNDA.n2308 GNDA.n2189 175.546
R1814 GNDA.n2232 GNDA.n2189 175.546
R1815 GNDA.n2241 GNDA.n2232 175.546
R1816 GNDA.n2241 GNDA.n2212 175.546
R1817 GNDA.n2246 GNDA.n2212 175.546
R1818 GNDA.n2246 GNDA.n470 175.546
R1819 GNDA.n2170 GNDA.n2135 175.546
R1820 GNDA.n2168 GNDA.n2167 175.546
R1821 GNDA.n2164 GNDA.n2163 175.546
R1822 GNDA.n2160 GNDA.n2159 175.546
R1823 GNDA.n2156 GNDA.n475 175.546
R1824 GNDA.n2178 GNDA.n475 175.546
R1825 GNDA.n992 GNDA.n991 175.546
R1826 GNDA.n997 GNDA.n994 175.546
R1827 GNDA.n1000 GNDA.n999 175.546
R1828 GNDA.n1005 GNDA.n1002 175.546
R1829 GNDA.n1008 GNDA.n1007 175.546
R1830 GNDA.n968 GNDA.n967 175.546
R1831 GNDA.n972 GNDA.n971 175.546
R1832 GNDA.n976 GNDA.n975 175.546
R1833 GNDA.n980 GNDA.n979 175.546
R1834 GNDA.n982 GNDA.n940 175.546
R1835 GNDA.n2125 GNDA.n2124 175.546
R1836 GNDA.n554 GNDA.n534 175.546
R1837 GNDA.n536 GNDA.n533 175.546
R1838 GNDA.n544 GNDA.n543 175.546
R1839 GNDA.n2062 GNDA.n517 175.546
R1840 GNDA.n960 GNDA.n959 175.546
R1841 GNDA.n956 GNDA.n955 175.546
R1842 GNDA.n952 GNDA.n951 175.546
R1843 GNDA.n948 GNDA.n947 175.546
R1844 GNDA.n944 GNDA.n943 175.546
R1845 GNDA.n1802 GNDA.n1064 175.546
R1846 GNDA.n1806 GNDA.n1064 175.546
R1847 GNDA.n1806 GNDA.n1062 175.546
R1848 GNDA.n1811 GNDA.n1062 175.546
R1849 GNDA.n1811 GNDA.n1060 175.546
R1850 GNDA.n1815 GNDA.n1060 175.546
R1851 GNDA.n1815 GNDA.n1059 175.546
R1852 GNDA.n1820 GNDA.n1059 175.546
R1853 GNDA.n1820 GNDA.n1057 175.546
R1854 GNDA.n1824 GNDA.n1057 175.546
R1855 GNDA.n1825 GNDA.n1824 175.546
R1856 GNDA.n1781 GNDA.n1780 175.546
R1857 GNDA.n1785 GNDA.n1784 175.546
R1858 GNDA.n1789 GNDA.n1788 175.546
R1859 GNDA.n1793 GNDA.n1792 175.546
R1860 GNDA.n1797 GNDA.n1796 175.546
R1861 GNDA.n1919 GNDA.n1918 175.546
R1862 GNDA.n1835 GNDA.n1834 175.546
R1863 GNDA.n1841 GNDA.n1840 175.546
R1864 GNDA.n1848 GNDA.n1847 175.546
R1865 GNDA.n1856 GNDA.n1855 175.546
R1866 GNDA.n1773 GNDA.n1772 175.546
R1867 GNDA.n1770 GNDA.n1750 175.546
R1868 GNDA.n1766 GNDA.n1764 175.546
R1869 GNDA.n1762 GNDA.n1757 175.546
R1870 GNDA.n2054 GNDA.n913 175.546
R1871 GNDA.n2040 GNDA.n2039 175.546
R1872 GNDA.n2036 GNDA.n2035 175.546
R1873 GNDA.n2033 GNDA.n996 175.546
R1874 GNDA.n2029 GNDA.n2027 175.546
R1875 GNDA.n2025 GNDA.n1004 175.546
R1876 GNDA.n1726 GNDA.n1725 175.546
R1877 GNDA.n1730 GNDA.n1729 175.546
R1878 GNDA.n1734 GNDA.n1733 175.546
R1879 GNDA.n1738 GNDA.n1737 175.546
R1880 GNDA.n1742 GNDA.n1741 175.546
R1881 GNDA.n2014 GNDA.n2013 175.546
R1882 GNDA.n1930 GNDA.n1929 175.546
R1883 GNDA.n1936 GNDA.n1935 175.546
R1884 GNDA.n1943 GNDA.n1942 175.546
R1885 GNDA.n1951 GNDA.n1950 175.546
R1886 GNDA.n1748 GNDA.n1747 175.546
R1887 GNDA.n1752 GNDA.n1751 175.546
R1888 GNDA.n1754 GNDA.n1753 175.546
R1889 GNDA.n1759 GNDA.n1758 175.546
R1890 GNDA.n2052 GNDA.n915 175.546
R1891 GNDA.n1662 GNDA.n1101 175.546
R1892 GNDA.n1662 GNDA.n1103 175.546
R1893 GNDA.n1658 GNDA.n1103 175.546
R1894 GNDA.n1658 GNDA.n1105 175.546
R1895 GNDA.n1654 GNDA.n1105 175.546
R1896 GNDA.n1654 GNDA.n1106 175.546
R1897 GNDA.n1650 GNDA.n1106 175.546
R1898 GNDA.n1650 GNDA.n1108 175.546
R1899 GNDA.n1646 GNDA.n1108 175.546
R1900 GNDA.n1646 GNDA.n1111 175.546
R1901 GNDA.n1641 GNDA.n1111 175.546
R1902 GNDA.n1686 GNDA.n1087 175.546
R1903 GNDA.n1686 GNDA.n1090 175.546
R1904 GNDA.n1682 GNDA.n1090 175.546
R1905 GNDA.n1682 GNDA.n1093 175.546
R1906 GNDA.n1678 GNDA.n1093 175.546
R1907 GNDA.n1678 GNDA.n1094 175.546
R1908 GNDA.n1674 GNDA.n1094 175.546
R1909 GNDA.n1674 GNDA.n1096 175.546
R1910 GNDA.n1670 GNDA.n1096 175.546
R1911 GNDA.n1670 GNDA.n1099 175.546
R1912 GNDA.n1666 GNDA.n1099 175.546
R1913 GNDA.n1605 GNDA.n1531 175.546
R1914 GNDA.n1609 GNDA.n1607 175.546
R1915 GNDA.n1620 GNDA.n1525 175.546
R1916 GNDA.n1624 GNDA.n1622 175.546
R1917 GNDA.n1635 GNDA.n1518 175.546
R1918 GNDA.n1692 GNDA.n1691 175.546
R1919 GNDA.n1692 GNDA.n1083 175.546
R1920 GNDA.n1698 GNDA.n1083 175.546
R1921 GNDA.n1698 GNDA.n1078 175.546
R1922 GNDA.n1704 GNDA.n1078 175.546
R1923 GNDA.n1706 GNDA.n1704 175.546
R1924 GNDA.n1707 GNDA.n1706 175.546
R1925 GNDA.n1707 GNDA.n1074 175.546
R1926 GNDA.n1713 GNDA.n1074 175.546
R1927 GNDA.n1713 GNDA.n1069 175.546
R1928 GNDA.n1719 GNDA.n1069 175.546
R1929 GNDA.n1397 GNDA.n1395 175.546
R1930 GNDA.n1403 GNDA.n1284 175.546
R1931 GNDA.n1407 GNDA.n1405 175.546
R1932 GNDA.n1417 GNDA.n1276 175.546
R1933 GNDA.n1420 GNDA.n1419 175.546
R1934 GNDA.n1330 GNDA.n1288 175.546
R1935 GNDA.n1330 GNDA.n1290 175.546
R1936 GNDA.n1326 GNDA.n1290 175.546
R1937 GNDA.n1326 GNDA.n1293 175.546
R1938 GNDA.n1322 GNDA.n1293 175.546
R1939 GNDA.n1322 GNDA.n1295 175.546
R1940 GNDA.n1318 GNDA.n1295 175.546
R1941 GNDA.n1318 GNDA.n1305 175.546
R1942 GNDA.n1314 GNDA.n1305 175.546
R1943 GNDA.n1314 GNDA.n1311 175.546
R1944 GNDA.n1311 GNDA.n1310 175.546
R1945 GNDA.n1268 GNDA.n1267 175.546
R1946 GNDA.n1184 GNDA.n1183 175.546
R1947 GNDA.n1190 GNDA.n1189 175.546
R1948 GNDA.n1197 GNDA.n1196 175.546
R1949 GNDA.n1205 GNDA.n1204 175.546
R1950 GNDA.n1694 GNDA.n1085 175.546
R1951 GNDA.n1695 GNDA.n1694 175.546
R1952 GNDA.n1695 GNDA.n1081 175.546
R1953 GNDA.n1701 GNDA.n1081 175.546
R1954 GNDA.n1702 GNDA.n1701 175.546
R1955 GNDA.n1702 GNDA.n1076 175.546
R1956 GNDA.n1709 GNDA.n1076 175.546
R1957 GNDA.n1710 GNDA.n1709 175.546
R1958 GNDA.n1710 GNDA.n1072 175.546
R1959 GNDA.n1716 GNDA.n1072 175.546
R1960 GNDA.n1717 GNDA.n1716 175.546
R1961 GNDA.n1411 GNDA.t209 172.876
R1962 GNDA.n1274 GNDA.t209 172.615
R1963 GNDA.n1449 GNDA.n1448 163.333
R1964 GNDA.n2250 GNDA.n2249 163.333
R1965 GNDA.n2066 GNDA.n2065 163.333
R1966 GNDA.n1955 GNDA.n1954 163.333
R1967 GNDA.n1860 GNDA.n1859 163.333
R1968 GNDA.n1209 GNDA.n1208 163.333
R1969 GNDA.n1631 GNDA.n1630 163.333
R1970 GNDA.n804 GNDA.n803 163.333
R1971 GNDA.n684 GNDA.n683 163.333
R1972 GNDA.n303 GNDA.n67 152
R1973 GNDA.n300 GNDA.n299 152
R1974 GNDA.n176 GNDA.n93 150
R1975 GNDA.n94 GNDA.n93 150
R1976 GNDA.n95 GNDA.n94 150
R1977 GNDA.n96 GNDA.n95 150
R1978 GNDA.n98 GNDA.n97 150
R1979 GNDA.n99 GNDA.n98 150
R1980 GNDA.n100 GNDA.n99 150
R1981 GNDA.n101 GNDA.n100 150
R1982 GNDA.n119 GNDA.n118 150
R1983 GNDA.n119 GNDA.n110 150
R1984 GNDA.n127 GNDA.n110 150
R1985 GNDA.n128 GNDA.n127 150
R1986 GNDA.n129 GNDA.n106 150
R1987 GNDA.n137 GNDA.n106 150
R1988 GNDA.n138 GNDA.n137 150
R1989 GNDA.n139 GNDA.n138 150
R1990 GNDA.n2538 GNDA.n2505 150
R1991 GNDA.n2506 GNDA.n2505 150
R1992 GNDA.n2507 GNDA.n2506 150
R1993 GNDA.n2508 GNDA.n2507 150
R1994 GNDA.n2510 GNDA.n2509 150
R1995 GNDA.n2511 GNDA.n2510 150
R1996 GNDA.n2512 GNDA.n2511 150
R1997 GNDA.n2513 GNDA.n2512 150
R1998 GNDA.n2498 GNDA.n2461 150
R1999 GNDA.n2462 GNDA.n2461 150
R2000 GNDA.n2463 GNDA.n2462 150
R2001 GNDA.n2464 GNDA.n2463 150
R2002 GNDA.n2466 GNDA.n2465 150
R2003 GNDA.n2467 GNDA.n2466 150
R2004 GNDA.n2468 GNDA.n2467 150
R2005 GNDA.n2469 GNDA.n2468 150
R2006 GNDA.n1481 GNDA.n1480 150
R2007 GNDA.n1477 GNDA.n1476 150
R2008 GNDA.n1473 GNDA.n1472 150
R2009 GNDA.n1469 GNDA.n1468 150
R2010 GNDA.n1465 GNDA.n1464 150
R2011 GNDA.n1461 GNDA.n1460 150
R2012 GNDA.n1457 GNDA.n1456 150
R2013 GNDA.n1453 GNDA.n1452 150
R2014 GNDA.n1510 GNDA.n1509 150
R2015 GNDA.n1502 GNDA.n1136 150
R2016 GNDA.n1434 GNDA.n1137 150
R2017 GNDA.n1441 GNDA.n1440 150
R2018 GNDA.n1499 GNDA.n1153 150
R2019 GNDA.n1495 GNDA.n1494 150
R2020 GNDA.n1491 GNDA.n1490 150
R2021 GNDA.n1487 GNDA.n1486 150
R2022 GNDA.n2282 GNDA.n2281 150
R2023 GNDA.n2278 GNDA.n2277 150
R2024 GNDA.n2274 GNDA.n2273 150
R2025 GNDA.n2270 GNDA.n2269 150
R2026 GNDA.n2266 GNDA.n2265 150
R2027 GNDA.n2262 GNDA.n2261 150
R2028 GNDA.n2258 GNDA.n2257 150
R2029 GNDA.n2254 GNDA.n2253 150
R2030 GNDA.n2316 GNDA.n2315 150
R2031 GNDA.n2303 GNDA.n2302 150
R2032 GNDA.n2305 GNDA.n2192 150
R2033 GNDA.n2238 GNDA.n2237 150
R2034 GNDA.n2300 GNDA.n2208 150
R2035 GNDA.n2296 GNDA.n2295 150
R2036 GNDA.n2292 GNDA.n2291 150
R2037 GNDA.n2288 GNDA.n2287 150
R2038 GNDA.n2098 GNDA.n2097 150
R2039 GNDA.n2094 GNDA.n2093 150
R2040 GNDA.n2090 GNDA.n2089 150
R2041 GNDA.n2086 GNDA.n2085 150
R2042 GNDA.n2082 GNDA.n2081 150
R2043 GNDA.n2078 GNDA.n2077 150
R2044 GNDA.n2074 GNDA.n2073 150
R2045 GNDA.n2070 GNDA.n2069 150
R2046 GNDA.n2121 GNDA.n497 150
R2047 GNDA.n551 GNDA.n498 150
R2048 GNDA.n548 GNDA.n547 150
R2049 GNDA.n540 GNDA.n539 150
R2050 GNDA.n2106 GNDA.n2105 150
R2051 GNDA.n2110 GNDA.n2109 150
R2052 GNDA.n2114 GNDA.n2113 150
R2053 GNDA.n2118 GNDA.n2117 150
R2054 GNDA.n1987 GNDA.n1986 150
R2055 GNDA.n1983 GNDA.n1982 150
R2056 GNDA.n1979 GNDA.n1978 150
R2057 GNDA.n1975 GNDA.n1974 150
R2058 GNDA.n1971 GNDA.n1970 150
R2059 GNDA.n1967 GNDA.n1966 150
R2060 GNDA.n1963 GNDA.n1962 150
R2061 GNDA.n1959 GNDA.n1958 150
R2062 GNDA.n2010 GNDA.n1015 150
R2063 GNDA.n1932 GNDA.n1016 150
R2064 GNDA.n1940 GNDA.n1939 150
R2065 GNDA.n1947 GNDA.n1946 150
R2066 GNDA.n1995 GNDA.n1994 150
R2067 GNDA.n1999 GNDA.n1998 150
R2068 GNDA.n2003 GNDA.n2002 150
R2069 GNDA.n2007 GNDA.n2006 150
R2070 GNDA.n1892 GNDA.n1891 150
R2071 GNDA.n1888 GNDA.n1887 150
R2072 GNDA.n1884 GNDA.n1883 150
R2073 GNDA.n1880 GNDA.n1879 150
R2074 GNDA.n1876 GNDA.n1875 150
R2075 GNDA.n1872 GNDA.n1871 150
R2076 GNDA.n1868 GNDA.n1867 150
R2077 GNDA.n1864 GNDA.n1863 150
R2078 GNDA.n1915 GNDA.n1036 150
R2079 GNDA.n1837 GNDA.n1037 150
R2080 GNDA.n1845 GNDA.n1844 150
R2081 GNDA.n1852 GNDA.n1851 150
R2082 GNDA.n1900 GNDA.n1899 150
R2083 GNDA.n1904 GNDA.n1903 150
R2084 GNDA.n1908 GNDA.n1907 150
R2085 GNDA.n1912 GNDA.n1911 150
R2086 GNDA.n1241 GNDA.n1240 150
R2087 GNDA.n1237 GNDA.n1236 150
R2088 GNDA.n1233 GNDA.n1232 150
R2089 GNDA.n1229 GNDA.n1228 150
R2090 GNDA.n1225 GNDA.n1224 150
R2091 GNDA.n1221 GNDA.n1220 150
R2092 GNDA.n1217 GNDA.n1216 150
R2093 GNDA.n1213 GNDA.n1212 150
R2094 GNDA.n1264 GNDA.n1160 150
R2095 GNDA.n1186 GNDA.n1161 150
R2096 GNDA.n1194 GNDA.n1193 150
R2097 GNDA.n1201 GNDA.n1200 150
R2098 GNDA.n1249 GNDA.n1248 150
R2099 GNDA.n1253 GNDA.n1252 150
R2100 GNDA.n1257 GNDA.n1256 150
R2101 GNDA.n1261 GNDA.n1260 150
R2102 GNDA.n1575 GNDA.n1573 150
R2103 GNDA.n1571 GNDA.n1539 150
R2104 GNDA.n1567 GNDA.n1565 150
R2105 GNDA.n1563 GNDA.n1541 150
R2106 GNDA.n1559 GNDA.n1557 150
R2107 GNDA.n1555 GNDA.n1543 150
R2108 GNDA.n1551 GNDA.n1550 150
R2109 GNDA.n1548 GNDA.n1546 150
R2110 GNDA.n1602 GNDA.n1600 150
R2111 GNDA.n1613 GNDA.n1527 150
R2112 GNDA.n1617 GNDA.n1615 150
R2113 GNDA.n1628 GNDA.n1522 150
R2114 GNDA.n1583 GNDA.n1581 150
R2115 GNDA.n1587 GNDA.n1535 150
R2116 GNDA.n1591 GNDA.n1589 150
R2117 GNDA.n1598 GNDA.n1533 150
R2118 GNDA.n836 GNDA.n835 150
R2119 GNDA.n832 GNDA.n831 150
R2120 GNDA.n828 GNDA.n827 150
R2121 GNDA.n824 GNDA.n823 150
R2122 GNDA.n820 GNDA.n819 150
R2123 GNDA.n816 GNDA.n815 150
R2124 GNDA.n812 GNDA.n811 150
R2125 GNDA.n808 GNDA.n807 150
R2126 GNDA.n871 GNDA.n870 150
R2127 GNDA.n858 GNDA.n857 150
R2128 GNDA.n860 GNDA.n759 150
R2129 GNDA.n792 GNDA.n791 150
R2130 GNDA.n855 GNDA.n775 150
R2131 GNDA.n851 GNDA.n850 150
R2132 GNDA.n847 GNDA.n846 150
R2133 GNDA.n843 GNDA.n842 150
R2134 GNDA.n716 GNDA.n715 150
R2135 GNDA.n712 GNDA.n711 150
R2136 GNDA.n708 GNDA.n707 150
R2137 GNDA.n704 GNDA.n703 150
R2138 GNDA.n700 GNDA.n699 150
R2139 GNDA.n696 GNDA.n695 150
R2140 GNDA.n692 GNDA.n691 150
R2141 GNDA.n688 GNDA.n687 150
R2142 GNDA.n2407 GNDA.n410 150
R2143 GNDA.n2397 GNDA.n2396 150
R2144 GNDA.n2410 GNDA.n391 150
R2145 GNDA.n673 GNDA.n392 150
R2146 GNDA.n724 GNDA.n723 150
R2147 GNDA.n728 GNDA.n727 150
R2148 GNDA.n732 GNDA.n731 150
R2149 GNDA.n734 GNDA.n409 150
R2150 GNDA.t116 GNDA.n337 148.466
R2151 GNDA.n337 GNDA.t36 148.466
R2152 GNDA.t308 GNDA.t64 147.84
R2153 GNDA.t13 GNDA.t126 144.321
R2154 GNDA.n2327 GNDA.n2326 139.077
R2155 GNDA.n2329 GNDA.n2328 139.077
R2156 GNDA.n2331 GNDA.n2330 139.077
R2157 GNDA.n2337 GNDA.n2336 139.077
R2158 GNDA.n2335 GNDA.n2334 139.077
R2159 GNDA.n2333 GNDA.n2332 139.077
R2160 GNDA.n416 GNDA.n415 139.077
R2161 GNDA.n2382 GNDA.n2381 139.077
R2162 GNDA.n2380 GNDA.n2379 139.077
R2163 GNDA.n376 GNDA.n375 139.077
R2164 GNDA.t33 GNDA.t151 139.041
R2165 GNDA.n2431 GNDA.t128 135.69
R2166 GNDA.n2218 GNDA.n2216 134.268
R2167 GNDA.n2226 GNDA.n2218 134.268
R2168 GNDA.n490 GNDA.n489 132.721
R2169 GNDA.n2436 GNDA.t264 130.001
R2170 GNDA.n2385 GNDA.t277 130.001
R2171 GNDA.n2376 GNDA.t255 130.001
R2172 GNDA.n2338 GNDA.t290 130.001
R2173 GNDA.n2343 GNDA.t216 130.001
R2174 GNDA.n2324 GNDA.t274 130.001
R2175 GNDA.n885 GNDA.n883 124.832
R2176 GNDA.n881 GNDA.n606 124.832
R2177 GNDA.n743 GNDA.n467 124.832
R2178 GNDA.n1425 GNDA.n1424 124.832
R2179 GNDA.n2347 GNDA.n2346 124.832
R2180 GNDA.n1010 GNDA.n557 124.832
R2181 GNDA.n2057 GNDA.n2056 124.832
R2182 GNDA.n2021 GNDA.n556 124.832
R2183 GNDA.n2050 GNDA.n558 124.832
R2184 GNDA.n1720 GNDA.n1719 124.832
R2185 GNDA.n1422 GNDA.n1273 124.832
R2186 GNDA.n1717 GNDA.n1066 124.832
R2187 GNDA.n378 GNDA.t34 115.948
R2188 GNDA.n1298 GNDA.t103 115.105
R2189 GNDA.n378 GNDA.t14 114.635
R2190 GNDA.n1299 GNDA.t97 114.635
R2191 GNDA.n277 GNDA.t211 103.665
R2192 GNDA.t222 GNDA.n17 103.665
R2193 GNDA.t254 GNDA.n417 101.942
R2194 GNDA.n2415 GNDA.n384 101.718
R2195 GNDA.n357 GNDA.n38 101.718
R2196 GNDA.n348 GNDA.n55 101.718
R2197 GNDA.n2451 GNDA.n31 101.718
R2198 GNDA.n2547 GNDA.n18 101.718
R2199 GNDA.n203 GNDA.n72 101.718
R2200 GNDA.n185 GNDA.n83 101.718
R2201 GNDA.n2495 GNDA.n25 101.718
R2202 GNDA.n2492 GNDA.n26 101.718
R2203 GNDA.n2488 GNDA.n27 101.718
R2204 GNDA.n2484 GNDA.n28 101.718
R2205 GNDA.n2480 GNDA.n29 101.718
R2206 GNDA.n2535 GNDA.n19 101.718
R2207 GNDA.n2532 GNDA.n20 101.718
R2208 GNDA.n2528 GNDA.n21 101.718
R2209 GNDA.n2524 GNDA.n22 101.718
R2210 GNDA.n2520 GNDA.n23 101.718
R2211 GNDA.n122 GNDA.n121 101.718
R2212 GNDA.n125 GNDA.n124 101.718
R2213 GNDA.n132 GNDA.n131 101.718
R2214 GNDA.n135 GNDA.n134 101.718
R2215 GNDA.n142 GNDA.n141 101.718
R2216 GNDA.n231 GNDA.n220 101.718
R2217 GNDA.n260 GNDA.n214 101.718
R2218 GNDA.n173 GNDA.n84 101.718
R2219 GNDA.n170 GNDA.n85 101.718
R2220 GNDA.n166 GNDA.n86 101.718
R2221 GNDA.n162 GNDA.n87 101.718
R2222 GNDA.n158 GNDA.n88 101.718
R2223 GNDA.n178 GNDA.n91 101.718
R2224 GNDA.n171 GNDA.n84 101.718
R2225 GNDA.n167 GNDA.n85 101.718
R2226 GNDA.n163 GNDA.n86 101.718
R2227 GNDA.n159 GNDA.n87 101.718
R2228 GNDA.n155 GNDA.n88 101.718
R2229 GNDA.n266 GNDA.n216 101.718
R2230 GNDA.n229 GNDA.n222 101.718
R2231 GNDA.n115 GNDA.n114 101.718
R2232 GNDA.n123 GNDA.n122 101.718
R2233 GNDA.n124 GNDA.n108 101.718
R2234 GNDA.n133 GNDA.n132 101.718
R2235 GNDA.n134 GNDA.n104 101.718
R2236 GNDA.n143 GNDA.n142 101.718
R2237 GNDA.n2540 GNDA.n2503 101.718
R2238 GNDA.n2533 GNDA.n19 101.718
R2239 GNDA.n2529 GNDA.n20 101.718
R2240 GNDA.n2525 GNDA.n21 101.718
R2241 GNDA.n2521 GNDA.n22 101.718
R2242 GNDA.n2517 GNDA.n23 101.718
R2243 GNDA.n2500 GNDA.n2459 101.718
R2244 GNDA.n2493 GNDA.n25 101.718
R2245 GNDA.n2489 GNDA.n26 101.718
R2246 GNDA.n2485 GNDA.n27 101.718
R2247 GNDA.n2481 GNDA.n28 101.718
R2248 GNDA.n2477 GNDA.n29 101.718
R2249 GNDA.n190 GNDA.n181 101.718
R2250 GNDA.n83 GNDA.n79 101.718
R2251 GNDA.n213 GNDA.n70 101.718
R2252 GNDA.n65 GNDA.n64 101.718
R2253 GNDA.n292 GNDA.n56 101.718
R2254 GNDA.n287 GNDA.n286 101.718
R2255 GNDA.n208 GNDA.n75 101.718
R2256 GNDA.n201 GNDA.n72 101.718
R2257 GNDA.n276 GNDA.n269 101.718
R2258 GNDA.n314 GNDA.n63 101.718
R2259 GNDA.n335 GNDA.n59 101.718
R2260 GNDA.n2552 GNDA.n2543 101.718
R2261 GNDA.n18 GNDA.n16 101.718
R2262 GNDA.n2456 GNDA.n2444 101.718
R2263 GNDA.n2449 GNDA.n31 101.718
R2264 GNDA.n325 GNDA.n324 101.718
R2265 GNDA.n346 GNDA.n339 101.718
R2266 GNDA.n363 GNDA.n40 101.718
R2267 GNDA.n2426 GNDA.n383 101.718
R2268 GNDA.n2215 GNDA.n2213 101.718
R2269 GNDA.n2222 GNDA.n2214 101.718
R2270 GNDA.n2221 GNDA.n2213 101.718
R2271 GNDA.n2048 GNDA.t209 47.6748
R2272 GNDA.n2374 GNDA.t209 47.6748
R2273 GNDA.n255 GNDA.n254 99.0842
R2274 GNDA.n253 GNDA.n252 99.0842
R2275 GNDA.n251 GNDA.n250 99.0842
R2276 GNDA.n249 GNDA.n248 99.0842
R2277 GNDA.n247 GNDA.n246 99.0842
R2278 GNDA.n245 GNDA.n244 99.0842
R2279 GNDA.n243 GNDA.n242 99.0842
R2280 GNDA.n241 GNDA.n240 99.0842
R2281 GNDA.n239 GNDA.n238 99.0842
R2282 GNDA.n237 GNDA.n236 99.0842
R2283 GNDA.n235 GNDA.n234 99.0842
R2284 GNDA.n353 GNDA.n352 99.0842
R2285 GNDA.n644 GNDA.t209 98.9756
R2286 GNDA.n745 GNDA.n744 98.8538
R2287 GNDA.n151 GNDA.n150 94.601
R2288 GNDA.n149 GNDA.n148 94.601
R2289 GNDA.n2471 GNDA.n2470 94.601
R2290 GNDA.n2473 GNDA.n2472 94.601
R2291 GNDA.n2388 GNDA.n2387 92.6754
R2292 GNDA.t92 GNDA.t31 92.1471
R2293 GNDA.t300 GNDA.t92 92.1471
R2294 GNDA.t313 GNDA.t300 92.1471
R2295 GNDA.t38 GNDA.t119 92.1471
R2296 GNDA.n2422 GNDA.n382 91.069
R2297 GNDA.n2417 GNDA.n382 91.069
R2298 GNDA.n2419 GNDA.n381 91.069
R2299 GNDA.n2420 GNDA.n2419 91.069
R2300 GNDA.n308 GNDA.n307 91.069
R2301 GNDA.n305 GNDA.n66 91.069
R2302 GNDA.n297 GNDA.n296 91.069
R2303 GNDA.n294 GNDA.n291 91.069
R2304 GNDA.n2224 GNDA.n2216 91.069
R2305 GNDA.n2226 GNDA.n2219 91.069
R2306 GNDA.t215 GNDA.n2244 90.616
R2307 GNDA.n210 GNDA.n69 90.4158
R2308 GNDA.n263 GNDA.n217 90.2704
R2309 GNDA.n259 GNDA.n217 90.2704
R2310 GNDA.n226 GNDA.n223 90.2704
R2311 GNDA.n223 GNDA.n219 90.2704
R2312 GNDA.n284 GNDA.n282 90.2704
R2313 GNDA.n273 GNDA.n270 90.2704
R2314 GNDA.n311 GNDA.n62 90.2704
R2315 GNDA.n332 GNDA.n60 90.2704
R2316 GNDA.n322 GNDA.n320 90.2704
R2317 GNDA.n343 GNDA.n340 90.2704
R2318 GNDA.n340 GNDA.n54 90.2704
R2319 GNDA.n360 GNDA.n41 90.2704
R2320 GNDA.n356 GNDA.n41 90.2704
R2321 GNDA.n1801 GNDA.t2 89.6052
R2322 GNDA.n1370 GNDA.n1344 88.5317
R2323 GNDA.n1371 GNDA.n1370 88.5317
R2324 GNDA.n1372 GNDA.n1371 88.5317
R2325 GNDA.n1372 GNDA.n1340 88.5317
R2326 GNDA.n1378 GNDA.n1340 88.5317
R2327 GNDA.n1380 GNDA.n1379 88.5317
R2328 GNDA.n1380 GNDA.n1336 88.5317
R2329 GNDA.n1387 GNDA.n1336 88.5317
R2330 GNDA.n1388 GNDA.n1387 88.5317
R2331 GNDA.n1389 GNDA.n1388 88.5317
R2332 GNDA.n1329 GNDA.n1291 88.5317
R2333 GNDA.n1329 GNDA.n1328 88.5317
R2334 GNDA.n1328 GNDA.n1327 88.5317
R2335 GNDA.n1327 GNDA.n1292 88.5317
R2336 GNDA.n1321 GNDA.n1292 88.5317
R2337 GNDA.n1320 GNDA.n1319 88.5317
R2338 GNDA.n1319 GNDA.n1304 88.5317
R2339 GNDA.n1313 GNDA.n1304 88.5317
R2340 GNDA.n1313 GNDA.n1312 88.5317
R2341 GNDA.n1312 GNDA.n1088 88.5317
R2342 GNDA.n1688 GNDA.n1687 88.5317
R2343 GNDA.n1687 GNDA.n1089 88.5317
R2344 GNDA.n1681 GNDA.n1089 88.5317
R2345 GNDA.n1681 GNDA.n1680 88.5317
R2346 GNDA.n1680 GNDA.n1679 88.5317
R2347 GNDA.n1673 GNDA.n1097 88.5317
R2348 GNDA.n1673 GNDA.n1672 88.5317
R2349 GNDA.n1672 GNDA.n1671 88.5317
R2350 GNDA.n1671 GNDA.n1098 88.5317
R2351 GNDA.n1665 GNDA.n1098 88.5317
R2352 GNDA.n191 GNDA.t38 88.3077
R2353 GNDA.t85 GNDA.n2438 85.4674
R2354 GNDA.t101 GNDA.t47 84.4682
R2355 GNDA.t62 GNDA.t89 84.4682
R2356 GNDA.t99 GNDA.t60 84.4682
R2357 GNDA.t95 GNDA.t48 84.4682
R2358 GNDA.t94 GNDA.t30 84.4682
R2359 GNDA.t211 GNDA.t87 84.4682
R2360 GNDA.t87 GNDA.t3 84.4682
R2361 GNDA.t3 GNDA.t68 84.4682
R2362 GNDA.t40 GNDA.t73 84.4682
R2363 GNDA.t149 GNDA.t130 84.4682
R2364 GNDA.t130 GNDA.t222 84.4682
R2365 GNDA.t113 GNDA.t136 84.4682
R2366 GNDA.t134 GNDA.t54 84.4682
R2367 GNDA.t76 GNDA.t133 84.4682
R2368 GNDA.t114 GNDA.t51 84.4682
R2369 GNDA.t298 GNDA.t299 84.4682
R2370 GNDA.n865 GNDA.t180 84.4377
R2371 GNDA.n1297 GNDA.n1296 84.306
R2372 GNDA.t12 GNDA.t139 82.3782
R2373 GNDA.t96 GNDA.t127 82.3782
R2374 GNDA.n1690 GNDA.n1689 80.9821
R2375 GNDA.t233 GNDA.t280 80.6288
R2376 GNDA.t270 GNDA.t257 80.6288
R2377 GNDA.t206 GNDA.t260 80.6288
R2378 GNDA.t247 GNDA.t227 80.6288
R2379 GNDA.n796 GNDA.t170 80.3188
R2380 GNDA.t106 GNDA.t251 76.7893
R2381 GNDA.t110 GNDA.t35 76.7893
R2382 GNDA.t304 GNDA.t283 76.7893
R2383 GNDA.n623 GNDA.n422 76.3222
R2384 GNDA.n627 GNDA.n423 76.3222
R2385 GNDA.n631 GNDA.n424 76.3222
R2386 GNDA.n635 GNDA.n425 76.3222
R2387 GNDA.n639 GNDA.n426 76.3222
R2388 GNDA.n643 GNDA.n427 76.3222
R2389 GNDA.n906 GNDA.n905 76.3222
R2390 GNDA.n903 GNDA.n585 76.3222
R2391 GNDA.n899 GNDA.n898 76.3222
R2392 GNDA.n892 GNDA.n592 76.3222
R2393 GNDA.n891 GNDA.n890 76.3222
R2394 GNDA.n884 GNDA.n600 76.3222
R2395 GNDA.n587 GNDA.n586 76.3222
R2396 GNDA.n590 GNDA.n589 76.3222
R2397 GNDA.n595 GNDA.n594 76.3222
R2398 GNDA.n598 GNDA.n597 76.3222
R2399 GNDA.n603 GNDA.n602 76.3222
R2400 GNDA.n606 GNDA.n605 76.3222
R2401 GNDA.n561 GNDA.n428 76.3222
R2402 GNDA.n565 GNDA.n429 76.3222
R2403 GNDA.n569 GNDA.n430 76.3222
R2404 GNDA.n573 GNDA.n431 76.3222
R2405 GNDA.n577 GNDA.n432 76.3222
R2406 GNDA.n581 GNDA.n433 76.3222
R2407 GNDA.n2368 GNDA.n2367 76.3222
R2408 GNDA.n2365 GNDA.n446 76.3222
R2409 GNDA.n2361 GNDA.n2360 76.3222
R2410 GNDA.n2354 GNDA.n453 76.3222
R2411 GNDA.n2353 GNDA.n2352 76.3222
R2412 GNDA.n466 GNDA.n461 76.3222
R2413 GNDA.n1286 GNDA.n1279 76.3222
R2414 GNDA.n1400 GNDA.n1280 76.3222
R2415 GNDA.n1282 GNDA.n1281 76.3222
R2416 GNDA.n1410 GNDA.n1278 76.3222
R2417 GNDA.n1414 GNDA.n1413 76.3222
R2418 GNDA.n1424 GNDA.n1155 76.3222
R2419 GNDA.n1516 GNDA.n1515 76.3222
R2420 GNDA.n1130 GNDA.n1124 76.3222
R2421 GNDA.n1505 GNDA.n1123 76.3222
R2422 GNDA.n1432 GNDA.n1122 76.3222
R2423 GNDA.n1436 GNDA.n1121 76.3222
R2424 GNDA.n1445 GNDA.n1120 76.3222
R2425 GNDA.n1365 GNDA.n477 76.3222
R2426 GNDA.n1362 GNDA.n478 76.3222
R2427 GNDA.n1358 GNDA.n479 76.3222
R2428 GNDA.n1354 GNDA.n480 76.3222
R2429 GNDA.n1350 GNDA.n481 76.3222
R2430 GNDA.n448 GNDA.n447 76.3222
R2431 GNDA.n451 GNDA.n450 76.3222
R2432 GNDA.n456 GNDA.n455 76.3222
R2433 GNDA.n459 GNDA.n458 76.3222
R2434 GNDA.n464 GNDA.n463 76.3222
R2435 GNDA.n2347 GNDA.n469 76.3222
R2436 GNDA.n2153 GNDA.n434 76.3222
R2437 GNDA.n2149 GNDA.n435 76.3222
R2438 GNDA.n2145 GNDA.n436 76.3222
R2439 GNDA.n2141 GNDA.n437 76.3222
R2440 GNDA.n2137 GNDA.n438 76.3222
R2441 GNDA.n2373 GNDA.n2372 76.3222
R2442 GNDA.n2175 GNDA.n2174 76.3222
R2443 GNDA.n2170 GNDA.n2134 76.3222
R2444 GNDA.n2167 GNDA.n2133 76.3222
R2445 GNDA.n2163 GNDA.n2132 76.3222
R2446 GNDA.n2159 GNDA.n2131 76.3222
R2447 GNDA.n2175 GNDA.n2135 76.3222
R2448 GNDA.n2168 GNDA.n2134 76.3222
R2449 GNDA.n2164 GNDA.n2133 76.3222
R2450 GNDA.n2160 GNDA.n2132 76.3222
R2451 GNDA.n2156 GNDA.n2131 76.3222
R2452 GNDA.n1363 GNDA.n477 76.3222
R2453 GNDA.n1359 GNDA.n478 76.3222
R2454 GNDA.n1355 GNDA.n479 76.3222
R2455 GNDA.n1351 GNDA.n480 76.3222
R2456 GNDA.n1347 GNDA.n481 76.3222
R2457 GNDA.n991 GNDA.n990 76.3222
R2458 GNDA.n994 GNDA.n993 76.3222
R2459 GNDA.n999 GNDA.n998 76.3222
R2460 GNDA.n1002 GNDA.n1001 76.3222
R2461 GNDA.n1007 GNDA.n1006 76.3222
R2462 GNDA.n1010 GNDA.n1009 76.3222
R2463 GNDA.n967 GNDA.n935 76.3222
R2464 GNDA.n971 GNDA.n936 76.3222
R2465 GNDA.n975 GNDA.n937 76.3222
R2466 GNDA.n979 GNDA.n938 76.3222
R2467 GNDA.n982 GNDA.n939 76.3222
R2468 GNDA.n2047 GNDA.n2046 76.3222
R2469 GNDA.n2129 GNDA.n491 76.3222
R2470 GNDA.n2124 GNDA.n495 76.3222
R2471 GNDA.n555 GNDA.n554 76.3222
R2472 GNDA.n536 GNDA.n532 76.3222
R2473 GNDA.n543 GNDA.n531 76.3222
R2474 GNDA.n2062 GNDA.n2061 76.3222
R2475 GNDA.n963 GNDA.n484 76.3222
R2476 GNDA.n959 GNDA.n485 76.3222
R2477 GNDA.n955 GNDA.n486 76.3222
R2478 GNDA.n951 GNDA.n487 76.3222
R2479 GNDA.n947 GNDA.n488 76.3222
R2480 GNDA.n943 GNDA.n489 76.3222
R2481 GNDA.n960 GNDA.n484 76.3222
R2482 GNDA.n956 GNDA.n485 76.3222
R2483 GNDA.n952 GNDA.n486 76.3222
R2484 GNDA.n948 GNDA.n487 76.3222
R2485 GNDA.n944 GNDA.n488 76.3222
R2486 GNDA.n1780 GNDA.n923 76.3222
R2487 GNDA.n1784 GNDA.n924 76.3222
R2488 GNDA.n1788 GNDA.n925 76.3222
R2489 GNDA.n1792 GNDA.n926 76.3222
R2490 GNDA.n1796 GNDA.n927 76.3222
R2491 GNDA.n1800 GNDA.n928 76.3222
R2492 GNDA.n910 GNDA.n524 76.3222
R2493 GNDA.n1918 GNDA.n523 76.3222
R2494 GNDA.n1835 GNDA.n522 76.3222
R2495 GNDA.n1841 GNDA.n521 76.3222
R2496 GNDA.n1847 GNDA.n520 76.3222
R2497 GNDA.n1856 GNDA.n519 76.3222
R2498 GNDA.n1776 GNDA.n1723 76.3222
R2499 GNDA.n1772 GNDA.n1771 76.3222
R2500 GNDA.n1765 GNDA.n1750 76.3222
R2501 GNDA.n1764 GNDA.n1763 76.3222
R2502 GNDA.n1757 GNDA.n1756 76.3222
R2503 GNDA.n2055 GNDA.n2054 76.3222
R2504 GNDA.n2042 GNDA.n2041 76.3222
R2505 GNDA.n2039 GNDA.n989 76.3222
R2506 GNDA.n2035 GNDA.n2034 76.3222
R2507 GNDA.n2028 GNDA.n996 76.3222
R2508 GNDA.n2027 GNDA.n2026 76.3222
R2509 GNDA.n2020 GNDA.n1004 76.3222
R2510 GNDA.n1725 GNDA.n929 76.3222
R2511 GNDA.n1729 GNDA.n930 76.3222
R2512 GNDA.n1733 GNDA.n931 76.3222
R2513 GNDA.n1737 GNDA.n932 76.3222
R2514 GNDA.n1741 GNDA.n933 76.3222
R2515 GNDA.n1745 GNDA.n934 76.3222
R2516 GNDA.n2017 GNDA.n530 76.3222
R2517 GNDA.n2013 GNDA.n529 76.3222
R2518 GNDA.n1930 GNDA.n528 76.3222
R2519 GNDA.n1936 GNDA.n527 76.3222
R2520 GNDA.n1942 GNDA.n526 76.3222
R2521 GNDA.n1951 GNDA.n525 76.3222
R2522 GNDA.n1747 GNDA.n916 76.3222
R2523 GNDA.n1751 GNDA.n917 76.3222
R2524 GNDA.n1753 GNDA.n918 76.3222
R2525 GNDA.n1758 GNDA.n919 76.3222
R2526 GNDA.n920 GNDA.n915 76.3222
R2527 GNDA.n2051 GNDA.n2050 76.3222
R2528 GNDA.n1530 GNDA.n1068 76.3222
R2529 GNDA.n1606 GNDA.n1605 76.3222
R2530 GNDA.n1609 GNDA.n1608 76.3222
R2531 GNDA.n1621 GNDA.n1620 76.3222
R2532 GNDA.n1624 GNDA.n1623 76.3222
R2533 GNDA.n1636 GNDA.n1635 76.3222
R2534 GNDA.n1394 GNDA.n1393 76.3222
R2535 GNDA.n1397 GNDA.n1396 76.3222
R2536 GNDA.n1404 GNDA.n1403 76.3222
R2537 GNDA.n1407 GNDA.n1406 76.3222
R2538 GNDA.n1418 GNDA.n1417 76.3222
R2539 GNDA.n1421 GNDA.n1420 76.3222
R2540 GNDA.n1272 GNDA.n1119 76.3222
R2541 GNDA.n1267 GNDA.n1118 76.3222
R2542 GNDA.n1184 GNDA.n1117 76.3222
R2543 GNDA.n1190 GNDA.n1116 76.3222
R2544 GNDA.n1196 GNDA.n1115 76.3222
R2545 GNDA.n1205 GNDA.n1114 76.3222
R2546 GNDA.n2052 GNDA.n2051 76.3222
R2547 GNDA.n1759 GNDA.n920 76.3222
R2548 GNDA.n1754 GNDA.n919 76.3222
R2549 GNDA.n1752 GNDA.n918 76.3222
R2550 GNDA.n1748 GNDA.n917 76.3222
R2551 GNDA.n1746 GNDA.n916 76.3222
R2552 GNDA.n1773 GNDA.n1723 76.3222
R2553 GNDA.n1771 GNDA.n1770 76.3222
R2554 GNDA.n1766 GNDA.n1765 76.3222
R2555 GNDA.n1763 GNDA.n1762 76.3222
R2556 GNDA.n1756 GNDA.n913 76.3222
R2557 GNDA.n2056 GNDA.n2055 76.3222
R2558 GNDA.n2047 GNDA.n940 76.3222
R2559 GNDA.n980 GNDA.n939 76.3222
R2560 GNDA.n976 GNDA.n938 76.3222
R2561 GNDA.n972 GNDA.n937 76.3222
R2562 GNDA.n968 GNDA.n936 76.3222
R2563 GNDA.n964 GNDA.n935 76.3222
R2564 GNDA.n1742 GNDA.n934 76.3222
R2565 GNDA.n1738 GNDA.n933 76.3222
R2566 GNDA.n1734 GNDA.n932 76.3222
R2567 GNDA.n1730 GNDA.n931 76.3222
R2568 GNDA.n1726 GNDA.n930 76.3222
R2569 GNDA.n988 GNDA.n929 76.3222
R2570 GNDA.n1797 GNDA.n928 76.3222
R2571 GNDA.n1793 GNDA.n927 76.3222
R2572 GNDA.n1789 GNDA.n926 76.3222
R2573 GNDA.n1785 GNDA.n925 76.3222
R2574 GNDA.n1781 GNDA.n924 76.3222
R2575 GNDA.n1777 GNDA.n923 76.3222
R2576 GNDA.n1516 GNDA.n1125 76.3222
R2577 GNDA.n1506 GNDA.n1124 76.3222
R2578 GNDA.n1431 GNDA.n1123 76.3222
R2579 GNDA.n1437 GNDA.n1122 76.3222
R2580 GNDA.n1444 GNDA.n1121 76.3222
R2581 GNDA.n1426 GNDA.n1120 76.3222
R2582 GNDA.n1268 GNDA.n1119 76.3222
R2583 GNDA.n1183 GNDA.n1118 76.3222
R2584 GNDA.n1189 GNDA.n1117 76.3222
R2585 GNDA.n1197 GNDA.n1116 76.3222
R2586 GNDA.n1204 GNDA.n1115 76.3222
R2587 GNDA.n1178 GNDA.n1114 76.3222
R2588 GNDA.n1531 GNDA.n1530 76.3222
R2589 GNDA.n1607 GNDA.n1606 76.3222
R2590 GNDA.n1608 GNDA.n1525 76.3222
R2591 GNDA.n1622 GNDA.n1621 76.3222
R2592 GNDA.n1623 GNDA.n1518 76.3222
R2593 GNDA.n1637 GNDA.n1636 76.3222
R2594 GNDA.n1412 GNDA.n1155 76.3222
R2595 GNDA.n1415 GNDA.n1414 76.3222
R2596 GNDA.n1410 GNDA.n1409 76.3222
R2597 GNDA.n1401 GNDA.n1281 76.3222
R2598 GNDA.n1287 GNDA.n1280 76.3222
R2599 GNDA.n1391 GNDA.n1279 76.3222
R2600 GNDA.n1395 GNDA.n1394 76.3222
R2601 GNDA.n1396 GNDA.n1284 76.3222
R2602 GNDA.n1405 GNDA.n1404 76.3222
R2603 GNDA.n1406 GNDA.n1276 76.3222
R2604 GNDA.n1419 GNDA.n1418 76.3222
R2605 GNDA.n1422 GNDA.n1421 76.3222
R2606 GNDA.n1009 GNDA.n1008 76.3222
R2607 GNDA.n1006 GNDA.n1005 76.3222
R2608 GNDA.n1001 GNDA.n1000 76.3222
R2609 GNDA.n998 GNDA.n997 76.3222
R2610 GNDA.n993 GNDA.n992 76.3222
R2611 GNDA.n990 GNDA.n941 76.3222
R2612 GNDA.n2041 GNDA.n2040 76.3222
R2613 GNDA.n2036 GNDA.n989 76.3222
R2614 GNDA.n2034 GNDA.n2033 76.3222
R2615 GNDA.n2029 GNDA.n2028 76.3222
R2616 GNDA.n2026 GNDA.n2025 76.3222
R2617 GNDA.n2021 GNDA.n2020 76.3222
R2618 GNDA.n469 GNDA.n465 76.3222
R2619 GNDA.n463 GNDA.n462 76.3222
R2620 GNDA.n458 GNDA.n457 76.3222
R2621 GNDA.n455 GNDA.n454 76.3222
R2622 GNDA.n450 GNDA.n449 76.3222
R2623 GNDA.n447 GNDA.n440 76.3222
R2624 GNDA.n2367 GNDA.n2366 76.3222
R2625 GNDA.n2362 GNDA.n446 76.3222
R2626 GNDA.n2360 GNDA.n2359 76.3222
R2627 GNDA.n2355 GNDA.n2354 76.3222
R2628 GNDA.n2352 GNDA.n2351 76.3222
R2629 GNDA.n467 GNDA.n466 76.3222
R2630 GNDA.n605 GNDA.n604 76.3222
R2631 GNDA.n602 GNDA.n601 76.3222
R2632 GNDA.n597 GNDA.n596 76.3222
R2633 GNDA.n594 GNDA.n593 76.3222
R2634 GNDA.n589 GNDA.n588 76.3222
R2635 GNDA.n586 GNDA.n582 76.3222
R2636 GNDA.n905 GNDA.n904 76.3222
R2637 GNDA.n900 GNDA.n585 76.3222
R2638 GNDA.n898 GNDA.n897 76.3222
R2639 GNDA.n893 GNDA.n892 76.3222
R2640 GNDA.n890 GNDA.n889 76.3222
R2641 GNDA.n885 GNDA.n884 76.3222
R2642 GNDA.n2373 GNDA.n439 76.3222
R2643 GNDA.n2140 GNDA.n438 76.3222
R2644 GNDA.n2144 GNDA.n437 76.3222
R2645 GNDA.n2148 GNDA.n436 76.3222
R2646 GNDA.n2152 GNDA.n435 76.3222
R2647 GNDA.n2136 GNDA.n434 76.3222
R2648 GNDA.n578 GNDA.n433 76.3222
R2649 GNDA.n574 GNDA.n432 76.3222
R2650 GNDA.n570 GNDA.n431 76.3222
R2651 GNDA.n566 GNDA.n430 76.3222
R2652 GNDA.n562 GNDA.n429 76.3222
R2653 GNDA.n445 GNDA.n428 76.3222
R2654 GNDA.n640 GNDA.n427 76.3222
R2655 GNDA.n636 GNDA.n426 76.3222
R2656 GNDA.n632 GNDA.n425 76.3222
R2657 GNDA.n628 GNDA.n424 76.3222
R2658 GNDA.n624 GNDA.n423 76.3222
R2659 GNDA.n584 GNDA.n422 76.3222
R2660 GNDA.n2125 GNDA.n491 76.3222
R2661 GNDA.n534 GNDA.n495 76.3222
R2662 GNDA.n555 GNDA.n533 76.3222
R2663 GNDA.n544 GNDA.n532 76.3222
R2664 GNDA.n531 GNDA.n517 76.3222
R2665 GNDA.n2061 GNDA.n518 76.3222
R2666 GNDA.n2014 GNDA.n530 76.3222
R2667 GNDA.n1929 GNDA.n529 76.3222
R2668 GNDA.n1935 GNDA.n528 76.3222
R2669 GNDA.n1943 GNDA.n527 76.3222
R2670 GNDA.n1950 GNDA.n526 76.3222
R2671 GNDA.n1924 GNDA.n525 76.3222
R2672 GNDA.n1919 GNDA.n524 76.3222
R2673 GNDA.n1834 GNDA.n523 76.3222
R2674 GNDA.n1840 GNDA.n522 76.3222
R2675 GNDA.n1848 GNDA.n521 76.3222
R2676 GNDA.n1855 GNDA.n520 76.3222
R2677 GNDA.n1829 GNDA.n519 76.3222
R2678 GNDA.t281 GNDA.n96 75.0005
R2679 GNDA.n97 GNDA.t281 75.0005
R2680 GNDA.t271 GNDA.n128 75.0005
R2681 GNDA.n129 GNDA.t271 75.0005
R2682 GNDA.n206 GNDA.t258 75.0005
R2683 GNDA.n77 GNDA.t258 75.0005
R2684 GNDA.n188 GNDA.t234 75.0005
R2685 GNDA.n183 GNDA.t234 75.0005
R2686 GNDA.n2550 GNDA.t207 75.0005
R2687 GNDA.n2545 GNDA.t207 75.0005
R2688 GNDA.n2454 GNDA.t228 75.0005
R2689 GNDA.n2446 GNDA.t228 75.0005
R2690 GNDA.t261 GNDA.n2508 75.0005
R2691 GNDA.n2509 GNDA.t261 75.0005
R2692 GNDA.t248 GNDA.n2464 75.0005
R2693 GNDA.n2465 GNDA.t248 75.0005
R2694 GNDA.n1468 GNDA.n1142 74.5978
R2695 GNDA.n1465 GNDA.n1142 74.5978
R2696 GNDA.n2269 GNDA.n2197 74.5978
R2697 GNDA.n2266 GNDA.n2197 74.5978
R2698 GNDA.n2085 GNDA.n504 74.5978
R2699 GNDA.n2082 GNDA.n504 74.5978
R2700 GNDA.n1974 GNDA.n1022 74.5978
R2701 GNDA.n1971 GNDA.n1022 74.5978
R2702 GNDA.n1879 GNDA.n1043 74.5978
R2703 GNDA.n1876 GNDA.n1043 74.5978
R2704 GNDA.n1228 GNDA.n1167 74.5978
R2705 GNDA.n1225 GNDA.n1167 74.5978
R2706 GNDA.n1558 GNDA.n1541 74.5978
R2707 GNDA.n1559 GNDA.n1558 74.5978
R2708 GNDA.n823 GNDA.n764 74.5978
R2709 GNDA.n820 GNDA.n764 74.5978
R2710 GNDA.n703 GNDA.n398 74.5978
R2711 GNDA.n700 GNDA.n398 74.5978
R2712 GNDA.n798 GNDA.t186 74.1404
R2713 GNDA.n336 GNDA.t81 72.9499
R2714 GNDA.n230 GNDA.t0 72.9499
R2715 GNDA.n755 GNDA.t182 70.0216
R2716 GNDA.n1510 GNDA.n1132 69.3109
R2717 GNDA.n1486 GNDA.n1132 69.3109
R2718 GNDA.n2316 GNDA.n2182 69.3109
R2719 GNDA.n2287 GNDA.n2182 69.3109
R2720 GNDA.n2119 GNDA.n497 69.3109
R2721 GNDA.n2119 GNDA.n2118 69.3109
R2722 GNDA.n2008 GNDA.n1015 69.3109
R2723 GNDA.n2008 GNDA.n2007 69.3109
R2724 GNDA.n1913 GNDA.n1036 69.3109
R2725 GNDA.n1913 GNDA.n1912 69.3109
R2726 GNDA.n1262 GNDA.n1160 69.3109
R2727 GNDA.n1262 GNDA.n1261 69.3109
R2728 GNDA.n1600 GNDA.n1599 69.3109
R2729 GNDA.n1599 GNDA.n1598 69.3109
R2730 GNDA.n871 GNDA.n751 69.3109
R2731 GNDA.n842 GNDA.n751 69.3109
R2732 GNDA.n2408 GNDA.n2407 69.3109
R2733 GNDA.n2408 GNDA.n409 69.3109
R2734 GNDA.t245 GNDA.n1500 65.8183
R2735 GNDA.t245 GNDA.n1151 65.8183
R2736 GNDA.t245 GNDA.n1150 65.8183
R2737 GNDA.t245 GNDA.n1149 65.8183
R2738 GNDA.t245 GNDA.n1140 65.8183
R2739 GNDA.t245 GNDA.n1147 65.8183
R2740 GNDA.t245 GNDA.n1138 65.8183
R2741 GNDA.t245 GNDA.n1148 65.8183
R2742 GNDA.t245 GNDA.n1146 65.8183
R2743 GNDA.t245 GNDA.n1145 65.8183
R2744 GNDA.t245 GNDA.n1144 65.8183
R2745 GNDA.t245 GNDA.n1143 65.8183
R2746 GNDA.t245 GNDA.n1141 65.8183
R2747 GNDA.t245 GNDA.n1139 65.8183
R2748 GNDA.n1501 GNDA.t245 65.8183
R2749 GNDA.t245 GNDA.n1133 65.8183
R2750 GNDA.t268 GNDA.n2301 65.8183
R2751 GNDA.t268 GNDA.n2206 65.8183
R2752 GNDA.t268 GNDA.n2205 65.8183
R2753 GNDA.t268 GNDA.n2204 65.8183
R2754 GNDA.t268 GNDA.n2195 65.8183
R2755 GNDA.t268 GNDA.n2202 65.8183
R2756 GNDA.t268 GNDA.n2193 65.8183
R2757 GNDA.t268 GNDA.n2203 65.8183
R2758 GNDA.t268 GNDA.n2201 65.8183
R2759 GNDA.t268 GNDA.n2200 65.8183
R2760 GNDA.t268 GNDA.n2199 65.8183
R2761 GNDA.t268 GNDA.n2198 65.8183
R2762 GNDA.t268 GNDA.n2196 65.8183
R2763 GNDA.t268 GNDA.n2194 65.8183
R2764 GNDA.n2304 GNDA.t268 65.8183
R2765 GNDA.t268 GNDA.n2183 65.8183
R2766 GNDA.t208 GNDA.n514 65.8183
R2767 GNDA.t208 GNDA.n513 65.8183
R2768 GNDA.t208 GNDA.n512 65.8183
R2769 GNDA.t208 GNDA.n511 65.8183
R2770 GNDA.t208 GNDA.n502 65.8183
R2771 GNDA.t208 GNDA.n509 65.8183
R2772 GNDA.t208 GNDA.n499 65.8183
R2773 GNDA.t208 GNDA.n510 65.8183
R2774 GNDA.t208 GNDA.n508 65.8183
R2775 GNDA.t208 GNDA.n507 65.8183
R2776 GNDA.t208 GNDA.n506 65.8183
R2777 GNDA.t208 GNDA.n505 65.8183
R2778 GNDA.t208 GNDA.n503 65.8183
R2779 GNDA.t208 GNDA.n501 65.8183
R2780 GNDA.t208 GNDA.n500 65.8183
R2781 GNDA.n2120 GNDA.t208 65.8183
R2782 GNDA.t241 GNDA.n1032 65.8183
R2783 GNDA.t241 GNDA.n1031 65.8183
R2784 GNDA.t241 GNDA.n1030 65.8183
R2785 GNDA.t241 GNDA.n1029 65.8183
R2786 GNDA.t241 GNDA.n1020 65.8183
R2787 GNDA.t241 GNDA.n1027 65.8183
R2788 GNDA.t241 GNDA.n1017 65.8183
R2789 GNDA.t241 GNDA.n1028 65.8183
R2790 GNDA.t241 GNDA.n1026 65.8183
R2791 GNDA.t241 GNDA.n1025 65.8183
R2792 GNDA.t241 GNDA.n1024 65.8183
R2793 GNDA.t241 GNDA.n1023 65.8183
R2794 GNDA.t241 GNDA.n1021 65.8183
R2795 GNDA.t241 GNDA.n1019 65.8183
R2796 GNDA.t241 GNDA.n1018 65.8183
R2797 GNDA.n2009 GNDA.t241 65.8183
R2798 GNDA.t278 GNDA.n1053 65.8183
R2799 GNDA.t278 GNDA.n1052 65.8183
R2800 GNDA.t278 GNDA.n1051 65.8183
R2801 GNDA.t278 GNDA.n1050 65.8183
R2802 GNDA.t278 GNDA.n1041 65.8183
R2803 GNDA.t278 GNDA.n1048 65.8183
R2804 GNDA.t278 GNDA.n1038 65.8183
R2805 GNDA.t278 GNDA.n1049 65.8183
R2806 GNDA.t278 GNDA.n1047 65.8183
R2807 GNDA.t278 GNDA.n1046 65.8183
R2808 GNDA.t278 GNDA.n1045 65.8183
R2809 GNDA.t278 GNDA.n1044 65.8183
R2810 GNDA.t278 GNDA.n1042 65.8183
R2811 GNDA.t278 GNDA.n1040 65.8183
R2812 GNDA.t278 GNDA.n1039 65.8183
R2813 GNDA.n1914 GNDA.t278 65.8183
R2814 GNDA.t213 GNDA.n1177 65.8183
R2815 GNDA.t213 GNDA.n1176 65.8183
R2816 GNDA.t213 GNDA.n1175 65.8183
R2817 GNDA.t213 GNDA.n1174 65.8183
R2818 GNDA.t213 GNDA.n1165 65.8183
R2819 GNDA.t213 GNDA.n1172 65.8183
R2820 GNDA.t213 GNDA.n1162 65.8183
R2821 GNDA.t213 GNDA.n1173 65.8183
R2822 GNDA.t213 GNDA.n1171 65.8183
R2823 GNDA.t213 GNDA.n1170 65.8183
R2824 GNDA.t213 GNDA.n1169 65.8183
R2825 GNDA.t213 GNDA.n1168 65.8183
R2826 GNDA.n1580 GNDA.t249 65.8183
R2827 GNDA.n1582 GNDA.t249 65.8183
R2828 GNDA.n1588 GNDA.t249 65.8183
R2829 GNDA.n1590 GNDA.t249 65.8183
R2830 GNDA.n1564 GNDA.t249 65.8183
R2831 GNDA.n1566 GNDA.t249 65.8183
R2832 GNDA.n1572 GNDA.t249 65.8183
R2833 GNDA.n1574 GNDA.t249 65.8183
R2834 GNDA.t249 GNDA.n1521 65.8183
R2835 GNDA.n1549 GNDA.t249 65.8183
R2836 GNDA.n1545 GNDA.t249 65.8183
R2837 GNDA.n1556 GNDA.t249 65.8183
R2838 GNDA.n1629 GNDA.t249 65.8183
R2839 GNDA.n1616 GNDA.t249 65.8183
R2840 GNDA.n1614 GNDA.t249 65.8183
R2841 GNDA.n1601 GNDA.t249 65.8183
R2842 GNDA.t213 GNDA.n1166 65.8183
R2843 GNDA.t213 GNDA.n1164 65.8183
R2844 GNDA.t213 GNDA.n1163 65.8183
R2845 GNDA.n1263 GNDA.t213 65.8183
R2846 GNDA.t244 GNDA.n856 65.8183
R2847 GNDA.t244 GNDA.n773 65.8183
R2848 GNDA.t244 GNDA.n772 65.8183
R2849 GNDA.t244 GNDA.n771 65.8183
R2850 GNDA.t244 GNDA.n762 65.8183
R2851 GNDA.t244 GNDA.n769 65.8183
R2852 GNDA.t244 GNDA.n760 65.8183
R2853 GNDA.t244 GNDA.n770 65.8183
R2854 GNDA.t244 GNDA.n768 65.8183
R2855 GNDA.t244 GNDA.n767 65.8183
R2856 GNDA.t244 GNDA.n766 65.8183
R2857 GNDA.t244 GNDA.n765 65.8183
R2858 GNDA.t244 GNDA.n763 65.8183
R2859 GNDA.t244 GNDA.n761 65.8183
R2860 GNDA.n859 GNDA.t244 65.8183
R2861 GNDA.t244 GNDA.n752 65.8183
R2862 GNDA.t217 GNDA.n408 65.8183
R2863 GNDA.t217 GNDA.n407 65.8183
R2864 GNDA.t217 GNDA.n406 65.8183
R2865 GNDA.t217 GNDA.n405 65.8183
R2866 GNDA.t217 GNDA.n396 65.8183
R2867 GNDA.t217 GNDA.n403 65.8183
R2868 GNDA.t217 GNDA.n394 65.8183
R2869 GNDA.t217 GNDA.n404 65.8183
R2870 GNDA.t217 GNDA.n402 65.8183
R2871 GNDA.t217 GNDA.n401 65.8183
R2872 GNDA.t217 GNDA.n400 65.8183
R2873 GNDA.t217 GNDA.n399 65.8183
R2874 GNDA.t217 GNDA.n397 65.8183
R2875 GNDA.n2409 GNDA.t217 65.8183
R2876 GNDA.t217 GNDA.n395 65.8183
R2877 GNDA.t217 GNDA.n393 65.8183
R2878 GNDA.t47 GNDA.t57 65.271
R2879 GNDA.t311 GNDA.t94 65.271
R2880 GNDA.t136 GNDA.t18 65.271
R2881 GNDA.t77 GNDA.t298 65.271
R2882 GNDA.n1827 GNDA.t209 65.0078
R2883 GNDA.t176 GNDA.n2188 63.8432
R2884 GNDA.n866 GNDA.t198 63.8432
R2885 GNDA.n2401 GNDA.t192 63.8432
R2886 GNDA.t16 GNDA.t91 62.9326
R2887 GNDA.t112 GNDA.t32 62.9326
R2888 GNDA.t32 GNDA.t120 62.9326
R2889 GNDA.t120 GNDA.t109 62.9326
R2890 GNDA.n2457 GNDA.n2442 61.4316
R2891 GNDA.n2231 GNDA.t178 59.7243
R2892 GNDA.n797 GNDA.t200 59.7243
R2893 GNDA.n678 GNDA.t190 59.7243
R2894 GNDA.n2322 GNDA.t124 58.6946
R2895 GNDA.n2310 GNDA.t125 58.6946
R2896 GNDA.t69 GNDA.n2242 58.6946
R2897 GNDA.t245 GNDA.n1132 57.8461
R2898 GNDA.t268 GNDA.n2182 57.8461
R2899 GNDA.t208 GNDA.n2119 57.8461
R2900 GNDA.t241 GNDA.n2008 57.8461
R2901 GNDA.t278 GNDA.n1913 57.8461
R2902 GNDA.n1599 GNDA.t249 57.8461
R2903 GNDA.t213 GNDA.n1262 57.8461
R2904 GNDA.t244 GNDA.n751 57.8461
R2905 GNDA.t217 GNDA.n2408 57.8461
R2906 GNDA.n179 GNDA.t233 57.5921
R2907 GNDA.t257 GNDA.n71 57.5921
R2908 GNDA.n267 GNDA.t7 57.5921
R2909 GNDA.n315 GNDA.t42 57.5921
R2910 GNDA.n2541 GNDA.t206 57.5921
R2911 GNDA.t227 GNDA.n2501 57.5921
R2912 GNDA.t301 GNDA.t166 56.6352
R2913 GNDA.n876 GNDA.t289 56.6352
R2914 GNDA.t118 GNDA.t162 56.6352
R2915 GNDA.n614 GNDA.n611 56.3995
R2916 GNDA.n1127 GNDA.n483 56.3995
R2917 GNDA.n2178 GNDA.n2177 56.3995
R2918 GNDA.n2177 GNDA.n472 56.3995
R2919 GNDA.n1126 GNDA.n483 56.3995
R2920 GNDA.n2130 GNDA.n490 56.3995
R2921 GNDA.n1825 GNDA.n1055 56.3995
R2922 GNDA.n1642 GNDA.n1641 56.3995
R2923 GNDA.n611 GNDA.n610 56.3995
R2924 GNDA.n1828 GNDA.n1055 56.3995
R2925 GNDA.n1642 GNDA.n1638 56.3995
R2926 GNDA.n2345 GNDA.n2344 55.6055
R2927 GNDA.t245 GNDA.n1142 55.2026
R2928 GNDA.t268 GNDA.n2197 55.2026
R2929 GNDA.t208 GNDA.n504 55.2026
R2930 GNDA.t241 GNDA.n1022 55.2026
R2931 GNDA.t278 GNDA.n1043 55.2026
R2932 GNDA.t213 GNDA.n1167 55.2026
R2933 GNDA.n1558 GNDA.t249 55.2026
R2934 GNDA.t244 GNDA.n764 55.2026
R2935 GNDA.t217 GNDA.n398 55.2026
R2936 GNDA.n879 GNDA.n878 54.5757
R2937 GNDA.n2386 GNDA.n414 54.5757
R2938 GNDA.t39 GNDA.n2402 54.5757
R2939 GNDA.n671 GNDA.t159 54.5757
R2940 GNDA.t314 GNDA.n374 54.5757
R2941 GNDA.t302 GNDA.t203 53.7527
R2942 GNDA.t155 GNDA.t105 53.7527
R2943 GNDA.t295 GNDA.t93 53.7527
R2944 GNDA.t79 GNDA.t83 53.7527
R2945 GNDA.t44 GNDA.t131 53.7527
R2946 GNDA.t4 GNDA.t104 53.7527
R2947 GNDA.t306 GNDA.t160 53.7527
R2948 GNDA.t238 GNDA.t46 53.7527
R2949 GNDA.t184 GNDA.n797 53.546
R2950 GNDA.n1483 GNDA.n1148 53.3664
R2951 GNDA.n1480 GNDA.n1138 53.3664
R2952 GNDA.n1476 GNDA.n1147 53.3664
R2953 GNDA.n1472 GNDA.n1140 53.3664
R2954 GNDA.n1461 GNDA.n1143 53.3664
R2955 GNDA.n1457 GNDA.n1144 53.3664
R2956 GNDA.n1453 GNDA.n1145 53.3664
R2957 GNDA.n1449 GNDA.n1146 53.3664
R2958 GNDA.n1509 GNDA.n1133 53.3664
R2959 GNDA.n1502 GNDA.n1501 53.3664
R2960 GNDA.n1434 GNDA.n1139 53.3664
R2961 GNDA.n1441 GNDA.n1141 53.3664
R2962 GNDA.n1500 GNDA.n1499 53.3664
R2963 GNDA.n1153 GNDA.n1151 53.3664
R2964 GNDA.n1494 GNDA.n1150 53.3664
R2965 GNDA.n1490 GNDA.n1149 53.3664
R2966 GNDA.n1500 GNDA.n1152 53.3664
R2967 GNDA.n1495 GNDA.n1151 53.3664
R2968 GNDA.n1491 GNDA.n1150 53.3664
R2969 GNDA.n1487 GNDA.n1149 53.3664
R2970 GNDA.n1469 GNDA.n1140 53.3664
R2971 GNDA.n1473 GNDA.n1147 53.3664
R2972 GNDA.n1477 GNDA.n1138 53.3664
R2973 GNDA.n1481 GNDA.n1148 53.3664
R2974 GNDA.n1452 GNDA.n1146 53.3664
R2975 GNDA.n1456 GNDA.n1145 53.3664
R2976 GNDA.n1460 GNDA.n1144 53.3664
R2977 GNDA.n1464 GNDA.n1143 53.3664
R2978 GNDA.n1448 GNDA.n1141 53.3664
R2979 GNDA.n1440 GNDA.n1139 53.3664
R2980 GNDA.n1501 GNDA.n1137 53.3664
R2981 GNDA.n1136 GNDA.n1133 53.3664
R2982 GNDA.n2284 GNDA.n2203 53.3664
R2983 GNDA.n2281 GNDA.n2193 53.3664
R2984 GNDA.n2277 GNDA.n2202 53.3664
R2985 GNDA.n2273 GNDA.n2195 53.3664
R2986 GNDA.n2262 GNDA.n2198 53.3664
R2987 GNDA.n2258 GNDA.n2199 53.3664
R2988 GNDA.n2254 GNDA.n2200 53.3664
R2989 GNDA.n2250 GNDA.n2201 53.3664
R2990 GNDA.n2315 GNDA.n2183 53.3664
R2991 GNDA.n2304 GNDA.n2303 53.3664
R2992 GNDA.n2194 GNDA.n2192 53.3664
R2993 GNDA.n2238 GNDA.n2196 53.3664
R2994 GNDA.n2301 GNDA.n2300 53.3664
R2995 GNDA.n2208 GNDA.n2206 53.3664
R2996 GNDA.n2295 GNDA.n2205 53.3664
R2997 GNDA.n2291 GNDA.n2204 53.3664
R2998 GNDA.n2301 GNDA.n2207 53.3664
R2999 GNDA.n2296 GNDA.n2206 53.3664
R3000 GNDA.n2292 GNDA.n2205 53.3664
R3001 GNDA.n2288 GNDA.n2204 53.3664
R3002 GNDA.n2270 GNDA.n2195 53.3664
R3003 GNDA.n2274 GNDA.n2202 53.3664
R3004 GNDA.n2278 GNDA.n2193 53.3664
R3005 GNDA.n2282 GNDA.n2203 53.3664
R3006 GNDA.n2253 GNDA.n2201 53.3664
R3007 GNDA.n2257 GNDA.n2200 53.3664
R3008 GNDA.n2261 GNDA.n2199 53.3664
R3009 GNDA.n2265 GNDA.n2198 53.3664
R3010 GNDA.n2249 GNDA.n2196 53.3664
R3011 GNDA.n2237 GNDA.n2194 53.3664
R3012 GNDA.n2305 GNDA.n2304 53.3664
R3013 GNDA.n2302 GNDA.n2183 53.3664
R3014 GNDA.n2101 GNDA.n510 53.3664
R3015 GNDA.n2097 GNDA.n499 53.3664
R3016 GNDA.n2093 GNDA.n509 53.3664
R3017 GNDA.n2089 GNDA.n502 53.3664
R3018 GNDA.n2078 GNDA.n505 53.3664
R3019 GNDA.n2074 GNDA.n506 53.3664
R3020 GNDA.n2070 GNDA.n507 53.3664
R3021 GNDA.n2066 GNDA.n508 53.3664
R3022 GNDA.n2121 GNDA.n2120 53.3664
R3023 GNDA.n551 GNDA.n500 53.3664
R3024 GNDA.n547 GNDA.n501 53.3664
R3025 GNDA.n540 GNDA.n503 53.3664
R3026 GNDA.n2105 GNDA.n514 53.3664
R3027 GNDA.n2106 GNDA.n513 53.3664
R3028 GNDA.n2110 GNDA.n512 53.3664
R3029 GNDA.n2114 GNDA.n511 53.3664
R3030 GNDA.n2102 GNDA.n514 53.3664
R3031 GNDA.n2109 GNDA.n513 53.3664
R3032 GNDA.n2113 GNDA.n512 53.3664
R3033 GNDA.n2117 GNDA.n511 53.3664
R3034 GNDA.n2086 GNDA.n502 53.3664
R3035 GNDA.n2090 GNDA.n509 53.3664
R3036 GNDA.n2094 GNDA.n499 53.3664
R3037 GNDA.n2098 GNDA.n510 53.3664
R3038 GNDA.n2069 GNDA.n508 53.3664
R3039 GNDA.n2073 GNDA.n507 53.3664
R3040 GNDA.n2077 GNDA.n506 53.3664
R3041 GNDA.n2081 GNDA.n505 53.3664
R3042 GNDA.n2065 GNDA.n503 53.3664
R3043 GNDA.n539 GNDA.n501 53.3664
R3044 GNDA.n548 GNDA.n500 53.3664
R3045 GNDA.n2120 GNDA.n498 53.3664
R3046 GNDA.n1990 GNDA.n1028 53.3664
R3047 GNDA.n1986 GNDA.n1017 53.3664
R3048 GNDA.n1982 GNDA.n1027 53.3664
R3049 GNDA.n1978 GNDA.n1020 53.3664
R3050 GNDA.n1967 GNDA.n1023 53.3664
R3051 GNDA.n1963 GNDA.n1024 53.3664
R3052 GNDA.n1959 GNDA.n1025 53.3664
R3053 GNDA.n1955 GNDA.n1026 53.3664
R3054 GNDA.n2010 GNDA.n2009 53.3664
R3055 GNDA.n1932 GNDA.n1018 53.3664
R3056 GNDA.n1940 GNDA.n1019 53.3664
R3057 GNDA.n1947 GNDA.n1021 53.3664
R3058 GNDA.n1994 GNDA.n1032 53.3664
R3059 GNDA.n1995 GNDA.n1031 53.3664
R3060 GNDA.n1999 GNDA.n1030 53.3664
R3061 GNDA.n2003 GNDA.n1029 53.3664
R3062 GNDA.n1991 GNDA.n1032 53.3664
R3063 GNDA.n1998 GNDA.n1031 53.3664
R3064 GNDA.n2002 GNDA.n1030 53.3664
R3065 GNDA.n2006 GNDA.n1029 53.3664
R3066 GNDA.n1975 GNDA.n1020 53.3664
R3067 GNDA.n1979 GNDA.n1027 53.3664
R3068 GNDA.n1983 GNDA.n1017 53.3664
R3069 GNDA.n1987 GNDA.n1028 53.3664
R3070 GNDA.n1958 GNDA.n1026 53.3664
R3071 GNDA.n1962 GNDA.n1025 53.3664
R3072 GNDA.n1966 GNDA.n1024 53.3664
R3073 GNDA.n1970 GNDA.n1023 53.3664
R3074 GNDA.n1954 GNDA.n1021 53.3664
R3075 GNDA.n1946 GNDA.n1019 53.3664
R3076 GNDA.n1939 GNDA.n1018 53.3664
R3077 GNDA.n2009 GNDA.n1016 53.3664
R3078 GNDA.n1895 GNDA.n1049 53.3664
R3079 GNDA.n1891 GNDA.n1038 53.3664
R3080 GNDA.n1887 GNDA.n1048 53.3664
R3081 GNDA.n1883 GNDA.n1041 53.3664
R3082 GNDA.n1872 GNDA.n1044 53.3664
R3083 GNDA.n1868 GNDA.n1045 53.3664
R3084 GNDA.n1864 GNDA.n1046 53.3664
R3085 GNDA.n1860 GNDA.n1047 53.3664
R3086 GNDA.n1915 GNDA.n1914 53.3664
R3087 GNDA.n1837 GNDA.n1039 53.3664
R3088 GNDA.n1845 GNDA.n1040 53.3664
R3089 GNDA.n1852 GNDA.n1042 53.3664
R3090 GNDA.n1899 GNDA.n1053 53.3664
R3091 GNDA.n1900 GNDA.n1052 53.3664
R3092 GNDA.n1904 GNDA.n1051 53.3664
R3093 GNDA.n1908 GNDA.n1050 53.3664
R3094 GNDA.n1896 GNDA.n1053 53.3664
R3095 GNDA.n1903 GNDA.n1052 53.3664
R3096 GNDA.n1907 GNDA.n1051 53.3664
R3097 GNDA.n1911 GNDA.n1050 53.3664
R3098 GNDA.n1880 GNDA.n1041 53.3664
R3099 GNDA.n1884 GNDA.n1048 53.3664
R3100 GNDA.n1888 GNDA.n1038 53.3664
R3101 GNDA.n1892 GNDA.n1049 53.3664
R3102 GNDA.n1863 GNDA.n1047 53.3664
R3103 GNDA.n1867 GNDA.n1046 53.3664
R3104 GNDA.n1871 GNDA.n1045 53.3664
R3105 GNDA.n1875 GNDA.n1044 53.3664
R3106 GNDA.n1859 GNDA.n1042 53.3664
R3107 GNDA.n1851 GNDA.n1040 53.3664
R3108 GNDA.n1844 GNDA.n1039 53.3664
R3109 GNDA.n1914 GNDA.n1037 53.3664
R3110 GNDA.n1244 GNDA.n1173 53.3664
R3111 GNDA.n1240 GNDA.n1162 53.3664
R3112 GNDA.n1236 GNDA.n1172 53.3664
R3113 GNDA.n1232 GNDA.n1165 53.3664
R3114 GNDA.n1221 GNDA.n1168 53.3664
R3115 GNDA.n1217 GNDA.n1169 53.3664
R3116 GNDA.n1213 GNDA.n1170 53.3664
R3117 GNDA.n1209 GNDA.n1171 53.3664
R3118 GNDA.n1264 GNDA.n1263 53.3664
R3119 GNDA.n1186 GNDA.n1163 53.3664
R3120 GNDA.n1194 GNDA.n1164 53.3664
R3121 GNDA.n1201 GNDA.n1166 53.3664
R3122 GNDA.n1248 GNDA.n1177 53.3664
R3123 GNDA.n1249 GNDA.n1176 53.3664
R3124 GNDA.n1253 GNDA.n1175 53.3664
R3125 GNDA.n1257 GNDA.n1174 53.3664
R3126 GNDA.n1245 GNDA.n1177 53.3664
R3127 GNDA.n1252 GNDA.n1176 53.3664
R3128 GNDA.n1256 GNDA.n1175 53.3664
R3129 GNDA.n1260 GNDA.n1174 53.3664
R3130 GNDA.n1229 GNDA.n1165 53.3664
R3131 GNDA.n1233 GNDA.n1172 53.3664
R3132 GNDA.n1237 GNDA.n1162 53.3664
R3133 GNDA.n1241 GNDA.n1173 53.3664
R3134 GNDA.n1212 GNDA.n1171 53.3664
R3135 GNDA.n1216 GNDA.n1170 53.3664
R3136 GNDA.n1220 GNDA.n1169 53.3664
R3137 GNDA.n1224 GNDA.n1168 53.3664
R3138 GNDA.n1574 GNDA.n1537 53.3664
R3139 GNDA.n1573 GNDA.n1572 53.3664
R3140 GNDA.n1566 GNDA.n1539 53.3664
R3141 GNDA.n1565 GNDA.n1564 53.3664
R3142 GNDA.n1556 GNDA.n1555 53.3664
R3143 GNDA.n1551 GNDA.n1545 53.3664
R3144 GNDA.n1549 GNDA.n1548 53.3664
R3145 GNDA.n1631 GNDA.n1521 53.3664
R3146 GNDA.n1602 GNDA.n1601 53.3664
R3147 GNDA.n1614 GNDA.n1613 53.3664
R3148 GNDA.n1617 GNDA.n1616 53.3664
R3149 GNDA.n1629 GNDA.n1628 53.3664
R3150 GNDA.n1581 GNDA.n1580 53.3664
R3151 GNDA.n1583 GNDA.n1582 53.3664
R3152 GNDA.n1588 GNDA.n1587 53.3664
R3153 GNDA.n1591 GNDA.n1590 53.3664
R3154 GNDA.n1580 GNDA.n1579 53.3664
R3155 GNDA.n1582 GNDA.n1535 53.3664
R3156 GNDA.n1589 GNDA.n1588 53.3664
R3157 GNDA.n1590 GNDA.n1533 53.3664
R3158 GNDA.n1564 GNDA.n1563 53.3664
R3159 GNDA.n1567 GNDA.n1566 53.3664
R3160 GNDA.n1572 GNDA.n1571 53.3664
R3161 GNDA.n1575 GNDA.n1574 53.3664
R3162 GNDA.n1546 GNDA.n1521 53.3664
R3163 GNDA.n1550 GNDA.n1549 53.3664
R3164 GNDA.n1545 GNDA.n1543 53.3664
R3165 GNDA.n1557 GNDA.n1556 53.3664
R3166 GNDA.n1630 GNDA.n1629 53.3664
R3167 GNDA.n1616 GNDA.n1522 53.3664
R3168 GNDA.n1615 GNDA.n1614 53.3664
R3169 GNDA.n1601 GNDA.n1527 53.3664
R3170 GNDA.n1208 GNDA.n1166 53.3664
R3171 GNDA.n1200 GNDA.n1164 53.3664
R3172 GNDA.n1193 GNDA.n1163 53.3664
R3173 GNDA.n1263 GNDA.n1161 53.3664
R3174 GNDA.n838 GNDA.n770 53.3664
R3175 GNDA.n835 GNDA.n760 53.3664
R3176 GNDA.n831 GNDA.n769 53.3664
R3177 GNDA.n827 GNDA.n762 53.3664
R3178 GNDA.n816 GNDA.n765 53.3664
R3179 GNDA.n812 GNDA.n766 53.3664
R3180 GNDA.n808 GNDA.n767 53.3664
R3181 GNDA.n804 GNDA.n768 53.3664
R3182 GNDA.n870 GNDA.n752 53.3664
R3183 GNDA.n859 GNDA.n858 53.3664
R3184 GNDA.n761 GNDA.n759 53.3664
R3185 GNDA.n791 GNDA.n763 53.3664
R3186 GNDA.n856 GNDA.n855 53.3664
R3187 GNDA.n775 GNDA.n773 53.3664
R3188 GNDA.n850 GNDA.n772 53.3664
R3189 GNDA.n846 GNDA.n771 53.3664
R3190 GNDA.n856 GNDA.n774 53.3664
R3191 GNDA.n851 GNDA.n773 53.3664
R3192 GNDA.n847 GNDA.n772 53.3664
R3193 GNDA.n843 GNDA.n771 53.3664
R3194 GNDA.n824 GNDA.n762 53.3664
R3195 GNDA.n828 GNDA.n769 53.3664
R3196 GNDA.n832 GNDA.n760 53.3664
R3197 GNDA.n836 GNDA.n770 53.3664
R3198 GNDA.n807 GNDA.n768 53.3664
R3199 GNDA.n811 GNDA.n767 53.3664
R3200 GNDA.n815 GNDA.n766 53.3664
R3201 GNDA.n819 GNDA.n765 53.3664
R3202 GNDA.n803 GNDA.n763 53.3664
R3203 GNDA.n792 GNDA.n761 53.3664
R3204 GNDA.n860 GNDA.n859 53.3664
R3205 GNDA.n857 GNDA.n752 53.3664
R3206 GNDA.n719 GNDA.n404 53.3664
R3207 GNDA.n715 GNDA.n394 53.3664
R3208 GNDA.n711 GNDA.n403 53.3664
R3209 GNDA.n707 GNDA.n396 53.3664
R3210 GNDA.n696 GNDA.n399 53.3664
R3211 GNDA.n692 GNDA.n400 53.3664
R3212 GNDA.n688 GNDA.n401 53.3664
R3213 GNDA.n684 GNDA.n402 53.3664
R3214 GNDA.n410 GNDA.n393 53.3664
R3215 GNDA.n2397 GNDA.n395 53.3664
R3216 GNDA.n2410 GNDA.n2409 53.3664
R3217 GNDA.n673 GNDA.n397 53.3664
R3218 GNDA.n723 GNDA.n408 53.3664
R3219 GNDA.n724 GNDA.n407 53.3664
R3220 GNDA.n728 GNDA.n406 53.3664
R3221 GNDA.n732 GNDA.n405 53.3664
R3222 GNDA.n720 GNDA.n408 53.3664
R3223 GNDA.n727 GNDA.n407 53.3664
R3224 GNDA.n731 GNDA.n406 53.3664
R3225 GNDA.n734 GNDA.n405 53.3664
R3226 GNDA.n704 GNDA.n396 53.3664
R3227 GNDA.n708 GNDA.n403 53.3664
R3228 GNDA.n712 GNDA.n394 53.3664
R3229 GNDA.n716 GNDA.n404 53.3664
R3230 GNDA.n687 GNDA.n402 53.3664
R3231 GNDA.n691 GNDA.n401 53.3664
R3232 GNDA.n695 GNDA.n400 53.3664
R3233 GNDA.n699 GNDA.n399 53.3664
R3234 GNDA.n683 GNDA.n397 53.3664
R3235 GNDA.n2409 GNDA.n392 53.3664
R3236 GNDA.n395 GNDA.n391 53.3664
R3237 GNDA.n2396 GNDA.n393 53.3664
R3238 GNDA.n1664 GNDA.n1663 52.7091
R3239 GNDA.n1663 GNDA.n1102 52.7091
R3240 GNDA.n1657 GNDA.n1102 52.7091
R3241 GNDA.n1657 GNDA.n1656 52.7091
R3242 GNDA.n1656 GNDA.n1655 52.7091
R3243 GNDA.n1649 GNDA.n1109 52.7091
R3244 GNDA.n1649 GNDA.n1648 52.7091
R3245 GNDA.n1648 GNDA.n1647 52.7091
R3246 GNDA.n1647 GNDA.n1110 52.7091
R3247 GNDA.n1640 GNDA.n1110 52.7091
R3248 GNDA.n1640 GNDA.n1639 52.7091
R3249 GNDA.n1801 GNDA.n1063 52.7091
R3250 GNDA.n1807 GNDA.n1063 52.7091
R3251 GNDA.n1808 GNDA.n1807 52.7091
R3252 GNDA.n1810 GNDA.n1808 52.7091
R3253 GNDA.n1810 GNDA.n1809 52.7091
R3254 GNDA.n1817 GNDA.n1816 52.7091
R3255 GNDA.n1819 GNDA.n1817 52.7091
R3256 GNDA.n1819 GNDA.n1818 52.7091
R3257 GNDA.n1818 GNDA.n1056 52.7091
R3258 GNDA.n1826 GNDA.n1056 52.7091
R3259 GNDA.n1827 GNDA.n1826 52.7091
R3260 GNDA.n644 GNDA.n620 52.7091
R3261 GNDA.n651 GNDA.n620 52.7091
R3262 GNDA.n652 GNDA.n651 52.7091
R3263 GNDA.n653 GNDA.n652 52.7091
R3264 GNDA.n653 GNDA.n386 52.7091
R3265 GNDA.n615 GNDA.n387 52.7091
R3266 GNDA.n661 GNDA.n615 52.7091
R3267 GNDA.n662 GNDA.n661 52.7091
R3268 GNDA.n665 GNDA.n662 52.7091
R3269 GNDA.n665 GNDA.n664 52.7091
R3270 GNDA.n664 GNDA.n663 52.7091
R3271 GNDA.t209 GNDA.n419 51.4866
R3272 GNDA.n2375 GNDA.t209 51.4866
R3273 GNDA.t89 GNDA.t22 49.9132
R3274 GNDA.t55 GNDA.t95 49.9132
R3275 GNDA.t54 GNDA.t317 49.9132
R3276 GNDA.t27 GNDA.t114 49.9132
R3277 GNDA.n866 GNDA.t172 49.4271
R3278 GNDA.t1 GNDA.n414 48.3974
R3279 GNDA.n2345 GNDA.t129 47.3677
R3280 GNDA.t9 GNDA.t273 46.338
R3281 GNDA.t263 GNDA.t15 46.338
R3282 GNDA.t209 GNDA.n1378 46.2335
R3283 GNDA.n1321 GNDA.t209 46.2335
R3284 GNDA.n1679 GNDA.t209 46.2335
R3285 GNDA.n191 GNDA.n179 46.0738
R3286 GNDA.n209 GNDA.n71 46.0738
R3287 GNDA.t7 GNDA.t286 46.0738
R3288 GNDA.t294 GNDA.t146 46.0738
R3289 GNDA.t98 GNDA.t121 46.0738
R3290 GNDA.t24 GNDA.t157 46.0738
R3291 GNDA.t17 GNDA.t71 46.0738
R3292 GNDA.t25 GNDA.t143 46.0738
R3293 GNDA.t6 GNDA.t315 46.0738
R3294 GNDA.t230 GNDA.t42 46.0738
R3295 GNDA.n2553 GNDA.n2541 46.0738
R3296 GNDA.n2501 GNDA.n2457 46.0738
R3297 GNDA.t273 GNDA.n2187 43.2488
R3298 GNDA.t172 GNDA.n755 43.2488
R3299 GNDA.n2402 GNDA.t188 43.2488
R3300 GNDA.n1379 GNDA.t209 42.2987
R3301 GNDA.t209 GNDA.n1320 42.2987
R3302 GNDA.n1097 GNDA.t209 42.2987
R3303 GNDA.t64 GNDA.t150 42.2405
R3304 GNDA.t150 GNDA.t13 42.2405
R3305 GNDA.t126 GNDA.t66 42.2405
R3306 GNDA.t66 GNDA.t33 42.2405
R3307 GNDA.n337 GNDA.t70 42.2344
R3308 GNDA.n864 GNDA.t50 42.2191
R3309 GNDA.t209 GNDA.t129 41.1894
R3310 GNDA.t209 GNDA.t1 41.1894
R3311 GNDA.t109 GNDA.t108 39.8575
R3312 GNDA.n2227 GNDA.n380 39.3903
R3313 GNDA.n2242 GNDA.t168 39.1299
R3314 GNDA.n787 GNDA.n786 39.1299
R3315 GNDA.n798 GNDA.t184 39.1299
R3316 GNDA.n679 GNDA.t263 39.1299
R3317 GNDA.t286 GNDA.t294 38.3949
R3318 GNDA.t146 GNDA.t98 38.3949
R3319 GNDA.t121 GNDA.t24 38.3949
R3320 GNDA.t157 GNDA.t17 38.3949
R3321 GNDA.t71 GNDA.t25 38.3949
R3322 GNDA.t143 GNDA.t6 38.3949
R3323 GNDA.t315 GNDA.t230 38.3949
R3324 GNDA.n744 GNDA.n419 38.1002
R3325 GNDA.n878 GNDA.n742 38.1002
R3326 GNDA.n2414 GNDA.t159 38.1002
R3327 GNDA.n679 GNDA.t314 38.1002
R3328 GNDA.n2375 GNDA.n417 37.0705
R3329 GNDA.t194 GNDA.t209 36.0408
R3330 GNDA.t209 GNDA.t174 36.0408
R3331 GNDA.n1655 GNDA.t209 35.7252
R3332 GNDA.n1809 GNDA.t209 35.7252
R3333 GNDA.t209 GNDA.n386 35.7252
R3334 GNDA.n2428 GNDA.n2427 35.3278
R3335 GNDA.n1639 GNDA.t65 35.1396
R3336 GNDA.t22 GNDA.t99 34.5555
R3337 GNDA.t60 GNDA.t55 34.5555
R3338 GNDA.t317 GNDA.t76 34.5555
R3339 GNDA.t133 GNDA.t27 34.5555
R3340 GNDA.n2187 GNDA.t124 33.9813
R3341 GNDA.t125 GNDA.n2309 33.9813
R3342 GNDA.n876 GNDA.n875 33.9813
R3343 GNDA.t178 GNDA.n2230 32.9516
R3344 GNDA.t200 GNDA.n796 32.9516
R3345 GNDA.t190 GNDA.n677 32.9516
R3346 GNDA.n2059 GNDA.t209 32.9056
R3347 GNDA.n1113 GNDA.t209 32.9056
R3348 GNDA.n2432 GNDA.n2431 32.3063
R3349 GNDA.t119 GNDA.t313 30.716
R3350 GNDA.t203 GNDA.t81 30.716
R3351 GNDA.t105 GNDA.t302 30.716
R3352 GNDA.t93 GNDA.t155 30.716
R3353 GNDA.t83 GNDA.t295 30.716
R3354 GNDA.t131 GNDA.t79 30.716
R3355 GNDA.t104 GNDA.t44 30.716
R3356 GNDA.t160 GNDA.t4 30.716
R3357 GNDA.t46 GNDA.t306 30.716
R3358 GNDA.t0 GNDA.t238 30.716
R3359 GNDA.n2561 GNDA.n0 29.8047
R3360 GNDA.t127 GNDA.n372 29.2831
R3361 GNDA.n2311 GNDA.t176 28.8327
R3362 GNDA.t198 GNDA.n865 28.8327
R3363 GNDA.t192 GNDA.n2391 28.8327
R3364 GNDA.n2311 GNDA.t301 27.803
R3365 GNDA.n2231 GNDA.t310 27.803
R3366 GNDA.n2244 GNDA.t11 27.803
R3367 GNDA.n1485 GNDA.n1484 27.5561
R3368 GNDA.n2286 GNDA.n2285 27.5561
R3369 GNDA.n2103 GNDA.n2100 27.5561
R3370 GNDA.n1992 GNDA.n1989 27.5561
R3371 GNDA.n1897 GNDA.n1894 27.5561
R3372 GNDA.n1246 GNDA.n1243 27.5561
R3373 GNDA.n1578 GNDA.n1577 27.5561
R3374 GNDA.n840 GNDA.n839 27.5561
R3375 GNDA.n721 GNDA.n718 27.5561
R3376 GNDA.t68 GNDA.n267 26.8766
R3377 GNDA.n315 GNDA.t106 26.8766
R3378 GNDA.t137 GNDA.t20 26.8766
R3379 GNDA.n1467 GNDA.n1466 26.6672
R3380 GNDA.n2268 GNDA.n2267 26.6672
R3381 GNDA.n2084 GNDA.n2083 26.6672
R3382 GNDA.n1973 GNDA.n1972 26.6672
R3383 GNDA.n1878 GNDA.n1877 26.6672
R3384 GNDA.n1227 GNDA.n1226 26.6672
R3385 GNDA.n1561 GNDA.n1560 26.6672
R3386 GNDA.n822 GNDA.n821 26.6672
R3387 GNDA.n702 GNDA.n701 26.6672
R3388 GNDA.t310 GNDA.t168 25.7435
R3389 GNDA.t188 GNDA.t309 25.7435
R3390 GNDA.n2218 GNDA.n2217 25.3679
R3391 GNDA.n290 GNDA.n289 24.991
R3392 GNDA.n280 GNDA.n279 24.7472
R3393 GNDA.n2561 GNDA.n2560 24.133
R3394 GNDA.n2326 GNDA.t177 24.0005
R3395 GNDA.n2326 GNDA.t167 24.0005
R3396 GNDA.n2328 GNDA.t195 24.0005
R3397 GNDA.n2328 GNDA.t179 24.0005
R3398 GNDA.n2330 GNDA.t169 24.0005
R3399 GNDA.n2330 GNDA.t197 24.0005
R3400 GNDA.n2336 GNDA.t183 24.0005
R3401 GNDA.n2336 GNDA.t173 24.0005
R3402 GNDA.n2334 GNDA.t199 24.0005
R3403 GNDA.n2334 GNDA.t181 24.0005
R3404 GNDA.n2332 GNDA.t171 24.0005
R3405 GNDA.n2332 GNDA.t201 24.0005
R3406 GNDA.n415 GNDA.t185 24.0005
R3407 GNDA.n415 GNDA.t187 24.0005
R3408 GNDA.n2381 GNDA.t165 24.0005
R3409 GNDA.n2381 GNDA.t189 24.0005
R3410 GNDA.n2379 GNDA.t193 24.0005
R3411 GNDA.n2379 GNDA.t175 24.0005
R3412 GNDA.n375 GNDA.t163 24.0005
R3413 GNDA.n375 GNDA.t191 24.0005
R3414 GNDA.n2387 GNDA.t145 23.6841
R3415 GNDA.t309 GNDA.n2401 23.6841
R3416 GNDA.n677 GNDA.t118 23.6841
R3417 GNDA.n309 GNDA.n303 23.6611
R3418 GNDA.n300 GNDA.n298 23.6611
R3419 GNDA.n146 GNDA.n145 22.8576
R3420 GNDA.n258 GNDA.n257 22.8576
R3421 GNDA.n233 GNDA.n232 22.8576
R3422 GNDA.n199 GNDA.n198 22.8576
R3423 GNDA.n194 GNDA.n193 22.8576
R3424 GNDA.n272 GNDA.n271 22.8576
R3425 GNDA.n318 GNDA.n317 22.8576
R3426 GNDA.n331 GNDA.n330 22.8576
R3427 GNDA.n328 GNDA.n327 22.8576
R3428 GNDA.n350 GNDA.n349 22.8576
R3429 GNDA.n355 GNDA.n354 22.8576
R3430 GNDA.n2556 GNDA.n2555 22.8576
R3431 GNDA.n2447 GNDA.n14 22.8576
R3432 GNDA.n2515 GNDA.n2514 22.8576
R3433 GNDA.n2475 GNDA.n2474 22.8576
R3434 GNDA.n153 GNDA.n152 22.8576
R3435 GNDA.n875 GNDA.t182 22.6544
R3436 GNDA.n2403 GNDA.t164 22.6544
R3437 GNDA.n2438 GNDA.t127 21.084
R3438 GNDA.n1300 GNDA.n1299 21.0192
R3439 GNDA.t91 GNDA.t112 20.9779
R3440 GNDA.n2325 GNDA.n2324 20.8233
R3441 GNDA.n2343 GNDA.n2342 20.8233
R3442 GNDA.n2339 GNDA.n2338 20.8233
R3443 GNDA.n2377 GNDA.n2376 20.8233
R3444 GNDA.n2385 GNDA.n2384 20.8233
R3445 GNDA.n2436 GNDA.n2435 20.8233
R3446 GNDA.n2229 GNDA.t209 20.5949
R3447 GNDA.t123 GNDA.n2229 20.5949
R3448 GNDA.n2344 GNDA.t11 20.5949
R3449 GNDA.t145 GNDA.n2386 20.5949
R3450 GNDA.n2425 GNDA.t148 20.5949
R3451 GNDA.n2425 GNDA.t209 20.5949
R3452 GNDA.n476 GNDA.t209 19.9378
R3453 GNDA.n51 GNDA.t100 19.7005
R3454 GNDA.n51 GNDA.t21 19.7005
R3455 GNDA.n49 GNDA.t8 19.7005
R3456 GNDA.n49 GNDA.t90 19.7005
R3457 GNDA.n47 GNDA.t63 19.7005
R3458 GNDA.n47 GNDA.t29 19.7005
R3459 GNDA.n45 GNDA.t102 19.7005
R3460 GNDA.n45 GNDA.t88 19.7005
R3461 GNDA.n43 GNDA.t61 19.7005
R3462 GNDA.n43 GNDA.t49 19.7005
R3463 GNDA.n42 GNDA.t84 19.7005
R3464 GNDA.n42 GNDA.t59 19.7005
R3465 GNDA.n12 GNDA.t161 19.7005
R3466 GNDA.n12 GNDA.t132 19.7005
R3467 GNDA.n10 GNDA.t141 19.7005
R3468 GNDA.n10 GNDA.t75 19.7005
R3469 GNDA.n8 GNDA.t140 19.7005
R3470 GNDA.n8 GNDA.t135 19.7005
R3471 GNDA.n6 GNDA.t297 19.7005
R3472 GNDA.n6 GNDA.t26 19.7005
R3473 GNDA.n4 GNDA.t142 19.7005
R3474 GNDA.n4 GNDA.t53 19.7005
R3475 GNDA.n3 GNDA.t52 19.7005
R3476 GNDA.n3 GNDA.t115 19.7005
R3477 GNDA.n1344 GNDA.t209 19.6741
R3478 GNDA.t57 GNDA.t62 19.1977
R3479 GNDA.t48 GNDA.t311 19.1977
R3480 GNDA.t18 GNDA.t134 19.1977
R3481 GNDA.t51 GNDA.t77 19.1977
R3482 GNDA.n301 GNDA.n290 19.0713
R3483 GNDA.n1302 GNDA.n1294 18.5605
R3484 GNDA.n2243 GNDA.t196 18.5355
R3485 GNDA.t186 GNDA.n742 18.5355
R3486 GNDA.n2442 GNDA.t16 18.3557
R3487 GNDA GNDA.n379 18.1546
R3488 GNDA.n197 GNDA.n194 18.1442
R3489 GNDA.n2557 GNDA.n14 18.1442
R3490 GNDA.n329 GNDA.n328 17.8005
R3491 GNDA.n1803 GNDA.n1799 17.5843
R3492 GNDA.n1667 GNDA.n1100 17.5843
R3493 GNDA.n646 GNDA.n642 17.5843
R3494 GNDA.t65 GNDA.t10 17.57
R3495 GNDA.n2323 GNDA.t209 17.5058
R3496 GNDA.n2438 GNDA.n2437 17.5058
R3497 GNDA.n1109 GNDA.t209 16.9844
R3498 GNDA.n1816 GNDA.t209 16.9844
R3499 GNDA.t209 GNDA.n387 16.9844
R3500 GNDA.n1367 GNDA.n1366 16.9379
R3501 GNDA.n2173 GNDA.n2155 16.9379
R3502 GNDA.n965 GNDA.n962 16.9379
R3503 GNDA.n1722 GNDA.n1721 16.7709
R3504 GNDA.n909 GNDA.n908 16.7709
R3505 GNDA.n2044 GNDA.n986 16.7709
R3506 GNDA.n2370 GNDA.n443 16.7709
R3507 GNDA.n2558 GNDA.n13 16.5057
R3508 GNDA.n210 GNDA.t212 16.0005
R3509 GNDA.n66 GNDA.t252 16.0005
R3510 GNDA.n307 GNDA.t231 16.0005
R3511 GNDA.n291 GNDA.t204 16.0005
R3512 GNDA.n296 GNDA.t284 16.0005
R3513 GNDA.n284 GNDA.t223 16.0005
R3514 GNDA.n270 GNDA.t225 16.0005
R3515 GNDA.n311 GNDA.t243 16.0005
R3516 GNDA.n60 GNDA.t220 16.0005
R3517 GNDA.n322 GNDA.t236 16.0005
R3518 GNDA.n1498 GNDA.n1485 16.0005
R3519 GNDA.n1498 GNDA.n1497 16.0005
R3520 GNDA.n1497 GNDA.n1496 16.0005
R3521 GNDA.n1496 GNDA.n1493 16.0005
R3522 GNDA.n1493 GNDA.n1492 16.0005
R3523 GNDA.n1492 GNDA.n1489 16.0005
R3524 GNDA.n1489 GNDA.n1488 16.0005
R3525 GNDA.n1488 GNDA.n1129 16.0005
R3526 GNDA.n1484 GNDA.n1482 16.0005
R3527 GNDA.n1482 GNDA.n1479 16.0005
R3528 GNDA.n1479 GNDA.n1478 16.0005
R3529 GNDA.n1478 GNDA.n1475 16.0005
R3530 GNDA.n1475 GNDA.n1474 16.0005
R3531 GNDA.n1474 GNDA.n1471 16.0005
R3532 GNDA.n1471 GNDA.n1470 16.0005
R3533 GNDA.n1470 GNDA.n1467 16.0005
R3534 GNDA.n1466 GNDA.n1463 16.0005
R3535 GNDA.n1463 GNDA.n1462 16.0005
R3536 GNDA.n1462 GNDA.n1459 16.0005
R3537 GNDA.n1459 GNDA.n1458 16.0005
R3538 GNDA.n1458 GNDA.n1455 16.0005
R3539 GNDA.n1455 GNDA.n1454 16.0005
R3540 GNDA.n1454 GNDA.n1451 16.0005
R3541 GNDA.n1451 GNDA.n1450 16.0005
R3542 GNDA.n2299 GNDA.n2286 16.0005
R3543 GNDA.n2299 GNDA.n2298 16.0005
R3544 GNDA.n2298 GNDA.n2297 16.0005
R3545 GNDA.n2297 GNDA.n2294 16.0005
R3546 GNDA.n2294 GNDA.n2293 16.0005
R3547 GNDA.n2293 GNDA.n2290 16.0005
R3548 GNDA.n2290 GNDA.n2289 16.0005
R3549 GNDA.n2289 GNDA.n2180 16.0005
R3550 GNDA.n2285 GNDA.n2283 16.0005
R3551 GNDA.n2283 GNDA.n2280 16.0005
R3552 GNDA.n2280 GNDA.n2279 16.0005
R3553 GNDA.n2279 GNDA.n2276 16.0005
R3554 GNDA.n2276 GNDA.n2275 16.0005
R3555 GNDA.n2275 GNDA.n2272 16.0005
R3556 GNDA.n2272 GNDA.n2271 16.0005
R3557 GNDA.n2271 GNDA.n2268 16.0005
R3558 GNDA.n2267 GNDA.n2264 16.0005
R3559 GNDA.n2264 GNDA.n2263 16.0005
R3560 GNDA.n2263 GNDA.n2260 16.0005
R3561 GNDA.n2260 GNDA.n2259 16.0005
R3562 GNDA.n2259 GNDA.n2256 16.0005
R3563 GNDA.n2256 GNDA.n2255 16.0005
R3564 GNDA.n2255 GNDA.n2252 16.0005
R3565 GNDA.n2252 GNDA.n2251 16.0005
R3566 GNDA.n2104 GNDA.n2103 16.0005
R3567 GNDA.n2107 GNDA.n2104 16.0005
R3568 GNDA.n2108 GNDA.n2107 16.0005
R3569 GNDA.n2111 GNDA.n2108 16.0005
R3570 GNDA.n2112 GNDA.n2111 16.0005
R3571 GNDA.n2115 GNDA.n2112 16.0005
R3572 GNDA.n2116 GNDA.n2115 16.0005
R3573 GNDA.n2116 GNDA.n493 16.0005
R3574 GNDA.n2100 GNDA.n2099 16.0005
R3575 GNDA.n2099 GNDA.n2096 16.0005
R3576 GNDA.n2096 GNDA.n2095 16.0005
R3577 GNDA.n2095 GNDA.n2092 16.0005
R3578 GNDA.n2092 GNDA.n2091 16.0005
R3579 GNDA.n2091 GNDA.n2088 16.0005
R3580 GNDA.n2088 GNDA.n2087 16.0005
R3581 GNDA.n2087 GNDA.n2084 16.0005
R3582 GNDA.n2083 GNDA.n2080 16.0005
R3583 GNDA.n2080 GNDA.n2079 16.0005
R3584 GNDA.n2079 GNDA.n2076 16.0005
R3585 GNDA.n2076 GNDA.n2075 16.0005
R3586 GNDA.n2075 GNDA.n2072 16.0005
R3587 GNDA.n2072 GNDA.n2071 16.0005
R3588 GNDA.n2071 GNDA.n2068 16.0005
R3589 GNDA.n2068 GNDA.n2067 16.0005
R3590 GNDA.n1993 GNDA.n1992 16.0005
R3591 GNDA.n1996 GNDA.n1993 16.0005
R3592 GNDA.n1997 GNDA.n1996 16.0005
R3593 GNDA.n2000 GNDA.n1997 16.0005
R3594 GNDA.n2001 GNDA.n2000 16.0005
R3595 GNDA.n2004 GNDA.n2001 16.0005
R3596 GNDA.n2005 GNDA.n2004 16.0005
R3597 GNDA.n2005 GNDA.n1012 16.0005
R3598 GNDA.n1989 GNDA.n1988 16.0005
R3599 GNDA.n1988 GNDA.n1985 16.0005
R3600 GNDA.n1985 GNDA.n1984 16.0005
R3601 GNDA.n1984 GNDA.n1981 16.0005
R3602 GNDA.n1981 GNDA.n1980 16.0005
R3603 GNDA.n1980 GNDA.n1977 16.0005
R3604 GNDA.n1977 GNDA.n1976 16.0005
R3605 GNDA.n1976 GNDA.n1973 16.0005
R3606 GNDA.n1972 GNDA.n1969 16.0005
R3607 GNDA.n1969 GNDA.n1968 16.0005
R3608 GNDA.n1968 GNDA.n1965 16.0005
R3609 GNDA.n1965 GNDA.n1964 16.0005
R3610 GNDA.n1964 GNDA.n1961 16.0005
R3611 GNDA.n1961 GNDA.n1960 16.0005
R3612 GNDA.n1960 GNDA.n1957 16.0005
R3613 GNDA.n1957 GNDA.n1956 16.0005
R3614 GNDA.n1898 GNDA.n1897 16.0005
R3615 GNDA.n1901 GNDA.n1898 16.0005
R3616 GNDA.n1902 GNDA.n1901 16.0005
R3617 GNDA.n1905 GNDA.n1902 16.0005
R3618 GNDA.n1906 GNDA.n1905 16.0005
R3619 GNDA.n1909 GNDA.n1906 16.0005
R3620 GNDA.n1910 GNDA.n1909 16.0005
R3621 GNDA.n1910 GNDA.n1033 16.0005
R3622 GNDA.n1894 GNDA.n1893 16.0005
R3623 GNDA.n1893 GNDA.n1890 16.0005
R3624 GNDA.n1890 GNDA.n1889 16.0005
R3625 GNDA.n1889 GNDA.n1886 16.0005
R3626 GNDA.n1886 GNDA.n1885 16.0005
R3627 GNDA.n1885 GNDA.n1882 16.0005
R3628 GNDA.n1882 GNDA.n1881 16.0005
R3629 GNDA.n1881 GNDA.n1878 16.0005
R3630 GNDA.n1877 GNDA.n1874 16.0005
R3631 GNDA.n1874 GNDA.n1873 16.0005
R3632 GNDA.n1873 GNDA.n1870 16.0005
R3633 GNDA.n1870 GNDA.n1869 16.0005
R3634 GNDA.n1869 GNDA.n1866 16.0005
R3635 GNDA.n1866 GNDA.n1865 16.0005
R3636 GNDA.n1865 GNDA.n1862 16.0005
R3637 GNDA.n1862 GNDA.n1861 16.0005
R3638 GNDA.n1247 GNDA.n1246 16.0005
R3639 GNDA.n1250 GNDA.n1247 16.0005
R3640 GNDA.n1251 GNDA.n1250 16.0005
R3641 GNDA.n1254 GNDA.n1251 16.0005
R3642 GNDA.n1255 GNDA.n1254 16.0005
R3643 GNDA.n1258 GNDA.n1255 16.0005
R3644 GNDA.n1259 GNDA.n1258 16.0005
R3645 GNDA.n1259 GNDA.n1157 16.0005
R3646 GNDA.n1243 GNDA.n1242 16.0005
R3647 GNDA.n1242 GNDA.n1239 16.0005
R3648 GNDA.n1239 GNDA.n1238 16.0005
R3649 GNDA.n1238 GNDA.n1235 16.0005
R3650 GNDA.n1235 GNDA.n1234 16.0005
R3651 GNDA.n1234 GNDA.n1231 16.0005
R3652 GNDA.n1231 GNDA.n1230 16.0005
R3653 GNDA.n1230 GNDA.n1227 16.0005
R3654 GNDA.n1226 GNDA.n1223 16.0005
R3655 GNDA.n1223 GNDA.n1222 16.0005
R3656 GNDA.n1222 GNDA.n1219 16.0005
R3657 GNDA.n1219 GNDA.n1218 16.0005
R3658 GNDA.n1218 GNDA.n1215 16.0005
R3659 GNDA.n1215 GNDA.n1214 16.0005
R3660 GNDA.n1214 GNDA.n1211 16.0005
R3661 GNDA.n1211 GNDA.n1210 16.0005
R3662 GNDA.n1578 GNDA.n1536 16.0005
R3663 GNDA.n1584 GNDA.n1536 16.0005
R3664 GNDA.n1585 GNDA.n1584 16.0005
R3665 GNDA.n1586 GNDA.n1585 16.0005
R3666 GNDA.n1586 GNDA.n1534 16.0005
R3667 GNDA.n1592 GNDA.n1534 16.0005
R3668 GNDA.n1593 GNDA.n1592 16.0005
R3669 GNDA.n1597 GNDA.n1593 16.0005
R3670 GNDA.n1577 GNDA.n1576 16.0005
R3671 GNDA.n1576 GNDA.n1538 16.0005
R3672 GNDA.n1570 GNDA.n1538 16.0005
R3673 GNDA.n1570 GNDA.n1569 16.0005
R3674 GNDA.n1569 GNDA.n1568 16.0005
R3675 GNDA.n1568 GNDA.n1540 16.0005
R3676 GNDA.n1562 GNDA.n1540 16.0005
R3677 GNDA.n1562 GNDA.n1561 16.0005
R3678 GNDA.n1560 GNDA.n1542 16.0005
R3679 GNDA.n1554 GNDA.n1542 16.0005
R3680 GNDA.n1554 GNDA.n1553 16.0005
R3681 GNDA.n1553 GNDA.n1552 16.0005
R3682 GNDA.n1552 GNDA.n1544 16.0005
R3683 GNDA.n1547 GNDA.n1544 16.0005
R3684 GNDA.n1547 GNDA.n1520 16.0005
R3685 GNDA.n1632 GNDA.n1520 16.0005
R3686 GNDA.n854 GNDA.n840 16.0005
R3687 GNDA.n854 GNDA.n853 16.0005
R3688 GNDA.n853 GNDA.n852 16.0005
R3689 GNDA.n852 GNDA.n849 16.0005
R3690 GNDA.n849 GNDA.n848 16.0005
R3691 GNDA.n848 GNDA.n845 16.0005
R3692 GNDA.n845 GNDA.n844 16.0005
R3693 GNDA.n844 GNDA.n841 16.0005
R3694 GNDA.n839 GNDA.n837 16.0005
R3695 GNDA.n837 GNDA.n834 16.0005
R3696 GNDA.n834 GNDA.n833 16.0005
R3697 GNDA.n833 GNDA.n830 16.0005
R3698 GNDA.n830 GNDA.n829 16.0005
R3699 GNDA.n829 GNDA.n826 16.0005
R3700 GNDA.n826 GNDA.n825 16.0005
R3701 GNDA.n825 GNDA.n822 16.0005
R3702 GNDA.n821 GNDA.n818 16.0005
R3703 GNDA.n818 GNDA.n817 16.0005
R3704 GNDA.n817 GNDA.n814 16.0005
R3705 GNDA.n814 GNDA.n813 16.0005
R3706 GNDA.n813 GNDA.n810 16.0005
R3707 GNDA.n810 GNDA.n809 16.0005
R3708 GNDA.n809 GNDA.n806 16.0005
R3709 GNDA.n806 GNDA.n805 16.0005
R3710 GNDA.n722 GNDA.n721 16.0005
R3711 GNDA.n725 GNDA.n722 16.0005
R3712 GNDA.n726 GNDA.n725 16.0005
R3713 GNDA.n729 GNDA.n726 16.0005
R3714 GNDA.n730 GNDA.n729 16.0005
R3715 GNDA.n733 GNDA.n730 16.0005
R3716 GNDA.n735 GNDA.n733 16.0005
R3717 GNDA.n736 GNDA.n735 16.0005
R3718 GNDA.n718 GNDA.n717 16.0005
R3719 GNDA.n717 GNDA.n714 16.0005
R3720 GNDA.n714 GNDA.n713 16.0005
R3721 GNDA.n713 GNDA.n710 16.0005
R3722 GNDA.n710 GNDA.n709 16.0005
R3723 GNDA.n709 GNDA.n706 16.0005
R3724 GNDA.n706 GNDA.n705 16.0005
R3725 GNDA.n705 GNDA.n702 16.0005
R3726 GNDA.n701 GNDA.n698 16.0005
R3727 GNDA.n698 GNDA.n697 16.0005
R3728 GNDA.n697 GNDA.n694 16.0005
R3729 GNDA.n694 GNDA.n693 16.0005
R3730 GNDA.n693 GNDA.n690 16.0005
R3731 GNDA.n690 GNDA.n689 16.0005
R3732 GNDA.n689 GNDA.n686 16.0005
R3733 GNDA.n686 GNDA.n685 16.0005
R3734 GNDA.n1301 GNDA.n1300 16.0005
R3735 GNDA.n1302 GNDA.n1301 16.0005
R3736 GNDA.t196 GNDA.t69 15.4463
R3737 GNDA.t164 GNDA.t39 15.4463
R3738 GNDA.n2474 GNDA.n2473 14.9255
R3739 GNDA.n152 GNDA.n151 14.9255
R3740 GNDA.n281 GNDA.n280 14.8213
R3741 GNDA.n303 GNDA.n302 14.8213
R3742 GNDA.n301 GNDA.n300 14.8213
R3743 GNDA.n2060 GNDA.n2059 14.555
R3744 GNDA.n1517 GNDA.n1113 14.555
R3745 GNDA.n2327 GNDA.n2325 14.363
R3746 GNDA.n354 GNDA.n353 14.363
R3747 GNDA.n235 GNDA.n233 14.0818
R3748 GNDA.n198 GNDA.n197 14.0193
R3749 GNDA.n2557 GNDA.n2556 14.0193
R3750 GNDA.n2342 GNDA.n2341 13.8005
R3751 GNDA.n2340 GNDA.n2339 13.8005
R3752 GNDA.n2378 GNDA.n2377 13.8005
R3753 GNDA.n2384 GNDA.n2383 13.8005
R3754 GNDA.n2435 GNDA.n2434 13.8005
R3755 GNDA.n147 GNDA.n146 13.8005
R3756 GNDA.n257 GNDA.n256 13.8005
R3757 GNDA.n271 GNDA.n61 13.8005
R3758 GNDA.n319 GNDA.n318 13.8005
R3759 GNDA.n330 GNDA.n329 13.8005
R3760 GNDA.n351 GNDA.n350 13.8005
R3761 GNDA.n2514 GNDA.n2 13.8005
R3762 GNDA.n2429 GNDA.n2428 12.7542
R3763 GNDA.n2309 GNDA.t194 12.3572
R3764 GNDA.t170 GNDA.n787 12.3572
R3765 GNDA.t162 GNDA.n671 12.3572
R3766 GNDA.t10 GNDA.t209 12.2992
R3767 GNDA.n877 GNDA.n380 12.2193
R3768 GNDA.n53 GNDA.n52 11.7557
R3769 GNDA.n1366 GNDA.n1364 11.6369
R3770 GNDA.n1364 GNDA.n1361 11.6369
R3771 GNDA.n1361 GNDA.n1360 11.6369
R3772 GNDA.n1360 GNDA.n1357 11.6369
R3773 GNDA.n1357 GNDA.n1356 11.6369
R3774 GNDA.n1356 GNDA.n1353 11.6369
R3775 GNDA.n1353 GNDA.n1352 11.6369
R3776 GNDA.n1352 GNDA.n1349 11.6369
R3777 GNDA.n1349 GNDA.n1348 11.6369
R3778 GNDA.n1348 GNDA.n1346 11.6369
R3779 GNDA.n2155 GNDA.n2154 11.6369
R3780 GNDA.n2154 GNDA.n2151 11.6369
R3781 GNDA.n2151 GNDA.n2150 11.6369
R3782 GNDA.n2150 GNDA.n2147 11.6369
R3783 GNDA.n2147 GNDA.n2146 11.6369
R3784 GNDA.n2146 GNDA.n2143 11.6369
R3785 GNDA.n2143 GNDA.n2142 11.6369
R3786 GNDA.n2142 GNDA.n2139 11.6369
R3787 GNDA.n2139 GNDA.n2138 11.6369
R3788 GNDA.n2138 GNDA.n441 11.6369
R3789 GNDA.n2371 GNDA.n441 11.6369
R3790 GNDA.n2173 GNDA.n2172 11.6369
R3791 GNDA.n2172 GNDA.n2171 11.6369
R3792 GNDA.n2171 GNDA.n2169 11.6369
R3793 GNDA.n2169 GNDA.n2166 11.6369
R3794 GNDA.n2166 GNDA.n2165 11.6369
R3795 GNDA.n2165 GNDA.n2162 11.6369
R3796 GNDA.n2162 GNDA.n2161 11.6369
R3797 GNDA.n2161 GNDA.n2158 11.6369
R3798 GNDA.n2158 GNDA.n2157 11.6369
R3799 GNDA.n2157 GNDA.n474 11.6369
R3800 GNDA.n962 GNDA.n961 11.6369
R3801 GNDA.n961 GNDA.n958 11.6369
R3802 GNDA.n958 GNDA.n957 11.6369
R3803 GNDA.n957 GNDA.n954 11.6369
R3804 GNDA.n954 GNDA.n953 11.6369
R3805 GNDA.n953 GNDA.n950 11.6369
R3806 GNDA.n950 GNDA.n949 11.6369
R3807 GNDA.n949 GNDA.n946 11.6369
R3808 GNDA.n946 GNDA.n945 11.6369
R3809 GNDA.n945 GNDA.n942 11.6369
R3810 GNDA.n966 GNDA.n965 11.6369
R3811 GNDA.n969 GNDA.n966 11.6369
R3812 GNDA.n970 GNDA.n969 11.6369
R3813 GNDA.n973 GNDA.n970 11.6369
R3814 GNDA.n974 GNDA.n973 11.6369
R3815 GNDA.n977 GNDA.n974 11.6369
R3816 GNDA.n978 GNDA.n977 11.6369
R3817 GNDA.n981 GNDA.n978 11.6369
R3818 GNDA.n983 GNDA.n981 11.6369
R3819 GNDA.n984 GNDA.n983 11.6369
R3820 GNDA.n2045 GNDA.n984 11.6369
R3821 GNDA.n1804 GNDA.n1803 11.6369
R3822 GNDA.n1805 GNDA.n1804 11.6369
R3823 GNDA.n1805 GNDA.n1061 11.6369
R3824 GNDA.n1812 GNDA.n1061 11.6369
R3825 GNDA.n1813 GNDA.n1812 11.6369
R3826 GNDA.n1814 GNDA.n1813 11.6369
R3827 GNDA.n1814 GNDA.n1058 11.6369
R3828 GNDA.n1821 GNDA.n1058 11.6369
R3829 GNDA.n1822 GNDA.n1821 11.6369
R3830 GNDA.n1823 GNDA.n1822 11.6369
R3831 GNDA.n1779 GNDA.n1778 11.6369
R3832 GNDA.n1782 GNDA.n1779 11.6369
R3833 GNDA.n1783 GNDA.n1782 11.6369
R3834 GNDA.n1786 GNDA.n1783 11.6369
R3835 GNDA.n1787 GNDA.n1786 11.6369
R3836 GNDA.n1790 GNDA.n1787 11.6369
R3837 GNDA.n1791 GNDA.n1790 11.6369
R3838 GNDA.n1794 GNDA.n1791 11.6369
R3839 GNDA.n1795 GNDA.n1794 11.6369
R3840 GNDA.n1798 GNDA.n1795 11.6369
R3841 GNDA.n1799 GNDA.n1798 11.6369
R3842 GNDA.n1724 GNDA.n985 11.6369
R3843 GNDA.n1727 GNDA.n1724 11.6369
R3844 GNDA.n1728 GNDA.n1727 11.6369
R3845 GNDA.n1731 GNDA.n1728 11.6369
R3846 GNDA.n1732 GNDA.n1731 11.6369
R3847 GNDA.n1735 GNDA.n1732 11.6369
R3848 GNDA.n1736 GNDA.n1735 11.6369
R3849 GNDA.n1739 GNDA.n1736 11.6369
R3850 GNDA.n1740 GNDA.n1739 11.6369
R3851 GNDA.n1743 GNDA.n1740 11.6369
R3852 GNDA.n1744 GNDA.n1743 11.6369
R3853 GNDA.n1685 GNDA.n1091 11.6369
R3854 GNDA.n1685 GNDA.n1684 11.6369
R3855 GNDA.n1684 GNDA.n1683 11.6369
R3856 GNDA.n1683 GNDA.n1092 11.6369
R3857 GNDA.n1677 GNDA.n1092 11.6369
R3858 GNDA.n1677 GNDA.n1676 11.6369
R3859 GNDA.n1676 GNDA.n1675 11.6369
R3860 GNDA.n1675 GNDA.n1095 11.6369
R3861 GNDA.n1669 GNDA.n1095 11.6369
R3862 GNDA.n1669 GNDA.n1668 11.6369
R3863 GNDA.n1668 GNDA.n1667 11.6369
R3864 GNDA.n1661 GNDA.n1100 11.6369
R3865 GNDA.n1661 GNDA.n1660 11.6369
R3866 GNDA.n1660 GNDA.n1659 11.6369
R3867 GNDA.n1659 GNDA.n1104 11.6369
R3868 GNDA.n1653 GNDA.n1104 11.6369
R3869 GNDA.n1653 GNDA.n1652 11.6369
R3870 GNDA.n1652 GNDA.n1651 11.6369
R3871 GNDA.n1651 GNDA.n1107 11.6369
R3872 GNDA.n1645 GNDA.n1107 11.6369
R3873 GNDA.n1645 GNDA.n1644 11.6369
R3874 GNDA.n647 GNDA.n646 11.6369
R3875 GNDA.n649 GNDA.n647 11.6369
R3876 GNDA.n649 GNDA.n648 11.6369
R3877 GNDA.n648 GNDA.n619 11.6369
R3878 GNDA.n619 GNDA.n617 11.6369
R3879 GNDA.n657 GNDA.n617 11.6369
R3880 GNDA.n658 GNDA.n657 11.6369
R3881 GNDA.n659 GNDA.n658 11.6369
R3882 GNDA.n659 GNDA.n612 11.6369
R3883 GNDA.n667 GNDA.n612 11.6369
R3884 GNDA.n622 GNDA.n559 11.6369
R3885 GNDA.n625 GNDA.n622 11.6369
R3886 GNDA.n626 GNDA.n625 11.6369
R3887 GNDA.n629 GNDA.n626 11.6369
R3888 GNDA.n630 GNDA.n629 11.6369
R3889 GNDA.n633 GNDA.n630 11.6369
R3890 GNDA.n634 GNDA.n633 11.6369
R3891 GNDA.n637 GNDA.n634 11.6369
R3892 GNDA.n638 GNDA.n637 11.6369
R3893 GNDA.n641 GNDA.n638 11.6369
R3894 GNDA.n642 GNDA.n641 11.6369
R3895 GNDA.n560 GNDA.n442 11.6369
R3896 GNDA.n563 GNDA.n560 11.6369
R3897 GNDA.n564 GNDA.n563 11.6369
R3898 GNDA.n567 GNDA.n564 11.6369
R3899 GNDA.n568 GNDA.n567 11.6369
R3900 GNDA.n571 GNDA.n568 11.6369
R3901 GNDA.n572 GNDA.n571 11.6369
R3902 GNDA.n575 GNDA.n572 11.6369
R3903 GNDA.n576 GNDA.n575 11.6369
R3904 GNDA.n579 GNDA.n576 11.6369
R3905 GNDA.n580 GNDA.n579 11.6369
R3906 GNDA.n1332 GNDA.n1331 11.6369
R3907 GNDA.n1331 GNDA.n1289 11.6369
R3908 GNDA.n1325 GNDA.n1289 11.6369
R3909 GNDA.n1325 GNDA.n1324 11.6369
R3910 GNDA.n1324 GNDA.n1323 11.6369
R3911 GNDA.n1317 GNDA.n1306 11.6369
R3912 GNDA.n1317 GNDA.n1316 11.6369
R3913 GNDA.n1316 GNDA.n1315 11.6369
R3914 GNDA.n1315 GNDA.n1307 11.6369
R3915 GNDA.n1309 GNDA.n1307 11.6369
R3916 GNDA.n1368 GNDA.n1367 11.6369
R3917 GNDA.n1368 GNDA.n1342 11.6369
R3918 GNDA.n1374 GNDA.n1342 11.6369
R3919 GNDA.n1375 GNDA.n1374 11.6369
R3920 GNDA.n1376 GNDA.n1375 11.6369
R3921 GNDA.n1376 GNDA.n1338 11.6369
R3922 GNDA.n1382 GNDA.n1338 11.6369
R3923 GNDA.n1383 GNDA.n1382 11.6369
R3924 GNDA.n1385 GNDA.n1383 11.6369
R3925 GNDA.n1385 GNDA.n1384 11.6369
R3926 GNDA.n1384 GNDA.n1335 11.6369
R3927 GNDA.t73 GNDA.n336 11.5188
R3928 GNDA.n230 GNDA.t149 11.5188
R3929 GNDA.n2434 GNDA.n2433 11.3792
R3930 GNDA.n2559 GNDA.n2558 10.2036
R3931 GNDA.n351 GNDA.n53 10.0943
R3932 GNDA.n377 GNDA.n0 9.75668
R3933 GNDA.n2226 GNDA.t152 9.6005
R3934 GNDA.n2216 GNDA.t154 9.6005
R3935 GNDA.n2419 GNDA.t86 9.6005
R3936 GNDA.n382 GNDA.t153 9.6005
R3937 GNDA.n217 GNDA.t287 9.6005
R3938 GNDA.n254 GNDA.t147 9.6005
R3939 GNDA.n254 GNDA.t122 9.6005
R3940 GNDA.n252 GNDA.t158 9.6005
R3941 GNDA.n252 GNDA.t72 9.6005
R3942 GNDA.n250 GNDA.t144 9.6005
R3943 GNDA.n250 GNDA.t316 9.6005
R3944 GNDA.n248 GNDA.t43 9.6005
R3945 GNDA.n248 GNDA.t107 9.6005
R3946 GNDA.n246 GNDA.t111 9.6005
R3947 GNDA.n246 GNDA.t138 9.6005
R3948 GNDA.n244 GNDA.t305 9.6005
R3949 GNDA.n244 GNDA.t41 9.6005
R3950 GNDA.n242 GNDA.t74 9.6005
R3951 GNDA.n242 GNDA.t82 9.6005
R3952 GNDA.n240 GNDA.t303 9.6005
R3953 GNDA.n240 GNDA.t156 9.6005
R3954 GNDA.n238 GNDA.t296 9.6005
R3955 GNDA.n238 GNDA.t80 9.6005
R3956 GNDA.n236 GNDA.t45 9.6005
R3957 GNDA.n236 GNDA.t5 9.6005
R3958 GNDA.n234 GNDA.t307 9.6005
R3959 GNDA.n234 GNDA.t239 9.6005
R3960 GNDA.n223 GNDA.t240 9.6005
R3961 GNDA.n340 GNDA.t293 9.6005
R3962 GNDA.n352 GNDA.t117 9.6005
R3963 GNDA.n352 GNDA.t37 9.6005
R3964 GNDA.n41 GNDA.t267 9.6005
R3965 GNDA.t2 GNDA.t209 9.37093
R3966 GNDA.n116 GNDA.n113 9.14336
R3967 GNDA.n120 GNDA.n113 9.14336
R3968 GNDA.n120 GNDA.n111 9.14336
R3969 GNDA.n126 GNDA.n111 9.14336
R3970 GNDA.n126 GNDA.n109 9.14336
R3971 GNDA.n130 GNDA.n109 9.14336
R3972 GNDA.n130 GNDA.n107 9.14336
R3973 GNDA.n136 GNDA.n107 9.14336
R3974 GNDA.n136 GNDA.n105 9.14336
R3975 GNDA.n140 GNDA.n105 9.14336
R3976 GNDA.n140 GNDA.n103 9.14336
R3977 GNDA.n265 GNDA.n264 9.14336
R3978 GNDA.n262 GNDA.n261 9.14336
R3979 GNDA.n228 GNDA.n227 9.14336
R3980 GNDA.n225 GNDA.n224 9.14336
R3981 GNDA.n285 GNDA.n283 9.14336
R3982 GNDA.n205 GNDA.n76 9.14336
R3983 GNDA.n205 GNDA.n204 9.14336
R3984 GNDA.n204 GNDA.n202 9.14336
R3985 GNDA.n187 GNDA.n182 9.14336
R3986 GNDA.n187 GNDA.n186 9.14336
R3987 GNDA.n186 GNDA.n184 9.14336
R3988 GNDA.n275 GNDA.n274 9.14336
R3989 GNDA.n313 GNDA.n312 9.14336
R3990 GNDA.n334 GNDA.n333 9.14336
R3991 GNDA.n323 GNDA.n321 9.14336
R3992 GNDA.n345 GNDA.n344 9.14336
R3993 GNDA.n342 GNDA.n341 9.14336
R3994 GNDA.n362 GNDA.n361 9.14336
R3995 GNDA.n359 GNDA.n358 9.14336
R3996 GNDA.n2549 GNDA.n2544 9.14336
R3997 GNDA.n2549 GNDA.n2548 9.14336
R3998 GNDA.n2548 GNDA.n2546 9.14336
R3999 GNDA.n2453 GNDA.n2445 9.14336
R4000 GNDA.n2453 GNDA.n2452 9.14336
R4001 GNDA.n2452 GNDA.n2450 9.14336
R4002 GNDA.n2537 GNDA.n2504 9.14336
R4003 GNDA.n2537 GNDA.n2536 9.14336
R4004 GNDA.n2536 GNDA.n2534 9.14336
R4005 GNDA.n2534 GNDA.n2531 9.14336
R4006 GNDA.n2531 GNDA.n2530 9.14336
R4007 GNDA.n2530 GNDA.n2527 9.14336
R4008 GNDA.n2527 GNDA.n2526 9.14336
R4009 GNDA.n2526 GNDA.n2523 9.14336
R4010 GNDA.n2523 GNDA.n2522 9.14336
R4011 GNDA.n2522 GNDA.n2519 9.14336
R4012 GNDA.n2519 GNDA.n2518 9.14336
R4013 GNDA.n2497 GNDA.n2460 9.14336
R4014 GNDA.n2497 GNDA.n2496 9.14336
R4015 GNDA.n2496 GNDA.n2494 9.14336
R4016 GNDA.n2494 GNDA.n2491 9.14336
R4017 GNDA.n2491 GNDA.n2490 9.14336
R4018 GNDA.n2490 GNDA.n2487 9.14336
R4019 GNDA.n2487 GNDA.n2486 9.14336
R4020 GNDA.n2486 GNDA.n2483 9.14336
R4021 GNDA.n2483 GNDA.n2482 9.14336
R4022 GNDA.n2482 GNDA.n2479 9.14336
R4023 GNDA.n2479 GNDA.n2478 9.14336
R4024 GNDA.n175 GNDA.n92 9.14336
R4025 GNDA.n175 GNDA.n174 9.14336
R4026 GNDA.n174 GNDA.n172 9.14336
R4027 GNDA.n172 GNDA.n169 9.14336
R4028 GNDA.n169 GNDA.n168 9.14336
R4029 GNDA.n168 GNDA.n165 9.14336
R4030 GNDA.n165 GNDA.n164 9.14336
R4031 GNDA.n164 GNDA.n161 9.14336
R4032 GNDA.n161 GNDA.n160 9.14336
R4033 GNDA.n160 GNDA.n157 9.14336
R4034 GNDA.n157 GNDA.n156 9.14336
R4035 GNDA.n2059 GNDA.n2058 8.60107
R4036 GNDA.n1113 GNDA.n1067 8.60107
R4037 GNDA.n212 GNDA.n211 8.53383
R4038 GNDA.t166 GNDA.n2310 8.23827
R4039 GNDA.t180 GNDA.n864 8.23827
R4040 GNDA.t174 GNDA.n2414 8.23827
R4041 GNDA.n2438 GNDA.n373 8.19962
R4042 GNDA.t251 GNDA.t110 7.67938
R4043 GNDA.t35 GNDA.t137 7.67938
R4044 GNDA.n337 GNDA.t20 7.67938
R4045 GNDA.t70 GNDA.t304 7.67938
R4046 GNDA.t283 GNDA.t40 7.67938
R4047 GNDA.n379 GNDA.n378 7.56675
R4048 GNDA.n1298 GNDA.n377 7.56675
R4049 GNDA.t139 GNDA.n2243 7.20855
R4050 GNDA.n2391 GNDA.t148 7.20855
R4051 GNDA.t15 GNDA.n678 7.20855
R4052 GNDA.n2437 GNDA.n374 7.20855
R4053 GNDA.n256 GNDA.n218 7.03175
R4054 GNDA.n2371 GNDA.n2370 6.72373
R4055 GNDA.n2045 GNDA.n2044 6.72373
R4056 GNDA.n1744 GNDA.n1722 6.72373
R4057 GNDA.n908 GNDA.n580 6.72373
R4058 GNDA.n1309 GNDA.n1308 6.72373
R4059 GNDA.n1335 GNDA.n1333 6.72373
R4060 GNDA.n2560 GNDA.n2559 6.28175
R4061 GNDA.n2560 GNDA.n1 6.28175
R4062 GNDA.n1778 GNDA.n1722 6.20656
R4063 GNDA.n2044 GNDA.n985 6.20656
R4064 GNDA.n1308 GNDA.n1091 6.20656
R4065 GNDA.n908 GNDA.n559 6.20656
R4066 GNDA.n2370 GNDA.n442 6.20656
R4067 GNDA.n1333 GNDA.n1332 6.20656
R4068 GNDA.t209 GNDA.t50 6.17883
R4069 GNDA.n1323 GNDA.n1294 6.07727
R4070 GNDA.n218 GNDA.n1 6.063
R4071 GNDA.n2227 GNDA.n2217 5.81868
R4072 GNDA.n2220 GNDA.n2217 5.81868
R4073 GNDA.n145 GNDA.n102 5.78934
R4074 GNDA.n200 GNDA.n199 5.78934
R4075 GNDA.n193 GNDA.n78 5.78934
R4076 GNDA.n2555 GNDA.n15 5.78934
R4077 GNDA.n2448 GNDA.n2447 5.78934
R4078 GNDA.n2516 GNDA.n2515 5.78934
R4079 GNDA.n2476 GNDA.n2475 5.78934
R4080 GNDA.n154 GNDA.n153 5.78934
R4081 GNDA.n379 GNDA.n0 5.737
R4082 GNDA.n1306 GNDA.n1294 5.5601
R4083 GNDA.n197 GNDA.n196 5.54068
R4084 GNDA.n2558 GNDA.n2557 5.54068
R4085 GNDA.n1450 GNDA.n1428 5.51161
R4086 GNDA.n2251 GNDA.n2210 5.51161
R4087 GNDA.n2067 GNDA.n515 5.51161
R4088 GNDA.n1956 GNDA.n1926 5.51161
R4089 GNDA.n1861 GNDA.n1831 5.51161
R4090 GNDA.n1210 GNDA.n1180 5.51161
R4091 GNDA.n1633 GNDA.n1632 5.51161
R4092 GNDA.n805 GNDA.n776 5.51161
R4093 GNDA.n685 GNDA.n607 5.51161
R4094 GNDA.n281 GNDA.n68 5.46925
R4095 GNDA.n195 GNDA.n61 5.46925
R4096 GNDA.n1830 GNDA.n1054 5.1717
R4097 GNDA.n1643 GNDA.n1112 5.1717
R4098 GNDA.n669 GNDA.n668 5.1717
R4099 GNDA.n786 GNDA.t209 5.14911
R4100 GNDA.t276 GNDA.t96 5.14911
R4101 GNDA.n52 GNDA.n50 5.063
R4102 GNDA.n13 GNDA.n11 5.063
R4103 GNDA.n1514 GNDA.n1128 4.9157
R4104 GNDA.n2320 GNDA.n2179 4.9157
R4105 GNDA.n2128 GNDA.n492 4.9157
R4106 GNDA.n264 GNDA.n263 4.46219
R4107 GNDA.n261 GNDA.n259 4.46219
R4108 GNDA.n263 GNDA.n262 4.46219
R4109 GNDA.n259 GNDA.n258 4.46219
R4110 GNDA.n227 GNDA.n226 4.46219
R4111 GNDA.n224 GNDA.n219 4.46219
R4112 GNDA.n226 GNDA.n225 4.46219
R4113 GNDA.n232 GNDA.n219 4.46219
R4114 GNDA.n283 GNDA.n282 4.46219
R4115 GNDA.n289 GNDA.n282 4.46219
R4116 GNDA.n274 GNDA.n273 4.46219
R4117 GNDA.n273 GNDA.n272 4.46219
R4118 GNDA.n312 GNDA.n62 4.46219
R4119 GNDA.n317 GNDA.n62 4.46219
R4120 GNDA.n333 GNDA.n332 4.46219
R4121 GNDA.n332 GNDA.n331 4.46219
R4122 GNDA.n321 GNDA.n320 4.46219
R4123 GNDA.n327 GNDA.n320 4.46219
R4124 GNDA.n344 GNDA.n343 4.46219
R4125 GNDA.n341 GNDA.n54 4.46219
R4126 GNDA.n343 GNDA.n342 4.46219
R4127 GNDA.n349 GNDA.n54 4.46219
R4128 GNDA.n361 GNDA.n360 4.46219
R4129 GNDA.n358 GNDA.n356 4.46219
R4130 GNDA.n360 GNDA.n359 4.46219
R4131 GNDA.n356 GNDA.n355 4.46219
R4132 GNDA.n1693 GNDA.n1086 4.26717
R4133 GNDA.n1693 GNDA.n1082 4.26717
R4134 GNDA.n1699 GNDA.n1082 4.26717
R4135 GNDA.n1700 GNDA.n1699 4.26717
R4136 GNDA.n1700 GNDA.n1079 4.26717
R4137 GNDA.n1079 GNDA.n1077 4.26717
R4138 GNDA.n1708 GNDA.n1077 4.26717
R4139 GNDA.n1708 GNDA.n1073 4.26717
R4140 GNDA.n1714 GNDA.n1073 4.26717
R4141 GNDA.n1715 GNDA.n1714 4.26717
R4142 GNDA.n1715 GNDA.n1070 4.26717
R4143 GNDA.n907 GNDA.n583 4.26717
R4144 GNDA.n902 GNDA.n583 4.26717
R4145 GNDA.n902 GNDA.n901 4.26717
R4146 GNDA.n901 GNDA.n591 4.26717
R4147 GNDA.n896 GNDA.n591 4.26717
R4148 GNDA.n896 GNDA.n895 4.26717
R4149 GNDA.n895 GNDA.n894 4.26717
R4150 GNDA.n894 GNDA.n599 4.26717
R4151 GNDA.n888 GNDA.n599 4.26717
R4152 GNDA.n888 GNDA.n887 4.26717
R4153 GNDA.n887 GNDA.n886 4.26717
R4154 GNDA.n1775 GNDA.n1774 4.26717
R4155 GNDA.n1774 GNDA.n1749 4.26717
R4156 GNDA.n1769 GNDA.n1749 4.26717
R4157 GNDA.n1769 GNDA.n1768 4.26717
R4158 GNDA.n1768 GNDA.n1767 4.26717
R4159 GNDA.n1767 GNDA.n1755 4.26717
R4160 GNDA.n1761 GNDA.n1755 4.26717
R4161 GNDA.n1761 GNDA.n1760 4.26717
R4162 GNDA.n1760 GNDA.n914 4.26717
R4163 GNDA.n2053 GNDA.n914 4.26717
R4164 GNDA.n2053 GNDA.n911 4.26717
R4165 GNDA.n1392 GNDA.n1285 4.26717
R4166 GNDA.n1398 GNDA.n1285 4.26717
R4167 GNDA.n1399 GNDA.n1398 4.26717
R4168 GNDA.n1402 GNDA.n1399 4.26717
R4169 GNDA.n1402 GNDA.n1283 4.26717
R4170 GNDA.n1408 GNDA.n1283 4.26717
R4171 GNDA.n1408 GNDA.n1277 4.26717
R4172 GNDA.n1416 GNDA.n1277 4.26717
R4173 GNDA.n1416 GNDA.n1275 4.26717
R4174 GNDA.n1275 GNDA.n1156 4.26717
R4175 GNDA.n1423 GNDA.n1156 4.26717
R4176 GNDA.n2043 GNDA.n987 4.26717
R4177 GNDA.n2038 GNDA.n987 4.26717
R4178 GNDA.n2038 GNDA.n2037 4.26717
R4179 GNDA.n2037 GNDA.n995 4.26717
R4180 GNDA.n2032 GNDA.n995 4.26717
R4181 GNDA.n2032 GNDA.n2031 4.26717
R4182 GNDA.n2031 GNDA.n2030 4.26717
R4183 GNDA.n2030 GNDA.n1003 4.26717
R4184 GNDA.n2024 GNDA.n1003 4.26717
R4185 GNDA.n2024 GNDA.n2023 4.26717
R4186 GNDA.n2023 GNDA.n2022 4.26717
R4187 GNDA.n2369 GNDA.n444 4.26717
R4188 GNDA.n2364 GNDA.n444 4.26717
R4189 GNDA.n2364 GNDA.n2363 4.26717
R4190 GNDA.n2363 GNDA.n452 4.26717
R4191 GNDA.n2358 GNDA.n452 4.26717
R4192 GNDA.n2358 GNDA.n2357 4.26717
R4193 GNDA.n2357 GNDA.n2356 4.26717
R4194 GNDA.n2356 GNDA.n460 4.26717
R4195 GNDA.n2350 GNDA.n460 4.26717
R4196 GNDA.n2350 GNDA.n2349 4.26717
R4197 GNDA.n2349 GNDA.n2348 4.26717
R4198 GNDA.n302 GNDA.n281 4.2505
R4199 GNDA GNDA.n2561 4.2117
R4200 GNDA.n211 GNDA.n69 4.17148
R4201 GNDA.n279 GNDA.n69 4.17148
R4202 GNDA.n2428 GNDA.n380 4.063
R4203 GNDA.n319 GNDA.n61 4.0005
R4204 GNDA.n1308 GNDA.n1086 3.93531
R4205 GNDA.n908 GNDA.n907 3.93531
R4206 GNDA.n1775 GNDA.n1722 3.93531
R4207 GNDA.n1392 GNDA.n1333 3.93531
R4208 GNDA.n2044 GNDA.n2043 3.93531
R4209 GNDA.n2370 GNDA.n2369 3.93531
R4210 GNDA.t280 GNDA.t101 3.83994
R4211 GNDA.t30 GNDA.t270 3.83994
R4212 GNDA.t260 GNDA.t113 3.83994
R4213 GNDA.t299 GNDA.t247 3.83994
R4214 GNDA.n1512 GNDA.n1511 3.7893
R4215 GNDA.n1508 GNDA.n1131 3.7893
R4216 GNDA.n1507 GNDA.n1134 3.7893
R4217 GNDA.n1504 GNDA.n1503 3.7893
R4218 GNDA.n1430 GNDA.n1135 3.7893
R4219 GNDA.n1439 GNDA.n1438 3.7893
R4220 GNDA.n1442 GNDA.n1429 3.7893
R4221 GNDA.n1447 GNDA.n1443 3.7893
R4222 GNDA.n2318 GNDA.n2317 3.7893
R4223 GNDA.n2314 GNDA.n2181 3.7893
R4224 GNDA.n2313 GNDA.n2184 3.7893
R4225 GNDA.n2191 GNDA.n2190 3.7893
R4226 GNDA.n2307 GNDA.n2306 3.7893
R4227 GNDA.n2236 GNDA.n2235 3.7893
R4228 GNDA.n2240 GNDA.n2239 3.7893
R4229 GNDA.n2248 GNDA.n2211 3.7893
R4230 GNDA.n2126 GNDA.n494 3.7893
R4231 GNDA.n2123 GNDA.n2122 3.7893
R4232 GNDA.n535 GNDA.n496 3.7893
R4233 GNDA.n553 GNDA.n552 3.7893
R4234 GNDA.n550 GNDA.n549 3.7893
R4235 GNDA.n545 GNDA.n538 3.7893
R4236 GNDA.n542 GNDA.n541 3.7893
R4237 GNDA.n2064 GNDA.n516 3.7893
R4238 GNDA.n2015 GNDA.n1013 3.7893
R4239 GNDA.n2012 GNDA.n2011 3.7893
R4240 GNDA.n1928 GNDA.n1014 3.7893
R4241 GNDA.n1933 GNDA.n1931 3.7893
R4242 GNDA.n1938 GNDA.n1934 3.7893
R4243 GNDA.n1945 GNDA.n1944 3.7893
R4244 GNDA.n1948 GNDA.n1927 3.7893
R4245 GNDA.n1953 GNDA.n1949 3.7893
R4246 GNDA.n1920 GNDA.n1034 3.7893
R4247 GNDA.n1917 GNDA.n1916 3.7893
R4248 GNDA.n1833 GNDA.n1035 3.7893
R4249 GNDA.n1838 GNDA.n1836 3.7893
R4250 GNDA.n1843 GNDA.n1839 3.7893
R4251 GNDA.n1850 GNDA.n1849 3.7893
R4252 GNDA.n1853 GNDA.n1832 3.7893
R4253 GNDA.n1858 GNDA.n1854 3.7893
R4254 GNDA.n1595 GNDA.n1532 3.7893
R4255 GNDA.n1604 GNDA.n1603 3.7893
R4256 GNDA.n1529 GNDA.n1528 3.7893
R4257 GNDA.n1612 GNDA.n1610 3.7893
R4258 GNDA.n1611 GNDA.n1526 3.7893
R4259 GNDA.n1524 GNDA.n1523 3.7893
R4260 GNDA.n1627 GNDA.n1625 3.7893
R4261 GNDA.n1626 GNDA.n1519 3.7893
R4262 GNDA.n1269 GNDA.n1158 3.7893
R4263 GNDA.n1266 GNDA.n1265 3.7893
R4264 GNDA.n1182 GNDA.n1159 3.7893
R4265 GNDA.n1187 GNDA.n1185 3.7893
R4266 GNDA.n1192 GNDA.n1188 3.7893
R4267 GNDA.n1199 GNDA.n1198 3.7893
R4268 GNDA.n1202 GNDA.n1181 3.7893
R4269 GNDA.n1207 GNDA.n1203 3.7893
R4270 GNDA.n873 GNDA.n872 3.7893
R4271 GNDA.n869 GNDA.n750 3.7893
R4272 GNDA.n868 GNDA.n753 3.7893
R4273 GNDA.n758 GNDA.n757 3.7893
R4274 GNDA.n862 GNDA.n861 3.7893
R4275 GNDA.n794 GNDA.n793 3.7893
R4276 GNDA.n790 GNDA.n777 3.7893
R4277 GNDA.n802 GNDA.n800 3.7893
R4278 GNDA.n2406 GNDA.n411 3.7893
R4279 GNDA.n2405 GNDA.n412 3.7893
R4280 GNDA.n2393 GNDA.n2392 3.7893
R4281 GNDA.n2399 GNDA.n2398 3.7893
R4282 GNDA.n2395 GNDA.n2394 3.7893
R4283 GNDA.n672 GNDA.n390 3.7893
R4284 GNDA.n675 GNDA.n674 3.7893
R4285 GNDA.n682 GNDA.n608 3.7893
R4286 GNDA.n1435 GNDA 3.7381
R4287 GNDA.n2234 GNDA 3.7381
R4288 GNDA.n546 GNDA 3.7381
R4289 GNDA.n1941 GNDA 3.7381
R4290 GNDA.n1846 GNDA 3.7381
R4291 GNDA GNDA.n1618 3.7381
R4292 GNDA.n1195 GNDA 3.7381
R4293 GNDA.n789 GNDA 3.7381
R4294 GNDA GNDA.n2411 3.7381
R4295 GNDA.n2433 GNDA.n377 3.51962
R4296 GNDA.n150 GNDA.t58 3.42907
R4297 GNDA.n150 GNDA.t23 3.42907
R4298 GNDA.n148 GNDA.t56 3.42907
R4299 GNDA.n148 GNDA.t312 3.42907
R4300 GNDA.n2470 GNDA.t19 3.42907
R4301 GNDA.n2470 GNDA.t318 3.42907
R4302 GNDA.n2472 GNDA.t28 3.42907
R4303 GNDA.n2472 GNDA.t78 3.42907
R4304 GNDA.n117 GNDA.n116 3.19754
R4305 GNDA.n103 GNDA.n102 3.19754
R4306 GNDA.n207 GNDA.n76 3.19754
R4307 GNDA.n202 GNDA.n200 3.19754
R4308 GNDA.n189 GNDA.n182 3.19754
R4309 GNDA.n184 GNDA.n78 3.19754
R4310 GNDA.n2551 GNDA.n2544 3.19754
R4311 GNDA.n2546 GNDA.n15 3.19754
R4312 GNDA.n2455 GNDA.n2445 3.19754
R4313 GNDA.n2450 GNDA.n2448 3.19754
R4314 GNDA.n2539 GNDA.n2504 3.19754
R4315 GNDA.n2518 GNDA.n2516 3.19754
R4316 GNDA.n2499 GNDA.n2460 3.19754
R4317 GNDA.n2478 GNDA.n2476 3.19754
R4318 GNDA.n177 GNDA.n92 3.19754
R4319 GNDA.n156 GNDA.n154 3.19754
R4320 GNDA.n2323 GNDA.n2322 3.08966
R4321 GNDA.n2188 GNDA.t9 3.08966
R4322 GNDA.n2230 GNDA.t123 3.08966
R4323 GNDA.n2245 GNDA.t12 3.08966
R4324 GNDA.n2403 GNDA.t127 3.08966
R4325 GNDA.n2421 GNDA.n381 2.86505
R4326 GNDA.n2422 GNDA.n2421 2.86505
R4327 GNDA.n2420 GNDA.n2416 2.86505
R4328 GNDA.n2417 GNDA.n2416 2.86505
R4329 GNDA.n2423 GNDA.n2422 2.86505
R4330 GNDA.n2418 GNDA.n2417 2.86505
R4331 GNDA.n2427 GNDA.n381 2.86505
R4332 GNDA.n2423 GNDA.n2420 2.86505
R4333 GNDA.n305 GNDA.n304 2.86505
R4334 GNDA.n308 GNDA.n304 2.86505
R4335 GNDA.n309 GNDA.n308 2.86505
R4336 GNDA.n306 GNDA.n305 2.86505
R4337 GNDA.n294 GNDA.n293 2.86505
R4338 GNDA.n297 GNDA.n293 2.86505
R4339 GNDA.n298 GNDA.n297 2.86505
R4340 GNDA.n295 GNDA.n294 2.86505
R4341 GNDA.n2223 GNDA.n2219 2.86505
R4342 GNDA.n2224 GNDA.n2223 2.86505
R4343 GNDA.n2225 GNDA.n2224 2.86505
R4344 GNDA.n2220 GNDA.n2219 2.86505
R4345 GNDA.n1514 GNDA.n1513 2.6629
R4346 GNDA.n1427 GNDA.n1154 2.6629
R4347 GNDA.n2320 GNDA.n2319 2.6629
R4348 GNDA.n2209 GNDA.n468 2.6629
R4349 GNDA.n2128 GNDA.n2127 2.6629
R4350 GNDA.n2019 GNDA.n1011 2.6629
R4351 GNDA.n2018 GNDA.n2016 2.6629
R4352 GNDA.n1925 GNDA.n1923 2.6629
R4353 GNDA.n1922 GNDA.n1921 2.6629
R4354 GNDA.n1596 GNDA.n1594 2.6629
R4355 GNDA.n1271 GNDA.n1270 2.6629
R4356 GNDA.n1179 GNDA.n1065 2.6629
R4357 GNDA.n749 GNDA.n748 2.6629
R4358 GNDA.n741 GNDA.n739 2.6629
R4359 GNDA.n738 GNDA.n737 2.6629
R4360 GNDA.n218 GNDA.n68 2.53175
R4361 GNDA.n195 GNDA.n53 2.5005
R4362 GNDA.n1428 GNDA.n1427 2.4581
R4363 GNDA.n2210 GNDA.n2209 2.4581
R4364 GNDA.n1011 GNDA.n515 2.4581
R4365 GNDA.n2019 GNDA.n2018 2.4581
R4366 GNDA.n1926 GNDA.n1925 2.4581
R4367 GNDA.n1923 GNDA.n1922 2.4581
R4368 GNDA.n1831 GNDA.n1830 2.4581
R4369 GNDA.n1594 GNDA.n1065 2.4581
R4370 GNDA.n1633 GNDA.n1112 2.4581
R4371 GNDA.n1271 GNDA.n1154 2.4581
R4372 GNDA.n1180 GNDA.n1179 2.4581
R4373 GNDA.n748 GNDA.n468 2.4581
R4374 GNDA.n776 GNDA.n741 2.4581
R4375 GNDA.n739 GNDA.n738 2.4581
R4376 GNDA.n669 GNDA.n607 2.4581
R4377 GNDA.n329 GNDA.n319 2.2505
R4378 GNDA.n1070 GNDA.n1065 2.18124
R4379 GNDA.n886 GNDA.n739 2.18124
R4380 GNDA.n1923 GNDA.n911 2.18124
R4381 GNDA.n1423 GNDA.n1154 2.18124
R4382 GNDA.n2022 GNDA.n2019 2.18124
R4383 GNDA.n2348 GNDA.n468 2.18124
R4384 GNDA.n1446 GNDA.n1428 2.1509
R4385 GNDA.n2247 GNDA.n2210 2.1509
R4386 GNDA.n2063 GNDA.n515 2.1509
R4387 GNDA.n1952 GNDA.n1926 2.1509
R4388 GNDA.n1857 GNDA.n1831 2.1509
R4389 GNDA.n1634 GNDA.n1633 2.1509
R4390 GNDA.n1206 GNDA.n1180 2.1509
R4391 GNDA.n801 GNDA.n776 2.1509
R4392 GNDA.n681 GNDA.n607 2.1509
R4393 GNDA.n1513 GNDA.n1129 2.13383
R4394 GNDA.n2319 GNDA.n2180 2.13383
R4395 GNDA.n2127 GNDA.n493 2.13383
R4396 GNDA.n2016 GNDA.n1012 2.13383
R4397 GNDA.n1921 GNDA.n1033 2.13383
R4398 GNDA.n1270 GNDA.n1157 2.13383
R4399 GNDA.n1597 GNDA.n1596 2.13383
R4400 GNDA.n841 GNDA.n749 2.13383
R4401 GNDA.n737 GNDA.n736 2.13383
R4402 GNDA.n2429 GNDA 2.09787
R4403 GNDA.n1721 GNDA.n1065 2.08643
R4404 GNDA.n882 GNDA.n739 2.08643
R4405 GNDA.n1923 GNDA.n909 2.08643
R4406 GNDA.n1154 GNDA.n986 2.08643
R4407 GNDA.n2019 GNDA.n443 2.08643
R4408 GNDA.n471 GNDA.n468 2.08643
R4409 GNDA.n2245 GNDA.t215 2.05994
R4410 GNDA.n745 GNDA.t289 2.05994
R4411 GNDA.n879 GNDA.t254 2.05994
R4412 GNDA.n2388 GNDA.t276 2.05994
R4413 GNDA.n196 GNDA.n195 2.0005
R4414 GNDA.n1513 GNDA.n1512 1.9461
R4415 GNDA.n2319 GNDA.n2318 1.9461
R4416 GNDA.n2127 GNDA.n2126 1.9461
R4417 GNDA.n2016 GNDA.n2015 1.9461
R4418 GNDA.n1921 GNDA.n1920 1.9461
R4419 GNDA.n1596 GNDA.n1595 1.9461
R4420 GNDA.n1270 GNDA.n1269 1.9461
R4421 GNDA.n873 GNDA.n749 1.9461
R4422 GNDA.n737 GNDA.n411 1.9461
R4423 GNDA.n1299 GNDA.n1298 1.90675
R4424 GNDA.t151 GNDA.n476 1.83728
R4425 GNDA.n302 GNDA.n301 1.7505
R4426 GNDA.n1346 GNDA.n1128 1.47392
R4427 GNDA.n2179 GNDA.n474 1.47392
R4428 GNDA.n942 GNDA.n492 1.47392
R4429 GNDA.n1823 GNDA.n1054 1.47392
R4430 GNDA.n1644 GNDA.n1643 1.47392
R4431 GNDA.n668 GNDA.n667 1.47392
R4432 GNDA.n196 GNDA.n68 1.35988
R4433 GNDA.n2559 GNDA.n2 1.28175
R4434 GNDA.n147 GNDA.n1 1.28175
R4435 GNDA.n2473 GNDA.n2471 1.1255
R4436 GNDA.n2471 GNDA.n2 1.1255
R4437 GNDA.n149 GNDA.n147 1.1255
R4438 GNDA.n151 GNDA.n149 1.1255
R4439 GNDA.n2383 GNDA.n2378 0.96925
R4440 GNDA.n2341 GNDA.n2340 0.96925
R4441 GNDA.n1511 GNDA.n1131 0.8197
R4442 GNDA.n1508 GNDA.n1507 0.8197
R4443 GNDA.n1504 GNDA.n1134 0.8197
R4444 GNDA.n1503 GNDA.n1135 0.8197
R4445 GNDA.n1438 GNDA.n1435 0.8197
R4446 GNDA.n1439 GNDA.n1429 0.8197
R4447 GNDA.n1443 GNDA.n1442 0.8197
R4448 GNDA.n1447 GNDA.n1446 0.8197
R4449 GNDA.n2317 GNDA.n2181 0.8197
R4450 GNDA.n2314 GNDA.n2313 0.8197
R4451 GNDA.n2190 GNDA.n2184 0.8197
R4452 GNDA.n2307 GNDA.n2191 0.8197
R4453 GNDA.n2235 GNDA.n2234 0.8197
R4454 GNDA.n2240 GNDA.n2236 0.8197
R4455 GNDA.n2239 GNDA.n2211 0.8197
R4456 GNDA.n2248 GNDA.n2247 0.8197
R4457 GNDA.n2123 GNDA.n494 0.8197
R4458 GNDA.n2122 GNDA.n496 0.8197
R4459 GNDA.n553 GNDA.n535 0.8197
R4460 GNDA.n552 GNDA.n550 0.8197
R4461 GNDA.n546 GNDA.n545 0.8197
R4462 GNDA.n542 GNDA.n538 0.8197
R4463 GNDA.n541 GNDA.n516 0.8197
R4464 GNDA.n2064 GNDA.n2063 0.8197
R4465 GNDA.n2012 GNDA.n1013 0.8197
R4466 GNDA.n2011 GNDA.n1014 0.8197
R4467 GNDA.n1931 GNDA.n1928 0.8197
R4468 GNDA.n1934 GNDA.n1933 0.8197
R4469 GNDA.n1944 GNDA.n1941 0.8197
R4470 GNDA.n1945 GNDA.n1927 0.8197
R4471 GNDA.n1949 GNDA.n1948 0.8197
R4472 GNDA.n1953 GNDA.n1952 0.8197
R4473 GNDA.n1917 GNDA.n1034 0.8197
R4474 GNDA.n1916 GNDA.n1035 0.8197
R4475 GNDA.n1836 GNDA.n1833 0.8197
R4476 GNDA.n1839 GNDA.n1838 0.8197
R4477 GNDA.n1849 GNDA.n1846 0.8197
R4478 GNDA.n1850 GNDA.n1832 0.8197
R4479 GNDA.n1854 GNDA.n1853 0.8197
R4480 GNDA.n1858 GNDA.n1857 0.8197
R4481 GNDA.n1604 GNDA.n1532 0.8197
R4482 GNDA.n1603 GNDA.n1529 0.8197
R4483 GNDA.n1610 GNDA.n1528 0.8197
R4484 GNDA.n1612 GNDA.n1611 0.8197
R4485 GNDA.n1618 GNDA.n1524 0.8197
R4486 GNDA.n1625 GNDA.n1523 0.8197
R4487 GNDA.n1627 GNDA.n1626 0.8197
R4488 GNDA.n1634 GNDA.n1519 0.8197
R4489 GNDA.n1266 GNDA.n1158 0.8197
R4490 GNDA.n1265 GNDA.n1159 0.8197
R4491 GNDA.n1185 GNDA.n1182 0.8197
R4492 GNDA.n1188 GNDA.n1187 0.8197
R4493 GNDA.n1198 GNDA.n1195 0.8197
R4494 GNDA.n1199 GNDA.n1181 0.8197
R4495 GNDA.n1203 GNDA.n1202 0.8197
R4496 GNDA.n1207 GNDA.n1206 0.8197
R4497 GNDA.n872 GNDA.n750 0.8197
R4498 GNDA.n869 GNDA.n868 0.8197
R4499 GNDA.n757 GNDA.n753 0.8197
R4500 GNDA.n862 GNDA.n758 0.8197
R4501 GNDA.n794 GNDA.n789 0.8197
R4502 GNDA.n793 GNDA.n790 0.8197
R4503 GNDA.n800 GNDA.n777 0.8197
R4504 GNDA.n802 GNDA.n801 0.8197
R4505 GNDA.n2406 GNDA.n2405 0.8197
R4506 GNDA.n2392 GNDA.n412 0.8197
R4507 GNDA.n2399 GNDA.n2393 0.8197
R4508 GNDA.n2398 GNDA.n2395 0.8197
R4509 GNDA.n2411 GNDA.n390 0.8197
R4510 GNDA.n675 GNDA.n672 0.8197
R4511 GNDA.n674 GNDA.n608 0.8197
R4512 GNDA.n682 GNDA.n681 0.8197
R4513 GNDA.n2176 GNDA.n476 0.575776
R4514 GNDA GNDA.n1430 0.5637
R4515 GNDA.n2306 GNDA 0.5637
R4516 GNDA.n549 GNDA 0.5637
R4517 GNDA.n1938 GNDA 0.5637
R4518 GNDA.n1843 GNDA 0.5637
R4519 GNDA.n1526 GNDA 0.5637
R4520 GNDA.n1192 GNDA 0.5637
R4521 GNDA.n861 GNDA 0.5637
R4522 GNDA.n2394 GNDA 0.5637
R4523 GNDA.n2434 GNDA.n376 0.563
R4524 GNDA.n2380 GNDA.n376 0.563
R4525 GNDA.n2382 GNDA.n2380 0.563
R4526 GNDA.n2383 GNDA.n2382 0.563
R4527 GNDA.n2378 GNDA.n416 0.563
R4528 GNDA.n2333 GNDA.n416 0.563
R4529 GNDA.n2335 GNDA.n2333 0.563
R4530 GNDA.n2337 GNDA.n2335 0.563
R4531 GNDA.n2340 GNDA.n2337 0.563
R4532 GNDA.n2341 GNDA.n2331 0.563
R4533 GNDA.n2331 GNDA.n2329 0.563
R4534 GNDA.n2329 GNDA.n2327 0.563
R4535 GNDA.n237 GNDA.n235 0.563
R4536 GNDA.n239 GNDA.n237 0.563
R4537 GNDA.n241 GNDA.n239 0.563
R4538 GNDA.n243 GNDA.n241 0.563
R4539 GNDA.n245 GNDA.n243 0.563
R4540 GNDA.n247 GNDA.n245 0.563
R4541 GNDA.n249 GNDA.n247 0.563
R4542 GNDA.n251 GNDA.n249 0.563
R4543 GNDA.n253 GNDA.n251 0.563
R4544 GNDA.n255 GNDA.n253 0.563
R4545 GNDA.n256 GNDA.n255 0.563
R4546 GNDA.n353 GNDA.n351 0.563
R4547 GNDA.n46 GNDA.n44 0.563
R4548 GNDA.n48 GNDA.n46 0.563
R4549 GNDA.n50 GNDA.n48 0.563
R4550 GNDA.n7 GNDA.n5 0.563
R4551 GNDA.n9 GNDA.n7 0.563
R4552 GNDA.n11 GNDA.n9 0.563
R4553 GNDA.n2432 GNDA.n2429 0.276625
R4554 GNDA.n1433 GNDA 0.2565
R4555 GNDA.n2233 GNDA 0.2565
R4556 GNDA.n537 GNDA 0.2565
R4557 GNDA GNDA.n1937 0.2565
R4558 GNDA GNDA.n1842 0.2565
R4559 GNDA.n1619 GNDA 0.2565
R4560 GNDA GNDA.n1191 0.2565
R4561 GNDA.n788 GNDA 0.2565
R4562 GNDA.n2412 GNDA 0.2565
R4563 GNDA.n2433 GNDA.n2432 0.22375
R4564 GNDA GNDA.n1433 0.0517
R4565 GNDA GNDA.n2233 0.0517
R4566 GNDA GNDA.n537 0.0517
R4567 GNDA.n1937 GNDA 0.0517
R4568 GNDA.n1842 GNDA 0.0517
R4569 GNDA.n1619 GNDA 0.0517
R4570 GNDA.n1191 GNDA 0.0517
R4571 GNDA GNDA.n788 0.0517
R4572 GNDA.n2412 GNDA 0.0517
R4573 VDDA.n345 VDDA.t290 1212.4
R4574 VDDA.n409 VDDA.t278 1212.4
R4575 VDDA.n105 VDDA.t306 1212.4
R4576 VDDA.n174 VDDA.t321 1212.4
R4577 VDDA.n418 VDDA.t295 905.125
R4578 VDDA.n417 VDDA.t305 905.125
R4579 VDDA.n202 VDDA.t330 794.668
R4580 VDDA.n206 VDDA.t327 794.668
R4581 VDDA.n186 VDDA.t284 794.668
R4582 VDDA.n231 VDDA.t369 794.668
R4583 VDDA.n526 VDDA.t341 708.125
R4584 VDDA.t341 VDDA.n482 708.125
R4585 VDDA.n503 VDDA.t277 708.125
R4586 VDDA.t277 VDDA.n485 708.125
R4587 VDDA.n415 VDDA.n414 682
R4588 VDDA.n548 VDDA.t373 676.966
R4589 VDDA.n418 VDDA.t294 672.274
R4590 VDDA.t303 VDDA.n417 672.274
R4591 VDDA.n505 VDDA.t300 660.001
R4592 VDDA.t340 VDDA.n527 657.76
R4593 VDDA.t276 VDDA.n504 657.76
R4594 VDDA.n430 VDDA.t324 652.076
R4595 VDDA.n464 VDDA.t354 652.076
R4596 VDDA.n246 VDDA.t287 652.076
R4597 VDDA.n279 VDDA.t360 652.076
R4598 VDDA.n11 VDDA.t318 652.076
R4599 VDDA.n44 VDDA.t272 652.076
R4600 VDDA.t364 VDDA.n625 645.231
R4601 VDDA.n626 VDDA.t343 645.231
R4602 VDDA.t313 VDDA.n594 643.038
R4603 VDDA.t337 VDDA.n547 643.038
R4604 VDDA.n595 VDDA.t310 643.038
R4605 VDDA.t282 VDDA.n633 643.037
R4606 VDDA.n634 VDDA.t358 643.037
R4607 VDDA.t349 VDDA.n611 643.037
R4608 VDDA.n612 VDDA.t270 643.037
R4609 VDDA.n309 VDDA.t345 624.725
R4610 VDDA.n72 VDDA.t351 624.725
R4611 VDDA.n319 VDDA.t333 601.867
R4612 VDDA.n84 VDDA.t366 601.867
R4613 VDDA.n380 VDDA.n323 587.407
R4614 VDDA.n388 VDDA.n387 587.407
R4615 VDDA.n374 VDDA.n373 587.407
R4616 VDDA.n354 VDDA.n353 587.407
R4617 VDDA.n134 VDDA.n106 587.407
R4618 VDDA.n119 VDDA.n115 587.407
R4619 VDDA.n145 VDDA.n88 587.407
R4620 VDDA.n153 VDDA.n152 587.407
R4621 VDDA.n573 VDDA.n541 587.407
R4622 VDDA.n569 VDDA.n568 587.407
R4623 VDDA.n586 VDDA.n585 587.407
R4624 VDDA.n580 VDDA.n535 587.407
R4625 VDDA.n463 VDDA.n423 585
R4626 VDDA.n445 VDDA.n444 585
R4627 VDDA.n404 VDDA.n380 585
R4628 VDDA.n403 VDDA.n381 585
R4629 VDDA.n402 VDDA.n382 585
R4630 VDDA.n399 VDDA.n383 585
R4631 VDDA.n398 VDDA.n384 585
R4632 VDDA.n395 VDDA.n385 585
R4633 VDDA.n394 VDDA.n386 585
R4634 VDDA.n391 VDDA.n387 585
R4635 VDDA.n373 VDDA.n372 585
R4636 VDDA.n369 VDDA.n347 585
R4637 VDDA.n368 VDDA.n348 585
R4638 VDDA.n365 VDDA.n349 585
R4639 VDDA.n364 VDDA.n350 585
R4640 VDDA.n361 VDDA.n351 585
R4641 VDDA.n360 VDDA.n352 585
R4642 VDDA.n357 VDDA.n353 585
R4643 VDDA.n278 VDDA.n237 585
R4644 VDDA.n260 VDDA.n259 585
R4645 VDDA.n219 VDDA.n218 585
R4646 VDDA.n216 VDDA.n215 585
R4647 VDDA.n230 VDDA.n179 585
R4648 VDDA.n201 VDDA.n188 585
R4649 VDDA.n169 VDDA.n145 585
R4650 VDDA.n168 VDDA.n146 585
R4651 VDDA.n167 VDDA.n147 585
R4652 VDDA.n164 VDDA.n148 585
R4653 VDDA.n163 VDDA.n149 585
R4654 VDDA.n160 VDDA.n150 585
R4655 VDDA.n159 VDDA.n151 585
R4656 VDDA.n156 VDDA.n152 585
R4657 VDDA.n132 VDDA.n106 585
R4658 VDDA.n131 VDDA.n130 585
R4659 VDDA.n129 VDDA.n109 585
R4660 VDDA.n128 VDDA.n127 585
R4661 VDDA.n126 VDDA.n125 585
R4662 VDDA.n124 VDDA.n114 585
R4663 VDDA.n123 VDDA.n122 585
R4664 VDDA.n121 VDDA.n115 585
R4665 VDDA.n43 VDDA.n2 585
R4666 VDDA.n25 VDDA.n24 585
R4667 VDDA.n585 VDDA.n584 585
R4668 VDDA.n583 VDDA.n580 585
R4669 VDDA.n571 VDDA.n541 585
R4670 VDDA.n570 VDDA.n569 585
R4671 VDDA.n528 VDDA.t316 540.818
R4672 VDDA.n317 VDDA.t335 464.281
R4673 VDDA.n314 VDDA.t335 464.281
R4674 VDDA.n308 VDDA.t347 464.281
R4675 VDDA.t347 VDDA.n307 464.281
R4676 VDDA.n71 VDDA.t353 464.281
R4677 VDDA.t353 VDDA.n70 464.281
R4678 VDDA.t368 VDDA.n63 464.281
R4679 VDDA.n79 VDDA.t368 464.281
R4680 VDDA.n416 VDDA.t302 447.226
R4681 VDDA.n419 VDDA.t293 447.226
R4682 VDDA.n593 VDDA.t312 419.108
R4683 VDDA.n596 VDDA.t309 419.108
R4684 VDDA.n546 VDDA.t336 413.084
R4685 VDDA.n549 VDDA.t372 413.084
R4686 VDDA.n632 VDDA.t281 409.067
R4687 VDDA.n635 VDDA.t357 409.067
R4688 VDDA.n624 VDDA.t363 409.067
R4689 VDDA.n627 VDDA.t342 409.067
R4690 VDDA.n610 VDDA.t348 409.067
R4691 VDDA.t15 VDDA.t340 407.144
R4692 VDDA.t203 VDDA.t15 407.144
R4693 VDDA.t394 VDDA.t203 407.144
R4694 VDDA.t182 VDDA.t394 407.144
R4695 VDDA.t201 VDDA.t182 407.144
R4696 VDDA.t129 VDDA.t201 407.144
R4697 VDDA.t404 VDDA.t129 407.144
R4698 VDDA.t33 VDDA.t404 407.144
R4699 VDDA.t36 VDDA.t33 407.144
R4700 VDDA.t180 VDDA.t36 407.144
R4701 VDDA.t86 VDDA.t180 407.144
R4702 VDDA.t402 VDDA.t86 407.144
R4703 VDDA.t156 VDDA.t402 407.144
R4704 VDDA.t381 VDDA.t156 407.144
R4705 VDDA.t44 VDDA.t381 407.144
R4706 VDDA.t379 VDDA.t44 407.144
R4707 VDDA.t84 VDDA.t379 407.144
R4708 VDDA.t176 VDDA.t84 407.144
R4709 VDDA.t316 VDDA.t176 407.144
R4710 VDDA.t396 VDDA.t276 407.144
R4711 VDDA.t166 VDDA.t396 407.144
R4712 VDDA.t42 VDDA.t166 407.144
R4713 VDDA.t178 VDDA.t42 407.144
R4714 VDDA.t160 VDDA.t178 407.144
R4715 VDDA.t174 VDDA.t160 407.144
R4716 VDDA.t154 VDDA.t174 407.144
R4717 VDDA.t400 VDDA.t154 407.144
R4718 VDDA.t205 VDDA.t400 407.144
R4719 VDDA.t17 VDDA.t205 407.144
R4720 VDDA.t186 VDDA.t17 407.144
R4721 VDDA.t64 VDDA.t186 407.144
R4722 VDDA.t411 VDDA.t64 407.144
R4723 VDDA.t413 VDDA.t411 407.144
R4724 VDDA.t383 VDDA.t413 407.144
R4725 VDDA.t158 VDDA.t383 407.144
R4726 VDDA.t184 VDDA.t158 407.144
R4727 VDDA.t398 VDDA.t184 407.144
R4728 VDDA.t300 VDDA.t398 407.144
R4729 VDDA.n613 VDDA.t269 390.322
R4730 VDDA.n526 VDDA.t339 379.582
R4731 VDDA.n503 VDDA.t275 379.582
R4732 VDDA.t315 VDDA.n529 379.277
R4733 VDDA.t30 VDDA.t313 373.214
R4734 VDDA.t218 VDDA.t30 373.214
R4735 VDDA.t310 VDDA.t218 373.214
R4736 VDDA.t153 VDDA.t337 373.214
R4737 VDDA.t32 VDDA.t153 373.214
R4738 VDDA.t373 VDDA.t32 373.214
R4739 VDDA.t8 VDDA.t282 373.214
R4740 VDDA.t4 VDDA.t8 373.214
R4741 VDDA.t151 VDDA.t4 373.214
R4742 VDDA.t13 VDDA.t151 373.214
R4743 VDDA.t358 VDDA.t13 373.214
R4744 VDDA.t90 VDDA.t364 373.214
R4745 VDDA.t377 VDDA.t90 373.214
R4746 VDDA.t199 VDDA.t377 373.214
R4747 VDDA.t6 VDDA.t199 373.214
R4748 VDDA.t88 VDDA.t6 373.214
R4749 VDDA.t46 VDDA.t88 373.214
R4750 VDDA.t164 VDDA.t46 373.214
R4751 VDDA.t111 VDDA.t164 373.214
R4752 VDDA.t212 VDDA.t111 373.214
R4753 VDDA.t216 VDDA.t212 373.214
R4754 VDDA.t343 VDDA.t216 373.214
R4755 VDDA.t21 VDDA.t349 373.214
R4756 VDDA.t145 VDDA.t21 373.214
R4757 VDDA.t214 VDDA.t145 373.214
R4758 VDDA.t48 VDDA.t214 373.214
R4759 VDDA.t270 VDDA.t48 373.214
R4760 VDDA.n566 VDDA.t296 360.868
R4761 VDDA.n591 VDDA.t266 360.868
R4762 VDDA.n530 VDDA.t315 358.858
R4763 VDDA.t339 VDDA.n525 358.858
R4764 VDDA.n506 VDDA.t299 358.858
R4765 VDDA.t275 VDDA.n502 358.858
R4766 VDDA.n625 VDDA.t365 354.154
R4767 VDDA.n626 VDDA.t344 354.154
R4768 VDDA.n505 VDDA.t301 354.065
R4769 VDDA.n595 VDDA.t311 354.065
R4770 VDDA.n594 VDDA.t314 354.063
R4771 VDDA.n547 VDDA.t338 354.063
R4772 VDDA.n481 VDDA.t317 351.793
R4773 VDDA.n548 VDDA.t374 347.224
R4774 VDDA.n607 VDDA.n606 345.127
R4775 VDDA.n609 VDDA.n608 345.127
R4776 VDDA.n603 VDDA.n602 344.7
R4777 VDDA.n630 VDDA.n629 344.7
R4778 VDDA.n479 VDDA.n478 341.675
R4779 VDDA.n509 VDDA.n508 341.675
R4780 VDDA.n511 VDDA.n510 341.675
R4781 VDDA.n513 VDDA.n512 341.675
R4782 VDDA.n515 VDDA.n514 341.675
R4783 VDDA.n517 VDDA.n516 341.675
R4784 VDDA.n519 VDDA.n518 341.675
R4785 VDDA.n521 VDDA.n520 341.675
R4786 VDDA.n523 VDDA.n522 341.675
R4787 VDDA.n484 VDDA.n483 341.675
R4788 VDDA.n487 VDDA.n486 341.675
R4789 VDDA.n489 VDDA.n488 341.675
R4790 VDDA.n491 VDDA.n490 341.675
R4791 VDDA.n493 VDDA.n492 341.675
R4792 VDDA.n495 VDDA.n494 341.675
R4793 VDDA.n497 VDDA.n496 341.675
R4794 VDDA.n499 VDDA.n498 341.675
R4795 VDDA.n501 VDDA.n500 341.675
R4796 VDDA.n605 VDDA.n604 339.272
R4797 VDDA.n616 VDDA.n615 339.272
R4798 VDDA.n618 VDDA.n617 339.272
R4799 VDDA.n620 VDDA.n619 339.272
R4800 VDDA.n622 VDDA.n621 339.272
R4801 VDDA.n599 VDDA.n598 334.772
R4802 VDDA.n611 VDDA.t350 332.267
R4803 VDDA.n612 VDDA.t271 332.267
R4804 VDDA.n633 VDDA.t283 332.084
R4805 VDDA.n634 VDDA.t359 332.084
R4806 VDDA.n218 VDDA.n210 291.053
R4807 VDDA.n218 VDDA.n217 291.053
R4808 VDDA.n215 VDDA.n208 291.053
R4809 VDDA.n215 VDDA.n214 291.053
R4810 VDDA.n451 VDDA.n423 290.233
R4811 VDDA.n457 VDDA.n423 290.233
R4812 VDDA.n452 VDDA.n423 290.233
R4813 VDDA.n444 VDDA.n432 290.233
R4814 VDDA.n444 VDDA.n437 290.233
R4815 VDDA.n444 VDDA.n442 290.233
R4816 VDDA.n266 VDDA.n237 290.233
R4817 VDDA.n272 VDDA.n237 290.233
R4818 VDDA.n267 VDDA.n237 290.233
R4819 VDDA.n259 VDDA.n248 290.233
R4820 VDDA.n259 VDDA.n253 290.233
R4821 VDDA.n259 VDDA.n258 290.233
R4822 VDDA.n223 VDDA.n179 290.233
R4823 VDDA.n224 VDDA.n179 290.233
R4824 VDDA.n193 VDDA.n188 290.233
R4825 VDDA.n197 VDDA.n188 290.233
R4826 VDDA.n31 VDDA.n2 290.233
R4827 VDDA.n37 VDDA.n2 290.233
R4828 VDDA.n32 VDDA.n2 290.233
R4829 VDDA.n24 VDDA.n13 290.233
R4830 VDDA.n24 VDDA.n18 290.233
R4831 VDDA.n24 VDDA.n23 290.233
R4832 VDDA.n312 VDDA.t334 267.188
R4833 VDDA.t346 VDDA.n311 267.188
R4834 VDDA.t352 VDDA.n74 267.188
R4835 VDDA.n81 VDDA.t367 267.188
R4836 VDDA.t294 VDDA.t207 259.091
R4837 VDDA.t207 VDDA.t303 259.091
R4838 VDDA.t109 VDDA.t297 251.471
R4839 VDDA.t131 VDDA.t109 251.471
R4840 VDDA.t101 VDDA.t131 251.471
R4841 VDDA.t93 VDDA.t101 251.471
R4842 VDDA.t24 VDDA.t93 251.471
R4843 VDDA.t409 VDDA.t24 251.471
R4844 VDDA.t105 VDDA.t409 251.471
R4845 VDDA.t28 VDDA.t105 251.471
R4846 VDDA.t26 VDDA.t28 251.471
R4847 VDDA.t107 VDDA.t26 251.471
R4848 VDDA.t96 VDDA.t107 251.471
R4849 VDDA.t98 VDDA.t96 251.471
R4850 VDDA.t0 VDDA.t98 251.471
R4851 VDDA.t388 VDDA.t0 251.471
R4852 VDDA.t406 VDDA.t388 251.471
R4853 VDDA.t81 VDDA.t406 251.471
R4854 VDDA.t267 VDDA.t81 251.471
R4855 VDDA.n381 VDDA.n380 246.25
R4856 VDDA.n382 VDDA.n381 246.25
R4857 VDDA.n383 VDDA.n382 246.25
R4858 VDDA.n385 VDDA.n384 246.25
R4859 VDDA.n386 VDDA.n385 246.25
R4860 VDDA.n387 VDDA.n386 246.25
R4861 VDDA.n373 VDDA.n347 246.25
R4862 VDDA.n348 VDDA.n347 246.25
R4863 VDDA.n349 VDDA.n348 246.25
R4864 VDDA.n351 VDDA.n350 246.25
R4865 VDDA.n352 VDDA.n351 246.25
R4866 VDDA.n353 VDDA.n352 246.25
R4867 VDDA.n130 VDDA.n106 246.25
R4868 VDDA.n130 VDDA.n129 246.25
R4869 VDDA.n129 VDDA.n128 246.25
R4870 VDDA.n125 VDDA.n124 246.25
R4871 VDDA.n124 VDDA.n123 246.25
R4872 VDDA.n123 VDDA.n115 246.25
R4873 VDDA.n146 VDDA.n145 246.25
R4874 VDDA.n147 VDDA.n146 246.25
R4875 VDDA.n148 VDDA.n147 246.25
R4876 VDDA.n150 VDDA.n149 246.25
R4877 VDDA.n151 VDDA.n150 246.25
R4878 VDDA.n152 VDDA.n151 246.25
R4879 VDDA.n307 VDDA.n302 243.698
R4880 VDDA.n70 VDDA.n65 243.698
R4881 VDDA.n587 VDDA.n586 243.698
R4882 VDDA.n452 VDDA.n449 242.903
R4883 VDDA.n442 VDDA.n428 242.903
R4884 VDDA.n267 VDDA.n264 242.903
R4885 VDDA.n258 VDDA.n242 242.903
R4886 VDDA.n224 VDDA.n182 242.903
R4887 VDDA.n198 VDDA.n197 242.903
R4888 VDDA.n32 VDDA.n29 242.903
R4889 VDDA.n23 VDDA.n7 242.903
R4890 VDDA.n463 VDDA.n462 238.367
R4891 VDDA.n408 VDDA.n407 238.367
R4892 VDDA.n310 VDDA.n309 238.367
R4893 VDDA.n278 VDDA.n277 238.367
R4894 VDDA.n220 VDDA.n219 238.367
R4895 VDDA.n230 VDDA.n229 238.367
R4896 VDDA.n216 VDDA.n183 238.367
R4897 VDDA.n173 VDDA.n172 238.367
R4898 VDDA.n73 VDDA.n72 238.367
R4899 VDDA.n43 VDDA.n42 238.367
R4900 VDDA.n529 VDDA.n528 238.367
R4901 VDDA.n528 VDDA.n480 238.367
R4902 VDDA.t297 VDDA.n575 237.5
R4903 VDDA.n588 VDDA.t267 237.5
R4904 VDDA.n228 VDDA.t370 221.121
R4905 VDDA.t285 VDDA.n221 221.121
R4906 VDDA.n221 VDDA.t328 221.121
R4907 VDDA.n199 VDDA.t331 221.121
R4908 VDDA.t334 VDDA.t192 217.708
R4909 VDDA.t192 VDDA.t210 217.708
R4910 VDDA.t210 VDDA.t113 217.708
R4911 VDDA.t113 VDDA.t209 217.708
R4912 VDDA.t209 VDDA.t197 217.708
R4913 VDDA.t197 VDDA.t385 217.708
R4914 VDDA.t385 VDDA.t35 217.708
R4915 VDDA.t35 VDDA.t211 217.708
R4916 VDDA.t211 VDDA.t70 217.708
R4917 VDDA.t70 VDDA.t69 217.708
R4918 VDDA.t69 VDDA.t346 217.708
R4919 VDDA.t72 VDDA.t352 217.708
R4920 VDDA.t76 VDDA.t72 217.708
R4921 VDDA.t63 VDDA.t76 217.708
R4922 VDDA.t150 VDDA.t63 217.708
R4923 VDDA.t124 VDDA.t150 217.708
R4924 VDDA.t80 VDDA.t124 217.708
R4925 VDDA.t38 VDDA.t80 217.708
R4926 VDDA.t10 VDDA.t38 217.708
R4927 VDDA.t128 VDDA.t10 217.708
R4928 VDDA.t148 VDDA.t128 217.708
R4929 VDDA.t367 VDDA.t148 217.708
R4930 VDDA.n178 VDDA.n177 213.186
R4931 VDDA.n204 VDDA.n203 213.186
R4932 VDDA.n388 VDDA.n329 190.333
R4933 VDDA.n354 VDDA.n335 190.333
R4934 VDDA.n314 VDDA.n313 190.333
R4935 VDDA.n153 VDDA.n142 190.333
R4936 VDDA.n119 VDDA.n95 190.333
R4937 VDDA.n80 VDDA.n79 190.333
R4938 VDDA.n574 VDDA.n573 190.333
R4939 VDDA.n425 VDDA.n424 185
R4940 VDDA.n460 VDDA.n459 185
R4941 VDDA.n461 VDDA.n460 185
R4942 VDDA.n458 VDDA.n450 185
R4943 VDDA.n456 VDDA.n455 185
R4944 VDDA.n454 VDDA.n453 185
R4945 VDDA.n446 VDDA.n445 185
R4946 VDDA.n447 VDDA.n446 185
R4947 VDDA.n431 VDDA.n429 185
R4948 VDDA.n434 VDDA.n433 185
R4949 VDDA.n436 VDDA.n435 185
R4950 VDDA.n439 VDDA.n438 185
R4951 VDDA.n441 VDDA.n440 185
R4952 VDDA.n379 VDDA.n324 185
R4953 VDDA.n405 VDDA.n404 185
R4954 VDDA.n406 VDDA.n405 185
R4955 VDDA.n403 VDDA.n378 185
R4956 VDDA.n402 VDDA.n401 185
R4957 VDDA.n400 VDDA.n399 185
R4958 VDDA.n398 VDDA.n397 185
R4959 VDDA.n396 VDDA.n395 185
R4960 VDDA.n394 VDDA.n393 185
R4961 VDDA.n392 VDDA.n391 185
R4962 VDDA.n390 VDDA.n389 185
R4963 VDDA.n406 VDDA.n329 185
R4964 VDDA.n376 VDDA.n375 185
R4965 VDDA.n377 VDDA.n376 185
R4966 VDDA.n346 VDDA.n336 185
R4967 VDDA.n372 VDDA.n371 185
R4968 VDDA.n370 VDDA.n369 185
R4969 VDDA.n368 VDDA.n367 185
R4970 VDDA.n366 VDDA.n365 185
R4971 VDDA.n364 VDDA.n363 185
R4972 VDDA.n362 VDDA.n361 185
R4973 VDDA.n360 VDDA.n359 185
R4974 VDDA.n358 VDDA.n357 185
R4975 VDDA.n356 VDDA.n355 185
R4976 VDDA.n377 VDDA.n335 185
R4977 VDDA.n304 VDDA.n303 185
R4978 VDDA.n306 VDDA.n305 185
R4979 VDDA.n318 VDDA.n298 185
R4980 VDDA.n312 VDDA.n298 185
R4981 VDDA.n316 VDDA.n299 185
R4982 VDDA.n315 VDDA.n300 185
R4983 VDDA.n313 VDDA.n312 185
R4984 VDDA.n239 VDDA.n238 185
R4985 VDDA.n275 VDDA.n274 185
R4986 VDDA.n276 VDDA.n275 185
R4987 VDDA.n273 VDDA.n265 185
R4988 VDDA.n271 VDDA.n270 185
R4989 VDDA.n269 VDDA.n268 185
R4990 VDDA.n261 VDDA.n260 185
R4991 VDDA.n262 VDDA.n261 185
R4992 VDDA.n247 VDDA.n243 185
R4993 VDDA.n250 VDDA.n249 185
R4994 VDDA.n252 VDDA.n251 185
R4995 VDDA.n255 VDDA.n254 185
R4996 VDDA.n257 VDDA.n256 185
R4997 VDDA.n181 VDDA.n180 185
R4998 VDDA.n227 VDDA.n226 185
R4999 VDDA.n228 VDDA.n227 185
R5000 VDDA.n225 VDDA.n222 185
R5001 VDDA.n209 VDDA.n185 185
R5002 VDDA.n213 VDDA.n184 185
R5003 VDDA.n221 VDDA.n184 185
R5004 VDDA.n212 VDDA.n211 185
R5005 VDDA.n201 VDDA.n200 185
R5006 VDDA.n200 VDDA.n199 185
R5007 VDDA.n190 VDDA.n189 185
R5008 VDDA.n195 VDDA.n194 185
R5009 VDDA.n196 VDDA.n192 185
R5010 VDDA.n144 VDDA.n89 185
R5011 VDDA.n170 VDDA.n169 185
R5012 VDDA.n171 VDDA.n170 185
R5013 VDDA.n168 VDDA.n143 185
R5014 VDDA.n167 VDDA.n166 185
R5015 VDDA.n165 VDDA.n164 185
R5016 VDDA.n163 VDDA.n162 185
R5017 VDDA.n161 VDDA.n160 185
R5018 VDDA.n159 VDDA.n158 185
R5019 VDDA.n157 VDDA.n156 185
R5020 VDDA.n155 VDDA.n154 185
R5021 VDDA.n171 VDDA.n142 185
R5022 VDDA.n136 VDDA.n135 185
R5023 VDDA.n137 VDDA.n136 185
R5024 VDDA.n133 VDDA.n96 185
R5025 VDDA.n132 VDDA.n107 185
R5026 VDDA.n131 VDDA.n108 185
R5027 VDDA.n110 VDDA.n109 185
R5028 VDDA.n127 VDDA.n111 185
R5029 VDDA.n126 VDDA.n112 185
R5030 VDDA.n114 VDDA.n113 185
R5031 VDDA.n122 VDDA.n116 185
R5032 VDDA.n121 VDDA.n117 185
R5033 VDDA.n120 VDDA.n118 185
R5034 VDDA.n137 VDDA.n95 185
R5035 VDDA.n67 VDDA.n66 185
R5036 VDDA.n69 VDDA.n68 185
R5037 VDDA.n83 VDDA.n82 185
R5038 VDDA.n82 VDDA.n81 185
R5039 VDDA.n77 VDDA.n64 185
R5040 VDDA.n78 VDDA.n76 185
R5041 VDDA.n81 VDDA.n80 185
R5042 VDDA.n4 VDDA.n3 185
R5043 VDDA.n40 VDDA.n39 185
R5044 VDDA.n41 VDDA.n40 185
R5045 VDDA.n38 VDDA.n30 185
R5046 VDDA.n36 VDDA.n35 185
R5047 VDDA.n34 VDDA.n33 185
R5048 VDDA.n26 VDDA.n25 185
R5049 VDDA.n27 VDDA.n26 185
R5050 VDDA.n12 VDDA.n8 185
R5051 VDDA.n15 VDDA.n14 185
R5052 VDDA.n17 VDDA.n16 185
R5053 VDDA.n20 VDDA.n19 185
R5054 VDDA.n22 VDDA.n21 185
R5055 VDDA.n579 VDDA.n578 185
R5056 VDDA.n584 VDDA.n577 185
R5057 VDDA.n588 VDDA.n577 185
R5058 VDDA.n583 VDDA.n582 185
R5059 VDDA.n581 VDDA.n536 185
R5060 VDDA.n590 VDDA.n589 185
R5061 VDDA.n589 VDDA.n588 185
R5062 VDDA.n575 VDDA.n574 185
R5063 VDDA.n572 VDDA.n540 185
R5064 VDDA.n571 VDDA.n542 185
R5065 VDDA.n570 VDDA.n543 185
R5066 VDDA.n545 VDDA.n544 185
R5067 VDDA.n567 VDDA.n539 185
R5068 VDDA.n575 VDDA.n539 185
R5069 VDDA.t370 VDDA.t170 180.173
R5070 VDDA.t170 VDDA.t190 180.173
R5071 VDDA.t190 VDDA.t188 180.173
R5072 VDDA.t188 VDDA.t376 180.173
R5073 VDDA.t376 VDDA.t285 180.173
R5074 VDDA.t375 VDDA.t328 180.173
R5075 VDDA.t172 VDDA.t375 180.173
R5076 VDDA.t162 VDDA.t172 180.173
R5077 VDDA.t171 VDDA.t162 180.173
R5078 VDDA.t331 VDDA.t171 180.173
R5079 VDDA.t325 VDDA.n447 170.513
R5080 VDDA.n461 VDDA.t355 170.513
R5081 VDDA.t288 VDDA.n262 170.513
R5082 VDDA.n276 VDDA.t361 170.513
R5083 VDDA.t319 VDDA.n27 170.513
R5084 VDDA.n41 VDDA.t273 170.513
R5085 VDDA.n534 VDDA.n533 168.435
R5086 VDDA.n552 VDDA.n551 168.435
R5087 VDDA.n554 VDDA.n553 168.435
R5088 VDDA.n556 VDDA.n555 168.435
R5089 VDDA.n558 VDDA.n557 168.435
R5090 VDDA.n560 VDDA.n559 168.435
R5091 VDDA.n562 VDDA.n561 168.435
R5092 VDDA.n564 VDDA.n563 168.435
R5093 VDDA.n443 VDDA.n422 159.803
R5094 VDDA.n236 VDDA.n235 159.803
R5095 VDDA.n245 VDDA.n244 159.803
R5096 VDDA.n281 VDDA.n280 159.803
R5097 VDDA.n283 VDDA.n282 159.803
R5098 VDDA.n1 VDDA.n0 159.803
R5099 VDDA.n10 VDDA.n9 159.803
R5100 VDDA.n46 VDDA.n45 159.803
R5101 VDDA.n48 VDDA.n47 159.803
R5102 VDDA.n286 VDDA.n285 155.303
R5103 VDDA.n51 VDDA.n50 155.303
R5104 VDDA.n460 VDDA.n425 150
R5105 VDDA.n460 VDDA.n450 150
R5106 VDDA.n455 VDDA.n454 150
R5107 VDDA.n446 VDDA.n429 150
R5108 VDDA.n435 VDDA.n434 150
R5109 VDDA.n440 VDDA.n439 150
R5110 VDDA.n405 VDDA.n324 150
R5111 VDDA.n405 VDDA.n378 150
R5112 VDDA.n401 VDDA.n400 150
R5113 VDDA.n397 VDDA.n396 150
R5114 VDDA.n393 VDDA.n392 150
R5115 VDDA.n389 VDDA.n329 150
R5116 VDDA.n376 VDDA.n336 150
R5117 VDDA.n371 VDDA.n370 150
R5118 VDDA.n367 VDDA.n366 150
R5119 VDDA.n363 VDDA.n362 150
R5120 VDDA.n359 VDDA.n358 150
R5121 VDDA.n355 VDDA.n335 150
R5122 VDDA.n305 VDDA.n303 150
R5123 VDDA.n299 VDDA.n298 150
R5124 VDDA.n313 VDDA.n300 150
R5125 VDDA.n275 VDDA.n239 150
R5126 VDDA.n275 VDDA.n265 150
R5127 VDDA.n270 VDDA.n269 150
R5128 VDDA.n261 VDDA.n243 150
R5129 VDDA.n251 VDDA.n250 150
R5130 VDDA.n256 VDDA.n255 150
R5131 VDDA.n185 VDDA.n184 150
R5132 VDDA.n211 VDDA.n184 150
R5133 VDDA.n227 VDDA.n181 150
R5134 VDDA.n227 VDDA.n222 150
R5135 VDDA.n200 VDDA.n190 150
R5136 VDDA.n194 VDDA.n192 150
R5137 VDDA.n170 VDDA.n89 150
R5138 VDDA.n170 VDDA.n143 150
R5139 VDDA.n166 VDDA.n165 150
R5140 VDDA.n162 VDDA.n161 150
R5141 VDDA.n158 VDDA.n157 150
R5142 VDDA.n154 VDDA.n142 150
R5143 VDDA.n136 VDDA.n96 150
R5144 VDDA.n108 VDDA.n107 150
R5145 VDDA.n111 VDDA.n110 150
R5146 VDDA.n113 VDDA.n112 150
R5147 VDDA.n117 VDDA.n116 150
R5148 VDDA.n118 VDDA.n95 150
R5149 VDDA.n68 VDDA.n66 150
R5150 VDDA.n82 VDDA.n64 150
R5151 VDDA.n80 VDDA.n76 150
R5152 VDDA.n40 VDDA.n4 150
R5153 VDDA.n40 VDDA.n30 150
R5154 VDDA.n35 VDDA.n34 150
R5155 VDDA.n26 VDDA.n8 150
R5156 VDDA.n16 VDDA.n15 150
R5157 VDDA.n21 VDDA.n20 150
R5158 VDDA.n578 VDDA.n577 150
R5159 VDDA.n582 VDDA.n577 150
R5160 VDDA.n589 VDDA.n536 150
R5161 VDDA.n574 VDDA.n540 150
R5162 VDDA.n543 VDDA.n542 150
R5163 VDDA.n544 VDDA.n539 150
R5164 VDDA.t248 VDDA.t325 146.155
R5165 VDDA.t355 VDDA.t248 146.155
R5166 VDDA.t232 VDDA.t288 146.155
R5167 VDDA.t228 VDDA.t232 146.155
R5168 VDDA.t236 VDDA.t228 146.155
R5169 VDDA.t246 VDDA.t236 146.155
R5170 VDDA.t256 VDDA.t246 146.155
R5171 VDDA.t226 VDDA.t256 146.155
R5172 VDDA.t224 VDDA.t226 146.155
R5173 VDDA.t230 VDDA.t224 146.155
R5174 VDDA.t238 VDDA.t230 146.155
R5175 VDDA.t250 VDDA.t238 146.155
R5176 VDDA.t361 VDDA.t250 146.155
R5177 VDDA.t244 VDDA.t319 146.155
R5178 VDDA.t240 VDDA.t244 146.155
R5179 VDDA.t252 VDDA.t240 146.155
R5180 VDDA.t258 VDDA.t252 146.155
R5181 VDDA.t220 VDDA.t258 146.155
R5182 VDDA.t222 VDDA.t220 146.155
R5183 VDDA.t234 VDDA.t222 146.155
R5184 VDDA.t242 VDDA.t234 146.155
R5185 VDDA.t254 VDDA.t242 146.155
R5186 VDDA.t260 VDDA.t254 146.155
R5187 VDDA.t273 VDDA.t260 146.155
R5188 VDDA.n322 VDDA.n321 145.429
R5189 VDDA.n338 VDDA.n337 145.429
R5190 VDDA.n340 VDDA.n339 145.429
R5191 VDDA.n342 VDDA.n341 145.429
R5192 VDDA.n344 VDDA.n343 145.429
R5193 VDDA.n87 VDDA.n86 145.429
R5194 VDDA.n98 VDDA.n97 145.429
R5195 VDDA.n100 VDDA.n99 145.429
R5196 VDDA.n102 VDDA.n101 145.429
R5197 VDDA.n104 VDDA.n103 145.429
R5198 VDDA.t280 VDDA.n383 123.126
R5199 VDDA.n384 VDDA.t280 123.126
R5200 VDDA.t292 VDDA.n349 123.126
R5201 VDDA.n350 VDDA.t292 123.126
R5202 VDDA.n128 VDDA.t308 123.126
R5203 VDDA.n125 VDDA.t308 123.126
R5204 VDDA.t323 VDDA.n148 123.126
R5205 VDDA.n149 VDDA.t323 123.126
R5206 VDDA.t298 VDDA.n541 123.126
R5207 VDDA.n569 VDDA.t298 123.126
R5208 VDDA.n585 VDDA.t268 123.126
R5209 VDDA.n580 VDDA.t268 123.126
R5210 VDDA.n406 VDDA.t279 100.195
R5211 VDDA.t291 VDDA.n377 100.195
R5212 VDDA.t307 VDDA.n137 100.195
R5213 VDDA.n171 VDDA.t322 100.195
R5214 VDDA.n289 VDDA.n287 97.4002
R5215 VDDA.n54 VDDA.n52 97.4002
R5216 VDDA.n297 VDDA.n296 96.8377
R5217 VDDA.n295 VDDA.n294 96.8377
R5218 VDDA.n293 VDDA.n292 96.8377
R5219 VDDA.n291 VDDA.n290 96.8377
R5220 VDDA.n289 VDDA.n288 96.8377
R5221 VDDA.n62 VDDA.n61 96.8377
R5222 VDDA.n60 VDDA.n59 96.8377
R5223 VDDA.n58 VDDA.n57 96.8377
R5224 VDDA.n56 VDDA.n55 96.8377
R5225 VDDA.n54 VDDA.n53 96.8377
R5226 VDDA.t279 VDDA.t57 81.6411
R5227 VDDA.t57 VDDA.t67 81.6411
R5228 VDDA.t67 VDDA.t55 81.6411
R5229 VDDA.t55 VDDA.t114 81.6411
R5230 VDDA.t114 VDDA.t53 81.6411
R5231 VDDA.t53 VDDA.t194 81.6411
R5232 VDDA.t194 VDDA.t19 81.6411
R5233 VDDA.t19 VDDA.t392 81.6411
R5234 VDDA.t392 VDDA.t117 81.6411
R5235 VDDA.t117 VDDA.t119 81.6411
R5236 VDDA.t119 VDDA.t291 81.6411
R5237 VDDA.t40 VDDA.t307 81.6411
R5238 VDDA.t137 VDDA.t40 81.6411
R5239 VDDA.t11 VDDA.t137 81.6411
R5240 VDDA.t73 VDDA.t11 81.6411
R5241 VDDA.t77 VDDA.t73 81.6411
R5242 VDDA.t59 VDDA.t77 81.6411
R5243 VDDA.t143 VDDA.t59 81.6411
R5244 VDDA.t135 VDDA.t143 81.6411
R5245 VDDA.t141 VDDA.t135 81.6411
R5246 VDDA.t125 VDDA.t141 81.6411
R5247 VDDA.t322 VDDA.t125 81.6411
R5248 VDDA.n462 VDDA.n461 65.8183
R5249 VDDA.n461 VDDA.n448 65.8183
R5250 VDDA.n461 VDDA.n449 65.8183
R5251 VDDA.n447 VDDA.n426 65.8183
R5252 VDDA.n447 VDDA.n427 65.8183
R5253 VDDA.n447 VDDA.n428 65.8183
R5254 VDDA.n407 VDDA.n406 65.8183
R5255 VDDA.n406 VDDA.n325 65.8183
R5256 VDDA.n406 VDDA.n326 65.8183
R5257 VDDA.n406 VDDA.n327 65.8183
R5258 VDDA.n406 VDDA.n328 65.8183
R5259 VDDA.n377 VDDA.n330 65.8183
R5260 VDDA.n377 VDDA.n331 65.8183
R5261 VDDA.n377 VDDA.n332 65.8183
R5262 VDDA.n377 VDDA.n333 65.8183
R5263 VDDA.n377 VDDA.n334 65.8183
R5264 VDDA.n311 VDDA.n310 65.8183
R5265 VDDA.n311 VDDA.n302 65.8183
R5266 VDDA.n312 VDDA.n301 65.8183
R5267 VDDA.n277 VDDA.n276 65.8183
R5268 VDDA.n276 VDDA.n263 65.8183
R5269 VDDA.n276 VDDA.n264 65.8183
R5270 VDDA.n262 VDDA.n240 65.8183
R5271 VDDA.n262 VDDA.n241 65.8183
R5272 VDDA.n262 VDDA.n242 65.8183
R5273 VDDA.n229 VDDA.n228 65.8183
R5274 VDDA.n228 VDDA.n182 65.8183
R5275 VDDA.n221 VDDA.n220 65.8183
R5276 VDDA.n221 VDDA.n183 65.8183
R5277 VDDA.n199 VDDA.n191 65.8183
R5278 VDDA.n199 VDDA.n198 65.8183
R5279 VDDA.n172 VDDA.n171 65.8183
R5280 VDDA.n171 VDDA.n138 65.8183
R5281 VDDA.n171 VDDA.n139 65.8183
R5282 VDDA.n171 VDDA.n140 65.8183
R5283 VDDA.n171 VDDA.n141 65.8183
R5284 VDDA.n137 VDDA.n90 65.8183
R5285 VDDA.n137 VDDA.n91 65.8183
R5286 VDDA.n137 VDDA.n92 65.8183
R5287 VDDA.n137 VDDA.n93 65.8183
R5288 VDDA.n137 VDDA.n94 65.8183
R5289 VDDA.n74 VDDA.n73 65.8183
R5290 VDDA.n74 VDDA.n65 65.8183
R5291 VDDA.n81 VDDA.n75 65.8183
R5292 VDDA.n42 VDDA.n41 65.8183
R5293 VDDA.n41 VDDA.n28 65.8183
R5294 VDDA.n41 VDDA.n29 65.8183
R5295 VDDA.n27 VDDA.n5 65.8183
R5296 VDDA.n27 VDDA.n6 65.8183
R5297 VDDA.n27 VDDA.n7 65.8183
R5298 VDDA.n588 VDDA.n587 65.8183
R5299 VDDA.n588 VDDA.n576 65.8183
R5300 VDDA.n575 VDDA.n537 65.8183
R5301 VDDA.n575 VDDA.n538 65.8183
R5302 VDDA.n475 VDDA.t417 59.5681
R5303 VDDA.n474 VDDA.t418 59.5681
R5304 VDDA.n450 VDDA.n448 53.3664
R5305 VDDA.n454 VDDA.n449 53.3664
R5306 VDDA.n462 VDDA.n425 53.3664
R5307 VDDA.n455 VDDA.n448 53.3664
R5308 VDDA.n429 VDDA.n426 53.3664
R5309 VDDA.n435 VDDA.n427 53.3664
R5310 VDDA.n440 VDDA.n428 53.3664
R5311 VDDA.n434 VDDA.n426 53.3664
R5312 VDDA.n439 VDDA.n427 53.3664
R5313 VDDA.n378 VDDA.n325 53.3664
R5314 VDDA.n400 VDDA.n326 53.3664
R5315 VDDA.n396 VDDA.n327 53.3664
R5316 VDDA.n392 VDDA.n328 53.3664
R5317 VDDA.n407 VDDA.n324 53.3664
R5318 VDDA.n401 VDDA.n325 53.3664
R5319 VDDA.n397 VDDA.n326 53.3664
R5320 VDDA.n393 VDDA.n327 53.3664
R5321 VDDA.n389 VDDA.n328 53.3664
R5322 VDDA.n336 VDDA.n330 53.3664
R5323 VDDA.n370 VDDA.n331 53.3664
R5324 VDDA.n366 VDDA.n332 53.3664
R5325 VDDA.n362 VDDA.n333 53.3664
R5326 VDDA.n358 VDDA.n334 53.3664
R5327 VDDA.n371 VDDA.n330 53.3664
R5328 VDDA.n367 VDDA.n331 53.3664
R5329 VDDA.n363 VDDA.n332 53.3664
R5330 VDDA.n359 VDDA.n333 53.3664
R5331 VDDA.n355 VDDA.n334 53.3664
R5332 VDDA.n310 VDDA.n303 53.3664
R5333 VDDA.n305 VDDA.n302 53.3664
R5334 VDDA.n301 VDDA.n299 53.3664
R5335 VDDA.n301 VDDA.n300 53.3664
R5336 VDDA.n265 VDDA.n263 53.3664
R5337 VDDA.n269 VDDA.n264 53.3664
R5338 VDDA.n277 VDDA.n239 53.3664
R5339 VDDA.n270 VDDA.n263 53.3664
R5340 VDDA.n243 VDDA.n240 53.3664
R5341 VDDA.n251 VDDA.n241 53.3664
R5342 VDDA.n256 VDDA.n242 53.3664
R5343 VDDA.n250 VDDA.n240 53.3664
R5344 VDDA.n255 VDDA.n241 53.3664
R5345 VDDA.n211 VDDA.n183 53.3664
R5346 VDDA.n222 VDDA.n182 53.3664
R5347 VDDA.n229 VDDA.n181 53.3664
R5348 VDDA.n220 VDDA.n185 53.3664
R5349 VDDA.n191 VDDA.n190 53.3664
R5350 VDDA.n198 VDDA.n192 53.3664
R5351 VDDA.n194 VDDA.n191 53.3664
R5352 VDDA.n143 VDDA.n138 53.3664
R5353 VDDA.n165 VDDA.n139 53.3664
R5354 VDDA.n161 VDDA.n140 53.3664
R5355 VDDA.n157 VDDA.n141 53.3664
R5356 VDDA.n172 VDDA.n89 53.3664
R5357 VDDA.n166 VDDA.n138 53.3664
R5358 VDDA.n162 VDDA.n139 53.3664
R5359 VDDA.n158 VDDA.n140 53.3664
R5360 VDDA.n154 VDDA.n141 53.3664
R5361 VDDA.n96 VDDA.n90 53.3664
R5362 VDDA.n108 VDDA.n91 53.3664
R5363 VDDA.n111 VDDA.n92 53.3664
R5364 VDDA.n113 VDDA.n93 53.3664
R5365 VDDA.n117 VDDA.n94 53.3664
R5366 VDDA.n107 VDDA.n90 53.3664
R5367 VDDA.n110 VDDA.n91 53.3664
R5368 VDDA.n112 VDDA.n92 53.3664
R5369 VDDA.n116 VDDA.n93 53.3664
R5370 VDDA.n118 VDDA.n94 53.3664
R5371 VDDA.n73 VDDA.n66 53.3664
R5372 VDDA.n68 VDDA.n65 53.3664
R5373 VDDA.n75 VDDA.n64 53.3664
R5374 VDDA.n76 VDDA.n75 53.3664
R5375 VDDA.n30 VDDA.n28 53.3664
R5376 VDDA.n34 VDDA.n29 53.3664
R5377 VDDA.n42 VDDA.n4 53.3664
R5378 VDDA.n35 VDDA.n28 53.3664
R5379 VDDA.n8 VDDA.n5 53.3664
R5380 VDDA.n16 VDDA.n6 53.3664
R5381 VDDA.n21 VDDA.n7 53.3664
R5382 VDDA.n15 VDDA.n5 53.3664
R5383 VDDA.n20 VDDA.n6 53.3664
R5384 VDDA.n582 VDDA.n576 53.3664
R5385 VDDA.n587 VDDA.n578 53.3664
R5386 VDDA.n576 VDDA.n536 53.3664
R5387 VDDA.n540 VDDA.n537 53.3664
R5388 VDDA.n543 VDDA.n538 53.3664
R5389 VDDA.n542 VDDA.n537 53.3664
R5390 VDDA.n544 VDDA.n538 53.3664
R5391 VDDA.n474 VDDA.t416 52.3888
R5392 VDDA.n231 VDDA.n230 51.6576
R5393 VDDA.n202 VDDA.n201 51.6576
R5394 VDDA.n476 VDDA.t415 48.9557
R5395 VDDA.n207 VDDA.n206 48.0005
R5396 VDDA.n207 VDDA.n186 48.0005
R5397 VDDA.n419 VDDA.n418 46.6291
R5398 VDDA.n417 VDDA.n416 46.6291
R5399 VDDA.n478 VDDA.t85 39.4005
R5400 VDDA.n478 VDDA.t177 39.4005
R5401 VDDA.n508 VDDA.t45 39.4005
R5402 VDDA.n508 VDDA.t380 39.4005
R5403 VDDA.n510 VDDA.t157 39.4005
R5404 VDDA.n510 VDDA.t382 39.4005
R5405 VDDA.n512 VDDA.t87 39.4005
R5406 VDDA.n512 VDDA.t403 39.4005
R5407 VDDA.n514 VDDA.t37 39.4005
R5408 VDDA.n514 VDDA.t181 39.4005
R5409 VDDA.n516 VDDA.t405 39.4005
R5410 VDDA.n516 VDDA.t34 39.4005
R5411 VDDA.n518 VDDA.t202 39.4005
R5412 VDDA.n518 VDDA.t130 39.4005
R5413 VDDA.n520 VDDA.t395 39.4005
R5414 VDDA.n520 VDDA.t183 39.4005
R5415 VDDA.n522 VDDA.t16 39.4005
R5416 VDDA.n522 VDDA.t204 39.4005
R5417 VDDA.n483 VDDA.t185 39.4005
R5418 VDDA.n483 VDDA.t399 39.4005
R5419 VDDA.n486 VDDA.t384 39.4005
R5420 VDDA.n486 VDDA.t159 39.4005
R5421 VDDA.n488 VDDA.t412 39.4005
R5422 VDDA.n488 VDDA.t414 39.4005
R5423 VDDA.n490 VDDA.t187 39.4005
R5424 VDDA.n490 VDDA.t65 39.4005
R5425 VDDA.n492 VDDA.t206 39.4005
R5426 VDDA.n492 VDDA.t18 39.4005
R5427 VDDA.n494 VDDA.t155 39.4005
R5428 VDDA.n494 VDDA.t401 39.4005
R5429 VDDA.n496 VDDA.t161 39.4005
R5430 VDDA.n496 VDDA.t175 39.4005
R5431 VDDA.n498 VDDA.t43 39.4005
R5432 VDDA.n498 VDDA.t179 39.4005
R5433 VDDA.n500 VDDA.t397 39.4005
R5434 VDDA.n500 VDDA.t167 39.4005
R5435 VDDA.n598 VDDA.t31 39.4005
R5436 VDDA.n598 VDDA.t219 39.4005
R5437 VDDA.n602 VDDA.t152 39.4005
R5438 VDDA.n602 VDDA.t14 39.4005
R5439 VDDA.n629 VDDA.t9 39.4005
R5440 VDDA.n629 VDDA.t5 39.4005
R5441 VDDA.n604 VDDA.t213 39.4005
R5442 VDDA.n604 VDDA.t217 39.4005
R5443 VDDA.n615 VDDA.t165 39.4005
R5444 VDDA.n615 VDDA.t112 39.4005
R5445 VDDA.n617 VDDA.t89 39.4005
R5446 VDDA.n617 VDDA.t47 39.4005
R5447 VDDA.n619 VDDA.t200 39.4005
R5448 VDDA.n619 VDDA.t7 39.4005
R5449 VDDA.n621 VDDA.t91 39.4005
R5450 VDDA.n621 VDDA.t378 39.4005
R5451 VDDA.n606 VDDA.t215 39.4005
R5452 VDDA.n606 VDDA.t49 39.4005
R5453 VDDA.n608 VDDA.t22 39.4005
R5454 VDDA.n608 VDDA.t146 39.4005
R5455 VDDA.n473 VDDA.n467 27.9413
R5456 VDDA.n635 VDDA.n634 27.2462
R5457 VDDA.n633 VDDA.n632 27.2462
R5458 VDDA.n613 VDDA.n612 27.2462
R5459 VDDA.n611 VDDA.n610 27.2462
R5460 VDDA.n594 VDDA.n593 25.087
R5461 VDDA.n596 VDDA.n595 25.087
R5462 VDDA.n627 VDDA.n626 25.0384
R5463 VDDA.n625 VDDA.n624 25.0384
R5464 VDDA.n547 VDDA.n546 22.9536
R5465 VDDA.n506 VDDA.n505 22.9536
R5466 VDDA.n464 VDDA.n463 22.8576
R5467 VDDA.n445 VDDA.n430 22.8576
R5468 VDDA.n409 VDDA.n408 22.8576
R5469 VDDA.n375 VDDA.n345 22.8576
R5470 VDDA.n319 VDDA.n318 22.8576
R5471 VDDA.n279 VDDA.n278 22.8576
R5472 VDDA.n260 VDDA.n246 22.8576
R5473 VDDA.n174 VDDA.n173 22.8576
R5474 VDDA.n135 VDDA.n105 22.8576
R5475 VDDA.n84 VDDA.n83 22.8576
R5476 VDDA.n44 VDDA.n43 22.8576
R5477 VDDA.n25 VDDA.n11 22.8576
R5478 VDDA.n591 VDDA.n590 22.8576
R5479 VDDA.n567 VDDA.n566 22.8576
R5480 VDDA.n414 VDDA.t208 21.8894
R5481 VDDA.n414 VDDA.t304 21.8894
R5482 VDDA.n467 VDDA.n466 20.883
R5483 VDDA.n530 VDDA.n480 20.7243
R5484 VDDA.n525 VDDA.n482 20.7243
R5485 VDDA.n502 VDDA.n485 20.7243
R5486 VDDA.n549 VDDA.n548 20.4312
R5487 VDDA.n473 VDDA.t3 19.9244
R5488 VDDA.n320 VDDA.n319 19.613
R5489 VDDA.n85 VDDA.n84 19.613
R5490 VDDA.n177 VDDA.t191 15.7605
R5491 VDDA.n177 VDDA.t189 15.7605
R5492 VDDA.n203 VDDA.t173 15.7605
R5493 VDDA.n203 VDDA.t163 15.7605
R5494 VDDA.n215 VDDA.t329 15.7605
R5495 VDDA.n218 VDDA.t286 15.7605
R5496 VDDA.n179 VDDA.t371 15.7605
R5497 VDDA.n188 VDDA.t332 15.7605
R5498 VDDA.n550 VDDA.n546 15.488
R5499 VDDA.n204 VDDA.n202 14.7224
R5500 VDDA.n502 VDDA.n501 14.6963
R5501 VDDA.n281 VDDA.n279 14.4255
R5502 VDDA.n246 VDDA.n245 14.4255
R5503 VDDA.n46 VDDA.n44 14.4255
R5504 VDDA.n11 VDDA.n10 14.4255
R5505 VDDA.n345 VDDA.n344 14.363
R5506 VDDA.n105 VDDA.n104 14.363
R5507 VDDA.n597 VDDA.n596 14.363
R5508 VDDA.n597 VDDA.n593 14.363
R5509 VDDA.n610 VDDA.n609 14.363
R5510 VDDA.n550 VDDA.n549 14.238
R5511 VDDA.n525 VDDA.n524 14.0713
R5512 VDDA.n531 VDDA.n530 14.0713
R5513 VDDA.n507 VDDA.n506 14.0713
R5514 VDDA.n430 VDDA.n422 14.0505
R5515 VDDA.n416 VDDA.n415 14.0505
R5516 VDDA.n465 VDDA.n464 13.8005
R5517 VDDA.n420 VDDA.n419 13.8005
R5518 VDDA.n410 VDDA.n409 13.8005
R5519 VDDA.n206 VDDA.n205 13.8005
R5520 VDDA.n187 VDDA.n186 13.8005
R5521 VDDA.n232 VDDA.n231 13.8005
R5522 VDDA.n175 VDDA.n174 13.8005
R5523 VDDA.n566 VDDA.n565 13.8005
R5524 VDDA.n592 VDDA.n591 13.8005
R5525 VDDA.n632 VDDA.n631 13.8005
R5526 VDDA.n624 VDDA.n623 13.8005
R5527 VDDA.n614 VDDA.n613 13.8005
R5528 VDDA.n628 VDDA.n627 13.8005
R5529 VDDA.n636 VDDA.n635 13.8005
R5530 VDDA.n533 VDDA.t407 13.1338
R5531 VDDA.n533 VDDA.t82 13.1338
R5532 VDDA.n551 VDDA.t1 13.1338
R5533 VDDA.n551 VDDA.t389 13.1338
R5534 VDDA.n553 VDDA.t97 13.1338
R5535 VDDA.n553 VDDA.t99 13.1338
R5536 VDDA.n555 VDDA.t27 13.1338
R5537 VDDA.n555 VDDA.t108 13.1338
R5538 VDDA.n557 VDDA.t106 13.1338
R5539 VDDA.n557 VDDA.t29 13.1338
R5540 VDDA.n559 VDDA.t25 13.1338
R5541 VDDA.n559 VDDA.t410 13.1338
R5542 VDDA.n561 VDDA.t102 13.1338
R5543 VDDA.n561 VDDA.t94 13.1338
R5544 VDDA.n563 VDDA.t110 13.1338
R5545 VDDA.n563 VDDA.t132 13.1338
R5546 VDDA.n637 VDDA.n636 11.4105
R5547 VDDA.t326 VDDA.n443 11.2576
R5548 VDDA.n443 VDDA.t249 11.2576
R5549 VDDA.n444 VDDA.t326 11.2576
R5550 VDDA.n423 VDDA.t356 11.2576
R5551 VDDA.n285 VDDA.t257 11.2576
R5552 VDDA.n285 VDDA.t227 11.2576
R5553 VDDA.n235 VDDA.t237 11.2576
R5554 VDDA.n235 VDDA.t247 11.2576
R5555 VDDA.n244 VDDA.t233 11.2576
R5556 VDDA.n244 VDDA.t229 11.2576
R5557 VDDA.n259 VDDA.t289 11.2576
R5558 VDDA.n237 VDDA.t362 11.2576
R5559 VDDA.n280 VDDA.t239 11.2576
R5560 VDDA.n280 VDDA.t251 11.2576
R5561 VDDA.n282 VDDA.t225 11.2576
R5562 VDDA.n282 VDDA.t231 11.2576
R5563 VDDA.n50 VDDA.t221 11.2576
R5564 VDDA.n50 VDDA.t223 11.2576
R5565 VDDA.n0 VDDA.t253 11.2576
R5566 VDDA.n0 VDDA.t259 11.2576
R5567 VDDA.n9 VDDA.t245 11.2576
R5568 VDDA.n9 VDDA.t241 11.2576
R5569 VDDA.n24 VDDA.t320 11.2576
R5570 VDDA.n2 VDDA.t274 11.2576
R5571 VDDA.n45 VDDA.t255 11.2576
R5572 VDDA.n45 VDDA.t261 11.2576
R5573 VDDA.n47 VDDA.t235 11.2576
R5574 VDDA.n47 VDDA.t243 11.2576
R5575 VDDA.n477 VDDA.n476 11.1572
R5576 VDDA.n320 VDDA.n297 10.8443
R5577 VDDA.n85 VDDA.n62 10.8443
R5578 VDDA.n601 VDDA.n600 9.7855
R5579 VDDA.n463 VDDA.n424 9.14336
R5580 VDDA.n459 VDDA.n458 9.14336
R5581 VDDA.n456 VDDA.n453 9.14336
R5582 VDDA.n445 VDDA.n431 9.14336
R5583 VDDA.n436 VDDA.n433 9.14336
R5584 VDDA.n441 VDDA.n438 9.14336
R5585 VDDA.n404 VDDA.n379 9.14336
R5586 VDDA.n404 VDDA.n403 9.14336
R5587 VDDA.n403 VDDA.n402 9.14336
R5588 VDDA.n402 VDDA.n399 9.14336
R5589 VDDA.n399 VDDA.n398 9.14336
R5590 VDDA.n398 VDDA.n395 9.14336
R5591 VDDA.n395 VDDA.n394 9.14336
R5592 VDDA.n394 VDDA.n391 9.14336
R5593 VDDA.n391 VDDA.n390 9.14336
R5594 VDDA.n372 VDDA.n346 9.14336
R5595 VDDA.n372 VDDA.n369 9.14336
R5596 VDDA.n369 VDDA.n368 9.14336
R5597 VDDA.n368 VDDA.n365 9.14336
R5598 VDDA.n365 VDDA.n364 9.14336
R5599 VDDA.n364 VDDA.n361 9.14336
R5600 VDDA.n361 VDDA.n360 9.14336
R5601 VDDA.n360 VDDA.n357 9.14336
R5602 VDDA.n357 VDDA.n356 9.14336
R5603 VDDA.n306 VDDA.n304 9.14336
R5604 VDDA.n316 VDDA.n315 9.14336
R5605 VDDA.n278 VDDA.n238 9.14336
R5606 VDDA.n274 VDDA.n273 9.14336
R5607 VDDA.n271 VDDA.n268 9.14336
R5608 VDDA.n260 VDDA.n247 9.14336
R5609 VDDA.n252 VDDA.n249 9.14336
R5610 VDDA.n257 VDDA.n254 9.14336
R5611 VDDA.n230 VDDA.n180 9.14336
R5612 VDDA.n226 VDDA.n225 9.14336
R5613 VDDA.n201 VDDA.n189 9.14336
R5614 VDDA.n196 VDDA.n195 9.14336
R5615 VDDA.n169 VDDA.n144 9.14336
R5616 VDDA.n169 VDDA.n168 9.14336
R5617 VDDA.n168 VDDA.n167 9.14336
R5618 VDDA.n167 VDDA.n164 9.14336
R5619 VDDA.n164 VDDA.n163 9.14336
R5620 VDDA.n163 VDDA.n160 9.14336
R5621 VDDA.n160 VDDA.n159 9.14336
R5622 VDDA.n159 VDDA.n156 9.14336
R5623 VDDA.n156 VDDA.n155 9.14336
R5624 VDDA.n133 VDDA.n132 9.14336
R5625 VDDA.n132 VDDA.n131 9.14336
R5626 VDDA.n131 VDDA.n109 9.14336
R5627 VDDA.n127 VDDA.n109 9.14336
R5628 VDDA.n127 VDDA.n126 9.14336
R5629 VDDA.n126 VDDA.n114 9.14336
R5630 VDDA.n122 VDDA.n114 9.14336
R5631 VDDA.n122 VDDA.n121 9.14336
R5632 VDDA.n121 VDDA.n120 9.14336
R5633 VDDA.n69 VDDA.n67 9.14336
R5634 VDDA.n78 VDDA.n77 9.14336
R5635 VDDA.n43 VDDA.n3 9.14336
R5636 VDDA.n39 VDDA.n38 9.14336
R5637 VDDA.n36 VDDA.n33 9.14336
R5638 VDDA.n25 VDDA.n12 9.14336
R5639 VDDA.n17 VDDA.n14 9.14336
R5640 VDDA.n22 VDDA.n19 9.14336
R5641 VDDA.n584 VDDA.n579 9.14336
R5642 VDDA.n584 VDDA.n583 9.14336
R5643 VDDA.n583 VDDA.n581 9.14336
R5644 VDDA.n572 VDDA.n571 9.14336
R5645 VDDA.n571 VDDA.n570 9.14336
R5646 VDDA.n570 VDDA.n545 9.14336
R5647 VDDA.n532 VDDA.n531 8.973
R5648 VDDA.n412 VDDA.n411 8.8755
R5649 VDDA.n234 VDDA.n233 8.28175
R5650 VDDA.n233 VDDA.n232 8.188
R5651 VDDA.n412 VDDA.n286 8.15675
R5652 VDDA.n234 VDDA.n51 8.15675
R5653 VDDA.n296 VDDA.t262 8.0005
R5654 VDDA.n296 VDDA.t168 8.0005
R5655 VDDA.n294 VDDA.t198 8.0005
R5656 VDDA.n294 VDDA.t196 8.0005
R5657 VDDA.n292 VDDA.t71 8.0005
R5658 VDDA.n292 VDDA.t116 8.0005
R5659 VDDA.n290 VDDA.t193 8.0005
R5660 VDDA.n290 VDDA.t169 8.0005
R5661 VDDA.n288 VDDA.t66 8.0005
R5662 VDDA.n288 VDDA.t386 8.0005
R5663 VDDA.n287 VDDA.t387 8.0005
R5664 VDDA.n287 VDDA.t263 8.0005
R5665 VDDA.n61 VDDA.t39 8.0005
R5666 VDDA.n61 VDDA.t265 8.0005
R5667 VDDA.n59 VDDA.t62 8.0005
R5668 VDDA.n59 VDDA.t139 8.0005
R5669 VDDA.n57 VDDA.t75 8.0005
R5670 VDDA.n57 VDDA.t140 8.0005
R5671 VDDA.n55 VDDA.t127 8.0005
R5672 VDDA.n55 VDDA.t147 8.0005
R5673 VDDA.n53 VDDA.t61 8.0005
R5674 VDDA.n53 VDDA.t79 8.0005
R5675 VDDA.n52 VDDA.t264 8.0005
R5676 VDDA.n52 VDDA.t149 8.0005
R5677 VDDA.n321 VDDA.t58 6.56717
R5678 VDDA.n321 VDDA.t68 6.56717
R5679 VDDA.n337 VDDA.t56 6.56717
R5680 VDDA.n337 VDDA.t115 6.56717
R5681 VDDA.n339 VDDA.t54 6.56717
R5682 VDDA.n339 VDDA.t195 6.56717
R5683 VDDA.n341 VDDA.t20 6.56717
R5684 VDDA.n341 VDDA.t393 6.56717
R5685 VDDA.n343 VDDA.t118 6.56717
R5686 VDDA.n343 VDDA.t120 6.56717
R5687 VDDA.n86 VDDA.t142 6.56717
R5688 VDDA.n86 VDDA.t126 6.56717
R5689 VDDA.n97 VDDA.t144 6.56717
R5690 VDDA.n97 VDDA.t136 6.56717
R5691 VDDA.n99 VDDA.t78 6.56717
R5692 VDDA.n99 VDDA.t60 6.56717
R5693 VDDA.n101 VDDA.t12 6.56717
R5694 VDDA.n101 VDDA.t74 6.56717
R5695 VDDA.n103 VDDA.t41 6.56717
R5696 VDDA.n103 VDDA.t138 6.56717
R5697 VDDA.n421 VDDA.n413 6.563
R5698 VDDA.n413 VDDA.n412 6.0005
R5699 VDDA.n413 VDDA.n234 6.0005
R5700 VDDA.n411 VDDA.n410 5.8755
R5701 VDDA.n176 VDDA.n175 5.8755
R5702 VDDA.n408 VDDA.n323 5.33286
R5703 VDDA.n375 VDDA.n374 5.33286
R5704 VDDA.n318 VDDA.n317 5.33286
R5705 VDDA.n309 VDDA.n308 5.33286
R5706 VDDA.n135 VDDA.n134 5.33286
R5707 VDDA.n173 VDDA.n88 5.33286
R5708 VDDA.n72 VDDA.n71 5.33286
R5709 VDDA.n83 VDDA.n63 5.33286
R5710 VDDA.n590 VDDA.n535 5.33286
R5711 VDDA.n568 VDDA.n567 5.33286
R5712 VDDA.n466 VDDA.n465 5.28175
R5713 VDDA.n421 VDDA.n420 5.28175
R5714 VDDA.n600 VDDA.n599 5.0005
R5715 VDDA.n411 VDDA.n320 4.96925
R5716 VDDA.n176 VDDA.n85 4.96925
R5717 VDDA.n477 VDDA.n473 4.5595
R5718 VDDA.n481 VDDA.n480 4.54311
R5719 VDDA.n529 VDDA.n481 4.54311
R5720 VDDA.n451 VDDA.n424 4.53698
R5721 VDDA.n458 VDDA.n457 4.53698
R5722 VDDA.n453 VDDA.n452 4.53698
R5723 VDDA.n459 VDDA.n451 4.53698
R5724 VDDA.n457 VDDA.n456 4.53698
R5725 VDDA.n432 VDDA.n431 4.53698
R5726 VDDA.n437 VDDA.n436 4.53698
R5727 VDDA.n442 VDDA.n441 4.53698
R5728 VDDA.n433 VDDA.n432 4.53698
R5729 VDDA.n438 VDDA.n437 4.53698
R5730 VDDA.n266 VDDA.n238 4.53698
R5731 VDDA.n273 VDDA.n272 4.53698
R5732 VDDA.n268 VDDA.n267 4.53698
R5733 VDDA.n274 VDDA.n266 4.53698
R5734 VDDA.n272 VDDA.n271 4.53698
R5735 VDDA.n248 VDDA.n247 4.53698
R5736 VDDA.n253 VDDA.n252 4.53698
R5737 VDDA.n258 VDDA.n257 4.53698
R5738 VDDA.n249 VDDA.n248 4.53698
R5739 VDDA.n254 VDDA.n253 4.53698
R5740 VDDA.n223 VDDA.n180 4.53698
R5741 VDDA.n225 VDDA.n224 4.53698
R5742 VDDA.n226 VDDA.n223 4.53698
R5743 VDDA.n193 VDDA.n189 4.53698
R5744 VDDA.n197 VDDA.n196 4.53698
R5745 VDDA.n195 VDDA.n193 4.53698
R5746 VDDA.n31 VDDA.n3 4.53698
R5747 VDDA.n38 VDDA.n37 4.53698
R5748 VDDA.n33 VDDA.n32 4.53698
R5749 VDDA.n39 VDDA.n31 4.53698
R5750 VDDA.n37 VDDA.n36 4.53698
R5751 VDDA.n13 VDDA.n12 4.53698
R5752 VDDA.n18 VDDA.n17 4.53698
R5753 VDDA.n23 VDDA.n22 4.53698
R5754 VDDA.n14 VDDA.n13 4.53698
R5755 VDDA.n19 VDDA.n18 4.53698
R5756 VDDA.n286 VDDA.n284 4.5005
R5757 VDDA.n51 VDDA.n49 4.5005
R5758 VDDA.n599 VDDA.n597 4.5005
R5759 VDDA.n527 VDDA.n482 4.48641
R5760 VDDA.n527 VDDA.n526 4.48641
R5761 VDDA.n504 VDDA.n485 4.48641
R5762 VDDA.n504 VDDA.n503 4.48641
R5763 VDDA.n475 VDDA.n474 4.12334
R5764 VDDA.n379 VDDA.n323 3.75335
R5765 VDDA.n390 VDDA.n388 3.75335
R5766 VDDA.n374 VDDA.n346 3.75335
R5767 VDDA.n356 VDDA.n354 3.75335
R5768 VDDA.n308 VDDA.n304 3.75335
R5769 VDDA.n307 VDDA.n306 3.75335
R5770 VDDA.n317 VDDA.n316 3.75335
R5771 VDDA.n315 VDDA.n314 3.75335
R5772 VDDA.n144 VDDA.n88 3.75335
R5773 VDDA.n155 VDDA.n153 3.75335
R5774 VDDA.n134 VDDA.n133 3.75335
R5775 VDDA.n120 VDDA.n119 3.75335
R5776 VDDA.n71 VDDA.n67 3.75335
R5777 VDDA.n70 VDDA.n69 3.75335
R5778 VDDA.n77 VDDA.n63 3.75335
R5779 VDDA.n79 VDDA.n78 3.75335
R5780 VDDA.n586 VDDA.n579 3.75335
R5781 VDDA.n581 VDDA.n535 3.75335
R5782 VDDA.n573 VDDA.n572 3.75335
R5783 VDDA.n568 VDDA.n545 3.75335
R5784 VDDA.n638 VDDA.n637 3.71013
R5785 VDDA.n476 VDDA.n475 3.43377
R5786 VDDA.n209 VDDA.n208 2.8957
R5787 VDDA.n210 VDDA.n209 2.8957
R5788 VDDA.n214 VDDA.n212 2.8957
R5789 VDDA.n217 VDDA.n212 2.8957
R5790 VDDA.n213 VDDA.n210 2.8957
R5791 VDDA.n217 VDDA.n216 2.8957
R5792 VDDA.n219 VDDA.n208 2.8957
R5793 VDDA.n214 VDDA.n213 2.8957
R5794 VDDA.n600 VDDA.n592 2.5005
R5795 VDDA.n219 VDDA.n207 2.32777
R5796 VDDA.n638 VDDA.n467 2.1343
R5797 VDDA VDDA.n638 2.0779
R5798 VDDA.n524 VDDA.n507 1.8755
R5799 VDDA.n565 VDDA.n550 1.84425
R5800 VDDA.n623 VDDA.n614 1.813
R5801 VDDA.n631 VDDA.n628 1.813
R5802 VDDA.n565 VDDA.n564 1.0005
R5803 VDDA.n564 VDDA.n562 1.0005
R5804 VDDA.n562 VDDA.n560 1.0005
R5805 VDDA.n560 VDDA.n558 1.0005
R5806 VDDA.n558 VDDA.n556 1.0005
R5807 VDDA.n556 VDDA.n554 1.0005
R5808 VDDA.n554 VDDA.n552 1.0005
R5809 VDDA.n552 VDDA.n534 1.0005
R5810 VDDA.n592 VDDA.n534 1.0005
R5811 VDDA.n466 VDDA.n421 0.938
R5812 VDDA.n205 VDDA.n204 0.922375
R5813 VDDA.n187 VDDA.n178 0.922375
R5814 VDDA.n232 VDDA.n178 0.922375
R5815 VDDA.n532 VDDA.n477 0.840625
R5816 VDDA.n601 VDDA.n532 0.74075
R5817 VDDA.n465 VDDA.n422 0.6255
R5818 VDDA.n420 VDDA.n415 0.6255
R5819 VDDA.n284 VDDA.n283 0.6255
R5820 VDDA.n283 VDDA.n281 0.6255
R5821 VDDA.n245 VDDA.n236 0.6255
R5822 VDDA.n284 VDDA.n236 0.6255
R5823 VDDA.n49 VDDA.n48 0.6255
R5824 VDDA.n48 VDDA.n46 0.6255
R5825 VDDA.n10 VDDA.n1 0.6255
R5826 VDDA.n49 VDDA.n1 0.6255
R5827 VDDA.n501 VDDA.n499 0.6255
R5828 VDDA.n499 VDDA.n497 0.6255
R5829 VDDA.n497 VDDA.n495 0.6255
R5830 VDDA.n495 VDDA.n493 0.6255
R5831 VDDA.n493 VDDA.n491 0.6255
R5832 VDDA.n491 VDDA.n489 0.6255
R5833 VDDA.n489 VDDA.n487 0.6255
R5834 VDDA.n487 VDDA.n484 0.6255
R5835 VDDA.n507 VDDA.n484 0.6255
R5836 VDDA.n524 VDDA.n523 0.6255
R5837 VDDA.n523 VDDA.n521 0.6255
R5838 VDDA.n521 VDDA.n519 0.6255
R5839 VDDA.n519 VDDA.n517 0.6255
R5840 VDDA.n517 VDDA.n515 0.6255
R5841 VDDA.n515 VDDA.n513 0.6255
R5842 VDDA.n513 VDDA.n511 0.6255
R5843 VDDA.n511 VDDA.n509 0.6255
R5844 VDDA.n509 VDDA.n479 0.6255
R5845 VDDA.n531 VDDA.n479 0.6255
R5846 VDDA.n344 VDDA.n342 0.563
R5847 VDDA.n342 VDDA.n340 0.563
R5848 VDDA.n340 VDDA.n338 0.563
R5849 VDDA.n338 VDDA.n322 0.563
R5850 VDDA.n410 VDDA.n322 0.563
R5851 VDDA.n291 VDDA.n289 0.563
R5852 VDDA.n293 VDDA.n291 0.563
R5853 VDDA.n295 VDDA.n293 0.563
R5854 VDDA.n297 VDDA.n295 0.563
R5855 VDDA.n104 VDDA.n102 0.563
R5856 VDDA.n102 VDDA.n100 0.563
R5857 VDDA.n100 VDDA.n98 0.563
R5858 VDDA.n98 VDDA.n87 0.563
R5859 VDDA.n175 VDDA.n87 0.563
R5860 VDDA.n56 VDDA.n54 0.563
R5861 VDDA.n58 VDDA.n56 0.563
R5862 VDDA.n60 VDDA.n58 0.563
R5863 VDDA.n62 VDDA.n60 0.563
R5864 VDDA.n609 VDDA.n607 0.563
R5865 VDDA.n614 VDDA.n607 0.563
R5866 VDDA.n623 VDDA.n622 0.563
R5867 VDDA.n622 VDDA.n620 0.563
R5868 VDDA.n620 VDDA.n618 0.563
R5869 VDDA.n618 VDDA.n616 0.563
R5870 VDDA.n616 VDDA.n605 0.563
R5871 VDDA.n628 VDDA.n605 0.563
R5872 VDDA.n631 VDDA.n630 0.563
R5873 VDDA.n630 VDDA.n603 0.563
R5874 VDDA.n636 VDDA.n603 0.563
R5875 VDDA.n233 VDDA.n176 0.46925
R5876 VDDA VDDA.n601 0.41175
R5877 VDDA.n205 VDDA.n187 0.3755
R5878 VDDA.t95 VDDA.t2 0.1603
R5879 VDDA.t123 VDDA.t100 0.1603
R5880 VDDA.t83 VDDA.t50 0.1603
R5881 VDDA.t408 VDDA.t104 0.1603
R5882 VDDA.t391 VDDA.t133 0.1603
R5883 VDDA.n469 VDDA.t134 0.159278
R5884 VDDA.n470 VDDA.t121 0.159278
R5885 VDDA.n471 VDDA.t52 0.159278
R5886 VDDA.n472 VDDA.t103 0.159278
R5887 VDDA.n472 VDDA.t390 0.1368
R5888 VDDA.n472 VDDA.t95 0.1368
R5889 VDDA.n471 VDDA.t51 0.1368
R5890 VDDA.n471 VDDA.t123 0.1368
R5891 VDDA.n470 VDDA.t23 0.1368
R5892 VDDA.n470 VDDA.t83 0.1368
R5893 VDDA.n469 VDDA.t92 0.1368
R5894 VDDA.n469 VDDA.t408 0.1368
R5895 VDDA.n468 VDDA.t122 0.1368
R5896 VDDA.n468 VDDA.t391 0.1368
R5897 VDDA.n637 VDDA 0.135625
R5898 VDDA.t134 VDDA.n468 0.00152174
R5899 VDDA.t121 VDDA.n469 0.00152174
R5900 VDDA.t52 VDDA.n470 0.00152174
R5901 VDDA.t103 VDDA.n471 0.00152174
R5902 VDDA.t3 VDDA.n472 0.00152174
R5903 bgr_0.V_TOP.n0 bgr_0.V_TOP.t29 369.534
R5904 bgr_0.V_TOP.n23 bgr_0.V_TOP.n21 339.961
R5905 bgr_0.V_TOP.n23 bgr_0.V_TOP.n22 339.272
R5906 bgr_0.V_TOP.n19 bgr_0.V_TOP.n18 339.272
R5907 bgr_0.V_TOP.n27 bgr_0.V_TOP.n26 339.272
R5908 bgr_0.V_TOP.n29 bgr_0.V_TOP.n28 339.272
R5909 bgr_0.V_TOP.n24 bgr_0.V_TOP.n20 334.772
R5910 bgr_0.V_TOP.n39 bgr_0.V_TOP.n38 224.934
R5911 bgr_0.V_TOP.n38 bgr_0.V_TOP.n37 224.934
R5912 bgr_0.V_TOP.n37 bgr_0.V_TOP.n36 224.934
R5913 bgr_0.V_TOP.n36 bgr_0.V_TOP.n35 224.934
R5914 bgr_0.V_TOP.n35 bgr_0.V_TOP.n34 224.934
R5915 bgr_0.V_TOP.n34 bgr_0.V_TOP.n33 224.934
R5916 bgr_0.V_TOP.n33 bgr_0.V_TOP.n32 224.934
R5917 bgr_0.V_TOP.n1 bgr_0.V_TOP.n0 224.934
R5918 bgr_0.V_TOP.n2 bgr_0.V_TOP.n1 224.934
R5919 bgr_0.V_TOP.n3 bgr_0.V_TOP.n2 224.934
R5920 bgr_0.V_TOP.n4 bgr_0.V_TOP.n3 224.934
R5921 bgr_0.V_TOP.n5 bgr_0.V_TOP.n4 224.934
R5922 bgr_0.V_TOP bgr_0.V_TOP.t48 214.222
R5923 bgr_0.V_TOP.n31 bgr_0.V_TOP.n30 163.175
R5924 bgr_0.V_TOP.n39 bgr_0.V_TOP.t24 144.601
R5925 bgr_0.V_TOP.n38 bgr_0.V_TOP.t33 144.601
R5926 bgr_0.V_TOP.n37 bgr_0.V_TOP.t39 144.601
R5927 bgr_0.V_TOP.n36 bgr_0.V_TOP.t16 144.601
R5928 bgr_0.V_TOP.n35 bgr_0.V_TOP.t15 144.601
R5929 bgr_0.V_TOP.n34 bgr_0.V_TOP.t28 144.601
R5930 bgr_0.V_TOP.n33 bgr_0.V_TOP.t38 144.601
R5931 bgr_0.V_TOP.n32 bgr_0.V_TOP.t14 144.601
R5932 bgr_0.V_TOP.n0 bgr_0.V_TOP.t30 144.601
R5933 bgr_0.V_TOP.n1 bgr_0.V_TOP.t18 144.601
R5934 bgr_0.V_TOP.n2 bgr_0.V_TOP.t46 144.601
R5935 bgr_0.V_TOP.n3 bgr_0.V_TOP.t37 144.601
R5936 bgr_0.V_TOP.n4 bgr_0.V_TOP.t26 144.601
R5937 bgr_0.V_TOP.n5 bgr_0.V_TOP.t27 144.601
R5938 bgr_0.V_TOP.n17 bgr_0.V_TOP.t12 108.424
R5939 bgr_0.V_TOP.n30 bgr_0.V_TOP.t5 95.4467
R5940 bgr_0.V_TOP bgr_0.V_TOP.n39 69.6227
R5941 bgr_0.V_TOP.n32 bgr_0.V_TOP.n31 69.6227
R5942 bgr_0.V_TOP.n31 bgr_0.V_TOP.n5 69.6227
R5943 bgr_0.V_TOP.n18 bgr_0.V_TOP.t6 39.4005
R5944 bgr_0.V_TOP.n18 bgr_0.V_TOP.t10 39.4005
R5945 bgr_0.V_TOP.n20 bgr_0.V_TOP.t4 39.4005
R5946 bgr_0.V_TOP.n20 bgr_0.V_TOP.t3 39.4005
R5947 bgr_0.V_TOP.n22 bgr_0.V_TOP.t0 39.4005
R5948 bgr_0.V_TOP.n22 bgr_0.V_TOP.t9 39.4005
R5949 bgr_0.V_TOP.n21 bgr_0.V_TOP.t8 39.4005
R5950 bgr_0.V_TOP.n21 bgr_0.V_TOP.t2 39.4005
R5951 bgr_0.V_TOP.n26 bgr_0.V_TOP.t1 39.4005
R5952 bgr_0.V_TOP.n26 bgr_0.V_TOP.t13 39.4005
R5953 bgr_0.V_TOP.n28 bgr_0.V_TOP.t11 39.4005
R5954 bgr_0.V_TOP.n28 bgr_0.V_TOP.t7 39.4005
R5955 bgr_0.V_TOP.n17 bgr_0.V_TOP.n16 37.1479
R5956 bgr_0.V_TOP.n19 bgr_0.V_TOP.n17 27.8371
R5957 bgr_0.V_TOP.n24 bgr_0.V_TOP.n23 8.313
R5958 bgr_0.V_TOP.n30 bgr_0.V_TOP.n29 5.188
R5959 bgr_0.V_TOP.n6 bgr_0.V_TOP.t31 4.8295
R5960 bgr_0.V_TOP.n7 bgr_0.V_TOP.t22 4.8295
R5961 bgr_0.V_TOP.n8 bgr_0.V_TOP.t20 4.8295
R5962 bgr_0.V_TOP.n9 bgr_0.V_TOP.t45 4.8295
R5963 bgr_0.V_TOP.n10 bgr_0.V_TOP.t42 4.8295
R5964 bgr_0.V_TOP.n11 bgr_0.V_TOP.t36 4.8295
R5965 bgr_0.V_TOP.n12 bgr_0.V_TOP.t17 4.8295
R5966 bgr_0.V_TOP.n13 bgr_0.V_TOP.t43 4.8295
R5967 bgr_0.V_TOP.n14 bgr_0.V_TOP.t34 4.8295
R5968 bgr_0.V_TOP.n6 bgr_0.V_TOP.t35 4.5005
R5969 bgr_0.V_TOP.n7 bgr_0.V_TOP.t32 4.5005
R5970 bgr_0.V_TOP.n8 bgr_0.V_TOP.t25 4.5005
R5971 bgr_0.V_TOP.n9 bgr_0.V_TOP.t21 4.5005
R5972 bgr_0.V_TOP.n10 bgr_0.V_TOP.t49 4.5005
R5973 bgr_0.V_TOP.n11 bgr_0.V_TOP.t44 4.5005
R5974 bgr_0.V_TOP.n12 bgr_0.V_TOP.t23 4.5005
R5975 bgr_0.V_TOP.n13 bgr_0.V_TOP.t19 4.5005
R5976 bgr_0.V_TOP.n16 bgr_0.V_TOP.t40 4.5005
R5977 bgr_0.V_TOP.n15 bgr_0.V_TOP.t47 4.5005
R5978 bgr_0.V_TOP.n14 bgr_0.V_TOP.t41 4.5005
R5979 bgr_0.V_TOP.n25 bgr_0.V_TOP.n24 4.5005
R5980 bgr_0.V_TOP.n29 bgr_0.V_TOP.n27 2.1255
R5981 bgr_0.V_TOP.n27 bgr_0.V_TOP.n25 2.1255
R5982 bgr_0.V_TOP.n25 bgr_0.V_TOP.n19 2.1255
R5983 bgr_0.V_TOP.n7 bgr_0.V_TOP.n6 0.3295
R5984 bgr_0.V_TOP.n9 bgr_0.V_TOP.n8 0.3295
R5985 bgr_0.V_TOP.n11 bgr_0.V_TOP.n10 0.3295
R5986 bgr_0.V_TOP.n13 bgr_0.V_TOP.n12 0.3295
R5987 bgr_0.V_TOP.n16 bgr_0.V_TOP.n15 0.3295
R5988 bgr_0.V_TOP.n15 bgr_0.V_TOP.n14 0.3295
R5989 bgr_0.V_TOP.n9 bgr_0.V_TOP.n7 0.2825
R5990 bgr_0.V_TOP.n11 bgr_0.V_TOP.n9 0.2825
R5991 bgr_0.V_TOP.n13 bgr_0.V_TOP.n11 0.2825
R5992 bgr_0.V_TOP.n14 bgr_0.V_TOP.n13 0.2825
R5993 VOUT-.n8 VOUT-.n0 149.19
R5994 VOUT-.n3 VOUT-.n1 149.19
R5995 VOUT-.n7 VOUT-.n6 148.626
R5996 VOUT-.n5 VOUT-.n4 148.626
R5997 VOUT-.n3 VOUT-.n2 148.626
R5998 VOUT-.n10 VOUT-.n9 144.126
R5999 VOUT-.n91 VOUT-.t3 112.184
R6000 VOUT-.n88 VOUT-.n86 98.9303
R6001 VOUT-.n90 VOUT-.n89 97.8053
R6002 VOUT-.n88 VOUT-.n87 97.8053
R6003 VOUT-.n85 VOUT-.n10 15.5682
R6004 VOUT-.n85 VOUT-.n84 11.5649
R6005 VOUT- VOUT-.n85 9.46925
R6006 VOUT-.n9 VOUT-.t11 6.56717
R6007 VOUT-.n9 VOUT-.t0 6.56717
R6008 VOUT-.n6 VOUT-.t7 6.56717
R6009 VOUT-.n6 VOUT-.t8 6.56717
R6010 VOUT-.n4 VOUT-.t4 6.56717
R6011 VOUT-.n4 VOUT-.t13 6.56717
R6012 VOUT-.n2 VOUT-.t10 6.56717
R6013 VOUT-.n2 VOUT-.t12 6.56717
R6014 VOUT-.n1 VOUT-.t9 6.56717
R6015 VOUT-.n1 VOUT-.t17 6.56717
R6016 VOUT-.n0 VOUT-.t16 6.56717
R6017 VOUT-.n0 VOUT-.t2 6.56717
R6018 VOUT-.n39 VOUT-.t68 4.8295
R6019 VOUT-.n47 VOUT-.t66 4.8295
R6020 VOUT-.n45 VOUT-.t115 4.8295
R6021 VOUT-.n43 VOUT-.t150 4.8295
R6022 VOUT-.n42 VOUT-.t132 4.8295
R6023 VOUT-.n41 VOUT-.t29 4.8295
R6024 VOUT-.n59 VOUT-.t125 4.8295
R6025 VOUT-.n60 VOUT-.t73 4.8295
R6026 VOUT-.n61 VOUT-.t23 4.8295
R6027 VOUT-.n62 VOUT-.t109 4.8295
R6028 VOUT-.n63 VOUT-.t76 4.8295
R6029 VOUT-.n64 VOUT-.t44 4.8295
R6030 VOUT-.n66 VOUT-.t37 4.8295
R6031 VOUT-.n67 VOUT-.t143 4.8295
R6032 VOUT-.n69 VOUT-.t70 4.8295
R6033 VOUT-.n70 VOUT-.t39 4.8295
R6034 VOUT-.n72 VOUT-.t32 4.8295
R6035 VOUT-.n73 VOUT-.t138 4.8295
R6036 VOUT-.n75 VOUT-.t131 4.8295
R6037 VOUT-.n76 VOUT-.t101 4.8295
R6038 VOUT-.n78 VOUT-.t28 4.8295
R6039 VOUT-.n79 VOUT-.t133 4.8295
R6040 VOUT-.n11 VOUT-.t26 4.8295
R6041 VOUT-.n13 VOUT-.t36 4.8295
R6042 VOUT-.n24 VOUT-.t140 4.8295
R6043 VOUT-.n25 VOUT-.t111 4.8295
R6044 VOUT-.n27 VOUT-.t41 4.8295
R6045 VOUT-.n28 VOUT-.t151 4.8295
R6046 VOUT-.n30 VOUT-.t80 4.8295
R6047 VOUT-.n31 VOUT-.t51 4.8295
R6048 VOUT-.n33 VOUT-.t49 4.8295
R6049 VOUT-.n34 VOUT-.t19 4.8295
R6050 VOUT-.n36 VOUT-.t85 4.8295
R6051 VOUT-.n37 VOUT-.t55 4.8295
R6052 VOUT-.n81 VOUT-.t124 4.8295
R6053 VOUT-.n49 VOUT-.t91 4.8154
R6054 VOUT-.n50 VOUT-.t69 4.8154
R6055 VOUT-.n51 VOUT-.t107 4.8154
R6056 VOUT-.n49 VOUT-.t31 4.806
R6057 VOUT-.n50 VOUT-.t149 4.806
R6058 VOUT-.n51 VOUT-.t50 4.806
R6059 VOUT-.n52 VOUT-.t144 4.806
R6060 VOUT-.n52 VOUT-.t83 4.806
R6061 VOUT-.n53 VOUT-.t120 4.806
R6062 VOUT-.n54 VOUT-.t104 4.806
R6063 VOUT-.n55 VOUT-.t137 4.806
R6064 VOUT-.n56 VOUT-.t35 4.806
R6065 VOUT-.n57 VOUT-.t156 4.806
R6066 VOUT-.n14 VOUT-.t71 4.806
R6067 VOUT-.n14 VOUT-.t113 4.806
R6068 VOUT-.n15 VOUT-.t114 4.806
R6069 VOUT-.n15 VOUT-.t24 4.806
R6070 VOUT-.n16 VOUT-.t65 4.806
R6071 VOUT-.n16 VOUT-.t62 4.806
R6072 VOUT-.n17 VOUT-.t154 4.806
R6073 VOUT-.n17 VOUT-.t95 4.806
R6074 VOUT-.n18 VOUT-.t105 4.806
R6075 VOUT-.n18 VOUT-.t126 4.806
R6076 VOUT-.n19 VOUT-.t141 4.806
R6077 VOUT-.n19 VOUT-.t38 4.806
R6078 VOUT-.n20 VOUT-.t92 4.806
R6079 VOUT-.n20 VOUT-.t74 4.806
R6080 VOUT-.n21 VOUT-.t42 4.806
R6081 VOUT-.n22 VOUT-.t82 4.806
R6082 VOUT-.n39 VOUT-.t86 4.5005
R6083 VOUT-.n40 VOUT-.t54 4.5005
R6084 VOUT-.n47 VOUT-.t77 4.5005
R6085 VOUT-.n48 VOUT-.t43 4.5005
R6086 VOUT-.n45 VOUT-.t58 4.5005
R6087 VOUT-.n46 VOUT-.t22 4.5005
R6088 VOUT-.n43 VOUT-.t94 4.5005
R6089 VOUT-.n44 VOUT-.t61 4.5005
R6090 VOUT-.n42 VOUT-.t99 4.5005
R6091 VOUT-.n41 VOUT-.t52 4.5005
R6092 VOUT-.n58 VOUT-.t155 4.5005
R6093 VOUT-.n57 VOUT-.t116 4.5005
R6094 VOUT-.n56 VOUT-.t136 4.5005
R6095 VOUT-.n55 VOUT-.t100 4.5005
R6096 VOUT-.n54 VOUT-.t64 4.5005
R6097 VOUT-.n53 VOUT-.t81 4.5005
R6098 VOUT-.n52 VOUT-.t45 4.5005
R6099 VOUT-.n51 VOUT-.t146 4.5005
R6100 VOUT-.n50 VOUT-.t108 4.5005
R6101 VOUT-.n49 VOUT-.t130 4.5005
R6102 VOUT-.n59 VOUT-.t152 4.5005
R6103 VOUT-.n60 VOUT-.t112 4.5005
R6104 VOUT-.n61 VOUT-.t47 4.5005
R6105 VOUT-.n62 VOUT-.t147 4.5005
R6106 VOUT-.n63 VOUT-.t27 4.5005
R6107 VOUT-.n65 VOUT-.t128 4.5005
R6108 VOUT-.n64 VOUT-.t97 4.5005
R6109 VOUT-.n66 VOUT-.t123 4.5005
R6110 VOUT-.n68 VOUT-.t88 4.5005
R6111 VOUT-.n67 VOUT-.t57 4.5005
R6112 VOUT-.n69 VOUT-.t20 4.5005
R6113 VOUT-.n71 VOUT-.t121 4.5005
R6114 VOUT-.n70 VOUT-.t87 4.5005
R6115 VOUT-.n72 VOUT-.t118 4.5005
R6116 VOUT-.n74 VOUT-.t84 4.5005
R6117 VOUT-.n73 VOUT-.t53 4.5005
R6118 VOUT-.n75 VOUT-.t79 4.5005
R6119 VOUT-.n77 VOUT-.t48 4.5005
R6120 VOUT-.n76 VOUT-.t153 4.5005
R6121 VOUT-.n78 VOUT-.t117 4.5005
R6122 VOUT-.n80 VOUT-.t78 4.5005
R6123 VOUT-.n79 VOUT-.t46 4.5005
R6124 VOUT-.n11 VOUT-.t119 4.5005
R6125 VOUT-.n12 VOUT-.t33 4.5005
R6126 VOUT-.n13 VOUT-.t122 4.5005
R6127 VOUT-.n23 VOUT-.t90 4.5005
R6128 VOUT-.n22 VOUT-.t56 4.5005
R6129 VOUT-.n21 VOUT-.t142 4.5005
R6130 VOUT-.n20 VOUT-.t110 4.5005
R6131 VOUT-.n19 VOUT-.t72 4.5005
R6132 VOUT-.n18 VOUT-.t25 4.5005
R6133 VOUT-.n17 VOUT-.t127 4.5005
R6134 VOUT-.n16 VOUT-.t93 4.5005
R6135 VOUT-.n15 VOUT-.t60 4.5005
R6136 VOUT-.n14 VOUT-.t148 4.5005
R6137 VOUT-.n24 VOUT-.t89 4.5005
R6138 VOUT-.n26 VOUT-.t59 4.5005
R6139 VOUT-.n25 VOUT-.t21 4.5005
R6140 VOUT-.n27 VOUT-.t129 4.5005
R6141 VOUT-.n29 VOUT-.t98 4.5005
R6142 VOUT-.n28 VOUT-.t63 4.5005
R6143 VOUT-.n30 VOUT-.t30 4.5005
R6144 VOUT-.n32 VOUT-.t134 4.5005
R6145 VOUT-.n31 VOUT-.t103 4.5005
R6146 VOUT-.n33 VOUT-.t135 4.5005
R6147 VOUT-.n35 VOUT-.t102 4.5005
R6148 VOUT-.n34 VOUT-.t67 4.5005
R6149 VOUT-.n36 VOUT-.t34 4.5005
R6150 VOUT-.n38 VOUT-.t139 4.5005
R6151 VOUT-.n37 VOUT-.t106 4.5005
R6152 VOUT-.n81 VOUT-.t75 4.5005
R6153 VOUT-.n82 VOUT-.t40 4.5005
R6154 VOUT-.n83 VOUT-.t145 4.5005
R6155 VOUT-.n84 VOUT-.t96 4.5005
R6156 VOUT-.n10 VOUT-.n8 4.5005
R6157 VOUT-.n89 VOUT-.t15 3.42907
R6158 VOUT-.n89 VOUT-.t6 3.42907
R6159 VOUT-.n87 VOUT-.t1 3.42907
R6160 VOUT-.n87 VOUT-.t5 3.42907
R6161 VOUT-.n86 VOUT-.t18 3.42907
R6162 VOUT-.n86 VOUT-.t14 3.42907
R6163 VOUT-.n91 VOUT-.n90 1.30519
R6164 VOUT- VOUT-.n91 1.24269
R6165 VOUT-.n90 VOUT-.n88 1.1255
R6166 VOUT-.n5 VOUT-.n3 0.563
R6167 VOUT-.n7 VOUT-.n5 0.563
R6168 VOUT-.n8 VOUT-.n7 0.563
R6169 VOUT-.n40 VOUT-.n39 0.3295
R6170 VOUT-.n48 VOUT-.n47 0.3295
R6171 VOUT-.n46 VOUT-.n45 0.3295
R6172 VOUT-.n44 VOUT-.n43 0.3295
R6173 VOUT-.n58 VOUT-.n41 0.3295
R6174 VOUT-.n58 VOUT-.n57 0.3295
R6175 VOUT-.n57 VOUT-.n56 0.3295
R6176 VOUT-.n56 VOUT-.n55 0.3295
R6177 VOUT-.n55 VOUT-.n54 0.3295
R6178 VOUT-.n54 VOUT-.n53 0.3295
R6179 VOUT-.n53 VOUT-.n52 0.3295
R6180 VOUT-.n52 VOUT-.n51 0.3295
R6181 VOUT-.n51 VOUT-.n50 0.3295
R6182 VOUT-.n50 VOUT-.n49 0.3295
R6183 VOUT-.n60 VOUT-.n59 0.3295
R6184 VOUT-.n62 VOUT-.n61 0.3295
R6185 VOUT-.n65 VOUT-.n63 0.3295
R6186 VOUT-.n65 VOUT-.n64 0.3295
R6187 VOUT-.n68 VOUT-.n66 0.3295
R6188 VOUT-.n68 VOUT-.n67 0.3295
R6189 VOUT-.n71 VOUT-.n69 0.3295
R6190 VOUT-.n71 VOUT-.n70 0.3295
R6191 VOUT-.n74 VOUT-.n72 0.3295
R6192 VOUT-.n74 VOUT-.n73 0.3295
R6193 VOUT-.n77 VOUT-.n75 0.3295
R6194 VOUT-.n77 VOUT-.n76 0.3295
R6195 VOUT-.n80 VOUT-.n78 0.3295
R6196 VOUT-.n80 VOUT-.n79 0.3295
R6197 VOUT-.n12 VOUT-.n11 0.3295
R6198 VOUT-.n23 VOUT-.n13 0.3295
R6199 VOUT-.n23 VOUT-.n22 0.3295
R6200 VOUT-.n22 VOUT-.n21 0.3295
R6201 VOUT-.n21 VOUT-.n20 0.3295
R6202 VOUT-.n20 VOUT-.n19 0.3295
R6203 VOUT-.n19 VOUT-.n18 0.3295
R6204 VOUT-.n18 VOUT-.n17 0.3295
R6205 VOUT-.n17 VOUT-.n16 0.3295
R6206 VOUT-.n16 VOUT-.n15 0.3295
R6207 VOUT-.n15 VOUT-.n14 0.3295
R6208 VOUT-.n26 VOUT-.n24 0.3295
R6209 VOUT-.n26 VOUT-.n25 0.3295
R6210 VOUT-.n29 VOUT-.n27 0.3295
R6211 VOUT-.n29 VOUT-.n28 0.3295
R6212 VOUT-.n32 VOUT-.n30 0.3295
R6213 VOUT-.n32 VOUT-.n31 0.3295
R6214 VOUT-.n35 VOUT-.n33 0.3295
R6215 VOUT-.n35 VOUT-.n34 0.3295
R6216 VOUT-.n38 VOUT-.n36 0.3295
R6217 VOUT-.n38 VOUT-.n37 0.3295
R6218 VOUT-.n82 VOUT-.n81 0.3295
R6219 VOUT-.n83 VOUT-.n82 0.3295
R6220 VOUT-.n84 VOUT-.n83 0.3295
R6221 VOUT-.n53 VOUT-.n48 0.306
R6222 VOUT-.n54 VOUT-.n46 0.306
R6223 VOUT-.n55 VOUT-.n44 0.306
R6224 VOUT-.n56 VOUT-.n42 0.306
R6225 VOUT-.n58 VOUT-.n40 0.2825
R6226 VOUT-.n60 VOUT-.n58 0.2825
R6227 VOUT-.n62 VOUT-.n60 0.2825
R6228 VOUT-.n65 VOUT-.n62 0.2825
R6229 VOUT-.n68 VOUT-.n65 0.2825
R6230 VOUT-.n71 VOUT-.n68 0.2825
R6231 VOUT-.n74 VOUT-.n71 0.2825
R6232 VOUT-.n77 VOUT-.n74 0.2825
R6233 VOUT-.n80 VOUT-.n77 0.2825
R6234 VOUT-.n23 VOUT-.n12 0.2825
R6235 VOUT-.n26 VOUT-.n23 0.2825
R6236 VOUT-.n29 VOUT-.n26 0.2825
R6237 VOUT-.n32 VOUT-.n29 0.2825
R6238 VOUT-.n35 VOUT-.n32 0.2825
R6239 VOUT-.n38 VOUT-.n35 0.2825
R6240 VOUT-.n82 VOUT-.n38 0.2825
R6241 VOUT-.n82 VOUT-.n80 0.2825
R6242 two_stage_opamp_dummy_magic_14_0.cap_res_X two_stage_opamp_dummy_magic_14_0.cap_res_X.t0 49.197
R6243 two_stage_opamp_dummy_magic_14_0.cap_res_X two_stage_opamp_dummy_magic_14_0.cap_res_X.t7 0.87
R6244 two_stage_opamp_dummy_magic_14_0.cap_res_X.t27 two_stage_opamp_dummy_magic_14_0.cap_res_X.t66 0.1603
R6245 two_stage_opamp_dummy_magic_14_0.cap_res_X.t49 two_stage_opamp_dummy_magic_14_0.cap_res_X.t88 0.1603
R6246 two_stage_opamp_dummy_magic_14_0.cap_res_X.t11 two_stage_opamp_dummy_magic_14_0.cap_res_X.t50 0.1603
R6247 two_stage_opamp_dummy_magic_14_0.cap_res_X.t112 two_stage_opamp_dummy_magic_14_0.cap_res_X.t13 0.1603
R6248 two_stage_opamp_dummy_magic_14_0.cap_res_X.t80 two_stage_opamp_dummy_magic_14_0.cap_res_X.t91 0.1603
R6249 two_stage_opamp_dummy_magic_14_0.cap_res_X.t114 two_stage_opamp_dummy_magic_14_0.cap_res_X.t80 0.1603
R6250 two_stage_opamp_dummy_magic_14_0.cap_res_X.t76 two_stage_opamp_dummy_magic_14_0.cap_res_X.t114 0.1603
R6251 two_stage_opamp_dummy_magic_14_0.cap_res_X.t99 two_stage_opamp_dummy_magic_14_0.cap_res_X.t42 0.1603
R6252 two_stage_opamp_dummy_magic_14_0.cap_res_X.t135 two_stage_opamp_dummy_magic_14_0.cap_res_X.t99 0.1603
R6253 two_stage_opamp_dummy_magic_14_0.cap_res_X.t93 two_stage_opamp_dummy_magic_14_0.cap_res_X.t135 0.1603
R6254 two_stage_opamp_dummy_magic_14_0.cap_res_X.t105 two_stage_opamp_dummy_magic_14_0.cap_res_X.t128 0.1603
R6255 two_stage_opamp_dummy_magic_14_0.cap_res_X.t71 two_stage_opamp_dummy_magic_14_0.cap_res_X.t89 0.1603
R6256 two_stage_opamp_dummy_magic_14_0.cap_res_X.t5 two_stage_opamp_dummy_magic_14_0.cap_res_X.t32 0.1603
R6257 two_stage_opamp_dummy_magic_14_0.cap_res_X.t110 two_stage_opamp_dummy_magic_14_0.cap_res_X.t134 0.1603
R6258 two_stage_opamp_dummy_magic_14_0.cap_res_X.t60 two_stage_opamp_dummy_magic_14_0.cap_res_X.t113 0.1603
R6259 two_stage_opamp_dummy_magic_14_0.cap_res_X.t130 two_stage_opamp_dummy_magic_14_0.cap_res_X.t81 0.1603
R6260 two_stage_opamp_dummy_magic_14_0.cap_res_X.t100 two_stage_opamp_dummy_magic_14_0.cap_res_X.t14 0.1603
R6261 two_stage_opamp_dummy_magic_14_0.cap_res_X.t34 two_stage_opamp_dummy_magic_14_0.cap_res_X.t120 0.1603
R6262 two_stage_opamp_dummy_magic_14_0.cap_res_X.t70 two_stage_opamp_dummy_magic_14_0.cap_res_X.t118 0.1603
R6263 two_stage_opamp_dummy_magic_14_0.cap_res_X.t137 two_stage_opamp_dummy_magic_14_0.cap_res_X.t87 0.1603
R6264 two_stage_opamp_dummy_magic_14_0.cap_res_X.t104 two_stage_opamp_dummy_magic_14_0.cap_res_X.t19 0.1603
R6265 two_stage_opamp_dummy_magic_14_0.cap_res_X.t39 two_stage_opamp_dummy_magic_14_0.cap_res_X.t125 0.1603
R6266 two_stage_opamp_dummy_magic_14_0.cap_res_X.t4 two_stage_opamp_dummy_magic_14_0.cap_res_X.t56 0.1603
R6267 two_stage_opamp_dummy_magic_14_0.cap_res_X.t78 two_stage_opamp_dummy_magic_14_0.cap_res_X.t26 0.1603
R6268 two_stage_opamp_dummy_magic_14_0.cap_res_X.t111 two_stage_opamp_dummy_magic_14_0.cap_res_X.t24 0.1603
R6269 two_stage_opamp_dummy_magic_14_0.cap_res_X.t40 two_stage_opamp_dummy_magic_14_0.cap_res_X.t129 0.1603
R6270 two_stage_opamp_dummy_magic_14_0.cap_res_X.t12 two_stage_opamp_dummy_magic_14_0.cap_res_X.t61 0.1603
R6271 two_stage_opamp_dummy_magic_14_0.cap_res_X.t82 two_stage_opamp_dummy_magic_14_0.cap_res_X.t33 0.1603
R6272 two_stage_opamp_dummy_magic_14_0.cap_res_X.t51 two_stage_opamp_dummy_magic_14_0.cap_res_X.t102 0.1603
R6273 two_stage_opamp_dummy_magic_14_0.cap_res_X.t123 two_stage_opamp_dummy_magic_14_0.cap_res_X.t72 0.1603
R6274 two_stage_opamp_dummy_magic_14_0.cap_res_X.t90 two_stage_opamp_dummy_magic_14_0.cap_res_X.t138 0.1603
R6275 two_stage_opamp_dummy_magic_14_0.cap_res_X.t22 two_stage_opamp_dummy_magic_14_0.cap_res_X.t108 0.1603
R6276 two_stage_opamp_dummy_magic_14_0.cap_res_X.t54 two_stage_opamp_dummy_magic_14_0.cap_res_X.t106 0.1603
R6277 two_stage_opamp_dummy_magic_14_0.cap_res_X.t127 two_stage_opamp_dummy_magic_14_0.cap_res_X.t77 0.1603
R6278 two_stage_opamp_dummy_magic_14_0.cap_res_X.t94 two_stage_opamp_dummy_magic_14_0.cap_res_X.t6 0.1603
R6279 two_stage_opamp_dummy_magic_14_0.cap_res_X.t28 two_stage_opamp_dummy_magic_14_0.cap_res_X.t116 0.1603
R6280 two_stage_opamp_dummy_magic_14_0.cap_res_X.t136 two_stage_opamp_dummy_magic_14_0.cap_res_X.t46 0.1603
R6281 two_stage_opamp_dummy_magic_14_0.cap_res_X.t68 two_stage_opamp_dummy_magic_14_0.cap_res_X.t17 0.1603
R6282 two_stage_opamp_dummy_magic_14_0.cap_res_X.t9 two_stage_opamp_dummy_magic_14_0.cap_res_X.t86 0.1603
R6283 two_stage_opamp_dummy_magic_14_0.cap_res_X.t97 two_stage_opamp_dummy_magic_14_0.cap_res_X.t43 0.1603
R6284 two_stage_opamp_dummy_magic_14_0.cap_res_X.t64 two_stage_opamp_dummy_magic_14_0.cap_res_X.t92 0.1603
R6285 two_stage_opamp_dummy_magic_14_0.cap_res_X.t30 two_stage_opamp_dummy_magic_14_0.cap_res_X.t3 0.1603
R6286 two_stage_opamp_dummy_magic_14_0.cap_res_X.t132 two_stage_opamp_dummy_magic_14_0.cap_res_X.t52 0.1603
R6287 two_stage_opamp_dummy_magic_14_0.cap_res_X.t85 two_stage_opamp_dummy_magic_14_0.cap_res_X.t16 0.1603
R6288 two_stage_opamp_dummy_magic_14_0.cap_res_X.t47 two_stage_opamp_dummy_magic_14_0.cap_res_X.t65 0.1603
R6289 two_stage_opamp_dummy_magic_14_0.cap_res_X.t15 two_stage_opamp_dummy_magic_14_0.cap_res_X.t115 0.1603
R6290 two_stage_opamp_dummy_magic_14_0.cap_res_X.t101 two_stage_opamp_dummy_magic_14_0.cap_res_X.t75 0.1603
R6291 two_stage_opamp_dummy_magic_14_0.cap_res_X.t35 two_stage_opamp_dummy_magic_14_0.cap_res_X.t121 0.1603
R6292 two_stage_opamp_dummy_magic_14_0.cap_res_X.t38 two_stage_opamp_dummy_magic_14_0.cap_res_X.t131 0.1603
R6293 two_stage_opamp_dummy_magic_14_0.cap_res_X.t58 two_stage_opamp_dummy_magic_14_0.cap_res_X.t25 0.1603
R6294 two_stage_opamp_dummy_magic_14_0.cap_res_X.t21 two_stage_opamp_dummy_magic_14_0.cap_res_X.t58 0.1603
R6295 two_stage_opamp_dummy_magic_14_0.cap_res_X.t96 two_stage_opamp_dummy_magic_14_0.cap_res_X.t57 0.1603
R6296 two_stage_opamp_dummy_magic_14_0.cap_res_X.t63 two_stage_opamp_dummy_magic_14_0.cap_res_X.t96 0.1603
R6297 two_stage_opamp_dummy_magic_14_0.cap_res_X.t7 two_stage_opamp_dummy_magic_14_0.cap_res_X.t63 0.1603
R6298 two_stage_opamp_dummy_magic_14_0.cap_res_X.n28 two_stage_opamp_dummy_magic_14_0.cap_res_X.t126 0.159278
R6299 two_stage_opamp_dummy_magic_14_0.cap_res_X.n29 two_stage_opamp_dummy_magic_14_0.cap_res_X.t8 0.159278
R6300 two_stage_opamp_dummy_magic_14_0.cap_res_X.n30 two_stage_opamp_dummy_magic_14_0.cap_res_X.t107 0.159278
R6301 two_stage_opamp_dummy_magic_14_0.cap_res_X.n31 two_stage_opamp_dummy_magic_14_0.cap_res_X.t74 0.159278
R6302 two_stage_opamp_dummy_magic_14_0.cap_res_X.n32 two_stage_opamp_dummy_magic_14_0.cap_res_X.t37 0.159278
R6303 two_stage_opamp_dummy_magic_14_0.cap_res_X.n33 two_stage_opamp_dummy_magic_14_0.cap_res_X.t53 0.159278
R6304 two_stage_opamp_dummy_magic_14_0.cap_res_X.n25 two_stage_opamp_dummy_magic_14_0.cap_res_X.t103 0.159278
R6305 two_stage_opamp_dummy_magic_14_0.cap_res_X.n0 two_stage_opamp_dummy_magic_14_0.cap_res_X.t44 0.159278
R6306 two_stage_opamp_dummy_magic_14_0.cap_res_X.n1 two_stage_opamp_dummy_magic_14_0.cap_res_X.t133 0.159278
R6307 two_stage_opamp_dummy_magic_14_0.cap_res_X.n2 two_stage_opamp_dummy_magic_14_0.cap_res_X.t95 0.159278
R6308 two_stage_opamp_dummy_magic_14_0.cap_res_X.n3 two_stage_opamp_dummy_magic_14_0.cap_res_X.t62 0.159278
R6309 two_stage_opamp_dummy_magic_14_0.cap_res_X.n4 two_stage_opamp_dummy_magic_14_0.cap_res_X.t31 0.159278
R6310 two_stage_opamp_dummy_magic_14_0.cap_res_X.n5 two_stage_opamp_dummy_magic_14_0.cap_res_X.t119 0.159278
R6311 two_stage_opamp_dummy_magic_14_0.cap_res_X.n6 two_stage_opamp_dummy_magic_14_0.cap_res_X.t83 0.159278
R6312 two_stage_opamp_dummy_magic_14_0.cap_res_X.t67 two_stage_opamp_dummy_magic_14_0.cap_res_X.n9 0.159278
R6313 two_stage_opamp_dummy_magic_14_0.cap_res_X.t98 two_stage_opamp_dummy_magic_14_0.cap_res_X.n10 0.159278
R6314 two_stage_opamp_dummy_magic_14_0.cap_res_X.t59 two_stage_opamp_dummy_magic_14_0.cap_res_X.n11 0.159278
R6315 two_stage_opamp_dummy_magic_14_0.cap_res_X.t23 two_stage_opamp_dummy_magic_14_0.cap_res_X.n12 0.159278
R6316 two_stage_opamp_dummy_magic_14_0.cap_res_X.t55 two_stage_opamp_dummy_magic_14_0.cap_res_X.n13 0.159278
R6317 two_stage_opamp_dummy_magic_14_0.cap_res_X.t18 two_stage_opamp_dummy_magic_14_0.cap_res_X.n14 0.159278
R6318 two_stage_opamp_dummy_magic_14_0.cap_res_X.t117 two_stage_opamp_dummy_magic_14_0.cap_res_X.n15 0.159278
R6319 two_stage_opamp_dummy_magic_14_0.cap_res_X.t79 two_stage_opamp_dummy_magic_14_0.cap_res_X.n16 0.159278
R6320 two_stage_opamp_dummy_magic_14_0.cap_res_X.t109 two_stage_opamp_dummy_magic_14_0.cap_res_X.n17 0.159278
R6321 two_stage_opamp_dummy_magic_14_0.cap_res_X.t73 two_stage_opamp_dummy_magic_14_0.cap_res_X.n18 0.159278
R6322 two_stage_opamp_dummy_magic_14_0.cap_res_X.t36 two_stage_opamp_dummy_magic_14_0.cap_res_X.n19 0.159278
R6323 two_stage_opamp_dummy_magic_14_0.cap_res_X.t69 two_stage_opamp_dummy_magic_14_0.cap_res_X.n20 0.159278
R6324 two_stage_opamp_dummy_magic_14_0.cap_res_X.t29 two_stage_opamp_dummy_magic_14_0.cap_res_X.n21 0.159278
R6325 two_stage_opamp_dummy_magic_14_0.cap_res_X.t10 two_stage_opamp_dummy_magic_14_0.cap_res_X.n22 0.159278
R6326 two_stage_opamp_dummy_magic_14_0.cap_res_X.t45 two_stage_opamp_dummy_magic_14_0.cap_res_X.n23 0.159278
R6327 two_stage_opamp_dummy_magic_14_0.cap_res_X.t2 two_stage_opamp_dummy_magic_14_0.cap_res_X.n24 0.159278
R6328 two_stage_opamp_dummy_magic_14_0.cap_res_X.n26 two_stage_opamp_dummy_magic_14_0.cap_res_X.t1 0.159278
R6329 two_stage_opamp_dummy_magic_14_0.cap_res_X.n27 two_stage_opamp_dummy_magic_14_0.cap_res_X.t122 0.159278
R6330 two_stage_opamp_dummy_magic_14_0.cap_res_X.n34 two_stage_opamp_dummy_magic_14_0.cap_res_X.t20 0.159278
R6331 two_stage_opamp_dummy_magic_14_0.cap_res_X.t103 two_stage_opamp_dummy_magic_14_0.cap_res_X.t71 0.137822
R6332 two_stage_opamp_dummy_magic_14_0.cap_res_X.n25 two_stage_opamp_dummy_magic_14_0.cap_res_X.t105 0.1368
R6333 two_stage_opamp_dummy_magic_14_0.cap_res_X.n24 two_stage_opamp_dummy_magic_14_0.cap_res_X.t84 0.1368
R6334 two_stage_opamp_dummy_magic_14_0.cap_res_X.n24 two_stage_opamp_dummy_magic_14_0.cap_res_X.t5 0.1368
R6335 two_stage_opamp_dummy_magic_14_0.cap_res_X.n23 two_stage_opamp_dummy_magic_14_0.cap_res_X.t48 0.1368
R6336 two_stage_opamp_dummy_magic_14_0.cap_res_X.n23 two_stage_opamp_dummy_magic_14_0.cap_res_X.t110 0.1368
R6337 two_stage_opamp_dummy_magic_14_0.cap_res_X.n22 two_stage_opamp_dummy_magic_14_0.cap_res_X.t60 0.1368
R6338 two_stage_opamp_dummy_magic_14_0.cap_res_X.n22 two_stage_opamp_dummy_magic_14_0.cap_res_X.t130 0.1368
R6339 two_stage_opamp_dummy_magic_14_0.cap_res_X.n21 two_stage_opamp_dummy_magic_14_0.cap_res_X.t100 0.1368
R6340 two_stage_opamp_dummy_magic_14_0.cap_res_X.n21 two_stage_opamp_dummy_magic_14_0.cap_res_X.t34 0.1368
R6341 two_stage_opamp_dummy_magic_14_0.cap_res_X.n20 two_stage_opamp_dummy_magic_14_0.cap_res_X.t70 0.1368
R6342 two_stage_opamp_dummy_magic_14_0.cap_res_X.n20 two_stage_opamp_dummy_magic_14_0.cap_res_X.t137 0.1368
R6343 two_stage_opamp_dummy_magic_14_0.cap_res_X.n19 two_stage_opamp_dummy_magic_14_0.cap_res_X.t104 0.1368
R6344 two_stage_opamp_dummy_magic_14_0.cap_res_X.n19 two_stage_opamp_dummy_magic_14_0.cap_res_X.t39 0.1368
R6345 two_stage_opamp_dummy_magic_14_0.cap_res_X.n18 two_stage_opamp_dummy_magic_14_0.cap_res_X.t4 0.1368
R6346 two_stage_opamp_dummy_magic_14_0.cap_res_X.n18 two_stage_opamp_dummy_magic_14_0.cap_res_X.t78 0.1368
R6347 two_stage_opamp_dummy_magic_14_0.cap_res_X.n17 two_stage_opamp_dummy_magic_14_0.cap_res_X.t111 0.1368
R6348 two_stage_opamp_dummy_magic_14_0.cap_res_X.n17 two_stage_opamp_dummy_magic_14_0.cap_res_X.t40 0.1368
R6349 two_stage_opamp_dummy_magic_14_0.cap_res_X.n16 two_stage_opamp_dummy_magic_14_0.cap_res_X.t12 0.1368
R6350 two_stage_opamp_dummy_magic_14_0.cap_res_X.n16 two_stage_opamp_dummy_magic_14_0.cap_res_X.t82 0.1368
R6351 two_stage_opamp_dummy_magic_14_0.cap_res_X.n15 two_stage_opamp_dummy_magic_14_0.cap_res_X.t51 0.1368
R6352 two_stage_opamp_dummy_magic_14_0.cap_res_X.n15 two_stage_opamp_dummy_magic_14_0.cap_res_X.t123 0.1368
R6353 two_stage_opamp_dummy_magic_14_0.cap_res_X.n14 two_stage_opamp_dummy_magic_14_0.cap_res_X.t90 0.1368
R6354 two_stage_opamp_dummy_magic_14_0.cap_res_X.n14 two_stage_opamp_dummy_magic_14_0.cap_res_X.t22 0.1368
R6355 two_stage_opamp_dummy_magic_14_0.cap_res_X.n13 two_stage_opamp_dummy_magic_14_0.cap_res_X.t54 0.1368
R6356 two_stage_opamp_dummy_magic_14_0.cap_res_X.n13 two_stage_opamp_dummy_magic_14_0.cap_res_X.t127 0.1368
R6357 two_stage_opamp_dummy_magic_14_0.cap_res_X.n12 two_stage_opamp_dummy_magic_14_0.cap_res_X.t94 0.1368
R6358 two_stage_opamp_dummy_magic_14_0.cap_res_X.n12 two_stage_opamp_dummy_magic_14_0.cap_res_X.t28 0.1368
R6359 two_stage_opamp_dummy_magic_14_0.cap_res_X.n11 two_stage_opamp_dummy_magic_14_0.cap_res_X.t136 0.1368
R6360 two_stage_opamp_dummy_magic_14_0.cap_res_X.n11 two_stage_opamp_dummy_magic_14_0.cap_res_X.t68 0.1368
R6361 two_stage_opamp_dummy_magic_14_0.cap_res_X.n10 two_stage_opamp_dummy_magic_14_0.cap_res_X.t35 0.1368
R6362 two_stage_opamp_dummy_magic_14_0.cap_res_X.n9 two_stage_opamp_dummy_magic_14_0.cap_res_X.t38 0.1368
R6363 two_stage_opamp_dummy_magic_14_0.cap_res_X.n29 two_stage_opamp_dummy_magic_14_0.cap_res_X.n28 0.1133
R6364 two_stage_opamp_dummy_magic_14_0.cap_res_X.n30 two_stage_opamp_dummy_magic_14_0.cap_res_X.n29 0.1133
R6365 two_stage_opamp_dummy_magic_14_0.cap_res_X.n31 two_stage_opamp_dummy_magic_14_0.cap_res_X.n30 0.1133
R6366 two_stage_opamp_dummy_magic_14_0.cap_res_X.n32 two_stage_opamp_dummy_magic_14_0.cap_res_X.n31 0.1133
R6367 two_stage_opamp_dummy_magic_14_0.cap_res_X.n33 two_stage_opamp_dummy_magic_14_0.cap_res_X.n32 0.1133
R6368 two_stage_opamp_dummy_magic_14_0.cap_res_X.n1 two_stage_opamp_dummy_magic_14_0.cap_res_X.n0 0.1133
R6369 two_stage_opamp_dummy_magic_14_0.cap_res_X.n2 two_stage_opamp_dummy_magic_14_0.cap_res_X.n1 0.1133
R6370 two_stage_opamp_dummy_magic_14_0.cap_res_X.n3 two_stage_opamp_dummy_magic_14_0.cap_res_X.n2 0.1133
R6371 two_stage_opamp_dummy_magic_14_0.cap_res_X.n4 two_stage_opamp_dummy_magic_14_0.cap_res_X.n3 0.1133
R6372 two_stage_opamp_dummy_magic_14_0.cap_res_X.n5 two_stage_opamp_dummy_magic_14_0.cap_res_X.n4 0.1133
R6373 two_stage_opamp_dummy_magic_14_0.cap_res_X.n6 two_stage_opamp_dummy_magic_14_0.cap_res_X.n5 0.1133
R6374 two_stage_opamp_dummy_magic_14_0.cap_res_X.n7 two_stage_opamp_dummy_magic_14_0.cap_res_X.n6 0.1133
R6375 two_stage_opamp_dummy_magic_14_0.cap_res_X.n8 two_stage_opamp_dummy_magic_14_0.cap_res_X.n7 0.1133
R6376 two_stage_opamp_dummy_magic_14_0.cap_res_X.n10 two_stage_opamp_dummy_magic_14_0.cap_res_X.n8 0.1133
R6377 two_stage_opamp_dummy_magic_14_0.cap_res_X.n26 two_stage_opamp_dummy_magic_14_0.cap_res_X.n25 0.1133
R6378 two_stage_opamp_dummy_magic_14_0.cap_res_X.n27 two_stage_opamp_dummy_magic_14_0.cap_res_X.n26 0.1133
R6379 two_stage_opamp_dummy_magic_14_0.cap_res_X.n34 two_stage_opamp_dummy_magic_14_0.cap_res_X.n27 0.1133
R6380 two_stage_opamp_dummy_magic_14_0.cap_res_X.n34 two_stage_opamp_dummy_magic_14_0.cap_res_X.n33 0.1133
R6381 two_stage_opamp_dummy_magic_14_0.cap_res_X.n28 two_stage_opamp_dummy_magic_14_0.cap_res_X.t27 0.00152174
R6382 two_stage_opamp_dummy_magic_14_0.cap_res_X.n29 two_stage_opamp_dummy_magic_14_0.cap_res_X.t49 0.00152174
R6383 two_stage_opamp_dummy_magic_14_0.cap_res_X.n30 two_stage_opamp_dummy_magic_14_0.cap_res_X.t11 0.00152174
R6384 two_stage_opamp_dummy_magic_14_0.cap_res_X.n31 two_stage_opamp_dummy_magic_14_0.cap_res_X.t112 0.00152174
R6385 two_stage_opamp_dummy_magic_14_0.cap_res_X.n32 two_stage_opamp_dummy_magic_14_0.cap_res_X.t76 0.00152174
R6386 two_stage_opamp_dummy_magic_14_0.cap_res_X.n33 two_stage_opamp_dummy_magic_14_0.cap_res_X.t93 0.00152174
R6387 two_stage_opamp_dummy_magic_14_0.cap_res_X.n0 two_stage_opamp_dummy_magic_14_0.cap_res_X.t9 0.00152174
R6388 two_stage_opamp_dummy_magic_14_0.cap_res_X.n1 two_stage_opamp_dummy_magic_14_0.cap_res_X.t97 0.00152174
R6389 two_stage_opamp_dummy_magic_14_0.cap_res_X.n2 two_stage_opamp_dummy_magic_14_0.cap_res_X.t64 0.00152174
R6390 two_stage_opamp_dummy_magic_14_0.cap_res_X.n3 two_stage_opamp_dummy_magic_14_0.cap_res_X.t30 0.00152174
R6391 two_stage_opamp_dummy_magic_14_0.cap_res_X.n4 two_stage_opamp_dummy_magic_14_0.cap_res_X.t132 0.00152174
R6392 two_stage_opamp_dummy_magic_14_0.cap_res_X.n5 two_stage_opamp_dummy_magic_14_0.cap_res_X.t85 0.00152174
R6393 two_stage_opamp_dummy_magic_14_0.cap_res_X.n6 two_stage_opamp_dummy_magic_14_0.cap_res_X.t47 0.00152174
R6394 two_stage_opamp_dummy_magic_14_0.cap_res_X.n7 two_stage_opamp_dummy_magic_14_0.cap_res_X.t15 0.00152174
R6395 two_stage_opamp_dummy_magic_14_0.cap_res_X.n8 two_stage_opamp_dummy_magic_14_0.cap_res_X.t101 0.00152174
R6396 two_stage_opamp_dummy_magic_14_0.cap_res_X.n9 two_stage_opamp_dummy_magic_14_0.cap_res_X.t124 0.00152174
R6397 two_stage_opamp_dummy_magic_14_0.cap_res_X.n10 two_stage_opamp_dummy_magic_14_0.cap_res_X.t67 0.00152174
R6398 two_stage_opamp_dummy_magic_14_0.cap_res_X.n11 two_stage_opamp_dummy_magic_14_0.cap_res_X.t98 0.00152174
R6399 two_stage_opamp_dummy_magic_14_0.cap_res_X.n12 two_stage_opamp_dummy_magic_14_0.cap_res_X.t59 0.00152174
R6400 two_stage_opamp_dummy_magic_14_0.cap_res_X.n13 two_stage_opamp_dummy_magic_14_0.cap_res_X.t23 0.00152174
R6401 two_stage_opamp_dummy_magic_14_0.cap_res_X.n14 two_stage_opamp_dummy_magic_14_0.cap_res_X.t55 0.00152174
R6402 two_stage_opamp_dummy_magic_14_0.cap_res_X.n15 two_stage_opamp_dummy_magic_14_0.cap_res_X.t18 0.00152174
R6403 two_stage_opamp_dummy_magic_14_0.cap_res_X.n16 two_stage_opamp_dummy_magic_14_0.cap_res_X.t117 0.00152174
R6404 two_stage_opamp_dummy_magic_14_0.cap_res_X.n17 two_stage_opamp_dummy_magic_14_0.cap_res_X.t79 0.00152174
R6405 two_stage_opamp_dummy_magic_14_0.cap_res_X.n18 two_stage_opamp_dummy_magic_14_0.cap_res_X.t109 0.00152174
R6406 two_stage_opamp_dummy_magic_14_0.cap_res_X.n19 two_stage_opamp_dummy_magic_14_0.cap_res_X.t73 0.00152174
R6407 two_stage_opamp_dummy_magic_14_0.cap_res_X.n20 two_stage_opamp_dummy_magic_14_0.cap_res_X.t36 0.00152174
R6408 two_stage_opamp_dummy_magic_14_0.cap_res_X.n21 two_stage_opamp_dummy_magic_14_0.cap_res_X.t69 0.00152174
R6409 two_stage_opamp_dummy_magic_14_0.cap_res_X.n22 two_stage_opamp_dummy_magic_14_0.cap_res_X.t29 0.00152174
R6410 two_stage_opamp_dummy_magic_14_0.cap_res_X.n23 two_stage_opamp_dummy_magic_14_0.cap_res_X.t10 0.00152174
R6411 two_stage_opamp_dummy_magic_14_0.cap_res_X.n24 two_stage_opamp_dummy_magic_14_0.cap_res_X.t45 0.00152174
R6412 two_stage_opamp_dummy_magic_14_0.cap_res_X.n25 two_stage_opamp_dummy_magic_14_0.cap_res_X.t2 0.00152174
R6413 two_stage_opamp_dummy_magic_14_0.cap_res_X.n26 two_stage_opamp_dummy_magic_14_0.cap_res_X.t41 0.00152174
R6414 two_stage_opamp_dummy_magic_14_0.cap_res_X.n27 two_stage_opamp_dummy_magic_14_0.cap_res_X.t21 0.00152174
R6415 two_stage_opamp_dummy_magic_14_0.cap_res_X.t57 two_stage_opamp_dummy_magic_14_0.cap_res_X.n34 0.00152174
R6416 VOUT+.n8 VOUT+.n6 149.19
R6417 VOUT+.n14 VOUT+.n13 149.19
R6418 VOUT+.n12 VOUT+.n11 148.626
R6419 VOUT+.n10 VOUT+.n9 148.626
R6420 VOUT+.n8 VOUT+.n7 148.626
R6421 VOUT+.n16 VOUT+.n15 144.126
R6422 VOUT+.n5 VOUT+.t0 112.184
R6423 VOUT+.n2 VOUT+.n0 98.9303
R6424 VOUT+.n4 VOUT+.n3 97.8053
R6425 VOUT+.n2 VOUT+.n1 97.8053
R6426 VOUT+.n91 VOUT+.n16 15.5682
R6427 VOUT+.n91 VOUT+.n90 11.5649
R6428 VOUT+ VOUT+.n91 9.2505
R6429 VOUT+.n15 VOUT+.t17 6.56717
R6430 VOUT+.n15 VOUT+.t9 6.56717
R6431 VOUT+.n13 VOUT+.t10 6.56717
R6432 VOUT+.n13 VOUT+.t16 6.56717
R6433 VOUT+.n11 VOUT+.t12 6.56717
R6434 VOUT+.n11 VOUT+.t1 6.56717
R6435 VOUT+.n9 VOUT+.t8 6.56717
R6436 VOUT+.n9 VOUT+.t4 6.56717
R6437 VOUT+.n7 VOUT+.t7 6.56717
R6438 VOUT+.n7 VOUT+.t5 6.56717
R6439 VOUT+.n6 VOUT+.t15 6.56717
R6440 VOUT+.n6 VOUT+.t6 6.56717
R6441 VOUT+.n45 VOUT+.t56 4.8295
R6442 VOUT+.n47 VOUT+.t105 4.8295
R6443 VOUT+.n48 VOUT+.t29 4.8295
R6444 VOUT+.n50 VOUT+.t60 4.8295
R6445 VOUT+.n52 VOUT+.t115 4.8295
R6446 VOUT+.n63 VOUT+.t20 4.8295
R6447 VOUT+.n66 VOUT+.t31 4.8295
R6448 VOUT+.n65 VOUT+.t121 4.8295
R6449 VOUT+.n68 VOUT+.t67 4.8295
R6450 VOUT+.n67 VOUT+.t152 4.8295
R6451 VOUT+.n69 VOUT+.t131 4.8295
R6452 VOUT+.n70 VOUT+.t118 4.8295
R6453 VOUT+.n72 VOUT+.t89 4.8295
R6454 VOUT+.n73 VOUT+.t76 4.8295
R6455 VOUT+.n75 VOUT+.t127 4.8295
R6456 VOUT+.n76 VOUT+.t110 4.8295
R6457 VOUT+.n78 VOUT+.t84 4.8295
R6458 VOUT+.n79 VOUT+.t68 4.8295
R6459 VOUT+.n81 VOUT+.t42 4.8295
R6460 VOUT+.n82 VOUT+.t30 4.8295
R6461 VOUT+.n84 VOUT+.t81 4.8295
R6462 VOUT+.n85 VOUT+.t64 4.8295
R6463 VOUT+.n17 VOUT+.t150 4.8295
R6464 VOUT+.n28 VOUT+.t75 4.8295
R6465 VOUT+.n30 VOUT+.t54 4.8295
R6466 VOUT+.n31 VOUT+.t34 4.8295
R6467 VOUT+.n33 VOUT+.t95 4.8295
R6468 VOUT+.n34 VOUT+.t79 4.8295
R6469 VOUT+.n36 VOUT+.t134 4.8295
R6470 VOUT+.n37 VOUT+.t122 4.8295
R6471 VOUT+.n39 VOUT+.t102 4.8295
R6472 VOUT+.n40 VOUT+.t82 4.8295
R6473 VOUT+.n42 VOUT+.t137 4.8295
R6474 VOUT+.n43 VOUT+.t126 4.8295
R6475 VOUT+.n87 VOUT+.t28 4.8295
R6476 VOUT+.n56 VOUT+.t57 4.8154
R6477 VOUT+.n55 VOUT+.t33 4.8154
R6478 VOUT+.n54 VOUT+.t77 4.8154
R6479 VOUT+.n62 VOUT+.t116 4.806
R6480 VOUT+.n61 VOUT+.t147 4.806
R6481 VOUT+.n60 VOUT+.t43 4.806
R6482 VOUT+.n59 VOUT+.t83 4.806
R6483 VOUT+.n58 VOUT+.t63 4.806
R6484 VOUT+.n57 VOUT+.t26 4.806
R6485 VOUT+.n57 VOUT+.t103 4.806
R6486 VOUT+.n56 VOUT+.t135 4.806
R6487 VOUT+.n55 VOUT+.t120 4.806
R6488 VOUT+.n54 VOUT+.t155 4.806
R6489 VOUT+.n27 VOUT+.t91 4.806
R6490 VOUT+.n26 VOUT+.t38 4.806
R6491 VOUT+.n25 VOUT+.t130 4.806
R6492 VOUT+.n25 VOUT+.t90 4.806
R6493 VOUT+.n24 VOUT+.t80 4.806
R6494 VOUT+.n24 VOUT+.t128 4.806
R6495 VOUT+.n23 VOUT+.t124 4.806
R6496 VOUT+.n23 VOUT+.t32 4.806
R6497 VOUT+.n22 VOUT+.t70 4.806
R6498 VOUT+.n22 VOUT+.t73 4.806
R6499 VOUT+.n21 VOUT+.t23 4.806
R6500 VOUT+.n21 VOUT+.t108 4.806
R6501 VOUT+.n20 VOUT+.t62 4.806
R6502 VOUT+.n20 VOUT+.t19 4.806
R6503 VOUT+.n19 VOUT+.t151 4.806
R6504 VOUT+.n19 VOUT+.t49 4.806
R6505 VOUT+.n46 VOUT+.t132 4.5005
R6506 VOUT+.n45 VOUT+.t96 4.5005
R6507 VOUT+.n47 VOUT+.t69 4.5005
R6508 VOUT+.n48 VOUT+.t139 4.5005
R6509 VOUT+.n49 VOUT+.t109 4.5005
R6510 VOUT+.n50 VOUT+.t37 4.5005
R6511 VOUT+.n51 VOUT+.t144 4.5005
R6512 VOUT+.n52 VOUT+.t21 4.5005
R6513 VOUT+.n53 VOUT+.t125 4.5005
R6514 VOUT+.n54 VOUT+.t119 4.5005
R6515 VOUT+.n55 VOUT+.t78 4.5005
R6516 VOUT+.n56 VOUT+.t97 4.5005
R6517 VOUT+.n57 VOUT+.t61 4.5005
R6518 VOUT+.n58 VOUT+.t27 4.5005
R6519 VOUT+.n59 VOUT+.t41 4.5005
R6520 VOUT+.n60 VOUT+.t145 4.5005
R6521 VOUT+.n61 VOUT+.t113 4.5005
R6522 VOUT+.n62 VOUT+.t72 4.5005
R6523 VOUT+.n64 VOUT+.t92 4.5005
R6524 VOUT+.n63 VOUT+.t55 4.5005
R6525 VOUT+.n66 VOUT+.t50 4.5005
R6526 VOUT+.n65 VOUT+.t156 4.5005
R6527 VOUT+.n68 VOUT+.t86 4.5005
R6528 VOUT+.n67 VOUT+.t47 4.5005
R6529 VOUT+.n69 VOUT+.t94 4.5005
R6530 VOUT+.n71 VOUT+.t39 4.5005
R6531 VOUT+.n70 VOUT+.t146 4.5005
R6532 VOUT+.n72 VOUT+.t53 4.5005
R6533 VOUT+.n74 VOUT+.t142 4.5005
R6534 VOUT+.n73 VOUT+.t112 4.5005
R6535 VOUT+.n75 VOUT+.t88 4.5005
R6536 VOUT+.n77 VOUT+.t35 4.5005
R6537 VOUT+.n76 VOUT+.t140 4.5005
R6538 VOUT+.n78 VOUT+.t46 4.5005
R6539 VOUT+.n80 VOUT+.t136 4.5005
R6540 VOUT+.n79 VOUT+.t104 4.5005
R6541 VOUT+.n81 VOUT+.t149 4.5005
R6542 VOUT+.n83 VOUT+.t99 4.5005
R6543 VOUT+.n82 VOUT+.t65 4.5005
R6544 VOUT+.n84 VOUT+.t40 4.5005
R6545 VOUT+.n86 VOUT+.t133 4.5005
R6546 VOUT+.n85 VOUT+.t98 4.5005
R6547 VOUT+.n18 VOUT+.t45 4.5005
R6548 VOUT+.n17 VOUT+.t101 4.5005
R6549 VOUT+.n19 VOUT+.t85 4.5005
R6550 VOUT+.n20 VOUT+.t48 4.5005
R6551 VOUT+.n21 VOUT+.t138 4.5005
R6552 VOUT+.n22 VOUT+.t107 4.5005
R6553 VOUT+.n23 VOUT+.t71 4.5005
R6554 VOUT+.n24 VOUT+.t25 4.5005
R6555 VOUT+.n25 VOUT+.t129 4.5005
R6556 VOUT+.n26 VOUT+.t87 4.5005
R6557 VOUT+.n27 VOUT+.t52 4.5005
R6558 VOUT+.n29 VOUT+.t141 4.5005
R6559 VOUT+.n28 VOUT+.t111 4.5005
R6560 VOUT+.n30 VOUT+.t24 4.5005
R6561 VOUT+.n32 VOUT+.t114 4.5005
R6562 VOUT+.n31 VOUT+.t74 4.5005
R6563 VOUT+.n33 VOUT+.t59 4.5005
R6564 VOUT+.n35 VOUT+.t148 4.5005
R6565 VOUT+.n34 VOUT+.t117 4.5005
R6566 VOUT+.n36 VOUT+.t100 4.5005
R6567 VOUT+.n38 VOUT+.t44 4.5005
R6568 VOUT+.n37 VOUT+.t153 4.5005
R6569 VOUT+.n39 VOUT+.t66 4.5005
R6570 VOUT+.n41 VOUT+.t154 4.5005
R6571 VOUT+.n40 VOUT+.t123 4.5005
R6572 VOUT+.n42 VOUT+.t106 4.5005
R6573 VOUT+.n44 VOUT+.t51 4.5005
R6574 VOUT+.n43 VOUT+.t22 4.5005
R6575 VOUT+.n90 VOUT+.t36 4.5005
R6576 VOUT+.n89 VOUT+.t143 4.5005
R6577 VOUT+.n88 VOUT+.t93 4.5005
R6578 VOUT+.n87 VOUT+.t58 4.5005
R6579 VOUT+.n16 VOUT+.n14 4.5005
R6580 VOUT+.n3 VOUT+.t11 3.42907
R6581 VOUT+.n3 VOUT+.t13 3.42907
R6582 VOUT+.n1 VOUT+.t18 3.42907
R6583 VOUT+.n1 VOUT+.t3 3.42907
R6584 VOUT+.n0 VOUT+.t14 3.42907
R6585 VOUT+.n0 VOUT+.t2 3.42907
R6586 VOUT+ VOUT+.n5 1.46144
R6587 VOUT+.n5 VOUT+.n4 1.30519
R6588 VOUT+.n4 VOUT+.n2 1.1255
R6589 VOUT+.n10 VOUT+.n8 0.563
R6590 VOUT+.n12 VOUT+.n10 0.563
R6591 VOUT+.n14 VOUT+.n12 0.563
R6592 VOUT+.n46 VOUT+.n45 0.3295
R6593 VOUT+.n49 VOUT+.n48 0.3295
R6594 VOUT+.n51 VOUT+.n50 0.3295
R6595 VOUT+.n53 VOUT+.n52 0.3295
R6596 VOUT+.n55 VOUT+.n54 0.3295
R6597 VOUT+.n56 VOUT+.n55 0.3295
R6598 VOUT+.n57 VOUT+.n56 0.3295
R6599 VOUT+.n58 VOUT+.n57 0.3295
R6600 VOUT+.n59 VOUT+.n58 0.3295
R6601 VOUT+.n60 VOUT+.n59 0.3295
R6602 VOUT+.n61 VOUT+.n60 0.3295
R6603 VOUT+.n62 VOUT+.n61 0.3295
R6604 VOUT+.n64 VOUT+.n62 0.3295
R6605 VOUT+.n64 VOUT+.n63 0.3295
R6606 VOUT+.n66 VOUT+.n65 0.3295
R6607 VOUT+.n68 VOUT+.n67 0.3295
R6608 VOUT+.n71 VOUT+.n69 0.3295
R6609 VOUT+.n71 VOUT+.n70 0.3295
R6610 VOUT+.n74 VOUT+.n72 0.3295
R6611 VOUT+.n74 VOUT+.n73 0.3295
R6612 VOUT+.n77 VOUT+.n75 0.3295
R6613 VOUT+.n77 VOUT+.n76 0.3295
R6614 VOUT+.n80 VOUT+.n78 0.3295
R6615 VOUT+.n80 VOUT+.n79 0.3295
R6616 VOUT+.n83 VOUT+.n81 0.3295
R6617 VOUT+.n83 VOUT+.n82 0.3295
R6618 VOUT+.n86 VOUT+.n84 0.3295
R6619 VOUT+.n86 VOUT+.n85 0.3295
R6620 VOUT+.n18 VOUT+.n17 0.3295
R6621 VOUT+.n20 VOUT+.n19 0.3295
R6622 VOUT+.n21 VOUT+.n20 0.3295
R6623 VOUT+.n22 VOUT+.n21 0.3295
R6624 VOUT+.n23 VOUT+.n22 0.3295
R6625 VOUT+.n24 VOUT+.n23 0.3295
R6626 VOUT+.n25 VOUT+.n24 0.3295
R6627 VOUT+.n26 VOUT+.n25 0.3295
R6628 VOUT+.n27 VOUT+.n26 0.3295
R6629 VOUT+.n29 VOUT+.n27 0.3295
R6630 VOUT+.n29 VOUT+.n28 0.3295
R6631 VOUT+.n32 VOUT+.n30 0.3295
R6632 VOUT+.n32 VOUT+.n31 0.3295
R6633 VOUT+.n35 VOUT+.n33 0.3295
R6634 VOUT+.n35 VOUT+.n34 0.3295
R6635 VOUT+.n38 VOUT+.n36 0.3295
R6636 VOUT+.n38 VOUT+.n37 0.3295
R6637 VOUT+.n41 VOUT+.n39 0.3295
R6638 VOUT+.n41 VOUT+.n40 0.3295
R6639 VOUT+.n44 VOUT+.n42 0.3295
R6640 VOUT+.n44 VOUT+.n43 0.3295
R6641 VOUT+.n90 VOUT+.n89 0.3295
R6642 VOUT+.n89 VOUT+.n88 0.3295
R6643 VOUT+.n88 VOUT+.n87 0.3295
R6644 VOUT+.n61 VOUT+.n47 0.306
R6645 VOUT+.n60 VOUT+.n49 0.306
R6646 VOUT+.n59 VOUT+.n51 0.306
R6647 VOUT+.n58 VOUT+.n53 0.306
R6648 VOUT+.n64 VOUT+.n46 0.2825
R6649 VOUT+.n66 VOUT+.n64 0.2825
R6650 VOUT+.n68 VOUT+.n66 0.2825
R6651 VOUT+.n71 VOUT+.n68 0.2825
R6652 VOUT+.n74 VOUT+.n71 0.2825
R6653 VOUT+.n77 VOUT+.n74 0.2825
R6654 VOUT+.n80 VOUT+.n77 0.2825
R6655 VOUT+.n83 VOUT+.n80 0.2825
R6656 VOUT+.n86 VOUT+.n83 0.2825
R6657 VOUT+.n29 VOUT+.n18 0.2825
R6658 VOUT+.n32 VOUT+.n29 0.2825
R6659 VOUT+.n35 VOUT+.n32 0.2825
R6660 VOUT+.n38 VOUT+.n35 0.2825
R6661 VOUT+.n41 VOUT+.n38 0.2825
R6662 VOUT+.n44 VOUT+.n41 0.2825
R6663 VOUT+.n88 VOUT+.n44 0.2825
R6664 VOUT+.n88 VOUT+.n86 0.2825
R6665 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t0 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t128 50.3211
R6666 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t102 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t137 0.1603
R6667 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t61 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t101 0.1603
R6668 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t1 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t36 0.1603
R6669 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t110 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t5 0.1603
R6670 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t11 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t39 0.1603
R6671 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t63 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t26 0.1603
R6672 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t45 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t81 0.1603
R6673 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t104 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t68 0.1603
R6674 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t17 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t47 0.1603
R6675 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t69 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t30 0.1603
R6676 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t53 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t89 0.1603
R6677 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t111 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t73 0.1603
R6678 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t92 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t127 0.1603
R6679 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t8 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t115 0.1603
R6680 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t59 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t93 0.1603
R6681 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t117 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t76 0.1603
R6682 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t99 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t129 0.1603
R6683 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t14 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t121 0.1603
R6684 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t135 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t31 0.1603
R6685 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t51 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t20 0.1603
R6686 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t34 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t75 0.1603
R6687 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t91 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t55 0.1603
R6688 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t4 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t35 0.1603
R6689 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t57 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t23 0.1603
R6690 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t40 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t78 0.1603
R6691 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t98 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t62 0.1603
R6692 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t83 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t123 0.1603
R6693 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t133 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t103 0.1603
R6694 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t46 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t82 0.1603
R6695 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t72 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t6 0.1603
R6696 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t109 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t95 0.1603
R6697 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t19 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t134 0.1603
R6698 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t50 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t87 0.1603
R6699 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t86 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t33 0.1603
R6700 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t132 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t77 0.1603
R6701 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t28 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t27 0.1603
R6702 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t70 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t119 0.1603
R6703 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t105 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t66 0.1603
R6704 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t56 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t7 0.1603
R6705 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t88 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t52 0.1603
R6706 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t44 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t88 0.1603
R6707 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t38 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t80 0.1603
R6708 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t79 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t124 0.1603
R6709 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t60 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t100 0.1603
R6710 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t96 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t131 0.1603
R6711 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t136 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t42 0.1603
R6712 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t32 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t136 0.1603
R6713 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t130 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t32 0.1603
R6714 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t120 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t97 0.1603
R6715 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t13 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t120 0.1603
R6716 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t116 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t13 0.1603
R6717 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t48 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t12 0.1603
R6718 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t18 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t48 0.1603
R6719 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t128 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t18 0.1603
R6720 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n31 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t25 0.159278
R6721 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n6 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t108 0.159278
R6722 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n7 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t138 0.159278
R6723 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n8 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t49 0.159278
R6724 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n9 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t84 0.159278
R6725 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n10 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t125 0.159278
R6726 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n11 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t29 0.159278
R6727 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n12 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t67 0.159278
R6728 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t16 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n15 0.159278
R6729 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t43 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n16 0.159278
R6730 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t9 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n17 0.159278
R6731 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t113 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n18 0.159278
R6732 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t3 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n19 0.159278
R6733 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t106 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n20 0.159278
R6734 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t64 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n21 0.159278
R6735 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t24 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n22 0.159278
R6736 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t58 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n23 0.159278
R6737 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t21 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n24 0.159278
R6738 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t122 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n25 0.159278
R6739 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t15 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n26 0.159278
R6740 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t118 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n27 0.159278
R6741 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t71 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n28 0.159278
R6742 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t107 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n29 0.159278
R6743 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t65 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n30 0.159278
R6744 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n32 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t41 0.159278
R6745 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n33 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t10 0.159278
R6746 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n0 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t2 0.159278
R6747 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n1 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t37 0.159278
R6748 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n2 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t22 0.159278
R6749 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n3 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t54 0.159278
R6750 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n4 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t94 0.159278
R6751 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n5 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t74 0.159278
R6752 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n34 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t114 0.159278
R6753 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t25 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t61 0.137822
R6754 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n31 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t102 0.1368
R6755 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n30 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t1 0.1368
R6756 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n30 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t126 0.1368
R6757 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n29 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t110 0.1368
R6758 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n29 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t90 0.1368
R6759 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n28 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t11 0.1368
R6760 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n28 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t63 0.1368
R6761 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n27 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t45 0.1368
R6762 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n27 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t104 0.1368
R6763 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n26 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t17 0.1368
R6764 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n26 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t69 0.1368
R6765 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n25 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t53 0.1368
R6766 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n25 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t111 0.1368
R6767 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n24 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t92 0.1368
R6768 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n24 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t8 0.1368
R6769 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n23 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t59 0.1368
R6770 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n23 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t117 0.1368
R6771 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n22 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t99 0.1368
R6772 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n22 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t14 0.1368
R6773 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n21 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t135 0.1368
R6774 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n21 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t51 0.1368
R6775 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n20 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t34 0.1368
R6776 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n20 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t91 0.1368
R6777 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n19 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t4 0.1368
R6778 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n19 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t57 0.1368
R6779 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n18 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t40 0.1368
R6780 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n18 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t98 0.1368
R6781 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n17 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t83 0.1368
R6782 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n17 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t133 0.1368
R6783 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n16 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t46 0.1368
R6784 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n15 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t56 0.1368
R6785 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n7 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n6 0.1133
R6786 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n8 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n7 0.1133
R6787 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n9 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n8 0.1133
R6788 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n10 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n9 0.1133
R6789 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n11 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n10 0.1133
R6790 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n12 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n11 0.1133
R6791 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n13 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n12 0.1133
R6792 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n14 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n13 0.1133
R6793 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n16 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n14 0.1133
R6794 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n32 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n31 0.1133
R6795 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n33 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n32 0.1133
R6796 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n1 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n0 0.1133
R6797 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n2 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n1 0.1133
R6798 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n3 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n2 0.1133
R6799 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n4 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n3 0.1133
R6800 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n5 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n4 0.1133
R6801 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n34 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n5 0.1133
R6802 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n34 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n33 0.1133
R6803 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n6 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t72 0.00152174
R6804 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n7 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t109 0.00152174
R6805 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n8 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t19 0.00152174
R6806 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n9 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t50 0.00152174
R6807 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n10 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t86 0.00152174
R6808 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n11 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t132 0.00152174
R6809 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n12 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t28 0.00152174
R6810 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n13 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t70 0.00152174
R6811 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n14 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t105 0.00152174
R6812 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n15 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t112 0.00152174
R6813 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n16 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t16 0.00152174
R6814 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n17 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t43 0.00152174
R6815 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n18 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t9 0.00152174
R6816 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n19 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t113 0.00152174
R6817 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n20 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t3 0.00152174
R6818 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n21 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t106 0.00152174
R6819 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n22 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t64 0.00152174
R6820 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n23 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t24 0.00152174
R6821 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n24 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t58 0.00152174
R6822 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n25 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t21 0.00152174
R6823 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n26 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t122 0.00152174
R6824 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n27 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t15 0.00152174
R6825 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n28 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t118 0.00152174
R6826 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n29 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t71 0.00152174
R6827 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n30 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t107 0.00152174
R6828 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n31 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t65 0.00152174
R6829 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n32 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t85 0.00152174
R6830 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n33 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t44 0.00152174
R6831 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n0 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t38 0.00152174
R6832 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n1 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t79 0.00152174
R6833 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n2 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t60 0.00152174
R6834 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n3 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t96 0.00152174
R6835 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n4 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t130 0.00152174
R6836 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n5 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t116 0.00152174
R6837 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t12 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n34 0.00152174
R6838 two_stage_opamp_dummy_magic_14_0.X.n47 two_stage_opamp_dummy_magic_14_0.X.t51 1172.87
R6839 two_stage_opamp_dummy_magic_14_0.X.n43 two_stage_opamp_dummy_magic_14_0.X.t27 1172.87
R6840 two_stage_opamp_dummy_magic_14_0.X.n50 two_stage_opamp_dummy_magic_14_0.X.t48 996.134
R6841 two_stage_opamp_dummy_magic_14_0.X.n49 two_stage_opamp_dummy_magic_14_0.X.t35 996.134
R6842 two_stage_opamp_dummy_magic_14_0.X.n48 two_stage_opamp_dummy_magic_14_0.X.t42 996.134
R6843 two_stage_opamp_dummy_magic_14_0.X.n47 two_stage_opamp_dummy_magic_14_0.X.t34 996.134
R6844 two_stage_opamp_dummy_magic_14_0.X.n43 two_stage_opamp_dummy_magic_14_0.X.t43 996.134
R6845 two_stage_opamp_dummy_magic_14_0.X.n44 two_stage_opamp_dummy_magic_14_0.X.t29 996.134
R6846 two_stage_opamp_dummy_magic_14_0.X.n45 two_stage_opamp_dummy_magic_14_0.X.t45 996.134
R6847 two_stage_opamp_dummy_magic_14_0.X.n46 two_stage_opamp_dummy_magic_14_0.X.t31 996.134
R6848 two_stage_opamp_dummy_magic_14_0.X.n25 two_stage_opamp_dummy_magic_14_0.X.t26 690.867
R6849 two_stage_opamp_dummy_magic_14_0.X.n20 two_stage_opamp_dummy_magic_14_0.X.t32 690.867
R6850 two_stage_opamp_dummy_magic_14_0.X.n16 two_stage_opamp_dummy_magic_14_0.X.t39 530.201
R6851 two_stage_opamp_dummy_magic_14_0.X.n11 two_stage_opamp_dummy_magic_14_0.X.t44 530.201
R6852 two_stage_opamp_dummy_magic_14_0.X.n25 two_stage_opamp_dummy_magic_14_0.X.t40 514.134
R6853 two_stage_opamp_dummy_magic_14_0.X.n26 two_stage_opamp_dummy_magic_14_0.X.t46 514.134
R6854 two_stage_opamp_dummy_magic_14_0.X.n27 two_stage_opamp_dummy_magic_14_0.X.t41 514.134
R6855 two_stage_opamp_dummy_magic_14_0.X.n24 two_stage_opamp_dummy_magic_14_0.X.t25 514.134
R6856 two_stage_opamp_dummy_magic_14_0.X.n23 two_stage_opamp_dummy_magic_14_0.X.t38 514.134
R6857 two_stage_opamp_dummy_magic_14_0.X.n22 two_stage_opamp_dummy_magic_14_0.X.t52 514.134
R6858 two_stage_opamp_dummy_magic_14_0.X.n21 two_stage_opamp_dummy_magic_14_0.X.t36 514.134
R6859 two_stage_opamp_dummy_magic_14_0.X.n20 two_stage_opamp_dummy_magic_14_0.X.t49 514.134
R6860 two_stage_opamp_dummy_magic_14_0.X.n18 two_stage_opamp_dummy_magic_14_0.X.t54 353.467
R6861 two_stage_opamp_dummy_magic_14_0.X.n17 two_stage_opamp_dummy_magic_14_0.X.t28 353.467
R6862 two_stage_opamp_dummy_magic_14_0.X.n16 two_stage_opamp_dummy_magic_14_0.X.t53 353.467
R6863 two_stage_opamp_dummy_magic_14_0.X.n11 two_stage_opamp_dummy_magic_14_0.X.t30 353.467
R6864 two_stage_opamp_dummy_magic_14_0.X.n12 two_stage_opamp_dummy_magic_14_0.X.t47 353.467
R6865 two_stage_opamp_dummy_magic_14_0.X.n13 two_stage_opamp_dummy_magic_14_0.X.t33 353.467
R6866 two_stage_opamp_dummy_magic_14_0.X.n14 two_stage_opamp_dummy_magic_14_0.X.t50 353.467
R6867 two_stage_opamp_dummy_magic_14_0.X.n15 two_stage_opamp_dummy_magic_14_0.X.t37 353.467
R6868 two_stage_opamp_dummy_magic_14_0.X.n50 two_stage_opamp_dummy_magic_14_0.X.n49 176.733
R6869 two_stage_opamp_dummy_magic_14_0.X.n49 two_stage_opamp_dummy_magic_14_0.X.n48 176.733
R6870 two_stage_opamp_dummy_magic_14_0.X.n48 two_stage_opamp_dummy_magic_14_0.X.n47 176.733
R6871 two_stage_opamp_dummy_magic_14_0.X.n44 two_stage_opamp_dummy_magic_14_0.X.n43 176.733
R6872 two_stage_opamp_dummy_magic_14_0.X.n45 two_stage_opamp_dummy_magic_14_0.X.n44 176.733
R6873 two_stage_opamp_dummy_magic_14_0.X.n46 two_stage_opamp_dummy_magic_14_0.X.n45 176.733
R6874 two_stage_opamp_dummy_magic_14_0.X.n18 two_stage_opamp_dummy_magic_14_0.X.n17 176.733
R6875 two_stage_opamp_dummy_magic_14_0.X.n17 two_stage_opamp_dummy_magic_14_0.X.n16 176.733
R6876 two_stage_opamp_dummy_magic_14_0.X.n12 two_stage_opamp_dummy_magic_14_0.X.n11 176.733
R6877 two_stage_opamp_dummy_magic_14_0.X.n13 two_stage_opamp_dummy_magic_14_0.X.n12 176.733
R6878 two_stage_opamp_dummy_magic_14_0.X.n14 two_stage_opamp_dummy_magic_14_0.X.n13 176.733
R6879 two_stage_opamp_dummy_magic_14_0.X.n15 two_stage_opamp_dummy_magic_14_0.X.n14 176.733
R6880 two_stage_opamp_dummy_magic_14_0.X.n27 two_stage_opamp_dummy_magic_14_0.X.n26 176.733
R6881 two_stage_opamp_dummy_magic_14_0.X.n26 two_stage_opamp_dummy_magic_14_0.X.n25 176.733
R6882 two_stage_opamp_dummy_magic_14_0.X.n21 two_stage_opamp_dummy_magic_14_0.X.n20 176.733
R6883 two_stage_opamp_dummy_magic_14_0.X.n22 two_stage_opamp_dummy_magic_14_0.X.n21 176.733
R6884 two_stage_opamp_dummy_magic_14_0.X.n23 two_stage_opamp_dummy_magic_14_0.X.n22 176.733
R6885 two_stage_opamp_dummy_magic_14_0.X.n24 two_stage_opamp_dummy_magic_14_0.X.n23 176.733
R6886 two_stage_opamp_dummy_magic_14_0.X.n52 two_stage_opamp_dummy_magic_14_0.X.n51 166.258
R6887 two_stage_opamp_dummy_magic_14_0.X.n2 two_stage_opamp_dummy_magic_14_0.X.n0 163.626
R6888 two_stage_opamp_dummy_magic_14_0.X.n8 two_stage_opamp_dummy_magic_14_0.X.n7 163.001
R6889 two_stage_opamp_dummy_magic_14_0.X.n6 two_stage_opamp_dummy_magic_14_0.X.n5 163.001
R6890 two_stage_opamp_dummy_magic_14_0.X.n4 two_stage_opamp_dummy_magic_14_0.X.n3 163.001
R6891 two_stage_opamp_dummy_magic_14_0.X.n2 two_stage_opamp_dummy_magic_14_0.X.n1 163.001
R6892 two_stage_opamp_dummy_magic_14_0.X.n29 two_stage_opamp_dummy_magic_14_0.X.n19 161.541
R6893 two_stage_opamp_dummy_magic_14_0.X.n29 two_stage_opamp_dummy_magic_14_0.X.n28 161.541
R6894 two_stage_opamp_dummy_magic_14_0.X.n10 two_stage_opamp_dummy_magic_14_0.X.n9 158.501
R6895 two_stage_opamp_dummy_magic_14_0.X.n32 two_stage_opamp_dummy_magic_14_0.X.n30 117.888
R6896 two_stage_opamp_dummy_magic_14_0.X.n40 two_stage_opamp_dummy_magic_14_0.X.n39 117.326
R6897 two_stage_opamp_dummy_magic_14_0.X.n38 two_stage_opamp_dummy_magic_14_0.X.n37 117.326
R6898 two_stage_opamp_dummy_magic_14_0.X.n36 two_stage_opamp_dummy_magic_14_0.X.n35 117.326
R6899 two_stage_opamp_dummy_magic_14_0.X.n34 two_stage_opamp_dummy_magic_14_0.X.n33 117.326
R6900 two_stage_opamp_dummy_magic_14_0.X.n32 two_stage_opamp_dummy_magic_14_0.X.n31 117.326
R6901 two_stage_opamp_dummy_magic_14_0.X.n19 two_stage_opamp_dummy_magic_14_0.X.n18 54.6272
R6902 two_stage_opamp_dummy_magic_14_0.X.n19 two_stage_opamp_dummy_magic_14_0.X.n15 54.6272
R6903 two_stage_opamp_dummy_magic_14_0.X.n28 two_stage_opamp_dummy_magic_14_0.X.n27 54.6272
R6904 two_stage_opamp_dummy_magic_14_0.X.n28 two_stage_opamp_dummy_magic_14_0.X.n24 54.6272
R6905 two_stage_opamp_dummy_magic_14_0.X.n51 two_stage_opamp_dummy_magic_14_0.X.n50 53.3126
R6906 two_stage_opamp_dummy_magic_14_0.X.n51 two_stage_opamp_dummy_magic_14_0.X.n46 53.3126
R6907 two_stage_opamp_dummy_magic_14_0.X.t8 two_stage_opamp_dummy_magic_14_0.X.n52 50.3023
R6908 two_stage_opamp_dummy_magic_14_0.X.n42 two_stage_opamp_dummy_magic_14_0.X.n10 16.8755
R6909 two_stage_opamp_dummy_magic_14_0.X.n39 two_stage_opamp_dummy_magic_14_0.X.t19 16.0005
R6910 two_stage_opamp_dummy_magic_14_0.X.n39 two_stage_opamp_dummy_magic_14_0.X.t10 16.0005
R6911 two_stage_opamp_dummy_magic_14_0.X.n37 two_stage_opamp_dummy_magic_14_0.X.t11 16.0005
R6912 two_stage_opamp_dummy_magic_14_0.X.n37 two_stage_opamp_dummy_magic_14_0.X.t18 16.0005
R6913 two_stage_opamp_dummy_magic_14_0.X.n35 two_stage_opamp_dummy_magic_14_0.X.t17 16.0005
R6914 two_stage_opamp_dummy_magic_14_0.X.n35 two_stage_opamp_dummy_magic_14_0.X.t21 16.0005
R6915 two_stage_opamp_dummy_magic_14_0.X.n33 two_stage_opamp_dummy_magic_14_0.X.t16 16.0005
R6916 two_stage_opamp_dummy_magic_14_0.X.n33 two_stage_opamp_dummy_magic_14_0.X.t4 16.0005
R6917 two_stage_opamp_dummy_magic_14_0.X.n31 two_stage_opamp_dummy_magic_14_0.X.t6 16.0005
R6918 two_stage_opamp_dummy_magic_14_0.X.n31 two_stage_opamp_dummy_magic_14_0.X.t9 16.0005
R6919 two_stage_opamp_dummy_magic_14_0.X.n30 two_stage_opamp_dummy_magic_14_0.X.t1 16.0005
R6920 two_stage_opamp_dummy_magic_14_0.X.n30 two_stage_opamp_dummy_magic_14_0.X.t20 16.0005
R6921 two_stage_opamp_dummy_magic_14_0.X.n41 two_stage_opamp_dummy_magic_14_0.X.n29 11.9693
R6922 two_stage_opamp_dummy_magic_14_0.X.n9 two_stage_opamp_dummy_magic_14_0.X.t7 11.2576
R6923 two_stage_opamp_dummy_magic_14_0.X.n9 two_stage_opamp_dummy_magic_14_0.X.t2 11.2576
R6924 two_stage_opamp_dummy_magic_14_0.X.n7 two_stage_opamp_dummy_magic_14_0.X.t13 11.2576
R6925 two_stage_opamp_dummy_magic_14_0.X.n7 two_stage_opamp_dummy_magic_14_0.X.t12 11.2576
R6926 two_stage_opamp_dummy_magic_14_0.X.n5 two_stage_opamp_dummy_magic_14_0.X.t3 11.2576
R6927 two_stage_opamp_dummy_magic_14_0.X.n5 two_stage_opamp_dummy_magic_14_0.X.t23 11.2576
R6928 two_stage_opamp_dummy_magic_14_0.X.n3 two_stage_opamp_dummy_magic_14_0.X.t0 11.2576
R6929 two_stage_opamp_dummy_magic_14_0.X.n3 two_stage_opamp_dummy_magic_14_0.X.t22 11.2576
R6930 two_stage_opamp_dummy_magic_14_0.X.n1 two_stage_opamp_dummy_magic_14_0.X.t15 11.2576
R6931 two_stage_opamp_dummy_magic_14_0.X.n1 two_stage_opamp_dummy_magic_14_0.X.t24 11.2576
R6932 two_stage_opamp_dummy_magic_14_0.X.n0 two_stage_opamp_dummy_magic_14_0.X.t14 11.2576
R6933 two_stage_opamp_dummy_magic_14_0.X.n0 two_stage_opamp_dummy_magic_14_0.X.t5 11.2576
R6934 two_stage_opamp_dummy_magic_14_0.X.n52 two_stage_opamp_dummy_magic_14_0.X.n42 7.09425
R6935 two_stage_opamp_dummy_magic_14_0.X.n41 two_stage_opamp_dummy_magic_14_0.X.n40 6.3755
R6936 two_stage_opamp_dummy_magic_14_0.X.n10 two_stage_opamp_dummy_magic_14_0.X.n8 5.1255
R6937 two_stage_opamp_dummy_magic_14_0.X.n42 two_stage_opamp_dummy_magic_14_0.X.n41 1.3755
R6938 two_stage_opamp_dummy_magic_14_0.X.n4 two_stage_opamp_dummy_magic_14_0.X.n2 0.6255
R6939 two_stage_opamp_dummy_magic_14_0.X.n6 two_stage_opamp_dummy_magic_14_0.X.n4 0.6255
R6940 two_stage_opamp_dummy_magic_14_0.X.n8 two_stage_opamp_dummy_magic_14_0.X.n6 0.6255
R6941 two_stage_opamp_dummy_magic_14_0.X.n34 two_stage_opamp_dummy_magic_14_0.X.n32 0.563
R6942 two_stage_opamp_dummy_magic_14_0.X.n36 two_stage_opamp_dummy_magic_14_0.X.n34 0.563
R6943 two_stage_opamp_dummy_magic_14_0.X.n38 two_stage_opamp_dummy_magic_14_0.X.n36 0.563
R6944 two_stage_opamp_dummy_magic_14_0.X.n40 two_stage_opamp_dummy_magic_14_0.X.n38 0.563
R6945 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.n2 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.n0 144.827
R6946 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.n2 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.n1 134.577
R6947 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.n12 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.t14 118.986
R6948 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.n5 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.n3 100.6
R6949 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.n11 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.n10 100.038
R6950 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.n9 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.n8 100.038
R6951 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.n7 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.n6 100.038
R6952 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.n5 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.n4 100.038
R6953 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.n13 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.n12 43.284
R6954 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.n13 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.n2 37.4067
R6955 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.n1 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.t10 24.0005
R6956 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.n1 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.t11 24.0005
R6957 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.n0 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.t12 24.0005
R6958 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.n0 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.t13 24.0005
R6959 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.n10 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.t7 8.0005
R6960 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.n10 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.t1 8.0005
R6961 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.n8 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.t6 8.0005
R6962 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.n8 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.t0 8.0005
R6963 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.n6 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.t5 8.0005
R6964 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.n6 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.t9 8.0005
R6965 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.n4 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.t3 8.0005
R6966 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.n4 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.t2 8.0005
R6967 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.n3 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.t4 8.0005
R6968 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.n3 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.t8 8.0005
R6969 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.n12 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.n11 5.6255
R6970 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.n7 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.n5 0.563
R6971 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.n9 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.n7 0.563
R6972 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.n11 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.n9 0.563
R6973 bgr_0.V_CMFB_S2 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.n13 0.047375
R6974 two_stage_opamp_dummy_magic_14_0.V_b_2nd_stage.n4 two_stage_opamp_dummy_magic_14_0.V_b_2nd_stage.t4 525.38
R6975 two_stage_opamp_dummy_magic_14_0.V_b_2nd_stage.n0 two_stage_opamp_dummy_magic_14_0.V_b_2nd_stage.t9 525.38
R6976 two_stage_opamp_dummy_magic_14_0.V_b_2nd_stage.n6 two_stage_opamp_dummy_magic_14_0.V_b_2nd_stage.t3 358.288
R6977 two_stage_opamp_dummy_magic_14_0.V_b_2nd_stage.n2 two_stage_opamp_dummy_magic_14_0.V_b_2nd_stage.t2 358.288
R6978 two_stage_opamp_dummy_magic_14_0.V_b_2nd_stage.n4 two_stage_opamp_dummy_magic_14_0.V_b_2nd_stage.t7 281.168
R6979 two_stage_opamp_dummy_magic_14_0.V_b_2nd_stage.n5 two_stage_opamp_dummy_magic_14_0.V_b_2nd_stage.t6 281.168
R6980 two_stage_opamp_dummy_magic_14_0.V_b_2nd_stage.n0 two_stage_opamp_dummy_magic_14_0.V_b_2nd_stage.t5 281.168
R6981 two_stage_opamp_dummy_magic_14_0.V_b_2nd_stage.n1 two_stage_opamp_dummy_magic_14_0.V_b_2nd_stage.t8 281.168
R6982 two_stage_opamp_dummy_magic_14_0.V_b_2nd_stage.n5 two_stage_opamp_dummy_magic_14_0.V_b_2nd_stage.n4 244.214
R6983 two_stage_opamp_dummy_magic_14_0.V_b_2nd_stage.n1 two_stage_opamp_dummy_magic_14_0.V_b_2nd_stage.n0 244.214
R6984 two_stage_opamp_dummy_magic_14_0.V_b_2nd_stage.n7 two_stage_opamp_dummy_magic_14_0.V_b_2nd_stage.n6 166.019
R6985 two_stage_opamp_dummy_magic_14_0.V_b_2nd_stage.n3 two_stage_opamp_dummy_magic_14_0.V_b_2nd_stage.n2 166.019
R6986 two_stage_opamp_dummy_magic_14_0.V_b_2nd_stage.n3 two_stage_opamp_dummy_magic_14_0.V_b_2nd_stage.t1 116.013
R6987 two_stage_opamp_dummy_magic_14_0.V_b_2nd_stage.t0 two_stage_opamp_dummy_magic_14_0.V_b_2nd_stage.n7 116.013
R6988 two_stage_opamp_dummy_magic_14_0.V_b_2nd_stage.n6 two_stage_opamp_dummy_magic_14_0.V_b_2nd_stage.n5 77.1205
R6989 two_stage_opamp_dummy_magic_14_0.V_b_2nd_stage.n2 two_stage_opamp_dummy_magic_14_0.V_b_2nd_stage.n1 77.1205
R6990 two_stage_opamp_dummy_magic_14_0.V_b_2nd_stage.n7 two_stage_opamp_dummy_magic_14_0.V_b_2nd_stage.n3 18.0005
R6991 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.n1 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.t11 688.859
R6992 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.n0 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.t8 651.343
R6993 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.n0 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.t9 647.968
R6994 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.n3 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.n2 514.134
R6995 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.n5 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.n4 214.056
R6996 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.n1 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.t7 174.726
R6997 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.n2 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.t13 174.726
R6998 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.n3 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.t10 174.726
R6999 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.n4 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.t12 174.726
R7000 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.n8 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.n6 173.591
R7001 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.n10 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.n9 169.216
R7002 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.n8 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.n7 169.216
R7003 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.n2 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.n1 128.534
R7004 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.n4 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.n3 128.534
R7005 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.n5 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.t4 126.049
R7006 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.n11 46.7438
R7007 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.n9 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.t0 13.1338
R7008 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.n9 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.t5 13.1338
R7009 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.n7 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.t3 13.1338
R7010 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.n7 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.t1 13.1338
R7011 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.n6 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.t6 13.1338
R7012 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.n6 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.t2 13.1338
R7013 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.n11 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.n10 10.0317
R7014 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.n10 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.n8 4.3755
R7015 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.n11 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.n5 3.03175
R7016 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.n0 1.53175
R7017 two_stage_opamp_dummy_magic_14_0.err_amp_out.n1 two_stage_opamp_dummy_magic_14_0.err_amp_out.t4 685.303
R7018 two_stage_opamp_dummy_magic_14_0.err_amp_out.n1 two_stage_opamp_dummy_magic_14_0.err_amp_out.n0 179.257
R7019 two_stage_opamp_dummy_magic_14_0.err_amp_out.n2 two_stage_opamp_dummy_magic_14_0.err_amp_out.n1 100.93
R7020 two_stage_opamp_dummy_magic_14_0.err_amp_out.n0 two_stage_opamp_dummy_magic_14_0.err_amp_out.t3 15.7605
R7021 two_stage_opamp_dummy_magic_14_0.err_amp_out.n0 two_stage_opamp_dummy_magic_14_0.err_amp_out.t0 15.7605
R7022 two_stage_opamp_dummy_magic_14_0.err_amp_out.n2 two_stage_opamp_dummy_magic_14_0.err_amp_out.t2 9.6005
R7023 two_stage_opamp_dummy_magic_14_0.err_amp_out.t1 two_stage_opamp_dummy_magic_14_0.err_amp_out.n2 9.6005
R7024 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n17 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t13 610.534
R7025 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n8 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t16 610.534
R7026 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n17 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t31 433.8
R7027 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n18 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t22 433.8
R7028 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n19 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t29 433.8
R7029 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n20 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t19 433.8
R7030 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n21 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t27 433.8
R7031 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n22 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t17 433.8
R7032 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n23 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t25 433.8
R7033 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n24 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t14 433.8
R7034 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n25 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t21 433.8
R7035 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n16 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t12 433.8
R7036 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n15 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t23 433.8
R7037 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n14 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t30 433.8
R7038 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n13 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t20 433.8
R7039 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n12 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t28 433.8
R7040 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n11 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t18 433.8
R7041 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n10 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t26 433.8
R7042 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n9 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t15 433.8
R7043 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n8 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t24 433.8
R7044 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n4 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n0 339.836
R7045 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n3 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n1 339.834
R7046 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n3 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n2 339.272
R7047 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n6 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n5 287.264
R7048 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n25 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n24 176.733
R7049 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n24 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n23 176.733
R7050 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n23 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n22 176.733
R7051 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n22 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n21 176.733
R7052 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n21 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n20 176.733
R7053 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n20 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n19 176.733
R7054 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n19 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n18 176.733
R7055 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n18 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n17 176.733
R7056 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n9 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n8 176.733
R7057 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n10 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n9 176.733
R7058 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n11 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n10 176.733
R7059 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n12 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n11 176.733
R7060 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n13 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n12 176.733
R7061 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n14 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n13 176.733
R7062 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n15 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n14 176.733
R7063 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n16 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n15 176.733
R7064 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n27 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n26 162.102
R7065 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n27 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n7 112.278
R7066 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n29 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n27 68.723
R7067 two_stage_opamp_dummy_magic_14_0.V_tail_gate two_stage_opamp_dummy_magic_14_0.V_tail_gate.n29 58.7539
R7068 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n26 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n25 54.6272
R7069 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n26 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n16 54.6272
R7070 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n29 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n28 53.2453
R7071 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n6 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n4 52.01
R7072 two_stage_opamp_dummy_magic_14_0.V_tail_gate two_stage_opamp_dummy_magic_14_0.V_tail_gate.n6 51.6642
R7073 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n5 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t0 39.4005
R7074 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n5 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t3 39.4005
R7075 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n2 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t2 39.4005
R7076 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n2 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t6 39.4005
R7077 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n1 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t5 39.4005
R7078 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n1 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t8 39.4005
R7079 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n0 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t11 39.4005
R7080 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n0 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t7 39.4005
R7081 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n28 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t9 16.0005
R7082 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n28 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t1 16.0005
R7083 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n7 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t4 16.0005
R7084 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n7 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t10 16.0005
R7085 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n4 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n3 0.563
R7086 two_stage_opamp_dummy_magic_14_0.V_source.n30 two_stage_opamp_dummy_magic_14_0.V_source.t5 217.776
R7087 two_stage_opamp_dummy_magic_14_0.V_source.n12 two_stage_opamp_dummy_magic_14_0.V_source.n10 114.469
R7088 two_stage_opamp_dummy_magic_14_0.V_source.n5 two_stage_opamp_dummy_magic_14_0.V_source.n3 114.469
R7089 two_stage_opamp_dummy_magic_14_0.V_source.n18 two_stage_opamp_dummy_magic_14_0.V_source.n17 113.906
R7090 two_stage_opamp_dummy_magic_14_0.V_source.n16 two_stage_opamp_dummy_magic_14_0.V_source.n15 113.906
R7091 two_stage_opamp_dummy_magic_14_0.V_source.n14 two_stage_opamp_dummy_magic_14_0.V_source.n13 113.906
R7092 two_stage_opamp_dummy_magic_14_0.V_source.n12 two_stage_opamp_dummy_magic_14_0.V_source.n11 113.906
R7093 two_stage_opamp_dummy_magic_14_0.V_source.n9 two_stage_opamp_dummy_magic_14_0.V_source.n8 113.906
R7094 two_stage_opamp_dummy_magic_14_0.V_source.n7 two_stage_opamp_dummy_magic_14_0.V_source.n6 113.906
R7095 two_stage_opamp_dummy_magic_14_0.V_source.n5 two_stage_opamp_dummy_magic_14_0.V_source.n4 113.906
R7096 two_stage_opamp_dummy_magic_14_0.V_source.n21 two_stage_opamp_dummy_magic_14_0.V_source.n20 109.406
R7097 two_stage_opamp_dummy_magic_14_0.V_source.n2 two_stage_opamp_dummy_magic_14_0.V_source.n0 102.941
R7098 two_stage_opamp_dummy_magic_14_0.V_source.n38 two_stage_opamp_dummy_magic_14_0.V_source.n37 102.285
R7099 two_stage_opamp_dummy_magic_14_0.V_source.n36 two_stage_opamp_dummy_magic_14_0.V_source.n35 102.284
R7100 two_stage_opamp_dummy_magic_14_0.V_source.n34 two_stage_opamp_dummy_magic_14_0.V_source.n33 102.284
R7101 two_stage_opamp_dummy_magic_14_0.V_source.n32 two_stage_opamp_dummy_magic_14_0.V_source.n31 102.284
R7102 two_stage_opamp_dummy_magic_14_0.V_source.n30 two_stage_opamp_dummy_magic_14_0.V_source.n29 102.284
R7103 two_stage_opamp_dummy_magic_14_0.V_source.n28 two_stage_opamp_dummy_magic_14_0.V_source.n27 102.284
R7104 two_stage_opamp_dummy_magic_14_0.V_source.n26 two_stage_opamp_dummy_magic_14_0.V_source.n25 102.284
R7105 two_stage_opamp_dummy_magic_14_0.V_source.n2 two_stage_opamp_dummy_magic_14_0.V_source.n1 102.284
R7106 two_stage_opamp_dummy_magic_14_0.V_source.n23 two_stage_opamp_dummy_magic_14_0.V_source.n22 97.7845
R7107 two_stage_opamp_dummy_magic_14_0.V_source.n20 two_stage_opamp_dummy_magic_14_0.V_source.t6 16.0005
R7108 two_stage_opamp_dummy_magic_14_0.V_source.n20 two_stage_opamp_dummy_magic_14_0.V_source.t8 16.0005
R7109 two_stage_opamp_dummy_magic_14_0.V_source.n17 two_stage_opamp_dummy_magic_14_0.V_source.t31 16.0005
R7110 two_stage_opamp_dummy_magic_14_0.V_source.n17 two_stage_opamp_dummy_magic_14_0.V_source.t36 16.0005
R7111 two_stage_opamp_dummy_magic_14_0.V_source.n15 two_stage_opamp_dummy_magic_14_0.V_source.t33 16.0005
R7112 two_stage_opamp_dummy_magic_14_0.V_source.n15 two_stage_opamp_dummy_magic_14_0.V_source.t10 16.0005
R7113 two_stage_opamp_dummy_magic_14_0.V_source.n13 two_stage_opamp_dummy_magic_14_0.V_source.t35 16.0005
R7114 two_stage_opamp_dummy_magic_14_0.V_source.n13 two_stage_opamp_dummy_magic_14_0.V_source.t34 16.0005
R7115 two_stage_opamp_dummy_magic_14_0.V_source.n11 two_stage_opamp_dummy_magic_14_0.V_source.t11 16.0005
R7116 two_stage_opamp_dummy_magic_14_0.V_source.n11 two_stage_opamp_dummy_magic_14_0.V_source.t0 16.0005
R7117 two_stage_opamp_dummy_magic_14_0.V_source.n10 two_stage_opamp_dummy_magic_14_0.V_source.t38 16.0005
R7118 two_stage_opamp_dummy_magic_14_0.V_source.n10 two_stage_opamp_dummy_magic_14_0.V_source.t32 16.0005
R7119 two_stage_opamp_dummy_magic_14_0.V_source.n8 two_stage_opamp_dummy_magic_14_0.V_source.t39 16.0005
R7120 two_stage_opamp_dummy_magic_14_0.V_source.n8 two_stage_opamp_dummy_magic_14_0.V_source.t4 16.0005
R7121 two_stage_opamp_dummy_magic_14_0.V_source.n6 two_stage_opamp_dummy_magic_14_0.V_source.t37 16.0005
R7122 two_stage_opamp_dummy_magic_14_0.V_source.n6 two_stage_opamp_dummy_magic_14_0.V_source.t9 16.0005
R7123 two_stage_opamp_dummy_magic_14_0.V_source.n4 two_stage_opamp_dummy_magic_14_0.V_source.t7 16.0005
R7124 two_stage_opamp_dummy_magic_14_0.V_source.n4 two_stage_opamp_dummy_magic_14_0.V_source.t3 16.0005
R7125 two_stage_opamp_dummy_magic_14_0.V_source.n3 two_stage_opamp_dummy_magic_14_0.V_source.t40 16.0005
R7126 two_stage_opamp_dummy_magic_14_0.V_source.n3 two_stage_opamp_dummy_magic_14_0.V_source.t2 16.0005
R7127 two_stage_opamp_dummy_magic_14_0.V_source.n35 two_stage_opamp_dummy_magic_14_0.V_source.t21 9.6005
R7128 two_stage_opamp_dummy_magic_14_0.V_source.n35 two_stage_opamp_dummy_magic_14_0.V_source.t28 9.6005
R7129 two_stage_opamp_dummy_magic_14_0.V_source.n33 two_stage_opamp_dummy_magic_14_0.V_source.t17 9.6005
R7130 two_stage_opamp_dummy_magic_14_0.V_source.n33 two_stage_opamp_dummy_magic_14_0.V_source.t25 9.6005
R7131 two_stage_opamp_dummy_magic_14_0.V_source.n31 two_stage_opamp_dummy_magic_14_0.V_source.t15 9.6005
R7132 two_stage_opamp_dummy_magic_14_0.V_source.n31 two_stage_opamp_dummy_magic_14_0.V_source.t23 9.6005
R7133 two_stage_opamp_dummy_magic_14_0.V_source.n29 two_stage_opamp_dummy_magic_14_0.V_source.t13 9.6005
R7134 two_stage_opamp_dummy_magic_14_0.V_source.n29 two_stage_opamp_dummy_magic_14_0.V_source.t20 9.6005
R7135 two_stage_opamp_dummy_magic_14_0.V_source.n27 two_stage_opamp_dummy_magic_14_0.V_source.t22 9.6005
R7136 two_stage_opamp_dummy_magic_14_0.V_source.n27 two_stage_opamp_dummy_magic_14_0.V_source.t12 9.6005
R7137 two_stage_opamp_dummy_magic_14_0.V_source.n25 two_stage_opamp_dummy_magic_14_0.V_source.t24 9.6005
R7138 two_stage_opamp_dummy_magic_14_0.V_source.n25 two_stage_opamp_dummy_magic_14_0.V_source.t14 9.6005
R7139 two_stage_opamp_dummy_magic_14_0.V_source.n22 two_stage_opamp_dummy_magic_14_0.V_source.t27 9.6005
R7140 two_stage_opamp_dummy_magic_14_0.V_source.n22 two_stage_opamp_dummy_magic_14_0.V_source.t16 9.6005
R7141 two_stage_opamp_dummy_magic_14_0.V_source.n1 two_stage_opamp_dummy_magic_14_0.V_source.t26 9.6005
R7142 two_stage_opamp_dummy_magic_14_0.V_source.n1 two_stage_opamp_dummy_magic_14_0.V_source.t18 9.6005
R7143 two_stage_opamp_dummy_magic_14_0.V_source.n0 two_stage_opamp_dummy_magic_14_0.V_source.t30 9.6005
R7144 two_stage_opamp_dummy_magic_14_0.V_source.n0 two_stage_opamp_dummy_magic_14_0.V_source.t1 9.6005
R7145 two_stage_opamp_dummy_magic_14_0.V_source.n38 two_stage_opamp_dummy_magic_14_0.V_source.t19 9.6005
R7146 two_stage_opamp_dummy_magic_14_0.V_source.t29 two_stage_opamp_dummy_magic_14_0.V_source.n38 9.6005
R7147 two_stage_opamp_dummy_magic_14_0.V_source.n21 two_stage_opamp_dummy_magic_14_0.V_source.n19 4.5005
R7148 two_stage_opamp_dummy_magic_14_0.V_source.n24 two_stage_opamp_dummy_magic_14_0.V_source.n23 4.5005
R7149 two_stage_opamp_dummy_magic_14_0.V_source.n19 two_stage_opamp_dummy_magic_14_0.V_source.n18 3.6255
R7150 two_stage_opamp_dummy_magic_14_0.V_source.n23 two_stage_opamp_dummy_magic_14_0.V_source.n21 1.61856
R7151 two_stage_opamp_dummy_magic_14_0.V_source.n32 two_stage_opamp_dummy_magic_14_0.V_source.n30 0.563
R7152 two_stage_opamp_dummy_magic_14_0.V_source.n34 two_stage_opamp_dummy_magic_14_0.V_source.n32 0.563
R7153 two_stage_opamp_dummy_magic_14_0.V_source.n36 two_stage_opamp_dummy_magic_14_0.V_source.n34 0.563
R7154 two_stage_opamp_dummy_magic_14_0.V_source.n37 two_stage_opamp_dummy_magic_14_0.V_source.n36 0.563
R7155 two_stage_opamp_dummy_magic_14_0.V_source.n14 two_stage_opamp_dummy_magic_14_0.V_source.n12 0.563
R7156 two_stage_opamp_dummy_magic_14_0.V_source.n16 two_stage_opamp_dummy_magic_14_0.V_source.n14 0.563
R7157 two_stage_opamp_dummy_magic_14_0.V_source.n18 two_stage_opamp_dummy_magic_14_0.V_source.n16 0.563
R7158 two_stage_opamp_dummy_magic_14_0.V_source.n7 two_stage_opamp_dummy_magic_14_0.V_source.n5 0.563
R7159 two_stage_opamp_dummy_magic_14_0.V_source.n9 two_stage_opamp_dummy_magic_14_0.V_source.n7 0.563
R7160 two_stage_opamp_dummy_magic_14_0.V_source.n19 two_stage_opamp_dummy_magic_14_0.V_source.n9 0.563
R7161 two_stage_opamp_dummy_magic_14_0.V_source.n24 two_stage_opamp_dummy_magic_14_0.V_source.n2 0.563
R7162 two_stage_opamp_dummy_magic_14_0.V_source.n26 two_stage_opamp_dummy_magic_14_0.V_source.n24 0.563
R7163 two_stage_opamp_dummy_magic_14_0.V_source.n28 two_stage_opamp_dummy_magic_14_0.V_source.n26 0.563
R7164 two_stage_opamp_dummy_magic_14_0.V_source.n37 two_stage_opamp_dummy_magic_14_0.V_source.n28 0.563
R7165 bgr_0.Vin+.n3 bgr_0.Vin+.n2 526.183
R7166 bgr_0.Vin+.n1 bgr_0.Vin+.n0 514.134
R7167 bgr_0.Vin+.n0 bgr_0.Vin+.t8 303.259
R7168 bgr_0.Vin+.n5 bgr_0.Vin+.n3 227.169
R7169 bgr_0.Vin+.n0 bgr_0.Vin+.t9 174.726
R7170 bgr_0.Vin+.n1 bgr_0.Vin+.t6 174.726
R7171 bgr_0.Vin+.n2 bgr_0.Vin+.t10 174.726
R7172 bgr_0.Vin+.n7 bgr_0.Vin+.n6 168.435
R7173 bgr_0.Vin+.n5 bgr_0.Vin+.n4 168.435
R7174 bgr_0.Vin+.n8 bgr_0.Vin+.t5 158.989
R7175 bgr_0.Vin+.n2 bgr_0.Vin+.n1 128.534
R7176 bgr_0.Vin+.t4 bgr_0.Vin+.n8 119.067
R7177 bgr_0.Vin+.n3 bgr_0.Vin+.t7 96.4005
R7178 bgr_0.Vin+.n8 bgr_0.Vin+.n7 35.0317
R7179 bgr_0.Vin+.n6 bgr_0.Vin+.t0 13.1338
R7180 bgr_0.Vin+.n6 bgr_0.Vin+.t3 13.1338
R7181 bgr_0.Vin+.n4 bgr_0.Vin+.t2 13.1338
R7182 bgr_0.Vin+.n4 bgr_0.Vin+.t1 13.1338
R7183 bgr_0.Vin+.n7 bgr_0.Vin+.n5 2.1255
R7184 two_stage_opamp_dummy_magic_14_0.VD3.n28 two_stage_opamp_dummy_magic_14_0.VD3.t6 652.076
R7185 two_stage_opamp_dummy_magic_14_0.VD3.n59 two_stage_opamp_dummy_magic_14_0.VD3.t9 652.076
R7186 two_stage_opamp_dummy_magic_14_0.VD3.n58 two_stage_opamp_dummy_magic_14_0.VD3.n11 585
R7187 two_stage_opamp_dummy_magic_14_0.VD3.n42 two_stage_opamp_dummy_magic_14_0.VD3.n29 585
R7188 two_stage_opamp_dummy_magic_14_0.VD3.n46 two_stage_opamp_dummy_magic_14_0.VD3.n11 290.233
R7189 two_stage_opamp_dummy_magic_14_0.VD3.n52 two_stage_opamp_dummy_magic_14_0.VD3.n11 290.233
R7190 two_stage_opamp_dummy_magic_14_0.VD3.n47 two_stage_opamp_dummy_magic_14_0.VD3.n11 290.233
R7191 two_stage_opamp_dummy_magic_14_0.VD3.n40 two_stage_opamp_dummy_magic_14_0.VD3.n29 290.233
R7192 two_stage_opamp_dummy_magic_14_0.VD3.n35 two_stage_opamp_dummy_magic_14_0.VD3.n29 290.233
R7193 two_stage_opamp_dummy_magic_14_0.VD3.n30 two_stage_opamp_dummy_magic_14_0.VD3.n29 290.233
R7194 two_stage_opamp_dummy_magic_14_0.VD3.n47 two_stage_opamp_dummy_magic_14_0.VD3.n15 242.903
R7195 two_stage_opamp_dummy_magic_14_0.VD3.n30 two_stage_opamp_dummy_magic_14_0.VD3.n18 242.903
R7196 two_stage_opamp_dummy_magic_14_0.VD3.n58 two_stage_opamp_dummy_magic_14_0.VD3.n57 238.367
R7197 two_stage_opamp_dummy_magic_14_0.VD3.n13 two_stage_opamp_dummy_magic_14_0.VD3.n12 185
R7198 two_stage_opamp_dummy_magic_14_0.VD3.n55 two_stage_opamp_dummy_magic_14_0.VD3.n54 185
R7199 two_stage_opamp_dummy_magic_14_0.VD3.n56 two_stage_opamp_dummy_magic_14_0.VD3.n55 185
R7200 two_stage_opamp_dummy_magic_14_0.VD3.n53 two_stage_opamp_dummy_magic_14_0.VD3.n45 185
R7201 two_stage_opamp_dummy_magic_14_0.VD3.n51 two_stage_opamp_dummy_magic_14_0.VD3.n50 185
R7202 two_stage_opamp_dummy_magic_14_0.VD3.n49 two_stage_opamp_dummy_magic_14_0.VD3.n48 185
R7203 two_stage_opamp_dummy_magic_14_0.VD3.n43 two_stage_opamp_dummy_magic_14_0.VD3.n42 185
R7204 two_stage_opamp_dummy_magic_14_0.VD3.n44 two_stage_opamp_dummy_magic_14_0.VD3.n43 185
R7205 two_stage_opamp_dummy_magic_14_0.VD3.n41 two_stage_opamp_dummy_magic_14_0.VD3.n19 185
R7206 two_stage_opamp_dummy_magic_14_0.VD3.n39 two_stage_opamp_dummy_magic_14_0.VD3.n38 185
R7207 two_stage_opamp_dummy_magic_14_0.VD3.n37 two_stage_opamp_dummy_magic_14_0.VD3.n36 185
R7208 two_stage_opamp_dummy_magic_14_0.VD3.n34 two_stage_opamp_dummy_magic_14_0.VD3.n33 185
R7209 two_stage_opamp_dummy_magic_14_0.VD3.n32 two_stage_opamp_dummy_magic_14_0.VD3.n31 185
R7210 two_stage_opamp_dummy_magic_14_0.VD3.n56 two_stage_opamp_dummy_magic_14_0.VD3.t10 170.513
R7211 two_stage_opamp_dummy_magic_14_0.VD3.t7 two_stage_opamp_dummy_magic_14_0.VD3.n44 170.513
R7212 two_stage_opamp_dummy_magic_14_0.VD3.n2 two_stage_opamp_dummy_magic_14_0.VD3.n0 163.626
R7213 two_stage_opamp_dummy_magic_14_0.VD3.n8 two_stage_opamp_dummy_magic_14_0.VD3.n7 163.001
R7214 two_stage_opamp_dummy_magic_14_0.VD3.n6 two_stage_opamp_dummy_magic_14_0.VD3.n5 163.001
R7215 two_stage_opamp_dummy_magic_14_0.VD3.n4 two_stage_opamp_dummy_magic_14_0.VD3.n3 163.001
R7216 two_stage_opamp_dummy_magic_14_0.VD3.n2 two_stage_opamp_dummy_magic_14_0.VD3.n1 163.001
R7217 two_stage_opamp_dummy_magic_14_0.VD3.n62 two_stage_opamp_dummy_magic_14_0.VD3.n61 162.999
R7218 two_stage_opamp_dummy_magic_14_0.VD3.n10 two_stage_opamp_dummy_magic_14_0.VD3.n9 159.803
R7219 two_stage_opamp_dummy_magic_14_0.VD3.n21 two_stage_opamp_dummy_magic_14_0.VD3.n20 159.803
R7220 two_stage_opamp_dummy_magic_14_0.VD3.n23 two_stage_opamp_dummy_magic_14_0.VD3.n22 159.803
R7221 two_stage_opamp_dummy_magic_14_0.VD3.n25 two_stage_opamp_dummy_magic_14_0.VD3.n24 159.803
R7222 two_stage_opamp_dummy_magic_14_0.VD3.n27 two_stage_opamp_dummy_magic_14_0.VD3.n26 159.803
R7223 two_stage_opamp_dummy_magic_14_0.VD3.n55 two_stage_opamp_dummy_magic_14_0.VD3.n13 150
R7224 two_stage_opamp_dummy_magic_14_0.VD3.n55 two_stage_opamp_dummy_magic_14_0.VD3.n45 150
R7225 two_stage_opamp_dummy_magic_14_0.VD3.n50 two_stage_opamp_dummy_magic_14_0.VD3.n49 150
R7226 two_stage_opamp_dummy_magic_14_0.VD3.n43 two_stage_opamp_dummy_magic_14_0.VD3.n19 150
R7227 two_stage_opamp_dummy_magic_14_0.VD3.n38 two_stage_opamp_dummy_magic_14_0.VD3.n37 150
R7228 two_stage_opamp_dummy_magic_14_0.VD3.n33 two_stage_opamp_dummy_magic_14_0.VD3.n32 150
R7229 two_stage_opamp_dummy_magic_14_0.VD3.t10 two_stage_opamp_dummy_magic_14_0.VD3.t2 146.155
R7230 two_stage_opamp_dummy_magic_14_0.VD3.t2 two_stage_opamp_dummy_magic_14_0.VD3.t14 146.155
R7231 two_stage_opamp_dummy_magic_14_0.VD3.t14 two_stage_opamp_dummy_magic_14_0.VD3.t12 146.155
R7232 two_stage_opamp_dummy_magic_14_0.VD3.t12 two_stage_opamp_dummy_magic_14_0.VD3.t4 146.155
R7233 two_stage_opamp_dummy_magic_14_0.VD3.t4 two_stage_opamp_dummy_magic_14_0.VD3.t34 146.155
R7234 two_stage_opamp_dummy_magic_14_0.VD3.t34 two_stage_opamp_dummy_magic_14_0.VD3.t0 146.155
R7235 two_stage_opamp_dummy_magic_14_0.VD3.t0 two_stage_opamp_dummy_magic_14_0.VD3.t32 146.155
R7236 two_stage_opamp_dummy_magic_14_0.VD3.t32 two_stage_opamp_dummy_magic_14_0.VD3.t18 146.155
R7237 two_stage_opamp_dummy_magic_14_0.VD3.t18 two_stage_opamp_dummy_magic_14_0.VD3.t36 146.155
R7238 two_stage_opamp_dummy_magic_14_0.VD3.t36 two_stage_opamp_dummy_magic_14_0.VD3.t16 146.155
R7239 two_stage_opamp_dummy_magic_14_0.VD3.t16 two_stage_opamp_dummy_magic_14_0.VD3.t7 146.155
R7240 two_stage_opamp_dummy_magic_14_0.VD3.n57 two_stage_opamp_dummy_magic_14_0.VD3.n56 65.8183
R7241 two_stage_opamp_dummy_magic_14_0.VD3.n56 two_stage_opamp_dummy_magic_14_0.VD3.n14 65.8183
R7242 two_stage_opamp_dummy_magic_14_0.VD3.n56 two_stage_opamp_dummy_magic_14_0.VD3.n15 65.8183
R7243 two_stage_opamp_dummy_magic_14_0.VD3.n44 two_stage_opamp_dummy_magic_14_0.VD3.n16 65.8183
R7244 two_stage_opamp_dummy_magic_14_0.VD3.n44 two_stage_opamp_dummy_magic_14_0.VD3.n17 65.8183
R7245 two_stage_opamp_dummy_magic_14_0.VD3.n44 two_stage_opamp_dummy_magic_14_0.VD3.n18 65.8183
R7246 two_stage_opamp_dummy_magic_14_0.VD3.n45 two_stage_opamp_dummy_magic_14_0.VD3.n14 53.3664
R7247 two_stage_opamp_dummy_magic_14_0.VD3.n49 two_stage_opamp_dummy_magic_14_0.VD3.n15 53.3664
R7248 two_stage_opamp_dummy_magic_14_0.VD3.n57 two_stage_opamp_dummy_magic_14_0.VD3.n13 53.3664
R7249 two_stage_opamp_dummy_magic_14_0.VD3.n50 two_stage_opamp_dummy_magic_14_0.VD3.n14 53.3664
R7250 two_stage_opamp_dummy_magic_14_0.VD3.n19 two_stage_opamp_dummy_magic_14_0.VD3.n16 53.3664
R7251 two_stage_opamp_dummy_magic_14_0.VD3.n37 two_stage_opamp_dummy_magic_14_0.VD3.n17 53.3664
R7252 two_stage_opamp_dummy_magic_14_0.VD3.n32 two_stage_opamp_dummy_magic_14_0.VD3.n18 53.3664
R7253 two_stage_opamp_dummy_magic_14_0.VD3.n38 two_stage_opamp_dummy_magic_14_0.VD3.n16 53.3664
R7254 two_stage_opamp_dummy_magic_14_0.VD3.n33 two_stage_opamp_dummy_magic_14_0.VD3.n17 53.3664
R7255 two_stage_opamp_dummy_magic_14_0.VD3.n59 two_stage_opamp_dummy_magic_14_0.VD3.n58 22.8576
R7256 two_stage_opamp_dummy_magic_14_0.VD3.n42 two_stage_opamp_dummy_magic_14_0.VD3.n28 22.8576
R7257 two_stage_opamp_dummy_magic_14_0.VD3.n28 two_stage_opamp_dummy_magic_14_0.VD3.n27 14.4255
R7258 two_stage_opamp_dummy_magic_14_0.VD3.n60 two_stage_opamp_dummy_magic_14_0.VD3.n59 13.8005
R7259 two_stage_opamp_dummy_magic_14_0.VD3.n61 two_stage_opamp_dummy_magic_14_0.VD3.n60 13.688
R7260 two_stage_opamp_dummy_magic_14_0.VD3.n9 two_stage_opamp_dummy_magic_14_0.VD3.t3 11.2576
R7261 two_stage_opamp_dummy_magic_14_0.VD3.n9 two_stage_opamp_dummy_magic_14_0.VD3.t15 11.2576
R7262 two_stage_opamp_dummy_magic_14_0.VD3.n20 two_stage_opamp_dummy_magic_14_0.VD3.t13 11.2576
R7263 two_stage_opamp_dummy_magic_14_0.VD3.n20 two_stage_opamp_dummy_magic_14_0.VD3.t5 11.2576
R7264 two_stage_opamp_dummy_magic_14_0.VD3.n22 two_stage_opamp_dummy_magic_14_0.VD3.t35 11.2576
R7265 two_stage_opamp_dummy_magic_14_0.VD3.n22 two_stage_opamp_dummy_magic_14_0.VD3.t1 11.2576
R7266 two_stage_opamp_dummy_magic_14_0.VD3.n24 two_stage_opamp_dummy_magic_14_0.VD3.t33 11.2576
R7267 two_stage_opamp_dummy_magic_14_0.VD3.n24 two_stage_opamp_dummy_magic_14_0.VD3.t19 11.2576
R7268 two_stage_opamp_dummy_magic_14_0.VD3.n26 two_stage_opamp_dummy_magic_14_0.VD3.t37 11.2576
R7269 two_stage_opamp_dummy_magic_14_0.VD3.n26 two_stage_opamp_dummy_magic_14_0.VD3.t17 11.2576
R7270 two_stage_opamp_dummy_magic_14_0.VD3.n11 two_stage_opamp_dummy_magic_14_0.VD3.t11 11.2576
R7271 two_stage_opamp_dummy_magic_14_0.VD3.n29 two_stage_opamp_dummy_magic_14_0.VD3.t8 11.2576
R7272 two_stage_opamp_dummy_magic_14_0.VD3.n7 two_stage_opamp_dummy_magic_14_0.VD3.t24 11.2576
R7273 two_stage_opamp_dummy_magic_14_0.VD3.n7 two_stage_opamp_dummy_magic_14_0.VD3.t27 11.2576
R7274 two_stage_opamp_dummy_magic_14_0.VD3.n5 two_stage_opamp_dummy_magic_14_0.VD3.t21 11.2576
R7275 two_stage_opamp_dummy_magic_14_0.VD3.n5 two_stage_opamp_dummy_magic_14_0.VD3.t22 11.2576
R7276 two_stage_opamp_dummy_magic_14_0.VD3.n3 two_stage_opamp_dummy_magic_14_0.VD3.t28 11.2576
R7277 two_stage_opamp_dummy_magic_14_0.VD3.n3 two_stage_opamp_dummy_magic_14_0.VD3.t20 11.2576
R7278 two_stage_opamp_dummy_magic_14_0.VD3.n1 two_stage_opamp_dummy_magic_14_0.VD3.t23 11.2576
R7279 two_stage_opamp_dummy_magic_14_0.VD3.n1 two_stage_opamp_dummy_magic_14_0.VD3.t26 11.2576
R7280 two_stage_opamp_dummy_magic_14_0.VD3.n0 two_stage_opamp_dummy_magic_14_0.VD3.t31 11.2576
R7281 two_stage_opamp_dummy_magic_14_0.VD3.n0 two_stage_opamp_dummy_magic_14_0.VD3.t25 11.2576
R7282 two_stage_opamp_dummy_magic_14_0.VD3.t29 two_stage_opamp_dummy_magic_14_0.VD3.n62 11.2576
R7283 two_stage_opamp_dummy_magic_14_0.VD3.n62 two_stage_opamp_dummy_magic_14_0.VD3.t30 11.2576
R7284 two_stage_opamp_dummy_magic_14_0.VD3.n58 two_stage_opamp_dummy_magic_14_0.VD3.n12 9.14336
R7285 two_stage_opamp_dummy_magic_14_0.VD3.n54 two_stage_opamp_dummy_magic_14_0.VD3.n53 9.14336
R7286 two_stage_opamp_dummy_magic_14_0.VD3.n51 two_stage_opamp_dummy_magic_14_0.VD3.n48 9.14336
R7287 two_stage_opamp_dummy_magic_14_0.VD3.n42 two_stage_opamp_dummy_magic_14_0.VD3.n41 9.14336
R7288 two_stage_opamp_dummy_magic_14_0.VD3.n39 two_stage_opamp_dummy_magic_14_0.VD3.n36 9.14336
R7289 two_stage_opamp_dummy_magic_14_0.VD3.n34 two_stage_opamp_dummy_magic_14_0.VD3.n31 9.14336
R7290 two_stage_opamp_dummy_magic_14_0.VD3.n46 two_stage_opamp_dummy_magic_14_0.VD3.n12 4.53698
R7291 two_stage_opamp_dummy_magic_14_0.VD3.n53 two_stage_opamp_dummy_magic_14_0.VD3.n52 4.53698
R7292 two_stage_opamp_dummy_magic_14_0.VD3.n48 two_stage_opamp_dummy_magic_14_0.VD3.n47 4.53698
R7293 two_stage_opamp_dummy_magic_14_0.VD3.n54 two_stage_opamp_dummy_magic_14_0.VD3.n46 4.53698
R7294 two_stage_opamp_dummy_magic_14_0.VD3.n52 two_stage_opamp_dummy_magic_14_0.VD3.n51 4.53698
R7295 two_stage_opamp_dummy_magic_14_0.VD3.n41 two_stage_opamp_dummy_magic_14_0.VD3.n40 4.53698
R7296 two_stage_opamp_dummy_magic_14_0.VD3.n36 two_stage_opamp_dummy_magic_14_0.VD3.n35 4.53698
R7297 two_stage_opamp_dummy_magic_14_0.VD3.n31 two_stage_opamp_dummy_magic_14_0.VD3.n30 4.53698
R7298 two_stage_opamp_dummy_magic_14_0.VD3.n40 two_stage_opamp_dummy_magic_14_0.VD3.n39 4.53698
R7299 two_stage_opamp_dummy_magic_14_0.VD3.n35 two_stage_opamp_dummy_magic_14_0.VD3.n34 4.53698
R7300 two_stage_opamp_dummy_magic_14_0.VD3.n27 two_stage_opamp_dummy_magic_14_0.VD3.n25 0.6255
R7301 two_stage_opamp_dummy_magic_14_0.VD3.n25 two_stage_opamp_dummy_magic_14_0.VD3.n23 0.6255
R7302 two_stage_opamp_dummy_magic_14_0.VD3.n23 two_stage_opamp_dummy_magic_14_0.VD3.n21 0.6255
R7303 two_stage_opamp_dummy_magic_14_0.VD3.n21 two_stage_opamp_dummy_magic_14_0.VD3.n10 0.6255
R7304 two_stage_opamp_dummy_magic_14_0.VD3.n60 two_stage_opamp_dummy_magic_14_0.VD3.n10 0.6255
R7305 two_stage_opamp_dummy_magic_14_0.VD3.n4 two_stage_opamp_dummy_magic_14_0.VD3.n2 0.6255
R7306 two_stage_opamp_dummy_magic_14_0.VD3.n6 two_stage_opamp_dummy_magic_14_0.VD3.n4 0.6255
R7307 two_stage_opamp_dummy_magic_14_0.VD3.n8 two_stage_opamp_dummy_magic_14_0.VD3.n6 0.6255
R7308 two_stage_opamp_dummy_magic_14_0.VD3.n61 two_stage_opamp_dummy_magic_14_0.VD3.n8 0.6255
R7309 bgr_0.V_mir1.n20 bgr_0.V_mir1.n19 325.473
R7310 bgr_0.V_mir1.n13 bgr_0.V_mir1.n12 325.473
R7311 bgr_0.V_mir1.n4 bgr_0.V_mir1.n3 325.473
R7312 bgr_0.V_mir1.n16 bgr_0.V_mir1.t19 310.488
R7313 bgr_0.V_mir1.n9 bgr_0.V_mir1.t21 310.488
R7314 bgr_0.V_mir1.n0 bgr_0.V_mir1.t20 310.488
R7315 bgr_0.V_mir1.n7 bgr_0.V_mir1.t2 278.312
R7316 bgr_0.V_mir1.n7 bgr_0.V_mir1.n6 228.939
R7317 bgr_0.V_mir1.n8 bgr_0.V_mir1.n5 224.439
R7318 bgr_0.V_mir1.n18 bgr_0.V_mir1.t9 184.097
R7319 bgr_0.V_mir1.n11 bgr_0.V_mir1.t5 184.097
R7320 bgr_0.V_mir1.n2 bgr_0.V_mir1.t3 184.097
R7321 bgr_0.V_mir1.n17 bgr_0.V_mir1.n16 167.094
R7322 bgr_0.V_mir1.n10 bgr_0.V_mir1.n9 167.094
R7323 bgr_0.V_mir1.n1 bgr_0.V_mir1.n0 167.094
R7324 bgr_0.V_mir1.n13 bgr_0.V_mir1.n11 152
R7325 bgr_0.V_mir1.n4 bgr_0.V_mir1.n2 152
R7326 bgr_0.V_mir1.n19 bgr_0.V_mir1.n18 152
R7327 bgr_0.V_mir1.n16 bgr_0.V_mir1.t22 120.501
R7328 bgr_0.V_mir1.n17 bgr_0.V_mir1.t13 120.501
R7329 bgr_0.V_mir1.n9 bgr_0.V_mir1.t17 120.501
R7330 bgr_0.V_mir1.n10 bgr_0.V_mir1.t11 120.501
R7331 bgr_0.V_mir1.n0 bgr_0.V_mir1.t18 120.501
R7332 bgr_0.V_mir1.n1 bgr_0.V_mir1.t7 120.501
R7333 bgr_0.V_mir1.n6 bgr_0.V_mir1.t16 48.0005
R7334 bgr_0.V_mir1.n6 bgr_0.V_mir1.t1 48.0005
R7335 bgr_0.V_mir1.n5 bgr_0.V_mir1.t0 48.0005
R7336 bgr_0.V_mir1.n5 bgr_0.V_mir1.t15 48.0005
R7337 bgr_0.V_mir1.n18 bgr_0.V_mir1.n17 40.7027
R7338 bgr_0.V_mir1.n11 bgr_0.V_mir1.n10 40.7027
R7339 bgr_0.V_mir1.n2 bgr_0.V_mir1.n1 40.7027
R7340 bgr_0.V_mir1.n12 bgr_0.V_mir1.t6 39.4005
R7341 bgr_0.V_mir1.n12 bgr_0.V_mir1.t12 39.4005
R7342 bgr_0.V_mir1.n3 bgr_0.V_mir1.t4 39.4005
R7343 bgr_0.V_mir1.n3 bgr_0.V_mir1.t8 39.4005
R7344 bgr_0.V_mir1.n20 bgr_0.V_mir1.t10 39.4005
R7345 bgr_0.V_mir1.t14 bgr_0.V_mir1.n20 39.4005
R7346 bgr_0.V_mir1.n15 bgr_0.V_mir1.n4 15.8005
R7347 bgr_0.V_mir1.n19 bgr_0.V_mir1.n15 15.8005
R7348 bgr_0.V_mir1.n14 bgr_0.V_mir1.n13 9.3005
R7349 bgr_0.V_mir1.n8 bgr_0.V_mir1.n7 5.8755
R7350 bgr_0.V_mir1.n15 bgr_0.V_mir1.n14 4.5005
R7351 bgr_0.V_mir1.n14 bgr_0.V_mir1.n8 0.78175
R7352 bgr_0.1st_Vout_1 bgr_0.1st_Vout_1.t13 354.854
R7353 bgr_0.1st_Vout_1.n5 bgr_0.1st_Vout_1.t21 346.8
R7354 bgr_0.1st_Vout_1.n20 bgr_0.1st_Vout_1.n19 339.522
R7355 bgr_0.1st_Vout_1.n7 bgr_0.1st_Vout_1.n6 339.522
R7356 bgr_0.1st_Vout_1.n15 bgr_0.1st_Vout_1.n14 335.022
R7357 bgr_0.1st_Vout_1.n11 bgr_0.1st_Vout_1.t9 275.909
R7358 bgr_0.1st_Vout_1.n11 bgr_0.1st_Vout_1.n10 227.909
R7359 bgr_0.1st_Vout_1.n13 bgr_0.1st_Vout_1.n12 222.034
R7360 bgr_0.1st_Vout_1.n17 bgr_0.1st_Vout_1.t22 184.097
R7361 bgr_0.1st_Vout_1.n17 bgr_0.1st_Vout_1.t32 184.097
R7362 bgr_0.1st_Vout_1.n8 bgr_0.1st_Vout_1.t16 184.097
R7363 bgr_0.1st_Vout_1.n8 bgr_0.1st_Vout_1.t36 184.097
R7364 bgr_0.1st_Vout_1.n18 bgr_0.1st_Vout_1.n17 166.05
R7365 bgr_0.1st_Vout_1.n9 bgr_0.1st_Vout_1.n8 166.05
R7366 bgr_0.1st_Vout_1.n5 bgr_0.1st_Vout_1.n4 54.2759
R7367 bgr_0.1st_Vout_1.n12 bgr_0.1st_Vout_1.t10 48.0005
R7368 bgr_0.1st_Vout_1.n12 bgr_0.1st_Vout_1.t7 48.0005
R7369 bgr_0.1st_Vout_1.n10 bgr_0.1st_Vout_1.t8 48.0005
R7370 bgr_0.1st_Vout_1.n10 bgr_0.1st_Vout_1.t6 48.0005
R7371 bgr_0.1st_Vout_1.n19 bgr_0.1st_Vout_1.t4 39.4005
R7372 bgr_0.1st_Vout_1.n19 bgr_0.1st_Vout_1.t2 39.4005
R7373 bgr_0.1st_Vout_1.n6 bgr_0.1st_Vout_1.t0 39.4005
R7374 bgr_0.1st_Vout_1.n6 bgr_0.1st_Vout_1.t3 39.4005
R7375 bgr_0.1st_Vout_1.n14 bgr_0.1st_Vout_1.t5 39.4005
R7376 bgr_0.1st_Vout_1.n14 bgr_0.1st_Vout_1.t1 39.4005
R7377 bgr_0.1st_Vout_1.n0 bgr_0.1st_Vout_1.t11 4.8295
R7378 bgr_0.1st_Vout_1.n0 bgr_0.1st_Vout_1.t29 4.8295
R7379 bgr_0.1st_Vout_1.n2 bgr_0.1st_Vout_1.t31 4.8295
R7380 bgr_0.1st_Vout_1.n1 bgr_0.1st_Vout_1.t20 4.8295
R7381 bgr_0.1st_Vout_1.n2 bgr_0.1st_Vout_1.t24 4.8295
R7382 bgr_0.1st_Vout_1.n2 bgr_0.1st_Vout_1.t14 4.8295
R7383 bgr_0.1st_Vout_1.n3 bgr_0.1st_Vout_1.t30 4.8295
R7384 bgr_0.1st_Vout_1.n3 bgr_0.1st_Vout_1.t18 4.8295
R7385 bgr_0.1st_Vout_1.n3 bgr_0.1st_Vout_1.t23 4.8295
R7386 bgr_0.1st_Vout_1.n0 bgr_0.1st_Vout_1.t15 4.5005
R7387 bgr_0.1st_Vout_1.n0 bgr_0.1st_Vout_1.t35 4.5005
R7388 bgr_0.1st_Vout_1.n2 bgr_0.1st_Vout_1.t34 4.5005
R7389 bgr_0.1st_Vout_1.n1 bgr_0.1st_Vout_1.t28 4.5005
R7390 bgr_0.1st_Vout_1.n2 bgr_0.1st_Vout_1.t27 4.5005
R7391 bgr_0.1st_Vout_1.n2 bgr_0.1st_Vout_1.t19 4.5005
R7392 bgr_0.1st_Vout_1.n3 bgr_0.1st_Vout_1.t33 4.5005
R7393 bgr_0.1st_Vout_1.n3 bgr_0.1st_Vout_1.t26 4.5005
R7394 bgr_0.1st_Vout_1.n3 bgr_0.1st_Vout_1.t25 4.5005
R7395 bgr_0.1st_Vout_1.n4 bgr_0.1st_Vout_1.t17 4.5005
R7396 bgr_0.1st_Vout_1.n4 bgr_0.1st_Vout_1.t12 4.5005
R7397 bgr_0.1st_Vout_1.n13 bgr_0.1st_Vout_1.n11 4.5005
R7398 bgr_0.1st_Vout_1.n16 bgr_0.1st_Vout_1.n15 4.5005
R7399 bgr_0.1st_Vout_1.n20 bgr_0.1st_Vout_1.n18 1.3755
R7400 bgr_0.1st_Vout_1.n16 bgr_0.1st_Vout_1.n9 1.3755
R7401 bgr_0.1st_Vout_1.n7 bgr_0.1st_Vout_1.n5 1.188
R7402 bgr_0.1st_Vout_1.n3 bgr_0.1st_Vout_1.n2 0.8935
R7403 bgr_0.1st_Vout_1.n2 bgr_0.1st_Vout_1.n0 0.8935
R7404 bgr_0.1st_Vout_1.n15 bgr_0.1st_Vout_1.n13 0.78175
R7405 bgr_0.1st_Vout_1.n4 bgr_0.1st_Vout_1.n3 0.6585
R7406 bgr_0.1st_Vout_1.n2 bgr_0.1st_Vout_1.n1 0.6585
R7407 bgr_0.1st_Vout_1.n18 bgr_0.1st_Vout_1.n16 0.6255
R7408 bgr_0.1st_Vout_1.n9 bgr_0.1st_Vout_1.n7 0.6255
R7409 bgr_0.1st_Vout_1 bgr_0.1st_Vout_1.n20 0.438
R7410 bgr_0.1st_Vout_2.n1 bgr_0.1st_Vout_2.t33 355.293
R7411 bgr_0.1st_Vout_2.n0 bgr_0.1st_Vout_2.t34 346.8
R7412 bgr_0.1st_Vout_2.n0 bgr_0.1st_Vout_2.n10 339.522
R7413 bgr_0.1st_Vout_2.n1 bgr_0.1st_Vout_2.n8 339.522
R7414 bgr_0.1st_Vout_2.n12 bgr_0.1st_Vout_2.n3 335.022
R7415 bgr_0.1st_Vout_2.n6 bgr_0.1st_Vout_2.t10 275.909
R7416 bgr_0.1st_Vout_2.n6 bgr_0.1st_Vout_2.n5 227.909
R7417 bgr_0.1st_Vout_2.n3 bgr_0.1st_Vout_2.n7 222.034
R7418 bgr_0.1st_Vout_2.n11 bgr_0.1st_Vout_2.t16 184.097
R7419 bgr_0.1st_Vout_2.n11 bgr_0.1st_Vout_2.t27 184.097
R7420 bgr_0.1st_Vout_2.n9 bgr_0.1st_Vout_2.t13 184.097
R7421 bgr_0.1st_Vout_2.n9 bgr_0.1st_Vout_2.t24 184.097
R7422 bgr_0.1st_Vout_2.n0 bgr_0.1st_Vout_2.n11 166.05
R7423 bgr_0.1st_Vout_2.n1 bgr_0.1st_Vout_2.n9 166.05
R7424 bgr_0.1st_Vout_2.n0 bgr_0.1st_Vout_2.n4 52.9634
R7425 bgr_0.1st_Vout_2.n7 bgr_0.1st_Vout_2.t6 48.0005
R7426 bgr_0.1st_Vout_2.n7 bgr_0.1st_Vout_2.t7 48.0005
R7427 bgr_0.1st_Vout_2.n5 bgr_0.1st_Vout_2.t5 48.0005
R7428 bgr_0.1st_Vout_2.n5 bgr_0.1st_Vout_2.t3 48.0005
R7429 bgr_0.1st_Vout_2.n10 bgr_0.1st_Vout_2.t8 39.4005
R7430 bgr_0.1st_Vout_2.n10 bgr_0.1st_Vout_2.t2 39.4005
R7431 bgr_0.1st_Vout_2.n8 bgr_0.1st_Vout_2.t4 39.4005
R7432 bgr_0.1st_Vout_2.n8 bgr_0.1st_Vout_2.t9 39.4005
R7433 bgr_0.1st_Vout_2.t0 bgr_0.1st_Vout_2.n12 39.4005
R7434 bgr_0.1st_Vout_2.n12 bgr_0.1st_Vout_2.t1 39.4005
R7435 bgr_0.1st_Vout_2.n3 bgr_0.1st_Vout_2.n1 5.28175
R7436 bgr_0.1st_Vout_2.n1 bgr_0.1st_Vout_2.n0 5.188
R7437 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.t17 4.8295
R7438 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.t35 4.8295
R7439 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.t11 4.8295
R7440 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.t26 4.8295
R7441 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.t30 4.8295
R7442 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.t19 4.8295
R7443 bgr_0.1st_Vout_2.n4 bgr_0.1st_Vout_2.t36 4.8295
R7444 bgr_0.1st_Vout_2.n4 bgr_0.1st_Vout_2.t25 4.8295
R7445 bgr_0.1st_Vout_2.n4 bgr_0.1st_Vout_2.t18 4.8295
R7446 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.t12 4.5005
R7447 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.t32 4.5005
R7448 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.t31 4.5005
R7449 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.t23 4.5005
R7450 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.t22 4.5005
R7451 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.t15 4.5005
R7452 bgr_0.1st_Vout_2.n4 bgr_0.1st_Vout_2.t29 4.5005
R7453 bgr_0.1st_Vout_2.n4 bgr_0.1st_Vout_2.t21 4.5005
R7454 bgr_0.1st_Vout_2.n4 bgr_0.1st_Vout_2.t28 4.5005
R7455 bgr_0.1st_Vout_2.n4 bgr_0.1st_Vout_2.t20 4.5005
R7456 bgr_0.1st_Vout_2.n4 bgr_0.1st_Vout_2.t14 4.5005
R7457 bgr_0.1st_Vout_2.n3 bgr_0.1st_Vout_2.n6 4.5005
R7458 bgr_0.1st_Vout_2.n4 bgr_0.1st_Vout_2.n2 3.1025
R7459 bgr_0.cap_res2.t20 bgr_0.cap_res2.t17 121.245
R7460 bgr_0.cap_res2.t12 bgr_0.cap_res2.t6 0.1603
R7461 bgr_0.cap_res2.t5 bgr_0.cap_res2.t0 0.1603
R7462 bgr_0.cap_res2.t10 bgr_0.cap_res2.t4 0.1603
R7463 bgr_0.cap_res2.t3 bgr_0.cap_res2.t19 0.1603
R7464 bgr_0.cap_res2.t18 bgr_0.cap_res2.t15 0.1603
R7465 bgr_0.cap_res2.n1 bgr_0.cap_res2.t2 0.159278
R7466 bgr_0.cap_res2.n2 bgr_0.cap_res2.t9 0.159278
R7467 bgr_0.cap_res2.n3 bgr_0.cap_res2.t16 0.159278
R7468 bgr_0.cap_res2.n4 bgr_0.cap_res2.t11 0.159278
R7469 bgr_0.cap_res2.n4 bgr_0.cap_res2.t14 0.1368
R7470 bgr_0.cap_res2.n4 bgr_0.cap_res2.t12 0.1368
R7471 bgr_0.cap_res2.n3 bgr_0.cap_res2.t8 0.1368
R7472 bgr_0.cap_res2.n3 bgr_0.cap_res2.t5 0.1368
R7473 bgr_0.cap_res2.n2 bgr_0.cap_res2.t13 0.1368
R7474 bgr_0.cap_res2.n2 bgr_0.cap_res2.t10 0.1368
R7475 bgr_0.cap_res2.n1 bgr_0.cap_res2.t7 0.1368
R7476 bgr_0.cap_res2.n1 bgr_0.cap_res2.t3 0.1368
R7477 bgr_0.cap_res2.n0 bgr_0.cap_res2.t1 0.1368
R7478 bgr_0.cap_res2.n0 bgr_0.cap_res2.t18 0.1368
R7479 bgr_0.cap_res2.t2 bgr_0.cap_res2.n0 0.00152174
R7480 bgr_0.cap_res2.t9 bgr_0.cap_res2.n1 0.00152174
R7481 bgr_0.cap_res2.t16 bgr_0.cap_res2.n2 0.00152174
R7482 bgr_0.cap_res2.t11 bgr_0.cap_res2.n3 0.00152174
R7483 bgr_0.cap_res2.t17 bgr_0.cap_res2.n4 0.00152174
R7484 two_stage_opamp_dummy_magic_14_0.Vb2.n25 two_stage_opamp_dummy_magic_14_0.Vb2.t31 650.273
R7485 two_stage_opamp_dummy_magic_14_0.Vb2.n27 two_stage_opamp_dummy_magic_14_0.Vb2.t0 650.273
R7486 two_stage_opamp_dummy_magic_14_0.Vb2.n4 two_stage_opamp_dummy_magic_14_0.Vb2.t12 611.739
R7487 two_stage_opamp_dummy_magic_14_0.Vb2.n0 two_stage_opamp_dummy_magic_14_0.Vb2.t22 611.739
R7488 two_stage_opamp_dummy_magic_14_0.Vb2.n13 two_stage_opamp_dummy_magic_14_0.Vb2.t13 611.739
R7489 two_stage_opamp_dummy_magic_14_0.Vb2.n9 two_stage_opamp_dummy_magic_14_0.Vb2.t23 611.739
R7490 two_stage_opamp_dummy_magic_14_0.Vb2.n28 two_stage_opamp_dummy_magic_14_0.Vb2.t27 445.423
R7491 two_stage_opamp_dummy_magic_14_0.Vb2.n4 two_stage_opamp_dummy_magic_14_0.Vb2.t17 421.75
R7492 two_stage_opamp_dummy_magic_14_0.Vb2.n5 two_stage_opamp_dummy_magic_14_0.Vb2.t24 421.75
R7493 two_stage_opamp_dummy_magic_14_0.Vb2.n6 two_stage_opamp_dummy_magic_14_0.Vb2.t28 421.75
R7494 two_stage_opamp_dummy_magic_14_0.Vb2.n7 two_stage_opamp_dummy_magic_14_0.Vb2.t29 421.75
R7495 two_stage_opamp_dummy_magic_14_0.Vb2.n0 two_stage_opamp_dummy_magic_14_0.Vb2.t26 421.75
R7496 two_stage_opamp_dummy_magic_14_0.Vb2.n1 two_stage_opamp_dummy_magic_14_0.Vb2.t19 421.75
R7497 two_stage_opamp_dummy_magic_14_0.Vb2.n2 two_stage_opamp_dummy_magic_14_0.Vb2.t14 421.75
R7498 two_stage_opamp_dummy_magic_14_0.Vb2.n3 two_stage_opamp_dummy_magic_14_0.Vb2.t32 421.75
R7499 two_stage_opamp_dummy_magic_14_0.Vb2.n13 two_stage_opamp_dummy_magic_14_0.Vb2.t18 421.75
R7500 two_stage_opamp_dummy_magic_14_0.Vb2.n14 two_stage_opamp_dummy_magic_14_0.Vb2.t25 421.75
R7501 two_stage_opamp_dummy_magic_14_0.Vb2.n15 two_stage_opamp_dummy_magic_14_0.Vb2.t21 421.75
R7502 two_stage_opamp_dummy_magic_14_0.Vb2.n16 two_stage_opamp_dummy_magic_14_0.Vb2.t30 421.75
R7503 two_stage_opamp_dummy_magic_14_0.Vb2.n9 two_stage_opamp_dummy_magic_14_0.Vb2.t16 421.75
R7504 two_stage_opamp_dummy_magic_14_0.Vb2.n10 two_stage_opamp_dummy_magic_14_0.Vb2.t20 421.75
R7505 two_stage_opamp_dummy_magic_14_0.Vb2.n11 two_stage_opamp_dummy_magic_14_0.Vb2.t15 421.75
R7506 two_stage_opamp_dummy_magic_14_0.Vb2.n12 two_stage_opamp_dummy_magic_14_0.Vb2.t11 421.75
R7507 two_stage_opamp_dummy_magic_14_0.Vb2.n30 two_stage_opamp_dummy_magic_14_0.Vb2.n17 169.352
R7508 two_stage_opamp_dummy_magic_14_0.Vb2.n5 two_stage_opamp_dummy_magic_14_0.Vb2.n4 167.094
R7509 two_stage_opamp_dummy_magic_14_0.Vb2.n6 two_stage_opamp_dummy_magic_14_0.Vb2.n5 167.094
R7510 two_stage_opamp_dummy_magic_14_0.Vb2.n7 two_stage_opamp_dummy_magic_14_0.Vb2.n6 167.094
R7511 two_stage_opamp_dummy_magic_14_0.Vb2.n1 two_stage_opamp_dummy_magic_14_0.Vb2.n0 167.094
R7512 two_stage_opamp_dummy_magic_14_0.Vb2.n2 two_stage_opamp_dummy_magic_14_0.Vb2.n1 167.094
R7513 two_stage_opamp_dummy_magic_14_0.Vb2.n3 two_stage_opamp_dummy_magic_14_0.Vb2.n2 167.094
R7514 two_stage_opamp_dummy_magic_14_0.Vb2.n14 two_stage_opamp_dummy_magic_14_0.Vb2.n13 167.094
R7515 two_stage_opamp_dummy_magic_14_0.Vb2.n15 two_stage_opamp_dummy_magic_14_0.Vb2.n14 167.094
R7516 two_stage_opamp_dummy_magic_14_0.Vb2.n16 two_stage_opamp_dummy_magic_14_0.Vb2.n15 167.094
R7517 two_stage_opamp_dummy_magic_14_0.Vb2.n10 two_stage_opamp_dummy_magic_14_0.Vb2.n9 167.094
R7518 two_stage_opamp_dummy_magic_14_0.Vb2.n11 two_stage_opamp_dummy_magic_14_0.Vb2.n10 167.094
R7519 two_stage_opamp_dummy_magic_14_0.Vb2.n12 two_stage_opamp_dummy_magic_14_0.Vb2.n11 167.094
R7520 two_stage_opamp_dummy_magic_14_0.Vb2 two_stage_opamp_dummy_magic_14_0.Vb2.n8 161.477
R7521 two_stage_opamp_dummy_magic_14_0.Vb2.n27 two_stage_opamp_dummy_magic_14_0.Vb2.n26 160.06
R7522 two_stage_opamp_dummy_magic_14_0.Vb2.n20 two_stage_opamp_dummy_magic_14_0.Vb2.n18 140.857
R7523 two_stage_opamp_dummy_magic_14_0.Vb2.n22 two_stage_opamp_dummy_magic_14_0.Vb2.n21 139.608
R7524 two_stage_opamp_dummy_magic_14_0.Vb2.n24 two_stage_opamp_dummy_magic_14_0.Vb2.n23 139.608
R7525 two_stage_opamp_dummy_magic_14_0.Vb2.n20 two_stage_opamp_dummy_magic_14_0.Vb2.n19 139.608
R7526 two_stage_opamp_dummy_magic_14_0.Vb2.n25 two_stage_opamp_dummy_magic_14_0.Vb2.n24 61.3349
R7527 two_stage_opamp_dummy_magic_14_0.Vb2.n8 two_stage_opamp_dummy_magic_14_0.Vb2.n7 49.8072
R7528 two_stage_opamp_dummy_magic_14_0.Vb2.n8 two_stage_opamp_dummy_magic_14_0.Vb2.n3 49.8072
R7529 two_stage_opamp_dummy_magic_14_0.Vb2.n17 two_stage_opamp_dummy_magic_14_0.Vb2.n16 49.8072
R7530 two_stage_opamp_dummy_magic_14_0.Vb2.n17 two_stage_opamp_dummy_magic_14_0.Vb2.n12 49.8072
R7531 two_stage_opamp_dummy_magic_14_0.Vb2.n18 two_stage_opamp_dummy_magic_14_0.Vb2.t7 24.0005
R7532 two_stage_opamp_dummy_magic_14_0.Vb2.n18 two_stage_opamp_dummy_magic_14_0.Vb2.t9 24.0005
R7533 two_stage_opamp_dummy_magic_14_0.Vb2.n21 two_stage_opamp_dummy_magic_14_0.Vb2.t5 24.0005
R7534 two_stage_opamp_dummy_magic_14_0.Vb2.n21 two_stage_opamp_dummy_magic_14_0.Vb2.t3 24.0005
R7535 two_stage_opamp_dummy_magic_14_0.Vb2.n23 two_stage_opamp_dummy_magic_14_0.Vb2.t10 24.0005
R7536 two_stage_opamp_dummy_magic_14_0.Vb2.n23 two_stage_opamp_dummy_magic_14_0.Vb2.t4 24.0005
R7537 two_stage_opamp_dummy_magic_14_0.Vb2.n19 two_stage_opamp_dummy_magic_14_0.Vb2.t6 24.0005
R7538 two_stage_opamp_dummy_magic_14_0.Vb2.n19 two_stage_opamp_dummy_magic_14_0.Vb2.t8 24.0005
R7539 two_stage_opamp_dummy_magic_14_0.Vb2.n30 two_stage_opamp_dummy_magic_14_0.Vb2.n29 12.8443
R7540 two_stage_opamp_dummy_magic_14_0.Vb2.n26 two_stage_opamp_dummy_magic_14_0.Vb2.t1 11.2576
R7541 two_stage_opamp_dummy_magic_14_0.Vb2.n26 two_stage_opamp_dummy_magic_14_0.Vb2.t2 11.2576
R7542 two_stage_opamp_dummy_magic_14_0.Vb2.n22 two_stage_opamp_dummy_magic_14_0.Vb2.n20 7.563
R7543 two_stage_opamp_dummy_magic_14_0.Vb2 two_stage_opamp_dummy_magic_14_0.Vb2.n30 7.2505
R7544 two_stage_opamp_dummy_magic_14_0.Vb2.n29 two_stage_opamp_dummy_magic_14_0.Vb2.n25 4.54113
R7545 two_stage_opamp_dummy_magic_14_0.Vb2.n28 two_stage_opamp_dummy_magic_14_0.Vb2.n27 2.84425
R7546 two_stage_opamp_dummy_magic_14_0.Vb2.n24 two_stage_opamp_dummy_magic_14_0.Vb2.n22 1.2505
R7547 two_stage_opamp_dummy_magic_14_0.Vb2.n29 two_stage_opamp_dummy_magic_14_0.Vb2.n28 0.928625
R7548 bgr_0.V_CUR_REF_REG.n4 bgr_0.V_CUR_REF_REG.n3 526.183
R7549 bgr_0.V_CUR_REF_REG.n2 bgr_0.V_CUR_REF_REG.n1 514.134
R7550 bgr_0.V_CUR_REF_REG.n5 bgr_0.V_CUR_REF_REG.n0 360.586
R7551 bgr_0.V_CUR_REF_REG.n1 bgr_0.V_CUR_REF_REG.t5 303.259
R7552 bgr_0.V_CUR_REF_REG.n5 bgr_0.V_CUR_REF_REG.n4 210.169
R7553 bgr_0.V_CUR_REF_REG.n1 bgr_0.V_CUR_REF_REG.t3 174.726
R7554 bgr_0.V_CUR_REF_REG.n2 bgr_0.V_CUR_REF_REG.t7 174.726
R7555 bgr_0.V_CUR_REF_REG.n3 bgr_0.V_CUR_REF_REG.t4 174.726
R7556 bgr_0.V_CUR_REF_REG.t0 bgr_0.V_CUR_REF_REG.n5 153.474
R7557 bgr_0.V_CUR_REF_REG.n3 bgr_0.V_CUR_REF_REG.n2 128.534
R7558 bgr_0.V_CUR_REF_REG.n4 bgr_0.V_CUR_REF_REG.t6 96.4005
R7559 bgr_0.V_CUR_REF_REG.n0 bgr_0.V_CUR_REF_REG.t1 39.4005
R7560 bgr_0.V_CUR_REF_REG.n0 bgr_0.V_CUR_REF_REG.t2 39.4005
R7561 bgr_0.V_p_2.n1 bgr_0.V_p_2.n2 229.562
R7562 bgr_0.V_p_2.n1 bgr_0.V_p_2.n5 228.939
R7563 bgr_0.V_p_2.n0 bgr_0.V_p_2.n4 228.939
R7564 bgr_0.V_p_2.n0 bgr_0.V_p_2.n3 228.939
R7565 bgr_0.V_p_2.n6 bgr_0.V_p_2.n1 228.938
R7566 bgr_0.V_p_2.n0 bgr_0.V_p_2.t10 98.7279
R7567 bgr_0.V_p_2.n5 bgr_0.V_p_2.t1 48.0005
R7568 bgr_0.V_p_2.n5 bgr_0.V_p_2.t5 48.0005
R7569 bgr_0.V_p_2.n4 bgr_0.V_p_2.t8 48.0005
R7570 bgr_0.V_p_2.n4 bgr_0.V_p_2.t0 48.0005
R7571 bgr_0.V_p_2.n3 bgr_0.V_p_2.t2 48.0005
R7572 bgr_0.V_p_2.n3 bgr_0.V_p_2.t6 48.0005
R7573 bgr_0.V_p_2.n2 bgr_0.V_p_2.t3 48.0005
R7574 bgr_0.V_p_2.n2 bgr_0.V_p_2.t7 48.0005
R7575 bgr_0.V_p_2.t9 bgr_0.V_p_2.n6 48.0005
R7576 bgr_0.V_p_2.n6 bgr_0.V_p_2.t4 48.0005
R7577 bgr_0.V_p_2.n1 bgr_0.V_p_2.n0 1.8755
R7578 a_7460_23988.t0 a_7460_23988.t1 178.133
R7579 two_stage_opamp_dummy_magic_14_0.V_err_gate.n2 two_stage_opamp_dummy_magic_14_0.V_err_gate.t6 479.322
R7580 two_stage_opamp_dummy_magic_14_0.V_err_gate.n2 two_stage_opamp_dummy_magic_14_0.V_err_gate.t8 479.322
R7581 two_stage_opamp_dummy_magic_14_0.V_err_gate.n6 two_stage_opamp_dummy_magic_14_0.V_err_gate.t9 479.322
R7582 two_stage_opamp_dummy_magic_14_0.V_err_gate.n6 two_stage_opamp_dummy_magic_14_0.V_err_gate.t7 479.322
R7583 two_stage_opamp_dummy_magic_14_0.V_err_gate.n3 two_stage_opamp_dummy_magic_14_0.V_err_gate.n1 178.625
R7584 two_stage_opamp_dummy_magic_14_0.V_err_gate.n5 two_stage_opamp_dummy_magic_14_0.V_err_gate.n4 177.987
R7585 two_stage_opamp_dummy_magic_14_0.V_err_gate two_stage_opamp_dummy_magic_14_0.V_err_gate.n0 175.013
R7586 two_stage_opamp_dummy_magic_14_0.V_err_gate.n3 two_stage_opamp_dummy_magic_14_0.V_err_gate.n2 165.8
R7587 two_stage_opamp_dummy_magic_14_0.V_err_gate two_stage_opamp_dummy_magic_14_0.V_err_gate.n6 165.8
R7588 two_stage_opamp_dummy_magic_14_0.V_err_gate.n0 two_stage_opamp_dummy_magic_14_0.V_err_gate.t1 24.0005
R7589 two_stage_opamp_dummy_magic_14_0.V_err_gate.n0 two_stage_opamp_dummy_magic_14_0.V_err_gate.t2 24.0005
R7590 two_stage_opamp_dummy_magic_14_0.V_err_gate.n4 two_stage_opamp_dummy_magic_14_0.V_err_gate.t3 15.7605
R7591 two_stage_opamp_dummy_magic_14_0.V_err_gate.n4 two_stage_opamp_dummy_magic_14_0.V_err_gate.t5 15.7605
R7592 two_stage_opamp_dummy_magic_14_0.V_err_gate.n1 two_stage_opamp_dummy_magic_14_0.V_err_gate.t0 15.7605
R7593 two_stage_opamp_dummy_magic_14_0.V_err_gate.n1 two_stage_opamp_dummy_magic_14_0.V_err_gate.t4 15.7605
R7594 two_stage_opamp_dummy_magic_14_0.V_err_gate two_stage_opamp_dummy_magic_14_0.V_err_gate.n5 1.76612
R7595 two_stage_opamp_dummy_magic_14_0.V_err_gate.n5 two_stage_opamp_dummy_magic_14_0.V_err_gate.n3 0.641125
R7596 two_stage_opamp_dummy_magic_14_0.V_err_mir_p two_stage_opamp_dummy_magic_14_0.V_err_mir_p.n0 187.315
R7597 two_stage_opamp_dummy_magic_14_0.V_err_mir_p two_stage_opamp_dummy_magic_14_0.V_err_mir_p.n1 177.755
R7598 two_stage_opamp_dummy_magic_14_0.V_err_mir_p.n0 two_stage_opamp_dummy_magic_14_0.V_err_mir_p.t3 15.7605
R7599 two_stage_opamp_dummy_magic_14_0.V_err_mir_p.n0 two_stage_opamp_dummy_magic_14_0.V_err_mir_p.t0 15.7605
R7600 two_stage_opamp_dummy_magic_14_0.V_err_mir_p.n1 two_stage_opamp_dummy_magic_14_0.V_err_mir_p.t1 15.7605
R7601 two_stage_opamp_dummy_magic_14_0.V_err_mir_p.n1 two_stage_opamp_dummy_magic_14_0.V_err_mir_p.t2 15.7605
R7602 two_stage_opamp_dummy_magic_14_0.Vb1.n17 two_stage_opamp_dummy_magic_14_0.Vb1.t11 449.868
R7603 two_stage_opamp_dummy_magic_14_0.Vb1.n13 two_stage_opamp_dummy_magic_14_0.Vb1.t15 449.868
R7604 two_stage_opamp_dummy_magic_14_0.Vb1.n8 two_stage_opamp_dummy_magic_14_0.Vb1.t10 449.868
R7605 two_stage_opamp_dummy_magic_14_0.Vb1.n4 two_stage_opamp_dummy_magic_14_0.Vb1.t14 449.868
R7606 two_stage_opamp_dummy_magic_14_0.Vb1.n2 two_stage_opamp_dummy_magic_14_0.Vb1.n0 339.961
R7607 two_stage_opamp_dummy_magic_14_0.Vb1.n2 two_stage_opamp_dummy_magic_14_0.Vb1.n1 339.272
R7608 two_stage_opamp_dummy_magic_14_0.Vb1.n17 two_stage_opamp_dummy_magic_14_0.Vb1.t20 273.134
R7609 two_stage_opamp_dummy_magic_14_0.Vb1.n18 two_stage_opamp_dummy_magic_14_0.Vb1.t9 273.134
R7610 two_stage_opamp_dummy_magic_14_0.Vb1.n19 two_stage_opamp_dummy_magic_14_0.Vb1.t18 273.134
R7611 two_stage_opamp_dummy_magic_14_0.Vb1.n20 two_stage_opamp_dummy_magic_14_0.Vb1.t6 273.134
R7612 two_stage_opamp_dummy_magic_14_0.Vb1.n16 two_stage_opamp_dummy_magic_14_0.Vb1.t23 273.134
R7613 two_stage_opamp_dummy_magic_14_0.Vb1.n15 two_stage_opamp_dummy_magic_14_0.Vb1.t7 273.134
R7614 two_stage_opamp_dummy_magic_14_0.Vb1.n14 two_stage_opamp_dummy_magic_14_0.Vb1.t16 273.134
R7615 two_stage_opamp_dummy_magic_14_0.Vb1.n13 two_stage_opamp_dummy_magic_14_0.Vb1.t25 273.134
R7616 two_stage_opamp_dummy_magic_14_0.Vb1.n8 two_stage_opamp_dummy_magic_14_0.Vb1.t19 273.134
R7617 two_stage_opamp_dummy_magic_14_0.Vb1.n9 two_stage_opamp_dummy_magic_14_0.Vb1.t8 273.134
R7618 two_stage_opamp_dummy_magic_14_0.Vb1.n10 two_stage_opamp_dummy_magic_14_0.Vb1.t17 273.134
R7619 two_stage_opamp_dummy_magic_14_0.Vb1.n11 two_stage_opamp_dummy_magic_14_0.Vb1.t13 273.134
R7620 two_stage_opamp_dummy_magic_14_0.Vb1.n7 two_stage_opamp_dummy_magic_14_0.Vb1.t22 273.134
R7621 two_stage_opamp_dummy_magic_14_0.Vb1.n6 two_stage_opamp_dummy_magic_14_0.Vb1.t12 273.134
R7622 two_stage_opamp_dummy_magic_14_0.Vb1.n5 two_stage_opamp_dummy_magic_14_0.Vb1.t21 273.134
R7623 two_stage_opamp_dummy_magic_14_0.Vb1.n4 two_stage_opamp_dummy_magic_14_0.Vb1.t24 273.134
R7624 two_stage_opamp_dummy_magic_14_0.Vb1.n20 two_stage_opamp_dummy_magic_14_0.Vb1.n19 176.733
R7625 two_stage_opamp_dummy_magic_14_0.Vb1.n19 two_stage_opamp_dummy_magic_14_0.Vb1.n18 176.733
R7626 two_stage_opamp_dummy_magic_14_0.Vb1.n18 two_stage_opamp_dummy_magic_14_0.Vb1.n17 176.733
R7627 two_stage_opamp_dummy_magic_14_0.Vb1.n14 two_stage_opamp_dummy_magic_14_0.Vb1.n13 176.733
R7628 two_stage_opamp_dummy_magic_14_0.Vb1.n15 two_stage_opamp_dummy_magic_14_0.Vb1.n14 176.733
R7629 two_stage_opamp_dummy_magic_14_0.Vb1.n16 two_stage_opamp_dummy_magic_14_0.Vb1.n15 176.733
R7630 two_stage_opamp_dummy_magic_14_0.Vb1.n11 two_stage_opamp_dummy_magic_14_0.Vb1.n10 176.733
R7631 two_stage_opamp_dummy_magic_14_0.Vb1.n10 two_stage_opamp_dummy_magic_14_0.Vb1.n9 176.733
R7632 two_stage_opamp_dummy_magic_14_0.Vb1.n9 two_stage_opamp_dummy_magic_14_0.Vb1.n8 176.733
R7633 two_stage_opamp_dummy_magic_14_0.Vb1.n5 two_stage_opamp_dummy_magic_14_0.Vb1.n4 176.733
R7634 two_stage_opamp_dummy_magic_14_0.Vb1.n6 two_stage_opamp_dummy_magic_14_0.Vb1.n5 176.733
R7635 two_stage_opamp_dummy_magic_14_0.Vb1.n7 two_stage_opamp_dummy_magic_14_0.Vb1.n6 176.733
R7636 two_stage_opamp_dummy_magic_14_0.Vb1.n3 two_stage_opamp_dummy_magic_14_0.Vb1.t2 175.553
R7637 two_stage_opamp_dummy_magic_14_0.Vb1.n22 two_stage_opamp_dummy_magic_14_0.Vb1.n12 172.207
R7638 two_stage_opamp_dummy_magic_14_0.Vb1.n22 two_stage_opamp_dummy_magic_14_0.Vb1.n21 165.8
R7639 two_stage_opamp_dummy_magic_14_0.Vb1.n3 two_stage_opamp_dummy_magic_14_0.Vb1.t1 62.3283
R7640 two_stage_opamp_dummy_magic_14_0.Vb1.n21 two_stage_opamp_dummy_magic_14_0.Vb1.n20 54.6272
R7641 two_stage_opamp_dummy_magic_14_0.Vb1.n21 two_stage_opamp_dummy_magic_14_0.Vb1.n16 54.6272
R7642 two_stage_opamp_dummy_magic_14_0.Vb1.n12 two_stage_opamp_dummy_magic_14_0.Vb1.n11 54.6272
R7643 two_stage_opamp_dummy_magic_14_0.Vb1.n12 two_stage_opamp_dummy_magic_14_0.Vb1.n7 54.6272
R7644 bgr_0.VB1_CUR_BIAS two_stage_opamp_dummy_magic_14_0.Vb1.n23 44.5005
R7645 two_stage_opamp_dummy_magic_14_0.Vb1.n1 two_stage_opamp_dummy_magic_14_0.Vb1.t3 39.4005
R7646 two_stage_opamp_dummy_magic_14_0.Vb1.n1 two_stage_opamp_dummy_magic_14_0.Vb1.t4 39.4005
R7647 two_stage_opamp_dummy_magic_14_0.Vb1.n0 two_stage_opamp_dummy_magic_14_0.Vb1.t5 39.4005
R7648 two_stage_opamp_dummy_magic_14_0.Vb1.n0 two_stage_opamp_dummy_magic_14_0.Vb1.t0 39.4005
R7649 two_stage_opamp_dummy_magic_14_0.Vb1.n23 two_stage_opamp_dummy_magic_14_0.Vb1.n3 21.8437
R7650 bgr_0.VB1_CUR_BIAS two_stage_opamp_dummy_magic_14_0.Vb1.n2 12.1255
R7651 two_stage_opamp_dummy_magic_14_0.Vb1.n23 two_stage_opamp_dummy_magic_14_0.Vb1.n22 6.92238
R7652 two_stage_opamp_dummy_magic_14_0.Y.n47 two_stage_opamp_dummy_magic_14_0.Y.t27 1172.87
R7653 two_stage_opamp_dummy_magic_14_0.Y.n43 two_stage_opamp_dummy_magic_14_0.Y.t33 1172.87
R7654 two_stage_opamp_dummy_magic_14_0.Y.n50 two_stage_opamp_dummy_magic_14_0.Y.t45 996.134
R7655 two_stage_opamp_dummy_magic_14_0.Y.n49 two_stage_opamp_dummy_magic_14_0.Y.t30 996.134
R7656 two_stage_opamp_dummy_magic_14_0.Y.n48 two_stage_opamp_dummy_magic_14_0.Y.t47 996.134
R7657 two_stage_opamp_dummy_magic_14_0.Y.n47 two_stage_opamp_dummy_magic_14_0.Y.t41 996.134
R7658 two_stage_opamp_dummy_magic_14_0.Y.n43 two_stage_opamp_dummy_magic_14_0.Y.t49 996.134
R7659 two_stage_opamp_dummy_magic_14_0.Y.n44 two_stage_opamp_dummy_magic_14_0.Y.t35 996.134
R7660 two_stage_opamp_dummy_magic_14_0.Y.n45 two_stage_opamp_dummy_magic_14_0.Y.t52 996.134
R7661 two_stage_opamp_dummy_magic_14_0.Y.n46 two_stage_opamp_dummy_magic_14_0.Y.t38 996.134
R7662 two_stage_opamp_dummy_magic_14_0.Y.n23 two_stage_opamp_dummy_magic_14_0.Y.t32 690.867
R7663 two_stage_opamp_dummy_magic_14_0.Y.n20 two_stage_opamp_dummy_magic_14_0.Y.t39 690.867
R7664 two_stage_opamp_dummy_magic_14_0.Y.n14 two_stage_opamp_dummy_magic_14_0.Y.t44 530.201
R7665 two_stage_opamp_dummy_magic_14_0.Y.n11 two_stage_opamp_dummy_magic_14_0.Y.t51 530.201
R7666 two_stage_opamp_dummy_magic_14_0.Y.n23 two_stage_opamp_dummy_magic_14_0.Y.t46 514.134
R7667 two_stage_opamp_dummy_magic_14_0.Y.n24 two_stage_opamp_dummy_magic_14_0.Y.t53 514.134
R7668 two_stage_opamp_dummy_magic_14_0.Y.n25 two_stage_opamp_dummy_magic_14_0.Y.t36 514.134
R7669 two_stage_opamp_dummy_magic_14_0.Y.n26 two_stage_opamp_dummy_magic_14_0.Y.t50 514.134
R7670 two_stage_opamp_dummy_magic_14_0.Y.n27 two_stage_opamp_dummy_magic_14_0.Y.t43 514.134
R7671 two_stage_opamp_dummy_magic_14_0.Y.n22 two_stage_opamp_dummy_magic_14_0.Y.t28 514.134
R7672 two_stage_opamp_dummy_magic_14_0.Y.n21 two_stage_opamp_dummy_magic_14_0.Y.t42 514.134
R7673 two_stage_opamp_dummy_magic_14_0.Y.n20 two_stage_opamp_dummy_magic_14_0.Y.t25 514.134
R7674 two_stage_opamp_dummy_magic_14_0.Y.n18 two_stage_opamp_dummy_magic_14_0.Y.t26 353.467
R7675 two_stage_opamp_dummy_magic_14_0.Y.n17 two_stage_opamp_dummy_magic_14_0.Y.t31 353.467
R7676 two_stage_opamp_dummy_magic_14_0.Y.n16 two_stage_opamp_dummy_magic_14_0.Y.t48 353.467
R7677 two_stage_opamp_dummy_magic_14_0.Y.n15 two_stage_opamp_dummy_magic_14_0.Y.t34 353.467
R7678 two_stage_opamp_dummy_magic_14_0.Y.n14 two_stage_opamp_dummy_magic_14_0.Y.t29 353.467
R7679 two_stage_opamp_dummy_magic_14_0.Y.n11 two_stage_opamp_dummy_magic_14_0.Y.t37 353.467
R7680 two_stage_opamp_dummy_magic_14_0.Y.n12 two_stage_opamp_dummy_magic_14_0.Y.t54 353.467
R7681 two_stage_opamp_dummy_magic_14_0.Y.n13 two_stage_opamp_dummy_magic_14_0.Y.t40 353.467
R7682 two_stage_opamp_dummy_magic_14_0.Y.n50 two_stage_opamp_dummy_magic_14_0.Y.n49 176.733
R7683 two_stage_opamp_dummy_magic_14_0.Y.n49 two_stage_opamp_dummy_magic_14_0.Y.n48 176.733
R7684 two_stage_opamp_dummy_magic_14_0.Y.n48 two_stage_opamp_dummy_magic_14_0.Y.n47 176.733
R7685 two_stage_opamp_dummy_magic_14_0.Y.n44 two_stage_opamp_dummy_magic_14_0.Y.n43 176.733
R7686 two_stage_opamp_dummy_magic_14_0.Y.n45 two_stage_opamp_dummy_magic_14_0.Y.n44 176.733
R7687 two_stage_opamp_dummy_magic_14_0.Y.n46 two_stage_opamp_dummy_magic_14_0.Y.n45 176.733
R7688 two_stage_opamp_dummy_magic_14_0.Y.n18 two_stage_opamp_dummy_magic_14_0.Y.n17 176.733
R7689 two_stage_opamp_dummy_magic_14_0.Y.n17 two_stage_opamp_dummy_magic_14_0.Y.n16 176.733
R7690 two_stage_opamp_dummy_magic_14_0.Y.n16 two_stage_opamp_dummy_magic_14_0.Y.n15 176.733
R7691 two_stage_opamp_dummy_magic_14_0.Y.n15 two_stage_opamp_dummy_magic_14_0.Y.n14 176.733
R7692 two_stage_opamp_dummy_magic_14_0.Y.n12 two_stage_opamp_dummy_magic_14_0.Y.n11 176.733
R7693 two_stage_opamp_dummy_magic_14_0.Y.n13 two_stage_opamp_dummy_magic_14_0.Y.n12 176.733
R7694 two_stage_opamp_dummy_magic_14_0.Y.n27 two_stage_opamp_dummy_magic_14_0.Y.n26 176.733
R7695 two_stage_opamp_dummy_magic_14_0.Y.n26 two_stage_opamp_dummy_magic_14_0.Y.n25 176.733
R7696 two_stage_opamp_dummy_magic_14_0.Y.n25 two_stage_opamp_dummy_magic_14_0.Y.n24 176.733
R7697 two_stage_opamp_dummy_magic_14_0.Y.n24 two_stage_opamp_dummy_magic_14_0.Y.n23 176.733
R7698 two_stage_opamp_dummy_magic_14_0.Y.n21 two_stage_opamp_dummy_magic_14_0.Y.n20 176.733
R7699 two_stage_opamp_dummy_magic_14_0.Y.n22 two_stage_opamp_dummy_magic_14_0.Y.n21 176.733
R7700 two_stage_opamp_dummy_magic_14_0.Y.n52 two_stage_opamp_dummy_magic_14_0.Y.n51 166.258
R7701 two_stage_opamp_dummy_magic_14_0.Y.n2 two_stage_opamp_dummy_magic_14_0.Y.n0 163.626
R7702 two_stage_opamp_dummy_magic_14_0.Y.n8 two_stage_opamp_dummy_magic_14_0.Y.n7 163.001
R7703 two_stage_opamp_dummy_magic_14_0.Y.n6 two_stage_opamp_dummy_magic_14_0.Y.n5 163.001
R7704 two_stage_opamp_dummy_magic_14_0.Y.n4 two_stage_opamp_dummy_magic_14_0.Y.n3 163.001
R7705 two_stage_opamp_dummy_magic_14_0.Y.n2 two_stage_opamp_dummy_magic_14_0.Y.n1 163.001
R7706 two_stage_opamp_dummy_magic_14_0.Y.n29 two_stage_opamp_dummy_magic_14_0.Y.n19 161.541
R7707 two_stage_opamp_dummy_magic_14_0.Y.n29 two_stage_opamp_dummy_magic_14_0.Y.n28 161.541
R7708 two_stage_opamp_dummy_magic_14_0.Y.n10 two_stage_opamp_dummy_magic_14_0.Y.n9 158.501
R7709 two_stage_opamp_dummy_magic_14_0.Y.n32 two_stage_opamp_dummy_magic_14_0.Y.n30 117.888
R7710 two_stage_opamp_dummy_magic_14_0.Y.n40 two_stage_opamp_dummy_magic_14_0.Y.n39 117.326
R7711 two_stage_opamp_dummy_magic_14_0.Y.n38 two_stage_opamp_dummy_magic_14_0.Y.n37 117.326
R7712 two_stage_opamp_dummy_magic_14_0.Y.n36 two_stage_opamp_dummy_magic_14_0.Y.n35 117.326
R7713 two_stage_opamp_dummy_magic_14_0.Y.n34 two_stage_opamp_dummy_magic_14_0.Y.n33 117.326
R7714 two_stage_opamp_dummy_magic_14_0.Y.n32 two_stage_opamp_dummy_magic_14_0.Y.n31 117.326
R7715 two_stage_opamp_dummy_magic_14_0.Y.n19 two_stage_opamp_dummy_magic_14_0.Y.n18 54.6272
R7716 two_stage_opamp_dummy_magic_14_0.Y.n19 two_stage_opamp_dummy_magic_14_0.Y.n13 54.6272
R7717 two_stage_opamp_dummy_magic_14_0.Y.n28 two_stage_opamp_dummy_magic_14_0.Y.n27 54.6272
R7718 two_stage_opamp_dummy_magic_14_0.Y.n28 two_stage_opamp_dummy_magic_14_0.Y.n22 54.6272
R7719 two_stage_opamp_dummy_magic_14_0.Y.n51 two_stage_opamp_dummy_magic_14_0.Y.n50 53.3126
R7720 two_stage_opamp_dummy_magic_14_0.Y.n51 two_stage_opamp_dummy_magic_14_0.Y.n46 53.3126
R7721 two_stage_opamp_dummy_magic_14_0.Y.t12 two_stage_opamp_dummy_magic_14_0.Y.n52 50.3031
R7722 two_stage_opamp_dummy_magic_14_0.Y.n42 two_stage_opamp_dummy_magic_14_0.Y.n10 16.8755
R7723 two_stage_opamp_dummy_magic_14_0.Y.n39 two_stage_opamp_dummy_magic_14_0.Y.t17 16.0005
R7724 two_stage_opamp_dummy_magic_14_0.Y.n39 two_stage_opamp_dummy_magic_14_0.Y.t24 16.0005
R7725 two_stage_opamp_dummy_magic_14_0.Y.n37 two_stage_opamp_dummy_magic_14_0.Y.t18 16.0005
R7726 two_stage_opamp_dummy_magic_14_0.Y.n37 two_stage_opamp_dummy_magic_14_0.Y.t19 16.0005
R7727 two_stage_opamp_dummy_magic_14_0.Y.n35 two_stage_opamp_dummy_magic_14_0.Y.t16 16.0005
R7728 two_stage_opamp_dummy_magic_14_0.Y.n35 two_stage_opamp_dummy_magic_14_0.Y.t22 16.0005
R7729 two_stage_opamp_dummy_magic_14_0.Y.n33 two_stage_opamp_dummy_magic_14_0.Y.t15 16.0005
R7730 two_stage_opamp_dummy_magic_14_0.Y.n33 two_stage_opamp_dummy_magic_14_0.Y.t20 16.0005
R7731 two_stage_opamp_dummy_magic_14_0.Y.n31 two_stage_opamp_dummy_magic_14_0.Y.t13 16.0005
R7732 two_stage_opamp_dummy_magic_14_0.Y.n31 two_stage_opamp_dummy_magic_14_0.Y.t14 16.0005
R7733 two_stage_opamp_dummy_magic_14_0.Y.n30 two_stage_opamp_dummy_magic_14_0.Y.t23 16.0005
R7734 two_stage_opamp_dummy_magic_14_0.Y.n30 two_stage_opamp_dummy_magic_14_0.Y.t21 16.0005
R7735 two_stage_opamp_dummy_magic_14_0.Y.n41 two_stage_opamp_dummy_magic_14_0.Y.n29 11.9693
R7736 two_stage_opamp_dummy_magic_14_0.Y.n9 two_stage_opamp_dummy_magic_14_0.Y.t7 11.2576
R7737 two_stage_opamp_dummy_magic_14_0.Y.n9 two_stage_opamp_dummy_magic_14_0.Y.t0 11.2576
R7738 two_stage_opamp_dummy_magic_14_0.Y.n7 two_stage_opamp_dummy_magic_14_0.Y.t3 11.2576
R7739 two_stage_opamp_dummy_magic_14_0.Y.n7 two_stage_opamp_dummy_magic_14_0.Y.t11 11.2576
R7740 two_stage_opamp_dummy_magic_14_0.Y.n5 two_stage_opamp_dummy_magic_14_0.Y.t4 11.2576
R7741 two_stage_opamp_dummy_magic_14_0.Y.n5 two_stage_opamp_dummy_magic_14_0.Y.t8 11.2576
R7742 two_stage_opamp_dummy_magic_14_0.Y.n3 two_stage_opamp_dummy_magic_14_0.Y.t5 11.2576
R7743 two_stage_opamp_dummy_magic_14_0.Y.n3 two_stage_opamp_dummy_magic_14_0.Y.t2 11.2576
R7744 two_stage_opamp_dummy_magic_14_0.Y.n1 two_stage_opamp_dummy_magic_14_0.Y.t10 11.2576
R7745 two_stage_opamp_dummy_magic_14_0.Y.n1 two_stage_opamp_dummy_magic_14_0.Y.t9 11.2576
R7746 two_stage_opamp_dummy_magic_14_0.Y.n0 two_stage_opamp_dummy_magic_14_0.Y.t1 11.2576
R7747 two_stage_opamp_dummy_magic_14_0.Y.n0 two_stage_opamp_dummy_magic_14_0.Y.t6 11.2576
R7748 two_stage_opamp_dummy_magic_14_0.Y.n52 two_stage_opamp_dummy_magic_14_0.Y.n42 7.09425
R7749 two_stage_opamp_dummy_magic_14_0.Y.n41 two_stage_opamp_dummy_magic_14_0.Y.n40 6.3755
R7750 two_stage_opamp_dummy_magic_14_0.Y.n10 two_stage_opamp_dummy_magic_14_0.Y.n8 5.1255
R7751 two_stage_opamp_dummy_magic_14_0.Y.n42 two_stage_opamp_dummy_magic_14_0.Y.n41 1.3755
R7752 two_stage_opamp_dummy_magic_14_0.Y.n4 two_stage_opamp_dummy_magic_14_0.Y.n2 0.6255
R7753 two_stage_opamp_dummy_magic_14_0.Y.n6 two_stage_opamp_dummy_magic_14_0.Y.n4 0.6255
R7754 two_stage_opamp_dummy_magic_14_0.Y.n8 two_stage_opamp_dummy_magic_14_0.Y.n6 0.6255
R7755 two_stage_opamp_dummy_magic_14_0.Y.n34 two_stage_opamp_dummy_magic_14_0.Y.n32 0.563
R7756 two_stage_opamp_dummy_magic_14_0.Y.n36 two_stage_opamp_dummy_magic_14_0.Y.n34 0.563
R7757 two_stage_opamp_dummy_magic_14_0.Y.n38 two_stage_opamp_dummy_magic_14_0.Y.n36 0.563
R7758 two_stage_opamp_dummy_magic_14_0.Y.n40 two_stage_opamp_dummy_magic_14_0.Y.n38 0.563
R7759 two_stage_opamp_dummy_magic_14_0.VD2.n16 two_stage_opamp_dummy_magic_14_0.VD2.n14 146.47
R7760 two_stage_opamp_dummy_magic_14_0.VD2.n11 two_stage_opamp_dummy_magic_14_0.VD2.n9 146.47
R7761 two_stage_opamp_dummy_magic_14_0.VD2.n18 two_stage_opamp_dummy_magic_14_0.VD2.n17 145.906
R7762 two_stage_opamp_dummy_magic_14_0.VD2.n16 two_stage_opamp_dummy_magic_14_0.VD2.n15 145.906
R7763 two_stage_opamp_dummy_magic_14_0.VD2.n13 two_stage_opamp_dummy_magic_14_0.VD2.n12 145.906
R7764 two_stage_opamp_dummy_magic_14_0.VD2.n11 two_stage_opamp_dummy_magic_14_0.VD2.n10 145.906
R7765 two_stage_opamp_dummy_magic_14_0.VD2.n6 two_stage_opamp_dummy_magic_14_0.VD2.n4 114.719
R7766 two_stage_opamp_dummy_magic_14_0.VD2.n3 two_stage_opamp_dummy_magic_14_0.VD2.n1 114.719
R7767 two_stage_opamp_dummy_magic_14_0.VD2.n6 two_stage_opamp_dummy_magic_14_0.VD2.n5 114.156
R7768 two_stage_opamp_dummy_magic_14_0.VD2.n3 two_stage_opamp_dummy_magic_14_0.VD2.n2 114.156
R7769 two_stage_opamp_dummy_magic_14_0.VD2.n8 two_stage_opamp_dummy_magic_14_0.VD2.n0 109.656
R7770 two_stage_opamp_dummy_magic_14_0.VD2.n5 two_stage_opamp_dummy_magic_14_0.VD2.t6 16.0005
R7771 two_stage_opamp_dummy_magic_14_0.VD2.n5 two_stage_opamp_dummy_magic_14_0.VD2.t10 16.0005
R7772 two_stage_opamp_dummy_magic_14_0.VD2.n4 two_stage_opamp_dummy_magic_14_0.VD2.t5 16.0005
R7773 two_stage_opamp_dummy_magic_14_0.VD2.n4 two_stage_opamp_dummy_magic_14_0.VD2.t9 16.0005
R7774 two_stage_opamp_dummy_magic_14_0.VD2.n2 two_stage_opamp_dummy_magic_14_0.VD2.t7 16.0005
R7775 two_stage_opamp_dummy_magic_14_0.VD2.n2 two_stage_opamp_dummy_magic_14_0.VD2.t11 16.0005
R7776 two_stage_opamp_dummy_magic_14_0.VD2.n1 two_stage_opamp_dummy_magic_14_0.VD2.t8 16.0005
R7777 two_stage_opamp_dummy_magic_14_0.VD2.n1 two_stage_opamp_dummy_magic_14_0.VD2.t3 16.0005
R7778 two_stage_opamp_dummy_magic_14_0.VD2.n17 two_stage_opamp_dummy_magic_14_0.VD2.t18 16.0005
R7779 two_stage_opamp_dummy_magic_14_0.VD2.n17 two_stage_opamp_dummy_magic_14_0.VD2.t2 16.0005
R7780 two_stage_opamp_dummy_magic_14_0.VD2.n15 two_stage_opamp_dummy_magic_14_0.VD2.t0 16.0005
R7781 two_stage_opamp_dummy_magic_14_0.VD2.n15 two_stage_opamp_dummy_magic_14_0.VD2.t21 16.0005
R7782 two_stage_opamp_dummy_magic_14_0.VD2.n14 two_stage_opamp_dummy_magic_14_0.VD2.t16 16.0005
R7783 two_stage_opamp_dummy_magic_14_0.VD2.n14 two_stage_opamp_dummy_magic_14_0.VD2.t14 16.0005
R7784 two_stage_opamp_dummy_magic_14_0.VD2.n12 two_stage_opamp_dummy_magic_14_0.VD2.t1 16.0005
R7785 two_stage_opamp_dummy_magic_14_0.VD2.n12 two_stage_opamp_dummy_magic_14_0.VD2.t19 16.0005
R7786 two_stage_opamp_dummy_magic_14_0.VD2.n10 two_stage_opamp_dummy_magic_14_0.VD2.t20 16.0005
R7787 two_stage_opamp_dummy_magic_14_0.VD2.n10 two_stage_opamp_dummy_magic_14_0.VD2.t17 16.0005
R7788 two_stage_opamp_dummy_magic_14_0.VD2.n9 two_stage_opamp_dummy_magic_14_0.VD2.t13 16.0005
R7789 two_stage_opamp_dummy_magic_14_0.VD2.n9 two_stage_opamp_dummy_magic_14_0.VD2.t15 16.0005
R7790 two_stage_opamp_dummy_magic_14_0.VD2.n0 two_stage_opamp_dummy_magic_14_0.VD2.t4 16.0005
R7791 two_stage_opamp_dummy_magic_14_0.VD2.n0 two_stage_opamp_dummy_magic_14_0.VD2.t12 16.0005
R7792 two_stage_opamp_dummy_magic_14_0.VD2 two_stage_opamp_dummy_magic_14_0.VD2.n19 4.64633
R7793 two_stage_opamp_dummy_magic_14_0.VD2.n8 two_stage_opamp_dummy_magic_14_0.VD2.n7 4.5005
R7794 two_stage_opamp_dummy_magic_14_0.VD2.n7 two_stage_opamp_dummy_magic_14_0.VD2.n6 0.563
R7795 two_stage_opamp_dummy_magic_14_0.VD2.n7 two_stage_opamp_dummy_magic_14_0.VD2.n3 0.563
R7796 two_stage_opamp_dummy_magic_14_0.VD2.n18 two_stage_opamp_dummy_magic_14_0.VD2.n16 0.563
R7797 two_stage_opamp_dummy_magic_14_0.VD2.n13 two_stage_opamp_dummy_magic_14_0.VD2.n11 0.563
R7798 two_stage_opamp_dummy_magic_14_0.VD2.n19 two_stage_opamp_dummy_magic_14_0.VD2.n18 0.234875
R7799 two_stage_opamp_dummy_magic_14_0.VD2.n19 two_stage_opamp_dummy_magic_14_0.VD2.n13 0.234875
R7800 two_stage_opamp_dummy_magic_14_0.VD2 two_stage_opamp_dummy_magic_14_0.VD2.n8 0.09425
R7801 bgr_0.PFET_GATE_10uA.n4 bgr_0.PFET_GATE_10uA.t13 369.534
R7802 bgr_0.PFET_GATE_10uA.n3 bgr_0.PFET_GATE_10uA.t12 369.534
R7803 bgr_0.PFET_GATE_10uA.n23 bgr_0.PFET_GATE_10uA.t29 369.534
R7804 bgr_0.PFET_GATE_10uA.n18 bgr_0.PFET_GATE_10uA.t17 369.534
R7805 bgr_0.PFET_GATE_10uA.n1 bgr_0.PFET_GATE_10uA.t21 369.534
R7806 bgr_0.PFET_GATE_10uA.n0 bgr_0.PFET_GATE_10uA.t20 369.534
R7807 bgr_0.PFET_GATE_10uA.n8 bgr_0.PFET_GATE_10uA.n6 341.397
R7808 bgr_0.PFET_GATE_10uA.n10 bgr_0.PFET_GATE_10uA.n9 339.272
R7809 bgr_0.PFET_GATE_10uA.n8 bgr_0.PFET_GATE_10uA.n7 339.272
R7810 bgr_0.PFET_GATE_10uA.n13 bgr_0.PFET_GATE_10uA.n12 334.772
R7811 bgr_0.PFET_GATE_10uA.n14 bgr_0.PFET_GATE_10uA.t14 238.322
R7812 bgr_0.PFET_GATE_10uA.n14 bgr_0.PFET_GATE_10uA.t27 238.322
R7813 bgr_0.PFET_GATE_10uA.n4 bgr_0.PFET_GATE_10uA.t26 192.8
R7814 bgr_0.PFET_GATE_10uA.n3 bgr_0.PFET_GATE_10uA.t19 192.8
R7815 bgr_0.PFET_GATE_10uA.n25 bgr_0.PFET_GATE_10uA.t16 192.8
R7816 bgr_0.PFET_GATE_10uA.n24 bgr_0.PFET_GATE_10uA.t23 192.8
R7817 bgr_0.PFET_GATE_10uA.n23 bgr_0.PFET_GATE_10uA.t22 192.8
R7818 bgr_0.PFET_GATE_10uA.n18 bgr_0.PFET_GATE_10uA.t24 192.8
R7819 bgr_0.PFET_GATE_10uA.n19 bgr_0.PFET_GATE_10uA.t10 192.8
R7820 bgr_0.PFET_GATE_10uA.n20 bgr_0.PFET_GATE_10uA.t18 192.8
R7821 bgr_0.PFET_GATE_10uA.n21 bgr_0.PFET_GATE_10uA.t25 192.8
R7822 bgr_0.PFET_GATE_10uA.n22 bgr_0.PFET_GATE_10uA.t11 192.8
R7823 bgr_0.PFET_GATE_10uA.n1 bgr_0.PFET_GATE_10uA.t15 192.8
R7824 bgr_0.PFET_GATE_10uA.n0 bgr_0.PFET_GATE_10uA.t28 192.8
R7825 bgr_0.PFET_GATE_10uA.n25 bgr_0.PFET_GATE_10uA.n24 176.733
R7826 bgr_0.PFET_GATE_10uA.n24 bgr_0.PFET_GATE_10uA.n23 176.733
R7827 bgr_0.PFET_GATE_10uA.n19 bgr_0.PFET_GATE_10uA.n18 176.733
R7828 bgr_0.PFET_GATE_10uA.n20 bgr_0.PFET_GATE_10uA.n19 176.733
R7829 bgr_0.PFET_GATE_10uA.n21 bgr_0.PFET_GATE_10uA.n20 176.733
R7830 bgr_0.PFET_GATE_10uA.n22 bgr_0.PFET_GATE_10uA.n21 176.733
R7831 bgr_0.PFET_GATE_10uA bgr_0.PFET_GATE_10uA.n2 171.321
R7832 bgr_0.PFET_GATE_10uA.n17 bgr_0.PFET_GATE_10uA.n5 168.166
R7833 bgr_0.PFET_GATE_10uA.n15 bgr_0.PFET_GATE_10uA.n14 167.519
R7834 bgr_0.PFET_GATE_10uA bgr_0.PFET_GATE_10uA.n26 166.071
R7835 bgr_0.PFET_GATE_10uA.n15 bgr_0.PFET_GATE_10uA.t6 137.48
R7836 bgr_0.PFET_GATE_10uA.n11 bgr_0.PFET_GATE_10uA.t7 100.635
R7837 bgr_0.PFET_GATE_10uA.n5 bgr_0.PFET_GATE_10uA.n4 56.2338
R7838 bgr_0.PFET_GATE_10uA.n5 bgr_0.PFET_GATE_10uA.n3 56.2338
R7839 bgr_0.PFET_GATE_10uA.n26 bgr_0.PFET_GATE_10uA.n25 56.2338
R7840 bgr_0.PFET_GATE_10uA.n26 bgr_0.PFET_GATE_10uA.n22 56.2338
R7841 bgr_0.PFET_GATE_10uA.n2 bgr_0.PFET_GATE_10uA.n1 56.2338
R7842 bgr_0.PFET_GATE_10uA.n2 bgr_0.PFET_GATE_10uA.n0 56.2338
R7843 bgr_0.PFET_GATE_10uA.n12 bgr_0.PFET_GATE_10uA.t9 39.4005
R7844 bgr_0.PFET_GATE_10uA.n12 bgr_0.PFET_GATE_10uA.t1 39.4005
R7845 bgr_0.PFET_GATE_10uA.n9 bgr_0.PFET_GATE_10uA.t3 39.4005
R7846 bgr_0.PFET_GATE_10uA.n9 bgr_0.PFET_GATE_10uA.t5 39.4005
R7847 bgr_0.PFET_GATE_10uA.n7 bgr_0.PFET_GATE_10uA.t2 39.4005
R7848 bgr_0.PFET_GATE_10uA.n7 bgr_0.PFET_GATE_10uA.t4 39.4005
R7849 bgr_0.PFET_GATE_10uA.n6 bgr_0.PFET_GATE_10uA.t0 39.4005
R7850 bgr_0.PFET_GATE_10uA.n6 bgr_0.PFET_GATE_10uA.t8 39.4005
R7851 bgr_0.PFET_GATE_10uA.n17 bgr_0.PFET_GATE_10uA.n16 27.5005
R7852 bgr_0.PFET_GATE_10uA.n16 bgr_0.PFET_GATE_10uA.n13 9.53175
R7853 bgr_0.PFET_GATE_10uA.n13 bgr_0.PFET_GATE_10uA.n11 4.5005
R7854 bgr_0.PFET_GATE_10uA bgr_0.PFET_GATE_10uA.n17 2.34425
R7855 bgr_0.PFET_GATE_10uA.n10 bgr_0.PFET_GATE_10uA.n8 2.1255
R7856 bgr_0.PFET_GATE_10uA.n11 bgr_0.PFET_GATE_10uA.n10 2.1255
R7857 bgr_0.PFET_GATE_10uA.n16 bgr_0.PFET_GATE_10uA.n15 1.688
R7858 VIN-.n9 VIN-.t1 490.075
R7859 VIN-.n4 VIN-.t3 449.868
R7860 VIN-.n0 VIN-.t6 449.868
R7861 VIN-.n4 VIN-.t8 273.134
R7862 VIN-.n5 VIN-.t2 273.134
R7863 VIN-.n6 VIN-.t7 273.134
R7864 VIN-.n7 VIN-.t5 273.134
R7865 VIN-.n3 VIN-.t10 273.134
R7866 VIN-.n2 VIN-.t4 273.134
R7867 VIN-.n1 VIN-.t9 273.134
R7868 VIN-.n0 VIN-.t0 273.134
R7869 VIN-.n7 VIN-.n6 176.733
R7870 VIN-.n6 VIN-.n5 176.733
R7871 VIN-.n5 VIN-.n4 176.733
R7872 VIN-.n1 VIN-.n0 176.733
R7873 VIN-.n2 VIN-.n1 176.733
R7874 VIN-.n3 VIN-.n2 176.733
R7875 VIN-.n9 VIN-.n8 165.8
R7876 VIN-.n8 VIN-.n7 56.2338
R7877 VIN-.n8 VIN-.n3 56.2338
R7878 VIN- VIN-.n9 2.14112
R7879 two_stage_opamp_dummy_magic_14_0.VD1.n3 two_stage_opamp_dummy_magic_14_0.VD1.n1 146.47
R7880 two_stage_opamp_dummy_magic_14_0.VD1.n18 two_stage_opamp_dummy_magic_14_0.VD1.n0 146.47
R7881 two_stage_opamp_dummy_magic_14_0.VD1.n17 two_stage_opamp_dummy_magic_14_0.VD1.n16 145.906
R7882 two_stage_opamp_dummy_magic_14_0.VD1.n5 two_stage_opamp_dummy_magic_14_0.VD1.n4 145.906
R7883 two_stage_opamp_dummy_magic_14_0.VD1.n3 two_stage_opamp_dummy_magic_14_0.VD1.n2 145.906
R7884 two_stage_opamp_dummy_magic_14_0.VD1.n19 two_stage_opamp_dummy_magic_14_0.VD1.n18 145.906
R7885 two_stage_opamp_dummy_magic_14_0.VD1.n12 two_stage_opamp_dummy_magic_14_0.VD1.n10 114.719
R7886 two_stage_opamp_dummy_magic_14_0.VD1.n9 two_stage_opamp_dummy_magic_14_0.VD1.n7 114.719
R7887 two_stage_opamp_dummy_magic_14_0.VD1.n12 two_stage_opamp_dummy_magic_14_0.VD1.n11 114.156
R7888 two_stage_opamp_dummy_magic_14_0.VD1.n9 two_stage_opamp_dummy_magic_14_0.VD1.n8 114.156
R7889 two_stage_opamp_dummy_magic_14_0.VD1.n14 two_stage_opamp_dummy_magic_14_0.VD1.n6 109.656
R7890 two_stage_opamp_dummy_magic_14_0.VD1.n16 two_stage_opamp_dummy_magic_14_0.VD1.t6 16.0005
R7891 two_stage_opamp_dummy_magic_14_0.VD1.n16 two_stage_opamp_dummy_magic_14_0.VD1.t0 16.0005
R7892 two_stage_opamp_dummy_magic_14_0.VD1.n11 two_stage_opamp_dummy_magic_14_0.VD1.t14 16.0005
R7893 two_stage_opamp_dummy_magic_14_0.VD1.n11 two_stage_opamp_dummy_magic_14_0.VD1.t19 16.0005
R7894 two_stage_opamp_dummy_magic_14_0.VD1.n10 two_stage_opamp_dummy_magic_14_0.VD1.t13 16.0005
R7895 two_stage_opamp_dummy_magic_14_0.VD1.n10 two_stage_opamp_dummy_magic_14_0.VD1.t18 16.0005
R7896 two_stage_opamp_dummy_magic_14_0.VD1.n8 two_stage_opamp_dummy_magic_14_0.VD1.t12 16.0005
R7897 two_stage_opamp_dummy_magic_14_0.VD1.n8 two_stage_opamp_dummy_magic_14_0.VD1.t17 16.0005
R7898 two_stage_opamp_dummy_magic_14_0.VD1.n7 two_stage_opamp_dummy_magic_14_0.VD1.t15 16.0005
R7899 two_stage_opamp_dummy_magic_14_0.VD1.n7 two_stage_opamp_dummy_magic_14_0.VD1.t10 16.0005
R7900 two_stage_opamp_dummy_magic_14_0.VD1.n6 two_stage_opamp_dummy_magic_14_0.VD1.t11 16.0005
R7901 two_stage_opamp_dummy_magic_14_0.VD1.n6 two_stage_opamp_dummy_magic_14_0.VD1.t16 16.0005
R7902 two_stage_opamp_dummy_magic_14_0.VD1.n4 two_stage_opamp_dummy_magic_14_0.VD1.t5 16.0005
R7903 two_stage_opamp_dummy_magic_14_0.VD1.n4 two_stage_opamp_dummy_magic_14_0.VD1.t3 16.0005
R7904 two_stage_opamp_dummy_magic_14_0.VD1.n2 two_stage_opamp_dummy_magic_14_0.VD1.t8 16.0005
R7905 two_stage_opamp_dummy_magic_14_0.VD1.n2 two_stage_opamp_dummy_magic_14_0.VD1.t2 16.0005
R7906 two_stage_opamp_dummy_magic_14_0.VD1.n1 two_stage_opamp_dummy_magic_14_0.VD1.t7 16.0005
R7907 two_stage_opamp_dummy_magic_14_0.VD1.n1 two_stage_opamp_dummy_magic_14_0.VD1.t21 16.0005
R7908 two_stage_opamp_dummy_magic_14_0.VD1.n0 two_stage_opamp_dummy_magic_14_0.VD1.t20 16.0005
R7909 two_stage_opamp_dummy_magic_14_0.VD1.n0 two_stage_opamp_dummy_magic_14_0.VD1.t4 16.0005
R7910 two_stage_opamp_dummy_magic_14_0.VD1.t9 two_stage_opamp_dummy_magic_14_0.VD1.n19 16.0005
R7911 two_stage_opamp_dummy_magic_14_0.VD1.n19 two_stage_opamp_dummy_magic_14_0.VD1.t1 16.0005
R7912 two_stage_opamp_dummy_magic_14_0.VD1.n15 two_stage_opamp_dummy_magic_14_0.VD1.n14 4.74008
R7913 two_stage_opamp_dummy_magic_14_0.VD1.n14 two_stage_opamp_dummy_magic_14_0.VD1.n13 4.5005
R7914 two_stage_opamp_dummy_magic_14_0.VD1.n13 two_stage_opamp_dummy_magic_14_0.VD1.n12 0.563
R7915 two_stage_opamp_dummy_magic_14_0.VD1.n13 two_stage_opamp_dummy_magic_14_0.VD1.n9 0.563
R7916 two_stage_opamp_dummy_magic_14_0.VD1.n5 two_stage_opamp_dummy_magic_14_0.VD1.n3 0.563
R7917 two_stage_opamp_dummy_magic_14_0.VD1.n18 two_stage_opamp_dummy_magic_14_0.VD1.n17 0.563
R7918 two_stage_opamp_dummy_magic_14_0.VD1.n15 two_stage_opamp_dummy_magic_14_0.VD1.n5 0.234875
R7919 two_stage_opamp_dummy_magic_14_0.VD1.n17 two_stage_opamp_dummy_magic_14_0.VD1.n15 0.234875
R7920 bgr_0.cap_res1.t20 bgr_0.cap_res1.t9 121.245
R7921 bgr_0.cap_res1.t15 bgr_0.cap_res1.t18 0.1603
R7922 bgr_0.cap_res1.t8 bgr_0.cap_res1.t14 0.1603
R7923 bgr_0.cap_res1.t13 bgr_0.cap_res1.t17 0.1603
R7924 bgr_0.cap_res1.t6 bgr_0.cap_res1.t12 0.1603
R7925 bgr_0.cap_res1.t0 bgr_0.cap_res1.t5 0.1603
R7926 bgr_0.cap_res1.n1 bgr_0.cap_res1.t16 0.159278
R7927 bgr_0.cap_res1.n2 bgr_0.cap_res1.t1 0.159278
R7928 bgr_0.cap_res1.n3 bgr_0.cap_res1.t7 0.159278
R7929 bgr_0.cap_res1.n4 bgr_0.cap_res1.t2 0.159278
R7930 bgr_0.cap_res1.n4 bgr_0.cap_res1.t15 0.1368
R7931 bgr_0.cap_res1.n4 bgr_0.cap_res1.t11 0.1368
R7932 bgr_0.cap_res1.n3 bgr_0.cap_res1.t8 0.1368
R7933 bgr_0.cap_res1.n3 bgr_0.cap_res1.t4 0.1368
R7934 bgr_0.cap_res1.n2 bgr_0.cap_res1.t13 0.1368
R7935 bgr_0.cap_res1.n2 bgr_0.cap_res1.t10 0.1368
R7936 bgr_0.cap_res1.n1 bgr_0.cap_res1.t6 0.1368
R7937 bgr_0.cap_res1.n1 bgr_0.cap_res1.t3 0.1368
R7938 bgr_0.cap_res1.n0 bgr_0.cap_res1.t0 0.1368
R7939 bgr_0.cap_res1.n0 bgr_0.cap_res1.t19 0.1368
R7940 bgr_0.cap_res1.t16 bgr_0.cap_res1.n0 0.00152174
R7941 bgr_0.cap_res1.t1 bgr_0.cap_res1.n1 0.00152174
R7942 bgr_0.cap_res1.t7 bgr_0.cap_res1.n2 0.00152174
R7943 bgr_0.cap_res1.t2 bgr_0.cap_res1.n3 0.00152174
R7944 bgr_0.cap_res1.t9 bgr_0.cap_res1.n4 0.00152174
R7945 bgr_0.V_mir2.n20 bgr_0.V_mir2.n19 325.473
R7946 bgr_0.V_mir2.n13 bgr_0.V_mir2.n12 325.473
R7947 bgr_0.V_mir2.n8 bgr_0.V_mir2.n7 325.473
R7948 bgr_0.V_mir2.n16 bgr_0.V_mir2.t21 310.488
R7949 bgr_0.V_mir2.n9 bgr_0.V_mir2.t22 310.488
R7950 bgr_0.V_mir2.n4 bgr_0.V_mir2.t20 310.488
R7951 bgr_0.V_mir2.n2 bgr_0.V_mir2.t14 278.312
R7952 bgr_0.V_mir2.n2 bgr_0.V_mir2.n1 228.939
R7953 bgr_0.V_mir2.n3 bgr_0.V_mir2.n0 224.439
R7954 bgr_0.V_mir2.n18 bgr_0.V_mir2.t10 184.097
R7955 bgr_0.V_mir2.n11 bgr_0.V_mir2.t8 184.097
R7956 bgr_0.V_mir2.n6 bgr_0.V_mir2.t0 184.097
R7957 bgr_0.V_mir2.n17 bgr_0.V_mir2.n16 167.094
R7958 bgr_0.V_mir2.n10 bgr_0.V_mir2.n9 167.094
R7959 bgr_0.V_mir2.n5 bgr_0.V_mir2.n4 167.094
R7960 bgr_0.V_mir2.n13 bgr_0.V_mir2.n11 152
R7961 bgr_0.V_mir2.n8 bgr_0.V_mir2.n6 152
R7962 bgr_0.V_mir2.n19 bgr_0.V_mir2.n18 152
R7963 bgr_0.V_mir2.n16 bgr_0.V_mir2.t19 120.501
R7964 bgr_0.V_mir2.n17 bgr_0.V_mir2.t6 120.501
R7965 bgr_0.V_mir2.n9 bgr_0.V_mir2.t18 120.501
R7966 bgr_0.V_mir2.n10 bgr_0.V_mir2.t2 120.501
R7967 bgr_0.V_mir2.n4 bgr_0.V_mir2.t17 120.501
R7968 bgr_0.V_mir2.n5 bgr_0.V_mir2.t4 120.501
R7969 bgr_0.V_mir2.n1 bgr_0.V_mir2.t16 48.0005
R7970 bgr_0.V_mir2.n1 bgr_0.V_mir2.t12 48.0005
R7971 bgr_0.V_mir2.n0 bgr_0.V_mir2.t15 48.0005
R7972 bgr_0.V_mir2.n0 bgr_0.V_mir2.t13 48.0005
R7973 bgr_0.V_mir2.n18 bgr_0.V_mir2.n17 40.7027
R7974 bgr_0.V_mir2.n11 bgr_0.V_mir2.n10 40.7027
R7975 bgr_0.V_mir2.n6 bgr_0.V_mir2.n5 40.7027
R7976 bgr_0.V_mir2.n12 bgr_0.V_mir2.t3 39.4005
R7977 bgr_0.V_mir2.n12 bgr_0.V_mir2.t9 39.4005
R7978 bgr_0.V_mir2.n7 bgr_0.V_mir2.t5 39.4005
R7979 bgr_0.V_mir2.n7 bgr_0.V_mir2.t1 39.4005
R7980 bgr_0.V_mir2.n20 bgr_0.V_mir2.t7 39.4005
R7981 bgr_0.V_mir2.t11 bgr_0.V_mir2.n20 39.4005
R7982 bgr_0.V_mir2.n14 bgr_0.V_mir2.n13 15.8005
R7983 bgr_0.V_mir2.n14 bgr_0.V_mir2.n8 15.8005
R7984 bgr_0.V_mir2.n19 bgr_0.V_mir2.n15 9.3005
R7985 bgr_0.V_mir2.n3 bgr_0.V_mir2.n2 5.8755
R7986 bgr_0.V_mir2.n15 bgr_0.V_mir2.n14 4.5005
R7987 bgr_0.V_mir2.n15 bgr_0.V_mir2.n3 0.78175
R7988 bgr_0.Vin-.n7 bgr_0.Vin-.t12 688.859
R7989 bgr_0.Vin-.n9 bgr_0.Vin-.n8 514.134
R7990 bgr_0.Vin-.n6 bgr_0.Vin-.n5 351.522
R7991 bgr_0.Vin-.n11 bgr_0.Vin-.n10 213.4
R7992 bgr_0.Vin-.n7 bgr_0.Vin-.t8 174.726
R7993 bgr_0.Vin-.n8 bgr_0.Vin-.t10 174.726
R7994 bgr_0.Vin-.n9 bgr_0.Vin-.t9 174.726
R7995 bgr_0.Vin-.n10 bgr_0.Vin-.t11 174.726
R7996 bgr_0.Vin-.n4 bgr_0.Vin-.n2 173.029
R7997 bgr_0.Vin-.n4 bgr_0.Vin-.n3 168.654
R7998 bgr_0.Vin-.n8 bgr_0.Vin-.n7 128.534
R7999 bgr_0.Vin-.n10 bgr_0.Vin-.n9 128.534
R8000 bgr_0.Vin-.n12 bgr_0.Vin-.t6 119.099
R8001 bgr_0.Vin-.n16 bgr_0.Vin-.n15 83.5719
R8002 bgr_0.Vin-.n1 bgr_0.Vin-.n0 83.5719
R8003 bgr_0.Vin-.n19 bgr_0.Vin-.n1 73.8495
R8004 bgr_0.Vin-.t7 bgr_0.Vin-.n14 65.0341
R8005 bgr_0.Vin-.n5 bgr_0.Vin-.t5 39.4005
R8006 bgr_0.Vin-.n5 bgr_0.Vin-.t4 39.4005
R8007 bgr_0.Vin-.n13 bgr_0.Vin-.n12 28.813
R8008 bgr_0.Vin-.n15 bgr_0.Vin-.n1 26.074
R8009 bgr_0.Vin-.n12 bgr_0.Vin-.n11 16.188
R8010 bgr_0.Vin-.n3 bgr_0.Vin-.t0 13.1338
R8011 bgr_0.Vin-.n3 bgr_0.Vin-.t2 13.1338
R8012 bgr_0.Vin-.n2 bgr_0.Vin-.t3 13.1338
R8013 bgr_0.Vin-.n2 bgr_0.Vin-.t1 13.1338
R8014 bgr_0.Vin-.n11 bgr_0.Vin-.n6 11.2193
R8015 bgr_0.Vin-.n6 bgr_0.Vin-.n4 3.8755
R8016 bgr_0.Vin-.n16 bgr_0.Vin-.n14 1.56483
R8017 bgr_0.Vin-.n18 bgr_0.Vin-.n17 1.5505
R8018 bgr_0.Vin-.n17 bgr_0.Vin-.n0 0.885803
R8019 bgr_0.Vin-.n17 bgr_0.Vin-.n16 0.77514
R8020 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_23.Emitter bgr_0.Vin-.n0 0.756696
R8021 bgr_0.Vin-.n19 bgr_0.Vin-.n18 0.711459
R8022 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_23.Emitter bgr_0.Vin-.n19 0.576566
R8023 bgr_0.Vin-.n14 bgr_0.Vin-.n13 0.531499
R8024 bgr_0.Vin-.n15 bgr_0.Vin-.t7 0.290206
R8025 bgr_0.Vin-.n18 bgr_0.Vin-.n13 0.00817857
R8026 bgr_0.V_p_1.n1 bgr_0.V_p_1.n5 229.562
R8027 bgr_0.V_p_1.n1 bgr_0.V_p_1.n4 228.939
R8028 bgr_0.V_p_1.n0 bgr_0.V_p_1.n3 228.939
R8029 bgr_0.V_p_1.n0 bgr_0.V_p_1.n2 228.939
R8030 bgr_0.V_p_1.n6 bgr_0.V_p_1.n1 228.938
R8031 bgr_0.V_p_1.n0 bgr_0.V_p_1.t10 98.7279
R8032 bgr_0.V_p_1.n5 bgr_0.V_p_1.t7 48.0005
R8033 bgr_0.V_p_1.n5 bgr_0.V_p_1.t0 48.0005
R8034 bgr_0.V_p_1.n4 bgr_0.V_p_1.t9 48.0005
R8035 bgr_0.V_p_1.n4 bgr_0.V_p_1.t2 48.0005
R8036 bgr_0.V_p_1.n3 bgr_0.V_p_1.t3 48.0005
R8037 bgr_0.V_p_1.n3 bgr_0.V_p_1.t5 48.0005
R8038 bgr_0.V_p_1.n2 bgr_0.V_p_1.t8 48.0005
R8039 bgr_0.V_p_1.n2 bgr_0.V_p_1.t1 48.0005
R8040 bgr_0.V_p_1.t4 bgr_0.V_p_1.n6 48.0005
R8041 bgr_0.V_p_1.n6 bgr_0.V_p_1.t6 48.0005
R8042 bgr_0.V_p_1.n1 bgr_0.V_p_1.n0 1.8755
R8043 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.n2 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.n0 144.827
R8044 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.n2 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.n1 134.577
R8045 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.n12 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.t10 118.986
R8046 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.n5 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.n3 100.6
R8047 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.n11 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.n10 100.038
R8048 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.n9 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.n8 100.038
R8049 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.n7 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.n6 100.038
R8050 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.n5 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.n4 100.038
R8051 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.n13 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.n12 43.284
R8052 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.n13 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.n2 37.4067
R8053 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.n1 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.t13 24.0005
R8054 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.n1 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.t11 24.0005
R8055 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.n0 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.t14 24.0005
R8056 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.n0 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.t12 24.0005
R8057 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.n10 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.t2 8.0005
R8058 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.n10 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.t7 8.0005
R8059 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.n8 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.t6 8.0005
R8060 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.n8 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.t0 8.0005
R8061 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.n6 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.t3 8.0005
R8062 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.n6 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.t1 8.0005
R8063 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.n4 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.t4 8.0005
R8064 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.n4 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.t8 8.0005
R8065 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.n3 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.t5 8.0005
R8066 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.n3 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.t9 8.0005
R8067 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.n12 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.n11 5.6255
R8068 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.n7 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.n5 0.563
R8069 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.n9 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.n7 0.563
R8070 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.n11 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.n9 0.563
R8071 bgr_0.V_CMFB_S4 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.n13 0.047375
R8072 VIN+.n9 VIN+.t8 490.072
R8073 VIN+.n4 VIN+.t4 449.868
R8074 VIN+.n0 VIN+.t5 449.868
R8075 VIN+.n4 VIN+.t9 273.134
R8076 VIN+.n5 VIN+.t3 273.134
R8077 VIN+.n6 VIN+.t7 273.134
R8078 VIN+.n7 VIN+.t1 273.134
R8079 VIN+.n3 VIN+.t10 273.134
R8080 VIN+.n2 VIN+.t2 273.134
R8081 VIN+.n1 VIN+.t6 273.134
R8082 VIN+.n0 VIN+.t0 273.134
R8083 VIN+.n7 VIN+.n6 176.733
R8084 VIN+.n6 VIN+.n5 176.733
R8085 VIN+.n5 VIN+.n4 176.733
R8086 VIN+.n1 VIN+.n0 176.733
R8087 VIN+.n2 VIN+.n1 176.733
R8088 VIN+.n3 VIN+.n2 176.733
R8089 VIN+.n9 VIN+.n8 165.8
R8090 VIN+.n8 VIN+.n7 56.2338
R8091 VIN+.n8 VIN+.n3 56.2338
R8092 VIN+ VIN+.n9 2.14112
R8093 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.n2 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.n0 345.264
R8094 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.n2 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.n1 344.7
R8095 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.n4 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.n3 292.5
R8096 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.n7 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.n5 209.251
R8097 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.n13 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.n12 208.689
R8098 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.n11 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.n10 208.689
R8099 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.n9 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.n8 208.689
R8100 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.n7 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.n6 208.689
R8101 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.n14 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.t10 120.305
R8102 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.n4 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.n2 52.763
R8103 bgr_0.V_CMFB_S3 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.n4 51.7297
R8104 bgr_0.V_CMFB_S3 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.n14 50.813
R8105 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.n3 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.t15 39.4005
R8106 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.n3 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.t14 39.4005
R8107 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.n1 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.t12 39.4005
R8108 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.n1 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.t11 39.4005
R8109 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.n0 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.t13 39.4005
R8110 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.n0 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.t16 39.4005
R8111 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.n12 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.t8 19.7005
R8112 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.n12 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.t3 19.7005
R8113 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.n10 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.t2 19.7005
R8114 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.n10 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.t6 19.7005
R8115 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.n8 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.t9 19.7005
R8116 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.n8 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.t7 19.7005
R8117 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.n6 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.t0 19.7005
R8118 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.n6 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.t4 19.7005
R8119 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.n5 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.t1 19.7005
R8120 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.n5 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.t5 19.7005
R8121 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.n14 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.n13 5.90675
R8122 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.n9 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.n7 0.563
R8123 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.n11 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.n9 0.563
R8124 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.n13 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.n11 0.563
R8125 two_stage_opamp_dummy_magic_14_0.VD4.n28 two_stage_opamp_dummy_magic_14_0.VD4.t23 652.076
R8126 two_stage_opamp_dummy_magic_14_0.VD4.n61 two_stage_opamp_dummy_magic_14_0.VD4.t20 652.076
R8127 two_stage_opamp_dummy_magic_14_0.VD4.n60 two_stage_opamp_dummy_magic_14_0.VD4.n13 585
R8128 two_stage_opamp_dummy_magic_14_0.VD4.n42 two_stage_opamp_dummy_magic_14_0.VD4.n41 585
R8129 two_stage_opamp_dummy_magic_14_0.VD4.n48 two_stage_opamp_dummy_magic_14_0.VD4.n13 290.233
R8130 two_stage_opamp_dummy_magic_14_0.VD4.n54 two_stage_opamp_dummy_magic_14_0.VD4.n13 290.233
R8131 two_stage_opamp_dummy_magic_14_0.VD4.n49 two_stage_opamp_dummy_magic_14_0.VD4.n13 290.233
R8132 two_stage_opamp_dummy_magic_14_0.VD4.n41 two_stage_opamp_dummy_magic_14_0.VD4.n30 290.233
R8133 two_stage_opamp_dummy_magic_14_0.VD4.n41 two_stage_opamp_dummy_magic_14_0.VD4.n35 290.233
R8134 two_stage_opamp_dummy_magic_14_0.VD4.n41 two_stage_opamp_dummy_magic_14_0.VD4.n40 290.233
R8135 two_stage_opamp_dummy_magic_14_0.VD4.n49 two_stage_opamp_dummy_magic_14_0.VD4.n46 242.903
R8136 two_stage_opamp_dummy_magic_14_0.VD4.n40 two_stage_opamp_dummy_magic_14_0.VD4.n18 242.903
R8137 two_stage_opamp_dummy_magic_14_0.VD4.n60 two_stage_opamp_dummy_magic_14_0.VD4.n59 238.367
R8138 two_stage_opamp_dummy_magic_14_0.VD4.n15 two_stage_opamp_dummy_magic_14_0.VD4.n14 185
R8139 two_stage_opamp_dummy_magic_14_0.VD4.n57 two_stage_opamp_dummy_magic_14_0.VD4.n56 185
R8140 two_stage_opamp_dummy_magic_14_0.VD4.n58 two_stage_opamp_dummy_magic_14_0.VD4.n57 185
R8141 two_stage_opamp_dummy_magic_14_0.VD4.n55 two_stage_opamp_dummy_magic_14_0.VD4.n47 185
R8142 two_stage_opamp_dummy_magic_14_0.VD4.n53 two_stage_opamp_dummy_magic_14_0.VD4.n52 185
R8143 two_stage_opamp_dummy_magic_14_0.VD4.n51 two_stage_opamp_dummy_magic_14_0.VD4.n50 185
R8144 two_stage_opamp_dummy_magic_14_0.VD4.n43 two_stage_opamp_dummy_magic_14_0.VD4.n42 185
R8145 two_stage_opamp_dummy_magic_14_0.VD4.n44 two_stage_opamp_dummy_magic_14_0.VD4.n43 185
R8146 two_stage_opamp_dummy_magic_14_0.VD4.n29 two_stage_opamp_dummy_magic_14_0.VD4.n19 185
R8147 two_stage_opamp_dummy_magic_14_0.VD4.n32 two_stage_opamp_dummy_magic_14_0.VD4.n31 185
R8148 two_stage_opamp_dummy_magic_14_0.VD4.n34 two_stage_opamp_dummy_magic_14_0.VD4.n33 185
R8149 two_stage_opamp_dummy_magic_14_0.VD4.n37 two_stage_opamp_dummy_magic_14_0.VD4.n36 185
R8150 two_stage_opamp_dummy_magic_14_0.VD4.n39 two_stage_opamp_dummy_magic_14_0.VD4.n38 185
R8151 two_stage_opamp_dummy_magic_14_0.VD4.t24 two_stage_opamp_dummy_magic_14_0.VD4.n44 170.513
R8152 two_stage_opamp_dummy_magic_14_0.VD4.n58 two_stage_opamp_dummy_magic_14_0.VD4.t21 170.513
R8153 two_stage_opamp_dummy_magic_14_0.VD4.n2 two_stage_opamp_dummy_magic_14_0.VD4.n0 163.626
R8154 two_stage_opamp_dummy_magic_14_0.VD4.n10 two_stage_opamp_dummy_magic_14_0.VD4.n9 163.001
R8155 two_stage_opamp_dummy_magic_14_0.VD4.n8 two_stage_opamp_dummy_magic_14_0.VD4.n7 163.001
R8156 two_stage_opamp_dummy_magic_14_0.VD4.n6 two_stage_opamp_dummy_magic_14_0.VD4.n5 163.001
R8157 two_stage_opamp_dummy_magic_14_0.VD4.n4 two_stage_opamp_dummy_magic_14_0.VD4.n3 163.001
R8158 two_stage_opamp_dummy_magic_14_0.VD4.n2 two_stage_opamp_dummy_magic_14_0.VD4.n1 163.001
R8159 two_stage_opamp_dummy_magic_14_0.VD4.n12 two_stage_opamp_dummy_magic_14_0.VD4.n11 159.804
R8160 two_stage_opamp_dummy_magic_14_0.VD4.n21 two_stage_opamp_dummy_magic_14_0.VD4.n20 159.803
R8161 two_stage_opamp_dummy_magic_14_0.VD4.n23 two_stage_opamp_dummy_magic_14_0.VD4.n22 159.803
R8162 two_stage_opamp_dummy_magic_14_0.VD4.n25 two_stage_opamp_dummy_magic_14_0.VD4.n24 159.803
R8163 two_stage_opamp_dummy_magic_14_0.VD4.n27 two_stage_opamp_dummy_magic_14_0.VD4.n26 159.803
R8164 two_stage_opamp_dummy_magic_14_0.VD4.n57 two_stage_opamp_dummy_magic_14_0.VD4.n15 150
R8165 two_stage_opamp_dummy_magic_14_0.VD4.n57 two_stage_opamp_dummy_magic_14_0.VD4.n47 150
R8166 two_stage_opamp_dummy_magic_14_0.VD4.n52 two_stage_opamp_dummy_magic_14_0.VD4.n51 150
R8167 two_stage_opamp_dummy_magic_14_0.VD4.n43 two_stage_opamp_dummy_magic_14_0.VD4.n19 150
R8168 two_stage_opamp_dummy_magic_14_0.VD4.n33 two_stage_opamp_dummy_magic_14_0.VD4.n32 150
R8169 two_stage_opamp_dummy_magic_14_0.VD4.n38 two_stage_opamp_dummy_magic_14_0.VD4.n37 150
R8170 two_stage_opamp_dummy_magic_14_0.VD4.t10 two_stage_opamp_dummy_magic_14_0.VD4.t24 146.155
R8171 two_stage_opamp_dummy_magic_14_0.VD4.t6 two_stage_opamp_dummy_magic_14_0.VD4.t10 146.155
R8172 two_stage_opamp_dummy_magic_14_0.VD4.t12 two_stage_opamp_dummy_magic_14_0.VD4.t6 146.155
R8173 two_stage_opamp_dummy_magic_14_0.VD4.t16 two_stage_opamp_dummy_magic_14_0.VD4.t12 146.155
R8174 two_stage_opamp_dummy_magic_14_0.VD4.t0 two_stage_opamp_dummy_magic_14_0.VD4.t16 146.155
R8175 two_stage_opamp_dummy_magic_14_0.VD4.t2 two_stage_opamp_dummy_magic_14_0.VD4.t0 146.155
R8176 two_stage_opamp_dummy_magic_14_0.VD4.t4 two_stage_opamp_dummy_magic_14_0.VD4.t2 146.155
R8177 two_stage_opamp_dummy_magic_14_0.VD4.t8 two_stage_opamp_dummy_magic_14_0.VD4.t4 146.155
R8178 two_stage_opamp_dummy_magic_14_0.VD4.t14 two_stage_opamp_dummy_magic_14_0.VD4.t8 146.155
R8179 two_stage_opamp_dummy_magic_14_0.VD4.t18 two_stage_opamp_dummy_magic_14_0.VD4.t14 146.155
R8180 two_stage_opamp_dummy_magic_14_0.VD4.t21 two_stage_opamp_dummy_magic_14_0.VD4.t18 146.155
R8181 two_stage_opamp_dummy_magic_14_0.VD4.n59 two_stage_opamp_dummy_magic_14_0.VD4.n58 65.8183
R8182 two_stage_opamp_dummy_magic_14_0.VD4.n58 two_stage_opamp_dummy_magic_14_0.VD4.n45 65.8183
R8183 two_stage_opamp_dummy_magic_14_0.VD4.n58 two_stage_opamp_dummy_magic_14_0.VD4.n46 65.8183
R8184 two_stage_opamp_dummy_magic_14_0.VD4.n44 two_stage_opamp_dummy_magic_14_0.VD4.n16 65.8183
R8185 two_stage_opamp_dummy_magic_14_0.VD4.n44 two_stage_opamp_dummy_magic_14_0.VD4.n17 65.8183
R8186 two_stage_opamp_dummy_magic_14_0.VD4.n44 two_stage_opamp_dummy_magic_14_0.VD4.n18 65.8183
R8187 two_stage_opamp_dummy_magic_14_0.VD4.n47 two_stage_opamp_dummy_magic_14_0.VD4.n45 53.3664
R8188 two_stage_opamp_dummy_magic_14_0.VD4.n51 two_stage_opamp_dummy_magic_14_0.VD4.n46 53.3664
R8189 two_stage_opamp_dummy_magic_14_0.VD4.n59 two_stage_opamp_dummy_magic_14_0.VD4.n15 53.3664
R8190 two_stage_opamp_dummy_magic_14_0.VD4.n52 two_stage_opamp_dummy_magic_14_0.VD4.n45 53.3664
R8191 two_stage_opamp_dummy_magic_14_0.VD4.n19 two_stage_opamp_dummy_magic_14_0.VD4.n16 53.3664
R8192 two_stage_opamp_dummy_magic_14_0.VD4.n33 two_stage_opamp_dummy_magic_14_0.VD4.n17 53.3664
R8193 two_stage_opamp_dummy_magic_14_0.VD4.n38 two_stage_opamp_dummy_magic_14_0.VD4.n18 53.3664
R8194 two_stage_opamp_dummy_magic_14_0.VD4.n32 two_stage_opamp_dummy_magic_14_0.VD4.n16 53.3664
R8195 two_stage_opamp_dummy_magic_14_0.VD4.n37 two_stage_opamp_dummy_magic_14_0.VD4.n17 53.3664
R8196 two_stage_opamp_dummy_magic_14_0.VD4.n61 two_stage_opamp_dummy_magic_14_0.VD4.n60 22.8576
R8197 two_stage_opamp_dummy_magic_14_0.VD4.n42 two_stage_opamp_dummy_magic_14_0.VD4.n28 22.8576
R8198 two_stage_opamp_dummy_magic_14_0.VD4.n28 two_stage_opamp_dummy_magic_14_0.VD4.n27 14.4255
R8199 two_stage_opamp_dummy_magic_14_0.VD4.n62 two_stage_opamp_dummy_magic_14_0.VD4.n61 13.8005
R8200 two_stage_opamp_dummy_magic_14_0.VD4.n20 two_stage_opamp_dummy_magic_14_0.VD4.t5 11.2576
R8201 two_stage_opamp_dummy_magic_14_0.VD4.n20 two_stage_opamp_dummy_magic_14_0.VD4.t9 11.2576
R8202 two_stage_opamp_dummy_magic_14_0.VD4.n22 two_stage_opamp_dummy_magic_14_0.VD4.t1 11.2576
R8203 two_stage_opamp_dummy_magic_14_0.VD4.n22 two_stage_opamp_dummy_magic_14_0.VD4.t3 11.2576
R8204 two_stage_opamp_dummy_magic_14_0.VD4.n24 two_stage_opamp_dummy_magic_14_0.VD4.t13 11.2576
R8205 two_stage_opamp_dummy_magic_14_0.VD4.n24 two_stage_opamp_dummy_magic_14_0.VD4.t17 11.2576
R8206 two_stage_opamp_dummy_magic_14_0.VD4.n26 two_stage_opamp_dummy_magic_14_0.VD4.t11 11.2576
R8207 two_stage_opamp_dummy_magic_14_0.VD4.n26 two_stage_opamp_dummy_magic_14_0.VD4.t7 11.2576
R8208 two_stage_opamp_dummy_magic_14_0.VD4.n41 two_stage_opamp_dummy_magic_14_0.VD4.t25 11.2576
R8209 two_stage_opamp_dummy_magic_14_0.VD4.n13 two_stage_opamp_dummy_magic_14_0.VD4.t22 11.2576
R8210 two_stage_opamp_dummy_magic_14_0.VD4.n9 two_stage_opamp_dummy_magic_14_0.VD4.t36 11.2576
R8211 two_stage_opamp_dummy_magic_14_0.VD4.n9 two_stage_opamp_dummy_magic_14_0.VD4.t30 11.2576
R8212 two_stage_opamp_dummy_magic_14_0.VD4.n7 two_stage_opamp_dummy_magic_14_0.VD4.t28 11.2576
R8213 two_stage_opamp_dummy_magic_14_0.VD4.n7 two_stage_opamp_dummy_magic_14_0.VD4.t31 11.2576
R8214 two_stage_opamp_dummy_magic_14_0.VD4.n5 two_stage_opamp_dummy_magic_14_0.VD4.t33 11.2576
R8215 two_stage_opamp_dummy_magic_14_0.VD4.n5 two_stage_opamp_dummy_magic_14_0.VD4.t35 11.2576
R8216 two_stage_opamp_dummy_magic_14_0.VD4.n3 two_stage_opamp_dummy_magic_14_0.VD4.t27 11.2576
R8217 two_stage_opamp_dummy_magic_14_0.VD4.n3 two_stage_opamp_dummy_magic_14_0.VD4.t26 11.2576
R8218 two_stage_opamp_dummy_magic_14_0.VD4.n1 two_stage_opamp_dummy_magic_14_0.VD4.t29 11.2576
R8219 two_stage_opamp_dummy_magic_14_0.VD4.n1 two_stage_opamp_dummy_magic_14_0.VD4.t32 11.2576
R8220 two_stage_opamp_dummy_magic_14_0.VD4.n0 two_stage_opamp_dummy_magic_14_0.VD4.t34 11.2576
R8221 two_stage_opamp_dummy_magic_14_0.VD4.n0 two_stage_opamp_dummy_magic_14_0.VD4.t37 11.2576
R8222 two_stage_opamp_dummy_magic_14_0.VD4.n11 two_stage_opamp_dummy_magic_14_0.VD4.t15 11.2576
R8223 two_stage_opamp_dummy_magic_14_0.VD4.n11 two_stage_opamp_dummy_magic_14_0.VD4.t19 11.2576
R8224 two_stage_opamp_dummy_magic_14_0.VD4.n60 two_stage_opamp_dummy_magic_14_0.VD4.n14 9.14336
R8225 two_stage_opamp_dummy_magic_14_0.VD4.n56 two_stage_opamp_dummy_magic_14_0.VD4.n55 9.14336
R8226 two_stage_opamp_dummy_magic_14_0.VD4.n53 two_stage_opamp_dummy_magic_14_0.VD4.n50 9.14336
R8227 two_stage_opamp_dummy_magic_14_0.VD4.n42 two_stage_opamp_dummy_magic_14_0.VD4.n29 9.14336
R8228 two_stage_opamp_dummy_magic_14_0.VD4.n34 two_stage_opamp_dummy_magic_14_0.VD4.n31 9.14336
R8229 two_stage_opamp_dummy_magic_14_0.VD4.n39 two_stage_opamp_dummy_magic_14_0.VD4.n36 9.14336
R8230 two_stage_opamp_dummy_magic_14_0.VD4.n63 two_stage_opamp_dummy_magic_14_0.VD4.n10 8.2505
R8231 two_stage_opamp_dummy_magic_14_0.VD4.n63 two_stage_opamp_dummy_magic_14_0.VD4.n62 5.3755
R8232 two_stage_opamp_dummy_magic_14_0.VD4.n48 two_stage_opamp_dummy_magic_14_0.VD4.n14 4.53698
R8233 two_stage_opamp_dummy_magic_14_0.VD4.n55 two_stage_opamp_dummy_magic_14_0.VD4.n54 4.53698
R8234 two_stage_opamp_dummy_magic_14_0.VD4.n50 two_stage_opamp_dummy_magic_14_0.VD4.n49 4.53698
R8235 two_stage_opamp_dummy_magic_14_0.VD4.n56 two_stage_opamp_dummy_magic_14_0.VD4.n48 4.53698
R8236 two_stage_opamp_dummy_magic_14_0.VD4.n54 two_stage_opamp_dummy_magic_14_0.VD4.n53 4.53698
R8237 two_stage_opamp_dummy_magic_14_0.VD4.n30 two_stage_opamp_dummy_magic_14_0.VD4.n29 4.53698
R8238 two_stage_opamp_dummy_magic_14_0.VD4.n35 two_stage_opamp_dummy_magic_14_0.VD4.n34 4.53698
R8239 two_stage_opamp_dummy_magic_14_0.VD4.n40 two_stage_opamp_dummy_magic_14_0.VD4.n39 4.53698
R8240 two_stage_opamp_dummy_magic_14_0.VD4.n31 two_stage_opamp_dummy_magic_14_0.VD4.n30 4.53698
R8241 two_stage_opamp_dummy_magic_14_0.VD4.n36 two_stage_opamp_dummy_magic_14_0.VD4.n35 4.53698
R8242 two_stage_opamp_dummy_magic_14_0.VD4.n4 two_stage_opamp_dummy_magic_14_0.VD4.n2 0.6255
R8243 two_stage_opamp_dummy_magic_14_0.VD4.n6 two_stage_opamp_dummy_magic_14_0.VD4.n4 0.6255
R8244 two_stage_opamp_dummy_magic_14_0.VD4.n8 two_stage_opamp_dummy_magic_14_0.VD4.n6 0.6255
R8245 two_stage_opamp_dummy_magic_14_0.VD4.n10 two_stage_opamp_dummy_magic_14_0.VD4.n8 0.6255
R8246 two_stage_opamp_dummy_magic_14_0.VD4.n62 two_stage_opamp_dummy_magic_14_0.VD4.n12 0.6255
R8247 two_stage_opamp_dummy_magic_14_0.VD4.n27 two_stage_opamp_dummy_magic_14_0.VD4.n25 0.6255
R8248 two_stage_opamp_dummy_magic_14_0.VD4.n25 two_stage_opamp_dummy_magic_14_0.VD4.n23 0.6255
R8249 two_stage_opamp_dummy_magic_14_0.VD4.n23 two_stage_opamp_dummy_magic_14_0.VD4.n21 0.6255
R8250 two_stage_opamp_dummy_magic_14_0.VD4.n21 two_stage_opamp_dummy_magic_14_0.VD4.n12 0.6255
R8251 two_stage_opamp_dummy_magic_14_0.VD4 two_stage_opamp_dummy_magic_14_0.VD4.n63 0.063
R8252 bgr_0.START_UP.n4 bgr_0.START_UP.t6 238.322
R8253 bgr_0.START_UP.n4 bgr_0.START_UP.t7 238.322
R8254 bgr_0.START_UP.n3 bgr_0.START_UP.n1 175.56
R8255 bgr_0.START_UP.n3 bgr_0.START_UP.n2 168.936
R8256 bgr_0.START_UP.n5 bgr_0.START_UP.n4 166.925
R8257 bgr_0.START_UP.n0 bgr_0.START_UP.t5 130.001
R8258 bgr_0.START_UP.n0 bgr_0.START_UP.t4 81.7074
R8259 bgr_0.START_UP bgr_0.START_UP.n0 36.9489
R8260 bgr_0.START_UP bgr_0.START_UP.n5 13.4693
R8261 bgr_0.START_UP.n1 bgr_0.START_UP.t0 13.1338
R8262 bgr_0.START_UP.n1 bgr_0.START_UP.t2 13.1338
R8263 bgr_0.START_UP.n2 bgr_0.START_UP.t1 13.1338
R8264 bgr_0.START_UP.n2 bgr_0.START_UP.t3 13.1338
R8265 bgr_0.START_UP.n5 bgr_0.START_UP.n3 4.21925
R8266 two_stage_opamp_dummy_magic_14_0.V_err_p.n1 two_stage_opamp_dummy_magic_14_0.V_err_p.n0 365.07
R8267 two_stage_opamp_dummy_magic_14_0.V_err_p.n0 two_stage_opamp_dummy_magic_14_0.V_err_p.t0 15.7605
R8268 two_stage_opamp_dummy_magic_14_0.V_err_p.n0 two_stage_opamp_dummy_magic_14_0.V_err_p.t3 15.7605
R8269 two_stage_opamp_dummy_magic_14_0.V_err_p.n1 two_stage_opamp_dummy_magic_14_0.V_err_p.t2 15.7605
R8270 two_stage_opamp_dummy_magic_14_0.V_err_p.t1 two_stage_opamp_dummy_magic_14_0.V_err_p.n1 15.7605
R8271 a_5980_2720.t0 a_5980_2720.t1 169.905
R8272 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n4 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.t2 652.076
R8273 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n14 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.t6 652.076
R8274 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n28 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n27 585
R8275 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n44 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n2 585
R8276 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n27 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n16 290.233
R8277 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n27 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n21 290.233
R8278 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n27 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n26 290.233
R8279 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n44 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n43 290.233
R8280 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n44 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n0 290.233
R8281 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n44 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n1 290.233
R8282 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n26 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n8 242.903
R8283 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n36 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n1 242.903
R8284 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n42 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n41 238.367
R8285 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n29 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n28 185
R8286 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n30 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n29 185
R8287 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n15 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n9 185
R8288 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n18 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n17 185
R8289 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n20 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n19 185
R8290 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n23 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n22 185
R8291 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n25 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n24 185
R8292 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n5 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n3 185
R8293 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n39 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n2 185
R8294 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n40 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n39 185
R8295 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n38 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n37 185
R8296 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n33 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n32 185
R8297 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n35 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n34 185
R8298 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.t7 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n30 170.513
R8299 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n40 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.t3 170.513
R8300 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n12 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n10 169.694
R8301 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n12 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n11 155.303
R8302 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n39 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n5 150
R8303 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n39 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n38 150
R8304 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n35 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n32 150
R8305 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n29 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n9 150
R8306 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n19 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n18 150
R8307 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n24 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n23 150
R8308 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.t0 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.t7 146.155
R8309 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.t3 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.t0 146.155
R8310 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n30 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n6 65.8183
R8311 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n30 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n7 65.8183
R8312 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n30 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n8 65.8183
R8313 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n41 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n40 65.8183
R8314 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n40 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n31 65.8183
R8315 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n40 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n36 65.8183
R8316 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n38 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n31 53.3664
R8317 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n36 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n35 53.3664
R8318 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n9 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n6 53.3664
R8319 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n19 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n7 53.3664
R8320 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n24 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n8 53.3664
R8321 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n18 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n6 53.3664
R8322 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n23 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n7 53.3664
R8323 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n41 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n5 53.3664
R8324 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n32 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n31 53.3664
R8325 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n28 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n14 22.8576
R8326 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n42 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n4 22.8576
R8327 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n14 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n13 14.4255
R8328 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n13 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n4 14.0505
R8329 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n11 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.t1 11.2576
R8330 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n11 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.t4 11.2576
R8331 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n10 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.t9 11.2576
R8332 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n10 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.t10 11.2576
R8333 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n27 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.t8 11.2576
R8334 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.t5 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n44 11.2576
R8335 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n28 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n15 9.14336
R8336 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n20 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n17 9.14336
R8337 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n25 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n22 9.14336
R8338 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n3 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n2 9.14336
R8339 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n37 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n2 9.14336
R8340 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n34 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n33 9.14336
R8341 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n16 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n15 4.53698
R8342 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n21 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n20 4.53698
R8343 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n26 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n25 4.53698
R8344 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n17 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n16 4.53698
R8345 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n22 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n21 4.53698
R8346 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n43 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n42 4.53698
R8347 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n37 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n0 4.53698
R8348 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n34 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n1 4.53698
R8349 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n43 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n3 4.53698
R8350 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n33 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n0 4.53698
R8351 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n13 two_stage_opamp_dummy_magic_14_0.Vb2_Vb3.n12 4.5005
R8352 a_14010_2720.t0 a_14010_2720.t1 169.905
R8353 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.n2 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.n0 344.837
R8354 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.n2 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.n1 344.274
R8355 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.n4 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.n3 292.5
R8356 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.n7 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.n5 209.251
R8357 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.n13 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.n12 208.689
R8358 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.n11 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.n10 208.689
R8359 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.n9 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.n8 208.689
R8360 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.n7 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.n6 208.689
R8361 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.n14 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.t16 120.305
R8362 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.n4 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.n2 52.3363
R8363 bgr_0.V_CMFB_S1 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.n4 52.1563
R8364 bgr_0.V_CMFB_S1 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.n14 50.813
R8365 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.n3 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.t11 39.4005
R8366 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.n3 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.t14 39.4005
R8367 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.n1 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.t10 39.4005
R8368 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.n1 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.t13 39.4005
R8369 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.n0 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.t15 39.4005
R8370 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.n0 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.t12 39.4005
R8371 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.n12 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.t4 19.7005
R8372 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.n12 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.t8 19.7005
R8373 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.n10 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.t3 19.7005
R8374 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.n10 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.t7 19.7005
R8375 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.n8 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.t2 19.7005
R8376 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.n8 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.t6 19.7005
R8377 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.n6 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.t0 19.7005
R8378 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.n6 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.t9 19.7005
R8379 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.n5 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.t1 19.7005
R8380 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.n5 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.t5 19.7005
R8381 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.n14 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.n13 5.90675
R8382 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.n9 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.n7 0.563
R8383 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.n11 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.n9 0.563
R8384 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.n13 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.n11 0.563
R8385 bgr_0.START_UP_NFET1 bgr_0.START_UP_NFET1.t0 141.653
R8386 two_stage_opamp_dummy_magic_14_0.err_amp_mir.n1 two_stage_opamp_dummy_magic_14_0.err_amp_mir.t5 554.301
R8387 two_stage_opamp_dummy_magic_14_0.err_amp_mir.n1 two_stage_opamp_dummy_magic_14_0.err_amp_mir.t0 442.837
R8388 two_stage_opamp_dummy_magic_14_0.err_amp_mir.n2 two_stage_opamp_dummy_magic_14_0.err_amp_mir.n0 193.744
R8389 two_stage_opamp_dummy_magic_14_0.err_amp_mir.n2 two_stage_opamp_dummy_magic_14_0.err_amp_mir.n1 173.088
R8390 two_stage_opamp_dummy_magic_14_0.err_amp_mir.n3 two_stage_opamp_dummy_magic_14_0.err_amp_mir.n2 86.8857
R8391 two_stage_opamp_dummy_magic_14_0.err_amp_mir.n0 two_stage_opamp_dummy_magic_14_0.err_amp_mir.t4 15.7605
R8392 two_stage_opamp_dummy_magic_14_0.err_amp_mir.n0 two_stage_opamp_dummy_magic_14_0.err_amp_mir.t3 15.7605
R8393 two_stage_opamp_dummy_magic_14_0.err_amp_mir.t1 two_stage_opamp_dummy_magic_14_0.err_amp_mir.n3 9.6005
R8394 two_stage_opamp_dummy_magic_14_0.err_amp_mir.n3 two_stage_opamp_dummy_magic_14_0.err_amp_mir.t2 9.6005
R8395 a_12530_23988.t0 a_12530_23988.t1 178.133
R8396 two_stage_opamp_dummy_magic_14_0.V_tot.n2 two_stage_opamp_dummy_magic_14_0.V_tot.t4 648.28
R8397 two_stage_opamp_dummy_magic_14_0.V_tot.n1 two_stage_opamp_dummy_magic_14_0.V_tot.t5 648.28
R8398 two_stage_opamp_dummy_magic_14_0.V_tot.n0 two_stage_opamp_dummy_magic_14_0.V_tot.t3 116.546
R8399 two_stage_opamp_dummy_magic_14_0.V_tot.n3 two_stage_opamp_dummy_magic_14_0.V_tot.t1 116.546
R8400 two_stage_opamp_dummy_magic_14_0.V_tot.n0 two_stage_opamp_dummy_magic_14_0.V_tot.t2 107.328
R8401 two_stage_opamp_dummy_magic_14_0.V_tot.t0 two_stage_opamp_dummy_magic_14_0.V_tot.n3 107.328
R8402 two_stage_opamp_dummy_magic_14_0.V_tot.n3 two_stage_opamp_dummy_magic_14_0.V_tot.n2 34.8494
R8403 two_stage_opamp_dummy_magic_14_0.V_tot.n1 two_stage_opamp_dummy_magic_14_0.V_tot.n0 34.8494
R8404 two_stage_opamp_dummy_magic_14_0.V_tot.n2 two_stage_opamp_dummy_magic_14_0.V_tot.n1 1.563
R8405 two_stage_opamp_dummy_magic_14_0.V_p_mir.n1 two_stage_opamp_dummy_magic_14_0.V_p_mir.n0 223.19
R8406 two_stage_opamp_dummy_magic_14_0.V_p_mir.n0 two_stage_opamp_dummy_magic_14_0.V_p_mir.t1 16.0005
R8407 two_stage_opamp_dummy_magic_14_0.V_p_mir.n0 two_stage_opamp_dummy_magic_14_0.V_p_mir.t0 16.0005
R8408 two_stage_opamp_dummy_magic_14_0.V_p_mir.t2 two_stage_opamp_dummy_magic_14_0.V_p_mir.n1 9.6005
R8409 two_stage_opamp_dummy_magic_14_0.V_p_mir.n1 two_stage_opamp_dummy_magic_14_0.V_p_mir.t3 9.6005
R8410 a_7580_22380.t0 a_7580_22380.t1 178.133
R8411 a_5700_5524.t0 a_5700_5524.t1 169.905
R8412 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n22 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t0 195.608
R8413 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n30 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n29 83.5719
R8414 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n28 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n27 83.5719
R8415 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n26 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n25 83.5719
R8416 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n104 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n103 83.5719
R8417 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n102 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n33 83.5719
R8418 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n101 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n100 83.5719
R8419 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n92 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n36 83.5719
R8420 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n85 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n37 83.5719
R8421 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n87 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n86 83.5719
R8422 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n79 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n41 83.5719
R8423 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n74 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n42 83.5719
R8424 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n66 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n65 83.5719
R8425 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n64 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n63 83.5719
R8426 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n62 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n61 83.5719
R8427 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n122 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n121 83.5719
R8428 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n120 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n119 83.5719
R8429 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n12 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n11 83.5719
R8430 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n130 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n129 83.5719
R8431 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n7 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n5 83.5719
R8432 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n135 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n4 83.5719
R8433 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n51 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n0 83.5719
R8434 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n52 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n50 83.5719
R8435 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n103 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n32 73.8495
R8436 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n116 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n11 73.8495
R8437 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n29 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n21 73.3165
R8438 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n94 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n36 73.3165
R8439 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n81 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n41 73.3165
R8440 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n67 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n66 73.3165
R8441 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n129 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n128 73.3165
R8442 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n51 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n1 73.3165
R8443 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n26 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n24 73.19
R8444 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n101 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n34 73.19
R8445 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n86 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n84 73.19
R8446 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n62 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n48 73.19
R8447 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n121 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n8 73.19
R8448 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n137 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n4 73.19
R8449 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n75 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t6 65.0299
R8450 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n53 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t3 65.0299
R8451 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n29 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n28 26.074
R8452 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n103 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n102 26.074
R8453 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n85 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n36 26.074
R8454 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n74 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n41 26.074
R8455 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n66 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n64 26.074
R8456 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n120 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n11 26.074
R8457 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n129 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n7 26.074
R8458 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n52 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n51 26.074
R8459 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t7 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n26 25.7843
R8460 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t8 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n101 25.7843
R8461 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n86 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t2 25.7843
R8462 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t5 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n62 25.7843
R8463 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n121 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t4 25.7843
R8464 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t1 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n4 25.7843
R8465 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n68 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n56 9.3005
R8466 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n56 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n46 9.3005
R8467 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n56 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 9.3005
R8468 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n72 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n56 9.3005
R8469 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n58 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n46 9.3005
R8470 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n58 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 9.3005
R8471 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n58 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n44 9.3005
R8472 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n72 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n58 9.3005
R8473 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n73 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n46 9.3005
R8474 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n73 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n45 9.3005
R8475 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n73 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 9.3005
R8476 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n73 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n44 9.3005
R8477 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n73 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n72 9.3005
R8478 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n72 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n60 9.3005
R8479 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n60 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n44 9.3005
R8480 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n60 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 9.3005
R8481 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n60 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n45 9.3005
R8482 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n72 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n55 9.3005
R8483 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n55 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n44 9.3005
R8484 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n55 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 9.3005
R8485 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n55 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n45 9.3005
R8486 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n68 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n55 9.3005
R8487 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n71 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n46 9.3005
R8488 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n71 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n45 9.3005
R8489 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n71 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 9.3005
R8490 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n72 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n71 9.3005
R8491 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n113 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n112 9.3005
R8492 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n112 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n111 9.3005
R8493 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n112 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 9.3005
R8494 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n112 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n14 9.3005
R8495 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n112 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n15 9.3005
R8496 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n111 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n109 9.3005
R8497 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n109 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 9.3005
R8498 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n109 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n14 9.3005
R8499 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n109 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n15 9.3005
R8500 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n111 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n108 9.3005
R8501 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n108 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 9.3005
R8502 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n108 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n14 9.3005
R8503 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n108 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n16 9.3005
R8504 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n108 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n15 9.3005
R8505 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n18 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n15 9.3005
R8506 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n18 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n16 9.3005
R8507 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n18 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n14 9.3005
R8508 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n18 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 9.3005
R8509 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n15 9.3005
R8510 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n16 9.3005
R8511 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n14 9.3005
R8512 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 9.3005
R8513 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n113 9.3005
R8514 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n111 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n110 9.3005
R8515 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n110 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 9.3005
R8516 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n110 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n14 9.3005
R8517 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n110 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n16 9.3005
R8518 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n110 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n15 9.3005
R8519 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n70 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n44 4.64654
R8520 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n57 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n45 4.64654
R8521 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n68 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n43 4.64654
R8522 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n59 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n46 4.64654
R8523 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n69 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n68 4.64654
R8524 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n23 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n16 4.64654
R8525 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n113 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n20 4.64654
R8526 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n111 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n13 4.64654
R8527 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n113 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n19 4.64654
R8528 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n96 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n34 2.36206
R8529 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n84 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n83 2.36206
R8530 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n125 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n8 2.36206
R8531 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n138 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n137 2.36206
R8532 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n95 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n94 2.19742
R8533 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n82 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n81 2.19742
R8534 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n128 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n126 2.19742
R8535 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n139 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n1 2.19742
R8536 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n75 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n42 1.56363
R8537 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n53 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n50 1.56363
R8538 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n141 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n140 1.5505
R8539 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n49 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n2 1.5505
R8540 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n127 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n6 1.5505
R8541 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n132 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n131 1.5505
R8542 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n134 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n133 1.5505
R8543 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n136 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n3 1.5505
R8544 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n118 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n117 1.5505
R8545 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n124 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n123 1.5505
R8546 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n10 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n9 1.5505
R8547 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n80 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n40 1.5505
R8548 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n78 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n77 1.5505
R8549 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n93 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n35 1.5505
R8550 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n91 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n90 1.5505
R8551 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n89 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n88 1.5505
R8552 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n39 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n38 1.5505
R8553 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n106 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n105 1.5505
R8554 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n99 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n31 1.5505
R8555 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n98 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n97 1.5505
R8556 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n25 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n16 1.25468
R8557 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n100 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n98 1.25468
R8558 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n87 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n39 1.25468
R8559 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n61 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n44 1.25468
R8560 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n123 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n122 1.25468
R8561 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n136 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n135 1.25468
R8562 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n111 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n21 1.19225
R8563 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n94 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n93 1.19225
R8564 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n81 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n80 1.19225
R8565 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n67 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n46 1.19225
R8566 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n128 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n127 1.19225
R8567 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n141 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n1 1.19225
R8568 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n27 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n14 1.07024
R8569 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n99 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n33 1.07024
R8570 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n88 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n37 1.07024
R8571 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n63 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 1.07024
R8572 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n119 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n10 1.07024
R8573 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n134 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n5 1.07024
R8574 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n24 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n16 1.0237
R8575 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n98 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n34 1.0237
R8576 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n84 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n39 1.0237
R8577 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n48 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n44 1.0237
R8578 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n123 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n8 1.0237
R8579 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n137 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n136 1.0237
R8580 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n30 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 0.885803
R8581 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n105 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n104 0.885803
R8582 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n92 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n91 0.885803
R8583 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n79 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n78 0.885803
R8584 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n65 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n45 0.885803
R8585 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n118 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n12 0.885803
R8586 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n131 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n130 0.885803
R8587 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n49 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n0 0.885803
R8588 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n24 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n15 0.812055
R8589 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n72 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n48 0.812055
R8590 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n27 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 0.77514
R8591 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n105 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n33 0.77514
R8592 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n91 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n37 0.77514
R8593 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n78 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n42 0.77514
R8594 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n63 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n45 0.77514
R8595 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n119 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n118 0.77514
R8596 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n131 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n5 0.77514
R8597 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n50 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n49 0.77514
R8598 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n30 0.756696
R8599 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n104 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.756696
R8600 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n92 0.756696
R8601 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n79 0.756696
R8602 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n65 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.756696
R8603 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n12 0.756696
R8604 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n130 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.756696
R8605 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n0 0.756696
R8606 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n117 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n116 0.711459
R8607 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n106 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n32 0.711459
R8608 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n113 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n21 0.647417
R8609 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n68 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n67 0.647417
R8610 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n25 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n14 0.590702
R8611 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n100 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n99 0.590702
R8612 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n88 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n87 0.590702
R8613 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n61 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 0.590702
R8614 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n122 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n10 0.590702
R8615 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n135 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n134 0.590702
R8616 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n32 0.576566
R8617 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n116 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.576566
R8618 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n54 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n53 0.530034
R8619 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n76 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n75 0.530034
R8620 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n28 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t7 0.290206
R8621 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n102 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t8 0.290206
R8622 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t2 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n85 0.290206
R8623 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t6 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n74 0.290206
R8624 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n64 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t5 0.290206
R8625 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t4 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n120 0.290206
R8626 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n7 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t1 0.290206
R8627 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t3 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n52 0.290206
R8628 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n111 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.203382
R8629 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n93 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.203382
R8630 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n80 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.203382
R8631 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n46 0.203382
R8632 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n127 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.203382
R8633 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n141 0.203382
R8634 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n139 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n138 0.154071
R8635 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n126 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n125 0.154071
R8636 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n83 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n82 0.154071
R8637 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n96 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n95 0.154071
R8638 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n76 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n73 0.137464
R8639 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n108 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n107 0.137464
R8640 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n55 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n54 0.134964
R8641 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n115 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 0.134964
R8642 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n140 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n2 0.0183571
R8643 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n140 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n139 0.0183571
R8644 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n138 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n3 0.0183571
R8645 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n133 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n3 0.0183571
R8646 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n133 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n132 0.0183571
R8647 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n132 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n6 0.0183571
R8648 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n126 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n6 0.0183571
R8649 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n125 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n124 0.0183571
R8650 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n124 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n9 0.0183571
R8651 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n77 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n40 0.0183571
R8652 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n82 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n40 0.0183571
R8653 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n83 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n38 0.0183571
R8654 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n89 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n38 0.0183571
R8655 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n90 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n89 0.0183571
R8656 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n90 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n35 0.0183571
R8657 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n95 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n35 0.0183571
R8658 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n97 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n96 0.0183571
R8659 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n97 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n31 0.0183571
R8660 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n115 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n9 0.0106786
R8661 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n107 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n31 0.0106786
R8662 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n110 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n22 0.0106786
R8663 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n60 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n59 0.00992001
R8664 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n71 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n69 0.00992001
R8665 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n70 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n56 0.00992001
R8666 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n58 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n57 0.00992001
R8667 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n73 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n43 0.00992001
R8668 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n57 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n56 0.00992001
R8669 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n58 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n43 0.00992001
R8670 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n69 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n60 0.00992001
R8671 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n59 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n55 0.00992001
R8672 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n71 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n70 0.00992001
R8673 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n18 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n13 0.00992001
R8674 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n110 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n19 0.00992001
R8675 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n109 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n23 0.00992001
R8676 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n108 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n20 0.00992001
R8677 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n112 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n23 0.00992001
R8678 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n109 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n20 0.00992001
R8679 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n19 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n18 0.00992001
R8680 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n13 0.00992001
R8681 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n54 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n2 0.00817857
R8682 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n117 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n115 0.00817857
R8683 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n77 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n76 0.00817857
R8684 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n107 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n106 0.00817857
R8685 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n112 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n22 0.00817857
R8686 a_5580_5524.t0 a_5580_5524.t1 262.248
R8687 a_12410_22380.t0 a_12410_22380.t1 178.133
R8688 a_13060_22630.t0 a_13060_22630.t1 178.133
R8689 a_6810_23838.t0 a_6810_23838.t1 178.133
R8690 a_6930_22664.t0 a_6930_22664.t1 178.133
R8691 two_stage_opamp_dummy_magic_14_0.Vb2_2.n32 two_stage_opamp_dummy_magic_14_0.Vb2_2.n31 692.967
R8692 two_stage_opamp_dummy_magic_14_0.Vb2_2.n34 two_stage_opamp_dummy_magic_14_0.Vb2_2.t4 652.076
R8693 two_stage_opamp_dummy_magic_14_0.Vb2_2.n30 two_stage_opamp_dummy_magic_14_0.Vb2_2.t7 652.076
R8694 two_stage_opamp_dummy_magic_14_0.Vb2_2.n36 two_stage_opamp_dummy_magic_14_0.Vb2_2.n0 587.407
R8695 two_stage_opamp_dummy_magic_14_0.Vb2_2.n41 two_stage_opamp_dummy_magic_14_0.Vb2_2.n2 587.407
R8696 two_stage_opamp_dummy_magic_14_0.Vb2_2.n29 two_stage_opamp_dummy_magic_14_0.Vb2_2.n11 585
R8697 two_stage_opamp_dummy_magic_14_0.Vb2_2.n3 two_stage_opamp_dummy_magic_14_0.Vb2_2.n0 585
R8698 two_stage_opamp_dummy_magic_14_0.Vb2_2.t6 two_stage_opamp_dummy_magic_14_0.Vb2_2.n44 585
R8699 two_stage_opamp_dummy_magic_14_0.Vb2_2.n43 two_stage_opamp_dummy_magic_14_0.Vb2_2.n2 585
R8700 two_stage_opamp_dummy_magic_14_0.Vb2_2.n17 two_stage_opamp_dummy_magic_14_0.Vb2_2.n11 290.233
R8701 two_stage_opamp_dummy_magic_14_0.Vb2_2.n23 two_stage_opamp_dummy_magic_14_0.Vb2_2.n11 290.233
R8702 two_stage_opamp_dummy_magic_14_0.Vb2_2.n18 two_stage_opamp_dummy_magic_14_0.Vb2_2.n11 290.233
R8703 two_stage_opamp_dummy_magic_14_0.Vb2_2.t6 two_stage_opamp_dummy_magic_14_0.Vb2_2.n0 246.25
R8704 two_stage_opamp_dummy_magic_14_0.Vb2_2.t6 two_stage_opamp_dummy_magic_14_0.Vb2_2.n2 246.25
R8705 two_stage_opamp_dummy_magic_14_0.Vb2_2.n41 two_stage_opamp_dummy_magic_14_0.Vb2_2.n40 243.698
R8706 two_stage_opamp_dummy_magic_14_0.Vb2_2.n18 two_stage_opamp_dummy_magic_14_0.Vb2_2.n15 242.903
R8707 two_stage_opamp_dummy_magic_14_0.Vb2_2.n29 two_stage_opamp_dummy_magic_14_0.Vb2_2.n28 238.367
R8708 two_stage_opamp_dummy_magic_14_0.Vb2_2.n13 two_stage_opamp_dummy_magic_14_0.Vb2_2.n12 185
R8709 two_stage_opamp_dummy_magic_14_0.Vb2_2.n26 two_stage_opamp_dummy_magic_14_0.Vb2_2.n25 185
R8710 two_stage_opamp_dummy_magic_14_0.Vb2_2.n27 two_stage_opamp_dummy_magic_14_0.Vb2_2.n26 185
R8711 two_stage_opamp_dummy_magic_14_0.Vb2_2.n24 two_stage_opamp_dummy_magic_14_0.Vb2_2.n16 185
R8712 two_stage_opamp_dummy_magic_14_0.Vb2_2.n22 two_stage_opamp_dummy_magic_14_0.Vb2_2.n21 185
R8713 two_stage_opamp_dummy_magic_14_0.Vb2_2.n20 two_stage_opamp_dummy_magic_14_0.Vb2_2.n19 185
R8714 two_stage_opamp_dummy_magic_14_0.Vb2_2.n38 two_stage_opamp_dummy_magic_14_0.Vb2_2.n37 185
R8715 two_stage_opamp_dummy_magic_14_0.Vb2_2.n39 two_stage_opamp_dummy_magic_14_0.Vb2_2.n38 185
R8716 two_stage_opamp_dummy_magic_14_0.Vb2_2.n35 two_stage_opamp_dummy_magic_14_0.Vb2_2.n10 185
R8717 two_stage_opamp_dummy_magic_14_0.Vb2_2.n7 two_stage_opamp_dummy_magic_14_0.Vb2_2.n3 185
R8718 two_stage_opamp_dummy_magic_14_0.Vb2_2.n44 two_stage_opamp_dummy_magic_14_0.Vb2_2.n4 185
R8719 two_stage_opamp_dummy_magic_14_0.Vb2_2.n43 two_stage_opamp_dummy_magic_14_0.Vb2_2.n5 185
R8720 two_stage_opamp_dummy_magic_14_0.Vb2_2.n42 two_stage_opamp_dummy_magic_14_0.Vb2_2.n6 185
R8721 two_stage_opamp_dummy_magic_14_0.Vb2_2.n39 two_stage_opamp_dummy_magic_14_0.Vb2_2.t5 170.513
R8722 two_stage_opamp_dummy_magic_14_0.Vb2_2.n27 two_stage_opamp_dummy_magic_14_0.Vb2_2.t8 170.513
R8723 two_stage_opamp_dummy_magic_14_0.Vb2_2.n32 two_stage_opamp_dummy_magic_14_0.Vb2_2.n1 155.304
R8724 two_stage_opamp_dummy_magic_14_0.Vb2_2.n26 two_stage_opamp_dummy_magic_14_0.Vb2_2.n13 150
R8725 two_stage_opamp_dummy_magic_14_0.Vb2_2.n26 two_stage_opamp_dummy_magic_14_0.Vb2_2.n16 150
R8726 two_stage_opamp_dummy_magic_14_0.Vb2_2.n21 two_stage_opamp_dummy_magic_14_0.Vb2_2.n20 150
R8727 two_stage_opamp_dummy_magic_14_0.Vb2_2.n38 two_stage_opamp_dummy_magic_14_0.Vb2_2.n10 150
R8728 two_stage_opamp_dummy_magic_14_0.Vb2_2.n7 two_stage_opamp_dummy_magic_14_0.Vb2_2.n4 150
R8729 two_stage_opamp_dummy_magic_14_0.Vb2_2.n6 two_stage_opamp_dummy_magic_14_0.Vb2_2.n5 150
R8730 two_stage_opamp_dummy_magic_14_0.Vb2_2.t0 two_stage_opamp_dummy_magic_14_0.Vb2_2.t5 146.155
R8731 two_stage_opamp_dummy_magic_14_0.Vb2_2.t8 two_stage_opamp_dummy_magic_14_0.Vb2_2.t0 146.155
R8732 two_stage_opamp_dummy_magic_14_0.Vb2_2.n28 two_stage_opamp_dummy_magic_14_0.Vb2_2.n27 65.8183
R8733 two_stage_opamp_dummy_magic_14_0.Vb2_2.n27 two_stage_opamp_dummy_magic_14_0.Vb2_2.n14 65.8183
R8734 two_stage_opamp_dummy_magic_14_0.Vb2_2.n27 two_stage_opamp_dummy_magic_14_0.Vb2_2.n15 65.8183
R8735 two_stage_opamp_dummy_magic_14_0.Vb2_2.n39 two_stage_opamp_dummy_magic_14_0.Vb2_2.n8 65.8183
R8736 two_stage_opamp_dummy_magic_14_0.Vb2_2.n39 two_stage_opamp_dummy_magic_14_0.Vb2_2.n9 65.8183
R8737 two_stage_opamp_dummy_magic_14_0.Vb2_2.n40 two_stage_opamp_dummy_magic_14_0.Vb2_2.n39 65.8183
R8738 two_stage_opamp_dummy_magic_14_0.Vb2_2.n16 two_stage_opamp_dummy_magic_14_0.Vb2_2.n14 53.3664
R8739 two_stage_opamp_dummy_magic_14_0.Vb2_2.n20 two_stage_opamp_dummy_magic_14_0.Vb2_2.n15 53.3664
R8740 two_stage_opamp_dummy_magic_14_0.Vb2_2.n28 two_stage_opamp_dummy_magic_14_0.Vb2_2.n13 53.3664
R8741 two_stage_opamp_dummy_magic_14_0.Vb2_2.n21 two_stage_opamp_dummy_magic_14_0.Vb2_2.n14 53.3664
R8742 two_stage_opamp_dummy_magic_14_0.Vb2_2.n10 two_stage_opamp_dummy_magic_14_0.Vb2_2.n8 53.3664
R8743 two_stage_opamp_dummy_magic_14_0.Vb2_2.n9 two_stage_opamp_dummy_magic_14_0.Vb2_2.n4 53.3664
R8744 two_stage_opamp_dummy_magic_14_0.Vb2_2.n40 two_stage_opamp_dummy_magic_14_0.Vb2_2.n6 53.3664
R8745 two_stage_opamp_dummy_magic_14_0.Vb2_2.n8 two_stage_opamp_dummy_magic_14_0.Vb2_2.n7 53.3664
R8746 two_stage_opamp_dummy_magic_14_0.Vb2_2.n9 two_stage_opamp_dummy_magic_14_0.Vb2_2.n5 53.3664
R8747 two_stage_opamp_dummy_magic_14_0.Vb2_2.n30 two_stage_opamp_dummy_magic_14_0.Vb2_2.n29 22.8576
R8748 two_stage_opamp_dummy_magic_14_0.Vb2_2.n37 two_stage_opamp_dummy_magic_14_0.Vb2_2.n34 22.8576
R8749 two_stage_opamp_dummy_magic_14_0.Vb2_2.n31 two_stage_opamp_dummy_magic_14_0.Vb2_2.t3 21.8894
R8750 two_stage_opamp_dummy_magic_14_0.Vb2_2.n31 two_stage_opamp_dummy_magic_14_0.Vb2_2.t2 21.8894
R8751 two_stage_opamp_dummy_magic_14_0.Vb2_2.n33 two_stage_opamp_dummy_magic_14_0.Vb2_2.n30 14.4255
R8752 two_stage_opamp_dummy_magic_14_0.Vb2_2.n34 two_stage_opamp_dummy_magic_14_0.Vb2_2.n33 14.0505
R8753 two_stage_opamp_dummy_magic_14_0.Vb2_2.n11 two_stage_opamp_dummy_magic_14_0.Vb2_2.t9 11.2576
R8754 two_stage_opamp_dummy_magic_14_0.Vb2_2.t6 two_stage_opamp_dummy_magic_14_0.Vb2_2.n1 11.2576
R8755 two_stage_opamp_dummy_magic_14_0.Vb2_2.n1 two_stage_opamp_dummy_magic_14_0.Vb2_2.t1 11.2576
R8756 two_stage_opamp_dummy_magic_14_0.Vb2_2.n29 two_stage_opamp_dummy_magic_14_0.Vb2_2.n12 9.14336
R8757 two_stage_opamp_dummy_magic_14_0.Vb2_2.n25 two_stage_opamp_dummy_magic_14_0.Vb2_2.n24 9.14336
R8758 two_stage_opamp_dummy_magic_14_0.Vb2_2.n22 two_stage_opamp_dummy_magic_14_0.Vb2_2.n19 9.14336
R8759 two_stage_opamp_dummy_magic_14_0.Vb2_2.n35 two_stage_opamp_dummy_magic_14_0.Vb2_2.n3 9.14336
R8760 two_stage_opamp_dummy_magic_14_0.Vb2_2.n44 two_stage_opamp_dummy_magic_14_0.Vb2_2.n3 9.14336
R8761 two_stage_opamp_dummy_magic_14_0.Vb2_2.n44 two_stage_opamp_dummy_magic_14_0.Vb2_2.n43 9.14336
R8762 two_stage_opamp_dummy_magic_14_0.Vb2_2.n43 two_stage_opamp_dummy_magic_14_0.Vb2_2.n42 9.14336
R8763 two_stage_opamp_dummy_magic_14_0.Vb2_2.n37 two_stage_opamp_dummy_magic_14_0.Vb2_2.n36 5.33286
R8764 two_stage_opamp_dummy_magic_14_0.Vb2_2.n17 two_stage_opamp_dummy_magic_14_0.Vb2_2.n12 4.53698
R8765 two_stage_opamp_dummy_magic_14_0.Vb2_2.n24 two_stage_opamp_dummy_magic_14_0.Vb2_2.n23 4.53698
R8766 two_stage_opamp_dummy_magic_14_0.Vb2_2.n19 two_stage_opamp_dummy_magic_14_0.Vb2_2.n18 4.53698
R8767 two_stage_opamp_dummy_magic_14_0.Vb2_2.n25 two_stage_opamp_dummy_magic_14_0.Vb2_2.n17 4.53698
R8768 two_stage_opamp_dummy_magic_14_0.Vb2_2.n23 two_stage_opamp_dummy_magic_14_0.Vb2_2.n22 4.53698
R8769 two_stage_opamp_dummy_magic_14_0.Vb2_2.n33 two_stage_opamp_dummy_magic_14_0.Vb2_2.n32 4.5005
R8770 two_stage_opamp_dummy_magic_14_0.Vb2_2.n36 two_stage_opamp_dummy_magic_14_0.Vb2_2.n35 3.75335
R8771 two_stage_opamp_dummy_magic_14_0.Vb2_2.n42 two_stage_opamp_dummy_magic_14_0.Vb2_2.n41 3.75335
R8772 a_13180_23838.t0 a_13180_23838.t1 178.133
R8773 a_14170_5524.t0 a_14170_5524.t1 262.248
R8774 a_14290_5524.t0 a_14290_5524.t1 169.905
C0 bgr_0.NFET_GATE_10uA bgr_0.START_UP_NFET1 0.351171f
C1 two_stage_opamp_dummy_magic_14_0.V_err_mir_p VDDA 0.671509f
C2 two_stage_opamp_dummy_magic_14_0.V_err_gate two_stage_opamp_dummy_magic_14_0.V_err_mir_p 0.429395f
C3 bgr_0.NFET_GATE_10uA two_stage_opamp_dummy_magic_14_0.Vb2 0.538556f
C4 bgr_0.START_UP_NFET1 VDDA 0.167059f
C5 two_stage_opamp_dummy_magic_14_0.Vb2 VDDA 1.44171f
C6 two_stage_opamp_dummy_magic_14_0.Vb2 two_stage_opamp_dummy_magic_14_0.V_err_gate 2.06924f
C7 two_stage_opamp_dummy_magic_14_0.cap_res_X VOUT+ 0.037134f
C8 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref VDDA 2.40167f
C9 two_stage_opamp_dummy_magic_14_0.V_err_gate two_stage_opamp_dummy_magic_14_0.V_err_amp_ref 0.804474f
C10 bgr_0.START_UP_NFET1 bgr_0.START_UP 0.145663f
C11 two_stage_opamp_dummy_magic_14_0.Vb2 bgr_0.START_UP 0.08188f
C12 bgr_0.START_UP two_stage_opamp_dummy_magic_14_0.V_err_amp_ref 1.36583f
C13 two_stage_opamp_dummy_magic_14_0.cap_res_X VOUT- 51.0174f
C14 two_stage_opamp_dummy_magic_14_0.Vb2 two_stage_opamp_dummy_magic_14_0.V_tail_gate 0.084214f
C15 VOUT+ VOUT- 0.397591f
C16 bgr_0.PFET_GATE_10uA two_stage_opamp_dummy_magic_14_0.cap_res_X 0.011459f
C17 two_stage_opamp_dummy_magic_14_0.VD4 VOUT+ 0.023279f
C18 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter VDDA 0.046803f
C19 bgr_0.V_TOP bgr_0.1st_Vout_1 2.47405f
C20 two_stage_opamp_dummy_magic_14_0.cap_res_X VDDA 0.39294f
C21 two_stage_opamp_dummy_magic_14_0.V_err_gate two_stage_opamp_dummy_magic_14_0.cap_res_X 0.333809f
C22 two_stage_opamp_dummy_magic_14_0.VD2 VIN+ 1.01398f
C23 VIN- li_11100_5020# 0.024834f
C24 VOUT+ VDDA 5.84806f
C25 two_stage_opamp_dummy_magic_14_0.Vb2 m1_10050_19490# 0.08176f
C26 two_stage_opamp_dummy_magic_14_0.V_tail_gate two_stage_opamp_dummy_magic_14_0.cap_res_X 0.245861f
C27 VOUT- VDDA 5.85106f
C28 two_stage_opamp_dummy_magic_14_0.V_err_gate VOUT- 0.040291f
C29 bgr_0.V_TOP two_stage_opamp_dummy_magic_14_0.Vb2 0.936691f
C30 bgr_0.V_TOP two_stage_opamp_dummy_magic_14_0.V_err_amp_ref 0.583702f
C31 two_stage_opamp_dummy_magic_14_0.Vb2 bgr_0.1st_Vout_1 0.042752f
C32 two_stage_opamp_dummy_magic_14_0.VD4 VDDA 4.39238f
C33 bgr_0.NFET_GATE_10uA bgr_0.PFET_GATE_10uA 0.012365f
C34 two_stage_opamp_dummy_magic_14_0.V_tail_gate two_stage_opamp_dummy_magic_14_0.VD2 0.023117f
C35 bgr_0.PFET_GATE_10uA VDDA 7.97055f
C36 two_stage_opamp_dummy_magic_14_0.V_tail_gate VOUT- 0.020352f
C37 VIN+ VIN- 0.141796f
C38 bgr_0.NFET_GATE_10uA VDDA 0.818988f
C39 bgr_0.NFET_GATE_10uA two_stage_opamp_dummy_magic_14_0.V_err_gate 3.50895f
C40 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter m1_10050_19490# 0.013969f
C41 two_stage_opamp_dummy_magic_14_0.V_err_gate VDDA 1.61242f
C42 bgr_0.PFET_GATE_10uA two_stage_opamp_dummy_magic_14_0.V_tail_gate 0.269369f
C43 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref two_stage_opamp_dummy_magic_14_0.V_err_mir_p 0.047419f
C44 bgr_0.NFET_GATE_10uA bgr_0.START_UP 1.64177f
C45 two_stage_opamp_dummy_magic_14_0.VD2 li_9020_5020# 0.073986f
C46 two_stage_opamp_dummy_magic_14_0.V_tail_gate VIN+ 0.055521f
C47 bgr_0.START_UP VDDA 1.09181f
C48 bgr_0.NFET_GATE_10uA two_stage_opamp_dummy_magic_14_0.V_tail_gate 0.038519f
C49 bgr_0.V_TOP bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.055802f
C50 two_stage_opamp_dummy_magic_14_0.V_tail_gate VDDA 3.41106f
C51 two_stage_opamp_dummy_magic_14_0.V_err_gate two_stage_opamp_dummy_magic_14_0.V_tail_gate 0.25337f
C52 two_stage_opamp_dummy_magic_14_0.V_tail_gate VIN- 0.15864f
C53 VIN+ li_9020_5020# 0.024834f
C54 m1_4880_3600# m2_4880_3600# 0.016063f
C55 bgr_0.V_TOP m2_10730_16580# 0.012f
C56 two_stage_opamp_dummy_magic_14_0.Vb2 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.01158f
C57 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.011335f
C58 two_stage_opamp_dummy_magic_14_0.Vb2 two_stage_opamp_dummy_magic_14_0.cap_res_X 0.615754f
C59 bgr_0.1st_Vout_1 m2_10730_16580# 0.075543f
C60 bgr_0.PFET_GATE_10uA m2_9370_16580# 0.012f
C61 bgr_0.V_TOP bgr_0.PFET_GATE_10uA 0.221314f
C62 two_stage_opamp_dummy_magic_14_0.V_err_gate m1_10050_19490# 0.091711f
C63 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref VOUT+ 0.041822f
C64 bgr_0.V_TOP bgr_0.NFET_GATE_10uA 0.052756f
C65 bgr_0.V_TOP VDDA 13.2374f
C66 bgr_0.NFET_GATE_10uA bgr_0.1st_Vout_1 0.03875f
C67 bgr_0.V_TOP two_stage_opamp_dummy_magic_14_0.V_err_gate 0.08195f
C68 bgr_0.1st_Vout_1 VDDA 0.896465f
C69 two_stage_opamp_dummy_magic_14_0.V_err_gate bgr_0.1st_Vout_1 0.041119f
C70 two_stage_opamp_dummy_magic_14_0.Vb2 VOUT- 0.058721f
C71 two_stage_opamp_dummy_magic_14_0.VD4 two_stage_opamp_dummy_magic_14_0.V_err_mir_p 0.0195f
C72 bgr_0.V_TOP bgr_0.START_UP 0.792764f
C73 two_stage_opamp_dummy_magic_14_0.Vb2 two_stage_opamp_dummy_magic_14_0.VD4 1.23597f
C74 bgr_0.START_UP bgr_0.1st_Vout_1 0.04354f
C75 two_stage_opamp_dummy_magic_14_0.VD4 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref 0.50647f
C76 bgr_0.START_UP_NFET1 bgr_0.PFET_GATE_10uA 0.0108f
C77 bgr_0.PFET_GATE_10uA two_stage_opamp_dummy_magic_14_0.V_err_amp_ref 1.69394f
C78 VIN- GNDA 1.44071f
C79 VIN+ GNDA 1.44759f
C80 VOUT- GNDA 15.84803f
C81 VOUT+ GNDA 15.878568f
C82 VDDA GNDA 0.121009p
C83 m2_4880_3600# GNDA 0.05269f $ **FLOATING
C84 m2_10730_16580# GNDA 0.0105f $ **FLOATING
C85 m2_9370_16580# GNDA 0.010002f $ **FLOATING
C86 m1_4880_3600# GNDA 0.059696f $ **FLOATING
C87 m1_10050_19490# GNDA 0.259273f $ **FLOATING
C88 li_11100_5020# GNDA 0.019798f $ **FLOATING
C89 li_9020_5020# GNDA 0.019798f $ **FLOATING
C90 two_stage_opamp_dummy_magic_14_0.VD2 GNDA 2.00032f
C91 two_stage_opamp_dummy_magic_14_0.cap_res_X GNDA 32.97633f
C92 two_stage_opamp_dummy_magic_14_0.V_err_mir_p GNDA 0.098639f
C93 two_stage_opamp_dummy_magic_14_0.V_tail_gate GNDA 8.759613f
C94 bgr_0.1st_Vout_1 GNDA 7.823503f
C95 bgr_0.START_UP GNDA 5.877827f
C96 bgr_0.START_UP_NFET1 GNDA 4.29564f
C97 two_stage_opamp_dummy_magic_14_0.V_err_gate GNDA 7.80031f
C98 two_stage_opamp_dummy_magic_14_0.Vb2 GNDA 7.393853f
C99 bgr_0.NFET_GATE_10uA GNDA 7.92412f
C100 bgr_0.V_TOP GNDA 9.96016f
C101 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter GNDA 17.8947f
C102 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref GNDA 6.84468f
C103 bgr_0.PFET_GATE_10uA GNDA 6.580853f
C104 two_stage_opamp_dummy_magic_14_0.VD4 GNDA 4.888977f
C105 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.t15 GNDA 0.01637f
C106 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.t12 GNDA 0.01637f
C107 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.n0 GNDA 0.041034f
C108 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.t10 GNDA 0.01637f
C109 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.t13 GNDA 0.01637f
C110 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.n1 GNDA 0.040818f
C111 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.n2 GNDA 0.362787f
C112 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.t11 GNDA 0.01637f
C113 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.t14 GNDA 0.01637f
C114 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.n3 GNDA 0.03274f
C115 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.n4 GNDA 0.060887f
C116 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.t16 GNDA 0.206157f
C117 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.t1 GNDA 0.03274f
C118 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.t5 GNDA 0.03274f
C119 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.n5 GNDA 0.097293f
C120 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.t0 GNDA 0.03274f
C121 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.t9 GNDA 0.03274f
C122 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.n6 GNDA 0.096862f
C123 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.n7 GNDA 0.331325f
C124 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.t2 GNDA 0.03274f
C125 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.t6 GNDA 0.03274f
C126 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.n8 GNDA 0.096862f
C127 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.n9 GNDA 0.171607f
C128 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.t3 GNDA 0.03274f
C129 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.t7 GNDA 0.03274f
C130 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.n10 GNDA 0.096862f
C131 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.n11 GNDA 0.171607f
C132 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.t4 GNDA 0.03274f
C133 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.t8 GNDA 0.03274f
C134 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.n12 GNDA 0.096862f
C135 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.n13 GNDA 0.239231f
C136 two_stage_opamp_dummy_magic_14_0.V_CMFB_S1.n14 GNDA 1.32734f
C137 bgr_0.V_CMFB_S1 GNDA 1.1041f
C138 bgr_0.START_UP.t4 GNDA 1.06745f
C139 bgr_0.START_UP.t5 GNDA 0.02806f
C140 bgr_0.START_UP.n0 GNDA 0.714928f
C141 bgr_0.START_UP.t0 GNDA 0.026778f
C142 bgr_0.START_UP.t2 GNDA 0.026778f
C143 bgr_0.START_UP.n1 GNDA 0.097147f
C144 bgr_0.START_UP.t1 GNDA 0.026778f
C145 bgr_0.START_UP.t3 GNDA 0.026778f
C146 bgr_0.START_UP.n2 GNDA 0.08937f
C147 bgr_0.START_UP.n3 GNDA 0.462855f
C148 bgr_0.START_UP.t7 GNDA 0.010062f
C149 bgr_0.START_UP.t6 GNDA 0.010062f
C150 bgr_0.START_UP.n4 GNDA 0.028407f
C151 bgr_0.START_UP.n5 GNDA 0.260836f
C152 two_stage_opamp_dummy_magic_14_0.VD4.t34 GNDA 0.030951f
C153 two_stage_opamp_dummy_magic_14_0.VD4.t37 GNDA 0.030951f
C154 two_stage_opamp_dummy_magic_14_0.VD4.n0 GNDA 0.108702f
C155 two_stage_opamp_dummy_magic_14_0.VD4.t29 GNDA 0.030951f
C156 two_stage_opamp_dummy_magic_14_0.VD4.t32 GNDA 0.030951f
C157 two_stage_opamp_dummy_magic_14_0.VD4.n1 GNDA 0.108329f
C158 two_stage_opamp_dummy_magic_14_0.VD4.n2 GNDA 0.202138f
C159 two_stage_opamp_dummy_magic_14_0.VD4.t27 GNDA 0.030951f
C160 two_stage_opamp_dummy_magic_14_0.VD4.t26 GNDA 0.030951f
C161 two_stage_opamp_dummy_magic_14_0.VD4.n3 GNDA 0.108329f
C162 two_stage_opamp_dummy_magic_14_0.VD4.n4 GNDA 0.104793f
C163 two_stage_opamp_dummy_magic_14_0.VD4.t33 GNDA 0.030951f
C164 two_stage_opamp_dummy_magic_14_0.VD4.t35 GNDA 0.030951f
C165 two_stage_opamp_dummy_magic_14_0.VD4.n5 GNDA 0.108329f
C166 two_stage_opamp_dummy_magic_14_0.VD4.n6 GNDA 0.104793f
C167 two_stage_opamp_dummy_magic_14_0.VD4.t28 GNDA 0.030951f
C168 two_stage_opamp_dummy_magic_14_0.VD4.t31 GNDA 0.030951f
C169 two_stage_opamp_dummy_magic_14_0.VD4.n7 GNDA 0.108329f
C170 two_stage_opamp_dummy_magic_14_0.VD4.n8 GNDA 0.104793f
C171 two_stage_opamp_dummy_magic_14_0.VD4.t36 GNDA 0.030951f
C172 two_stage_opamp_dummy_magic_14_0.VD4.t30 GNDA 0.030951f
C173 two_stage_opamp_dummy_magic_14_0.VD4.n9 GNDA 0.108329f
C174 two_stage_opamp_dummy_magic_14_0.VD4.n10 GNDA 0.153987f
C175 two_stage_opamp_dummy_magic_14_0.VD4.t15 GNDA 0.030951f
C176 two_stage_opamp_dummy_magic_14_0.VD4.t19 GNDA 0.030951f
C177 two_stage_opamp_dummy_magic_14_0.VD4.n11 GNDA 0.10726f
C178 two_stage_opamp_dummy_magic_14_0.VD4.n12 GNDA 0.104977f
C179 two_stage_opamp_dummy_magic_14_0.VD4.t22 GNDA 0.030951f
C180 two_stage_opamp_dummy_magic_14_0.VD4.n13 GNDA 0.092854f
C181 two_stage_opamp_dummy_magic_14_0.VD4.n14 GNDA 0.030951f
C182 two_stage_opamp_dummy_magic_14_0.VD4.n15 GNDA 0.017686f
C183 two_stage_opamp_dummy_magic_14_0.VD4.n18 GNDA 0.014321f
C184 two_stage_opamp_dummy_magic_14_0.VD4.n19 GNDA 0.017686f
C185 two_stage_opamp_dummy_magic_14_0.VD4.t23 GNDA 0.054268f
C186 two_stage_opamp_dummy_magic_14_0.VD4.t5 GNDA 0.030951f
C187 two_stage_opamp_dummy_magic_14_0.VD4.t9 GNDA 0.030951f
C188 two_stage_opamp_dummy_magic_14_0.VD4.n20 GNDA 0.10726f
C189 two_stage_opamp_dummy_magic_14_0.VD4.n21 GNDA 0.104977f
C190 two_stage_opamp_dummy_magic_14_0.VD4.t1 GNDA 0.030951f
C191 two_stage_opamp_dummy_magic_14_0.VD4.t3 GNDA 0.030951f
C192 two_stage_opamp_dummy_magic_14_0.VD4.n22 GNDA 0.10726f
C193 two_stage_opamp_dummy_magic_14_0.VD4.n23 GNDA 0.104977f
C194 two_stage_opamp_dummy_magic_14_0.VD4.t13 GNDA 0.030951f
C195 two_stage_opamp_dummy_magic_14_0.VD4.t17 GNDA 0.030951f
C196 two_stage_opamp_dummy_magic_14_0.VD4.n24 GNDA 0.10726f
C197 two_stage_opamp_dummy_magic_14_0.VD4.n25 GNDA 0.104977f
C198 two_stage_opamp_dummy_magic_14_0.VD4.t11 GNDA 0.030951f
C199 two_stage_opamp_dummy_magic_14_0.VD4.t7 GNDA 0.030951f
C200 two_stage_opamp_dummy_magic_14_0.VD4.n26 GNDA 0.10726f
C201 two_stage_opamp_dummy_magic_14_0.VD4.n27 GNDA 0.134403f
C202 two_stage_opamp_dummy_magic_14_0.VD4.n28 GNDA 0.046089f
C203 two_stage_opamp_dummy_magic_14_0.VD4.n29 GNDA 0.030951f
C204 two_stage_opamp_dummy_magic_14_0.VD4.n31 GNDA 0.030951f
C205 two_stage_opamp_dummy_magic_14_0.VD4.n32 GNDA 0.017686f
C206 two_stage_opamp_dummy_magic_14_0.VD4.n33 GNDA 0.017686f
C207 two_stage_opamp_dummy_magic_14_0.VD4.n34 GNDA 0.030951f
C208 two_stage_opamp_dummy_magic_14_0.VD4.n36 GNDA 0.030951f
C209 two_stage_opamp_dummy_magic_14_0.VD4.n37 GNDA 0.017686f
C210 two_stage_opamp_dummy_magic_14_0.VD4.n38 GNDA 0.017686f
C211 two_stage_opamp_dummy_magic_14_0.VD4.n39 GNDA 0.030951f
C212 two_stage_opamp_dummy_magic_14_0.VD4.n40 GNDA 0.031222f
C213 two_stage_opamp_dummy_magic_14_0.VD4.t25 GNDA 0.030951f
C214 two_stage_opamp_dummy_magic_14_0.VD4.n41 GNDA 0.092854f
C215 two_stage_opamp_dummy_magic_14_0.VD4.n42 GNDA 0.029837f
C216 two_stage_opamp_dummy_magic_14_0.VD4.n43 GNDA 0.017686f
C217 two_stage_opamp_dummy_magic_14_0.VD4.n44 GNDA 0.258664f
C218 two_stage_opamp_dummy_magic_14_0.VD4.t24 GNDA 0.224175f
C219 two_stage_opamp_dummy_magic_14_0.VD4.t10 GNDA 0.206931f
C220 two_stage_opamp_dummy_magic_14_0.VD4.t6 GNDA 0.206931f
C221 two_stage_opamp_dummy_magic_14_0.VD4.t12 GNDA 0.206931f
C222 two_stage_opamp_dummy_magic_14_0.VD4.t16 GNDA 0.206931f
C223 two_stage_opamp_dummy_magic_14_0.VD4.t0 GNDA 0.206931f
C224 two_stage_opamp_dummy_magic_14_0.VD4.t2 GNDA 0.206931f
C225 two_stage_opamp_dummy_magic_14_0.VD4.t4 GNDA 0.206931f
C226 two_stage_opamp_dummy_magic_14_0.VD4.t8 GNDA 0.206931f
C227 two_stage_opamp_dummy_magic_14_0.VD4.t14 GNDA 0.206931f
C228 two_stage_opamp_dummy_magic_14_0.VD4.t18 GNDA 0.206931f
C229 two_stage_opamp_dummy_magic_14_0.VD4.t21 GNDA 0.224175f
C230 two_stage_opamp_dummy_magic_14_0.VD4.n46 GNDA 0.014321f
C231 two_stage_opamp_dummy_magic_14_0.VD4.n47 GNDA 0.017686f
C232 two_stage_opamp_dummy_magic_14_0.VD4.n49 GNDA 0.031222f
C233 two_stage_opamp_dummy_magic_14_0.VD4.n50 GNDA 0.030951f
C234 two_stage_opamp_dummy_magic_14_0.VD4.n51 GNDA 0.017686f
C235 two_stage_opamp_dummy_magic_14_0.VD4.n52 GNDA 0.017686f
C236 two_stage_opamp_dummy_magic_14_0.VD4.n53 GNDA 0.030951f
C237 two_stage_opamp_dummy_magic_14_0.VD4.n55 GNDA 0.030951f
C238 two_stage_opamp_dummy_magic_14_0.VD4.n56 GNDA 0.030951f
C239 two_stage_opamp_dummy_magic_14_0.VD4.n57 GNDA 0.017686f
C240 two_stage_opamp_dummy_magic_14_0.VD4.n58 GNDA 0.258664f
C241 two_stage_opamp_dummy_magic_14_0.VD4.n59 GNDA 0.013727f
C242 two_stage_opamp_dummy_magic_14_0.VD4.n60 GNDA 0.033797f
C243 two_stage_opamp_dummy_magic_14_0.VD4.t20 GNDA 0.054268f
C244 two_stage_opamp_dummy_magic_14_0.VD4.n61 GNDA 0.044756f
C245 two_stage_opamp_dummy_magic_14_0.VD4.n62 GNDA 0.062101f
C246 two_stage_opamp_dummy_magic_14_0.VD4.n63 GNDA 0.087485f
C247 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.t13 GNDA 0.01637f
C248 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.t16 GNDA 0.01637f
C249 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.n0 GNDA 0.041052f
C250 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.t12 GNDA 0.01637f
C251 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.t11 GNDA 0.01637f
C252 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.n1 GNDA 0.040835f
C253 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.n2 GNDA 0.363013f
C254 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.t15 GNDA 0.01637f
C255 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.t14 GNDA 0.01637f
C256 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.n3 GNDA 0.03274f
C257 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.n4 GNDA 0.060861f
C258 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.t10 GNDA 0.206157f
C259 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.t1 GNDA 0.03274f
C260 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.t5 GNDA 0.03274f
C261 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.n5 GNDA 0.097293f
C262 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.t0 GNDA 0.03274f
C263 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.t4 GNDA 0.03274f
C264 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.n6 GNDA 0.096862f
C265 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.n7 GNDA 0.331325f
C266 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.t9 GNDA 0.03274f
C267 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.t7 GNDA 0.03274f
C268 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.n8 GNDA 0.096862f
C269 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.n9 GNDA 0.171607f
C270 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.t2 GNDA 0.03274f
C271 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.t6 GNDA 0.03274f
C272 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.n10 GNDA 0.096862f
C273 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.n11 GNDA 0.171607f
C274 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.t8 GNDA 0.03274f
C275 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.t3 GNDA 0.03274f
C276 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.n12 GNDA 0.096862f
C277 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.n13 GNDA 0.239231f
C278 two_stage_opamp_dummy_magic_14_0.V_CMFB_S3.n14 GNDA 1.32734f
C279 bgr_0.V_CMFB_S3 GNDA 1.10386f
C280 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.t14 GNDA 0.020156f
C281 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.t12 GNDA 0.020156f
C282 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.n0 GNDA 0.073261f
C283 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.t13 GNDA 0.020156f
C284 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.t11 GNDA 0.020156f
C285 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.n1 GNDA 0.060879f
C286 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.n2 GNDA 1.18743f
C287 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.t10 GNDA 0.247627f
C288 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.t5 GNDA 0.060467f
C289 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.t9 GNDA 0.060467f
C290 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.n3 GNDA 0.252232f
C291 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.t4 GNDA 0.060467f
C292 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.t8 GNDA 0.060467f
C293 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.n4 GNDA 0.251304f
C294 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.n5 GNDA 0.345024f
C295 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.t3 GNDA 0.060467f
C296 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.t1 GNDA 0.060467f
C297 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.n6 GNDA 0.251304f
C298 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.n7 GNDA 0.18003f
C299 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.t6 GNDA 0.060467f
C300 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.t0 GNDA 0.060467f
C301 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.n8 GNDA 0.251304f
C302 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.n9 GNDA 0.18003f
C303 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.t2 GNDA 0.060467f
C304 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.t7 GNDA 0.060467f
C305 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.n10 GNDA 0.251304f
C306 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.n11 GNDA 0.249769f
C307 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.n12 GNDA 1.34239f
C308 two_stage_opamp_dummy_magic_14_0.V_CMFB_S4.n13 GNDA 1.98073f
C309 bgr_0.V_CMFB_S4 GNDA 0.010078f
C310 bgr_0.Vin-.n0 GNDA 0.069747f
C311 bgr_0.Vin-.n1 GNDA 0.316148f
C312 bgr_0.Vin-.t3 GNDA 0.027101f
C313 bgr_0.Vin-.t1 GNDA 0.027101f
C314 bgr_0.Vin-.n2 GNDA 0.094346f
C315 bgr_0.Vin-.t0 GNDA 0.027101f
C316 bgr_0.Vin-.t2 GNDA 0.027101f
C317 bgr_0.Vin-.n3 GNDA 0.090091f
C318 bgr_0.Vin-.n4 GNDA 0.386489f
C319 bgr_0.Vin-.n5 GNDA 0.027681f
C320 bgr_0.Vin-.n6 GNDA 0.366254f
C321 bgr_0.Vin-.t12 GNDA 0.022346f
C322 bgr_0.Vin-.n7 GNDA 0.026209f
C323 bgr_0.Vin-.n8 GNDA 0.021455f
C324 bgr_0.Vin-.n9 GNDA 0.021455f
C325 bgr_0.Vin-.n10 GNDA 0.036491f
C326 bgr_0.Vin-.n11 GNDA 0.497932f
C327 bgr_0.Vin-.t6 GNDA 0.117924f
C328 bgr_0.Vin-.n12 GNDA 0.655831f
C329 bgr_0.Vin-.n13 GNDA 1.07297f
C330 bgr_0.Vin-.n14 GNDA 0.471323f
C331 bgr_0.Vin-.t7 GNDA 0.261631f
C332 bgr_0.Vin-.n15 GNDA 0.069875f
C333 bgr_0.Vin-.n16 GNDA 0.119593f
C334 bgr_0.Vin-.n17 GNDA 0.07053f
C335 bgr_0.Vin-.n18 GNDA 0.579028f
C336 bgr_0.Vin-.n19 GNDA 0.358216f
C337 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_23.Emitter GNDA 0.086538f
C338 bgr_0.V_mir2.t7 GNDA 0.019293f
C339 bgr_0.V_mir2.n0 GNDA 0.025223f
C340 bgr_0.V_mir2.t14 GNDA 0.041163f
C341 bgr_0.V_mir2.n1 GNDA 0.027381f
C342 bgr_0.V_mir2.n2 GNDA 0.451535f
C343 bgr_0.V_mir2.n3 GNDA 0.146338f
C344 bgr_0.V_mir2.t4 GNDA 0.023151f
C345 bgr_0.V_mir2.t17 GNDA 0.023151f
C346 bgr_0.V_mir2.t20 GNDA 0.037369f
C347 bgr_0.V_mir2.n4 GNDA 0.041731f
C348 bgr_0.V_mir2.n5 GNDA 0.028507f
C349 bgr_0.V_mir2.t0 GNDA 0.02939f
C350 bgr_0.V_mir2.n6 GNDA 0.044354f
C351 bgr_0.V_mir2.t5 GNDA 0.019293f
C352 bgr_0.V_mir2.t1 GNDA 0.019293f
C353 bgr_0.V_mir2.n7 GNDA 0.044166f
C354 bgr_0.V_mir2.n8 GNDA 0.109943f
C355 bgr_0.V_mir2.t2 GNDA 0.023151f
C356 bgr_0.V_mir2.t18 GNDA 0.023151f
C357 bgr_0.V_mir2.t22 GNDA 0.037369f
C358 bgr_0.V_mir2.n9 GNDA 0.041731f
C359 bgr_0.V_mir2.n10 GNDA 0.028507f
C360 bgr_0.V_mir2.t8 GNDA 0.02939f
C361 bgr_0.V_mir2.n11 GNDA 0.044354f
C362 bgr_0.V_mir2.t3 GNDA 0.019293f
C363 bgr_0.V_mir2.t9 GNDA 0.019293f
C364 bgr_0.V_mir2.n12 GNDA 0.044166f
C365 bgr_0.V_mir2.n13 GNDA 0.111042f
C366 bgr_0.V_mir2.n14 GNDA 0.381359f
C367 bgr_0.V_mir2.n15 GNDA 0.051125f
C368 bgr_0.V_mir2.t6 GNDA 0.023151f
C369 bgr_0.V_mir2.t19 GNDA 0.023151f
C370 bgr_0.V_mir2.t21 GNDA 0.037369f
C371 bgr_0.V_mir2.n16 GNDA 0.041731f
C372 bgr_0.V_mir2.n17 GNDA 0.028507f
C373 bgr_0.V_mir2.t10 GNDA 0.02939f
C374 bgr_0.V_mir2.n18 GNDA 0.044354f
C375 bgr_0.V_mir2.n19 GNDA 0.085095f
C376 bgr_0.V_mir2.n20 GNDA 0.044166f
C377 bgr_0.V_mir2.t11 GNDA 0.019293f
C378 bgr_0.cap_res1.t11 GNDA 0.331712f
C379 bgr_0.cap_res1.t18 GNDA 0.349187f
C380 bgr_0.cap_res1.t15 GNDA 0.350452f
C381 bgr_0.cap_res1.t4 GNDA 0.331712f
C382 bgr_0.cap_res1.t14 GNDA 0.349187f
C383 bgr_0.cap_res1.t8 GNDA 0.350452f
C384 bgr_0.cap_res1.t10 GNDA 0.331712f
C385 bgr_0.cap_res1.t17 GNDA 0.349187f
C386 bgr_0.cap_res1.t13 GNDA 0.350452f
C387 bgr_0.cap_res1.t3 GNDA 0.331712f
C388 bgr_0.cap_res1.t12 GNDA 0.349187f
C389 bgr_0.cap_res1.t6 GNDA 0.350452f
C390 bgr_0.cap_res1.t19 GNDA 0.331712f
C391 bgr_0.cap_res1.t5 GNDA 0.349187f
C392 bgr_0.cap_res1.t0 GNDA 0.350452f
C393 bgr_0.cap_res1.n0 GNDA 0.23406f
C394 bgr_0.cap_res1.t16 GNDA 0.186395f
C395 bgr_0.cap_res1.n1 GNDA 0.253961f
C396 bgr_0.cap_res1.t1 GNDA 0.186395f
C397 bgr_0.cap_res1.n2 GNDA 0.253961f
C398 bgr_0.cap_res1.t7 GNDA 0.186395f
C399 bgr_0.cap_res1.n3 GNDA 0.253961f
C400 bgr_0.cap_res1.t2 GNDA 0.186395f
C401 bgr_0.cap_res1.n4 GNDA 0.253961f
C402 bgr_0.cap_res1.t9 GNDA 0.363549f
C403 bgr_0.cap_res1.t20 GNDA 0.08421f
C404 bgr_0.PFET_GATE_10uA.t28 GNDA 0.020856f
C405 bgr_0.PFET_GATE_10uA.t20 GNDA 0.030831f
C406 bgr_0.PFET_GATE_10uA.n0 GNDA 0.033972f
C407 bgr_0.PFET_GATE_10uA.t15 GNDA 0.020856f
C408 bgr_0.PFET_GATE_10uA.t21 GNDA 0.030831f
C409 bgr_0.PFET_GATE_10uA.n1 GNDA 0.033972f
C410 bgr_0.PFET_GATE_10uA.n2 GNDA 0.040878f
C411 bgr_0.PFET_GATE_10uA.t19 GNDA 0.020856f
C412 bgr_0.PFET_GATE_10uA.t12 GNDA 0.030831f
C413 bgr_0.PFET_GATE_10uA.n3 GNDA 0.033972f
C414 bgr_0.PFET_GATE_10uA.t26 GNDA 0.020856f
C415 bgr_0.PFET_GATE_10uA.t13 GNDA 0.030831f
C416 bgr_0.PFET_GATE_10uA.n4 GNDA 0.033972f
C417 bgr_0.PFET_GATE_10uA.n5 GNDA 0.034081f
C418 bgr_0.PFET_GATE_10uA.t7 GNDA 0.312465f
C419 bgr_0.PFET_GATE_10uA.t0 GNDA 0.021391f
C420 bgr_0.PFET_GATE_10uA.t8 GNDA 0.021391f
C421 bgr_0.PFET_GATE_10uA.n6 GNDA 0.054673f
C422 bgr_0.PFET_GATE_10uA.t2 GNDA 0.021391f
C423 bgr_0.PFET_GATE_10uA.t4 GNDA 0.021391f
C424 bgr_0.PFET_GATE_10uA.n7 GNDA 0.05326f
C425 bgr_0.PFET_GATE_10uA.n8 GNDA 0.520952f
C426 bgr_0.PFET_GATE_10uA.t3 GNDA 0.021391f
C427 bgr_0.PFET_GATE_10uA.t5 GNDA 0.021391f
C428 bgr_0.PFET_GATE_10uA.n9 GNDA 0.05326f
C429 bgr_0.PFET_GATE_10uA.n10 GNDA 0.295408f
C430 bgr_0.PFET_GATE_10uA.n11 GNDA 0.603055f
C431 bgr_0.PFET_GATE_10uA.t9 GNDA 0.021391f
C432 bgr_0.PFET_GATE_10uA.t1 GNDA 0.021391f
C433 bgr_0.PFET_GATE_10uA.n12 GNDA 0.05159f
C434 bgr_0.PFET_GATE_10uA.n13 GNDA 0.275411f
C435 bgr_0.PFET_GATE_10uA.t6 GNDA 0.464967f
C436 bgr_0.PFET_GATE_10uA.t27 GNDA 0.024114f
C437 bgr_0.PFET_GATE_10uA.t14 GNDA 0.024114f
C438 bgr_0.PFET_GATE_10uA.n14 GNDA 0.069715f
C439 bgr_0.PFET_GATE_10uA.n15 GNDA 1.91969f
C440 bgr_0.PFET_GATE_10uA.n16 GNDA 0.771508f
C441 bgr_0.PFET_GATE_10uA.n17 GNDA 0.759224f
C442 bgr_0.PFET_GATE_10uA.t11 GNDA 0.020856f
C443 bgr_0.PFET_GATE_10uA.t25 GNDA 0.020856f
C444 bgr_0.PFET_GATE_10uA.t18 GNDA 0.020856f
C445 bgr_0.PFET_GATE_10uA.t10 GNDA 0.020856f
C446 bgr_0.PFET_GATE_10uA.t24 GNDA 0.020856f
C447 bgr_0.PFET_GATE_10uA.t17 GNDA 0.030831f
C448 bgr_0.PFET_GATE_10uA.n18 GNDA 0.038154f
C449 bgr_0.PFET_GATE_10uA.n19 GNDA 0.027273f
C450 bgr_0.PFET_GATE_10uA.n20 GNDA 0.027273f
C451 bgr_0.PFET_GATE_10uA.n21 GNDA 0.027273f
C452 bgr_0.PFET_GATE_10uA.n22 GNDA 0.023091f
C453 bgr_0.PFET_GATE_10uA.t16 GNDA 0.020856f
C454 bgr_0.PFET_GATE_10uA.t23 GNDA 0.020856f
C455 bgr_0.PFET_GATE_10uA.t22 GNDA 0.020856f
C456 bgr_0.PFET_GATE_10uA.t29 GNDA 0.030831f
C457 bgr_0.PFET_GATE_10uA.n23 GNDA 0.038154f
C458 bgr_0.PFET_GATE_10uA.n24 GNDA 0.027273f
C459 bgr_0.PFET_GATE_10uA.n25 GNDA 0.023091f
C460 bgr_0.PFET_GATE_10uA.n26 GNDA 0.031695f
C461 two_stage_opamp_dummy_magic_14_0.Y.t1 GNDA 0.030836f
C462 two_stage_opamp_dummy_magic_14_0.Y.t6 GNDA 0.030836f
C463 two_stage_opamp_dummy_magic_14_0.Y.n0 GNDA 0.108297f
C464 two_stage_opamp_dummy_magic_14_0.Y.t10 GNDA 0.030836f
C465 two_stage_opamp_dummy_magic_14_0.Y.t9 GNDA 0.030836f
C466 two_stage_opamp_dummy_magic_14_0.Y.n1 GNDA 0.107926f
C467 two_stage_opamp_dummy_magic_14_0.Y.n2 GNDA 0.201386f
C468 two_stage_opamp_dummy_magic_14_0.Y.t5 GNDA 0.030836f
C469 two_stage_opamp_dummy_magic_14_0.Y.t2 GNDA 0.030836f
C470 two_stage_opamp_dummy_magic_14_0.Y.n3 GNDA 0.107926f
C471 two_stage_opamp_dummy_magic_14_0.Y.n4 GNDA 0.104403f
C472 two_stage_opamp_dummy_magic_14_0.Y.t4 GNDA 0.030836f
C473 two_stage_opamp_dummy_magic_14_0.Y.t8 GNDA 0.030836f
C474 two_stage_opamp_dummy_magic_14_0.Y.n5 GNDA 0.107926f
C475 two_stage_opamp_dummy_magic_14_0.Y.n6 GNDA 0.104403f
C476 two_stage_opamp_dummy_magic_14_0.Y.t3 GNDA 0.030836f
C477 two_stage_opamp_dummy_magic_14_0.Y.t11 GNDA 0.030836f
C478 two_stage_opamp_dummy_magic_14_0.Y.n7 GNDA 0.107926f
C479 two_stage_opamp_dummy_magic_14_0.Y.n8 GNDA 0.122969f
C480 two_stage_opamp_dummy_magic_14_0.Y.t7 GNDA 0.030836f
C481 two_stage_opamp_dummy_magic_14_0.Y.t0 GNDA 0.030836f
C482 two_stage_opamp_dummy_magic_14_0.Y.n9 GNDA 0.105762f
C483 two_stage_opamp_dummy_magic_14_0.Y.n10 GNDA 0.180803f
C484 two_stage_opamp_dummy_magic_14_0.Y.t40 GNDA 0.018502f
C485 two_stage_opamp_dummy_magic_14_0.Y.t54 GNDA 0.018502f
C486 two_stage_opamp_dummy_magic_14_0.Y.t37 GNDA 0.018502f
C487 two_stage_opamp_dummy_magic_14_0.Y.t51 GNDA 0.022466f
C488 two_stage_opamp_dummy_magic_14_0.Y.n11 GNDA 0.022466f
C489 two_stage_opamp_dummy_magic_14_0.Y.n12 GNDA 0.014537f
C490 two_stage_opamp_dummy_magic_14_0.Y.n13 GNDA 0.012822f
C491 two_stage_opamp_dummy_magic_14_0.Y.t26 GNDA 0.018502f
C492 two_stage_opamp_dummy_magic_14_0.Y.t31 GNDA 0.018502f
C493 two_stage_opamp_dummy_magic_14_0.Y.t48 GNDA 0.018502f
C494 two_stage_opamp_dummy_magic_14_0.Y.t34 GNDA 0.018502f
C495 two_stage_opamp_dummy_magic_14_0.Y.t29 GNDA 0.018502f
C496 two_stage_opamp_dummy_magic_14_0.Y.t44 GNDA 0.022466f
C497 two_stage_opamp_dummy_magic_14_0.Y.n14 GNDA 0.022466f
C498 two_stage_opamp_dummy_magic_14_0.Y.n15 GNDA 0.014537f
C499 two_stage_opamp_dummy_magic_14_0.Y.n16 GNDA 0.014537f
C500 two_stage_opamp_dummy_magic_14_0.Y.n17 GNDA 0.014537f
C501 two_stage_opamp_dummy_magic_14_0.Y.n18 GNDA 0.012822f
C502 two_stage_opamp_dummy_magic_14_0.Y.n19 GNDA 0.013323f
C503 two_stage_opamp_dummy_magic_14_0.Y.t28 GNDA 0.028413f
C504 two_stage_opamp_dummy_magic_14_0.Y.t42 GNDA 0.028413f
C505 two_stage_opamp_dummy_magic_14_0.Y.t25 GNDA 0.028413f
C506 two_stage_opamp_dummy_magic_14_0.Y.t39 GNDA 0.032301f
C507 two_stage_opamp_dummy_magic_14_0.Y.n20 GNDA 0.029151f
C508 two_stage_opamp_dummy_magic_14_0.Y.n21 GNDA 0.017841f
C509 two_stage_opamp_dummy_magic_14_0.Y.n22 GNDA 0.016126f
C510 two_stage_opamp_dummy_magic_14_0.Y.t43 GNDA 0.028413f
C511 two_stage_opamp_dummy_magic_14_0.Y.t50 GNDA 0.028413f
C512 two_stage_opamp_dummy_magic_14_0.Y.t36 GNDA 0.028413f
C513 two_stage_opamp_dummy_magic_14_0.Y.t53 GNDA 0.028413f
C514 two_stage_opamp_dummy_magic_14_0.Y.t46 GNDA 0.028413f
C515 two_stage_opamp_dummy_magic_14_0.Y.t32 GNDA 0.032301f
C516 two_stage_opamp_dummy_magic_14_0.Y.n23 GNDA 0.029151f
C517 two_stage_opamp_dummy_magic_14_0.Y.n24 GNDA 0.017841f
C518 two_stage_opamp_dummy_magic_14_0.Y.n25 GNDA 0.017841f
C519 two_stage_opamp_dummy_magic_14_0.Y.n26 GNDA 0.017841f
C520 two_stage_opamp_dummy_magic_14_0.Y.n27 GNDA 0.016126f
C521 two_stage_opamp_dummy_magic_14_0.Y.n28 GNDA 0.013323f
C522 two_stage_opamp_dummy_magic_14_0.Y.n29 GNDA 0.108435f
C523 two_stage_opamp_dummy_magic_14_0.Y.t23 GNDA 0.013215f
C524 two_stage_opamp_dummy_magic_14_0.Y.t21 GNDA 0.013215f
C525 two_stage_opamp_dummy_magic_14_0.Y.n30 GNDA 0.048379f
C526 two_stage_opamp_dummy_magic_14_0.Y.t13 GNDA 0.013215f
C527 two_stage_opamp_dummy_magic_14_0.Y.t14 GNDA 0.013215f
C528 two_stage_opamp_dummy_magic_14_0.Y.n31 GNDA 0.047973f
C529 two_stage_opamp_dummy_magic_14_0.Y.n32 GNDA 0.175886f
C530 two_stage_opamp_dummy_magic_14_0.Y.t15 GNDA 0.013215f
C531 two_stage_opamp_dummy_magic_14_0.Y.t20 GNDA 0.013215f
C532 two_stage_opamp_dummy_magic_14_0.Y.n33 GNDA 0.047973f
C533 two_stage_opamp_dummy_magic_14_0.Y.n34 GNDA 0.091229f
C534 two_stage_opamp_dummy_magic_14_0.Y.t16 GNDA 0.013215f
C535 two_stage_opamp_dummy_magic_14_0.Y.t22 GNDA 0.013215f
C536 two_stage_opamp_dummy_magic_14_0.Y.n35 GNDA 0.047973f
C537 two_stage_opamp_dummy_magic_14_0.Y.n36 GNDA 0.091229f
C538 two_stage_opamp_dummy_magic_14_0.Y.t18 GNDA 0.013215f
C539 two_stage_opamp_dummy_magic_14_0.Y.t19 GNDA 0.013215f
C540 two_stage_opamp_dummy_magic_14_0.Y.n37 GNDA 0.047973f
C541 two_stage_opamp_dummy_magic_14_0.Y.n38 GNDA 0.091229f
C542 two_stage_opamp_dummy_magic_14_0.Y.t17 GNDA 0.013215f
C543 two_stage_opamp_dummy_magic_14_0.Y.t24 GNDA 0.013215f
C544 two_stage_opamp_dummy_magic_14_0.Y.n39 GNDA 0.047973f
C545 two_stage_opamp_dummy_magic_14_0.Y.n40 GNDA 0.137095f
C546 two_stage_opamp_dummy_magic_14_0.Y.n41 GNDA 0.114012f
C547 two_stage_opamp_dummy_magic_14_0.Y.n42 GNDA 0.217579f
C548 two_stage_opamp_dummy_magic_14_0.Y.t38 GNDA 0.058148f
C549 two_stage_opamp_dummy_magic_14_0.Y.t52 GNDA 0.058148f
C550 two_stage_opamp_dummy_magic_14_0.Y.t35 GNDA 0.058148f
C551 two_stage_opamp_dummy_magic_14_0.Y.t49 GNDA 0.058148f
C552 two_stage_opamp_dummy_magic_14_0.Y.t33 GNDA 0.061932f
C553 two_stage_opamp_dummy_magic_14_0.Y.n43 GNDA 0.049078f
C554 two_stage_opamp_dummy_magic_14_0.Y.n44 GNDA 0.027753f
C555 two_stage_opamp_dummy_magic_14_0.Y.n45 GNDA 0.027753f
C556 two_stage_opamp_dummy_magic_14_0.Y.n46 GNDA 0.026044f
C557 two_stage_opamp_dummy_magic_14_0.Y.t45 GNDA 0.058148f
C558 two_stage_opamp_dummy_magic_14_0.Y.t30 GNDA 0.058148f
C559 two_stage_opamp_dummy_magic_14_0.Y.t47 GNDA 0.058148f
C560 two_stage_opamp_dummy_magic_14_0.Y.t41 GNDA 0.058148f
C561 two_stage_opamp_dummy_magic_14_0.Y.t27 GNDA 0.061932f
C562 two_stage_opamp_dummy_magic_14_0.Y.n47 GNDA 0.049078f
C563 two_stage_opamp_dummy_magic_14_0.Y.n48 GNDA 0.027753f
C564 two_stage_opamp_dummy_magic_14_0.Y.n49 GNDA 0.027753f
C565 two_stage_opamp_dummy_magic_14_0.Y.n50 GNDA 0.026044f
C566 two_stage_opamp_dummy_magic_14_0.Y.n51 GNDA 0.015843f
C567 two_stage_opamp_dummy_magic_14_0.Y.n52 GNDA 0.500074f
C568 two_stage_opamp_dummy_magic_14_0.Y.t12 GNDA 0.428359f
C569 two_stage_opamp_dummy_magic_14_0.Vb1.n0 GNDA 0.01994f
C570 two_stage_opamp_dummy_magic_14_0.Vb1.n1 GNDA 0.019806f
C571 two_stage_opamp_dummy_magic_14_0.Vb1.n2 GNDA 0.217486f
C572 two_stage_opamp_dummy_magic_14_0.Vb1.t1 GNDA 0.226679f
C573 two_stage_opamp_dummy_magic_14_0.Vb1.t2 GNDA 0.036499f
C574 two_stage_opamp_dummy_magic_14_0.Vb1.n3 GNDA 0.325297f
C575 two_stage_opamp_dummy_magic_14_0.Vb1.t22 GNDA 0.01223f
C576 two_stage_opamp_dummy_magic_14_0.Vb1.t12 GNDA 0.01223f
C577 two_stage_opamp_dummy_magic_14_0.Vb1.t21 GNDA 0.01223f
C578 two_stage_opamp_dummy_magic_14_0.Vb1.t24 GNDA 0.01223f
C579 two_stage_opamp_dummy_magic_14_0.Vb1.t14 GNDA 0.015863f
C580 two_stage_opamp_dummy_magic_14_0.Vb1.n4 GNDA 0.017248f
C581 two_stage_opamp_dummy_magic_14_0.Vb1.n5 GNDA 0.011634f
C582 two_stage_opamp_dummy_magic_14_0.Vb1.n6 GNDA 0.011634f
C583 two_stage_opamp_dummy_magic_14_0.Vb1.n7 GNDA 0.010085f
C584 two_stage_opamp_dummy_magic_14_0.Vb1.t13 GNDA 0.01223f
C585 two_stage_opamp_dummy_magic_14_0.Vb1.t17 GNDA 0.01223f
C586 two_stage_opamp_dummy_magic_14_0.Vb1.t8 GNDA 0.01223f
C587 two_stage_opamp_dummy_magic_14_0.Vb1.t19 GNDA 0.01223f
C588 two_stage_opamp_dummy_magic_14_0.Vb1.t10 GNDA 0.015863f
C589 two_stage_opamp_dummy_magic_14_0.Vb1.n8 GNDA 0.017248f
C590 two_stage_opamp_dummy_magic_14_0.Vb1.n9 GNDA 0.011634f
C591 two_stage_opamp_dummy_magic_14_0.Vb1.n10 GNDA 0.011634f
C592 two_stage_opamp_dummy_magic_14_0.Vb1.n11 GNDA 0.010085f
C593 two_stage_opamp_dummy_magic_14_0.Vb1.n12 GNDA 0.016518f
C594 two_stage_opamp_dummy_magic_14_0.Vb1.t23 GNDA 0.01223f
C595 two_stage_opamp_dummy_magic_14_0.Vb1.t7 GNDA 0.01223f
C596 two_stage_opamp_dummy_magic_14_0.Vb1.t16 GNDA 0.01223f
C597 two_stage_opamp_dummy_magic_14_0.Vb1.t25 GNDA 0.01223f
C598 two_stage_opamp_dummy_magic_14_0.Vb1.t15 GNDA 0.015863f
C599 two_stage_opamp_dummy_magic_14_0.Vb1.n13 GNDA 0.017248f
C600 two_stage_opamp_dummy_magic_14_0.Vb1.n14 GNDA 0.011634f
C601 two_stage_opamp_dummy_magic_14_0.Vb1.n15 GNDA 0.011634f
C602 two_stage_opamp_dummy_magic_14_0.Vb1.n16 GNDA 0.010085f
C603 two_stage_opamp_dummy_magic_14_0.Vb1.t6 GNDA 0.01223f
C604 two_stage_opamp_dummy_magic_14_0.Vb1.t18 GNDA 0.01223f
C605 two_stage_opamp_dummy_magic_14_0.Vb1.t9 GNDA 0.01223f
C606 two_stage_opamp_dummy_magic_14_0.Vb1.t20 GNDA 0.01223f
C607 two_stage_opamp_dummy_magic_14_0.Vb1.t11 GNDA 0.015863f
C608 two_stage_opamp_dummy_magic_14_0.Vb1.n17 GNDA 0.017248f
C609 two_stage_opamp_dummy_magic_14_0.Vb1.n18 GNDA 0.011634f
C610 two_stage_opamp_dummy_magic_14_0.Vb1.n19 GNDA 0.011634f
C611 two_stage_opamp_dummy_magic_14_0.Vb1.n20 GNDA 0.010085f
C612 two_stage_opamp_dummy_magic_14_0.Vb1.n21 GNDA 0.012503f
C613 two_stage_opamp_dummy_magic_14_0.Vb1.n22 GNDA 0.268752f
C614 two_stage_opamp_dummy_magic_14_0.Vb1.n23 GNDA 0.707133f
C615 bgr_0.VB1_CUR_BIAS GNDA 0.456038f
C616 two_stage_opamp_dummy_magic_14_0.V_err_gate.t1 GNDA 0.019171f
C617 two_stage_opamp_dummy_magic_14_0.V_err_gate.t2 GNDA 0.019171f
C618 two_stage_opamp_dummy_magic_14_0.V_err_gate.n0 GNDA 0.291518f
C619 two_stage_opamp_dummy_magic_14_0.V_err_gate.t0 GNDA 0.047929f
C620 two_stage_opamp_dummy_magic_14_0.V_err_gate.t4 GNDA 0.047929f
C621 two_stage_opamp_dummy_magic_14_0.V_err_gate.n1 GNDA 0.14684f
C622 two_stage_opamp_dummy_magic_14_0.V_err_gate.t8 GNDA 0.05352f
C623 two_stage_opamp_dummy_magic_14_0.V_err_gate.t6 GNDA 0.05352f
C624 two_stage_opamp_dummy_magic_14_0.V_err_gate.n2 GNDA 0.080392f
C625 two_stage_opamp_dummy_magic_14_0.V_err_gate.n3 GNDA 0.296704f
C626 two_stage_opamp_dummy_magic_14_0.V_err_gate.t3 GNDA 0.047929f
C627 two_stage_opamp_dummy_magic_14_0.V_err_gate.t5 GNDA 0.047929f
C628 two_stage_opamp_dummy_magic_14_0.V_err_gate.n4 GNDA 0.146204f
C629 two_stage_opamp_dummy_magic_14_0.V_err_gate.n5 GNDA 0.22702f
C630 two_stage_opamp_dummy_magic_14_0.V_err_gate.t7 GNDA 0.05352f
C631 two_stage_opamp_dummy_magic_14_0.V_err_gate.t9 GNDA 0.05352f
C632 two_stage_opamp_dummy_magic_14_0.V_err_gate.n6 GNDA 0.080392f
C633 two_stage_opamp_dummy_magic_14_0.Vb2.t32 GNDA 0.043632f
C634 two_stage_opamp_dummy_magic_14_0.Vb2.t14 GNDA 0.043632f
C635 two_stage_opamp_dummy_magic_14_0.Vb2.t19 GNDA 0.043632f
C636 two_stage_opamp_dummy_magic_14_0.Vb2.t26 GNDA 0.043632f
C637 two_stage_opamp_dummy_magic_14_0.Vb2.t22 GNDA 0.050351f
C638 two_stage_opamp_dummy_magic_14_0.Vb2.n0 GNDA 0.04088f
C639 two_stage_opamp_dummy_magic_14_0.Vb2.n1 GNDA 0.025122f
C640 two_stage_opamp_dummy_magic_14_0.Vb2.n2 GNDA 0.025122f
C641 two_stage_opamp_dummy_magic_14_0.Vb2.n3 GNDA 0.023309f
C642 two_stage_opamp_dummy_magic_14_0.Vb2.t29 GNDA 0.043632f
C643 two_stage_opamp_dummy_magic_14_0.Vb2.t28 GNDA 0.043632f
C644 two_stage_opamp_dummy_magic_14_0.Vb2.t24 GNDA 0.043632f
C645 two_stage_opamp_dummy_magic_14_0.Vb2.t17 GNDA 0.043632f
C646 two_stage_opamp_dummy_magic_14_0.Vb2.t12 GNDA 0.050351f
C647 two_stage_opamp_dummy_magic_14_0.Vb2.n4 GNDA 0.04088f
C648 two_stage_opamp_dummy_magic_14_0.Vb2.n5 GNDA 0.025122f
C649 two_stage_opamp_dummy_magic_14_0.Vb2.n6 GNDA 0.025122f
C650 two_stage_opamp_dummy_magic_14_0.Vb2.n7 GNDA 0.023309f
C651 two_stage_opamp_dummy_magic_14_0.Vb2.n8 GNDA 0.013512f
C652 two_stage_opamp_dummy_magic_14_0.Vb2.t11 GNDA 0.043632f
C653 two_stage_opamp_dummy_magic_14_0.Vb2.t15 GNDA 0.043632f
C654 two_stage_opamp_dummy_magic_14_0.Vb2.t20 GNDA 0.043632f
C655 two_stage_opamp_dummy_magic_14_0.Vb2.t16 GNDA 0.043632f
C656 two_stage_opamp_dummy_magic_14_0.Vb2.t23 GNDA 0.050351f
C657 two_stage_opamp_dummy_magic_14_0.Vb2.n9 GNDA 0.04088f
C658 two_stage_opamp_dummy_magic_14_0.Vb2.n10 GNDA 0.025122f
C659 two_stage_opamp_dummy_magic_14_0.Vb2.n11 GNDA 0.025122f
C660 two_stage_opamp_dummy_magic_14_0.Vb2.n12 GNDA 0.023309f
C661 two_stage_opamp_dummy_magic_14_0.Vb2.t30 GNDA 0.043632f
C662 two_stage_opamp_dummy_magic_14_0.Vb2.t21 GNDA 0.043632f
C663 two_stage_opamp_dummy_magic_14_0.Vb2.t25 GNDA 0.043632f
C664 two_stage_opamp_dummy_magic_14_0.Vb2.t18 GNDA 0.043632f
C665 two_stage_opamp_dummy_magic_14_0.Vb2.t13 GNDA 0.050351f
C666 two_stage_opamp_dummy_magic_14_0.Vb2.n13 GNDA 0.04088f
C667 two_stage_opamp_dummy_magic_14_0.Vb2.n14 GNDA 0.025122f
C668 two_stage_opamp_dummy_magic_14_0.Vb2.n15 GNDA 0.025122f
C669 two_stage_opamp_dummy_magic_14_0.Vb2.n16 GNDA 0.023309f
C670 two_stage_opamp_dummy_magic_14_0.Vb2.n17 GNDA 0.016397f
C671 two_stage_opamp_dummy_magic_14_0.Vb2.n18 GNDA 0.03003f
C672 two_stage_opamp_dummy_magic_14_0.Vb2.n19 GNDA 0.029147f
C673 two_stage_opamp_dummy_magic_14_0.Vb2.n20 GNDA 0.303104f
C674 two_stage_opamp_dummy_magic_14_0.Vb2.n21 GNDA 0.029147f
C675 two_stage_opamp_dummy_magic_14_0.Vb2.n22 GNDA 0.204441f
C676 two_stage_opamp_dummy_magic_14_0.Vb2.n23 GNDA 0.029147f
C677 two_stage_opamp_dummy_magic_14_0.Vb2.n24 GNDA 0.808923f
C678 two_stage_opamp_dummy_magic_14_0.Vb2.t31 GNDA 0.053353f
C679 two_stage_opamp_dummy_magic_14_0.Vb2.n25 GNDA 0.723168f
C680 two_stage_opamp_dummy_magic_14_0.Vb2.t1 GNDA 0.030851f
C681 two_stage_opamp_dummy_magic_14_0.Vb2.t2 GNDA 0.030851f
C682 two_stage_opamp_dummy_magic_14_0.Vb2.n26 GNDA 0.107063f
C683 two_stage_opamp_dummy_magic_14_0.Vb2.t0 GNDA 0.053353f
C684 two_stage_opamp_dummy_magic_14_0.Vb2.n27 GNDA 0.18525f
C685 two_stage_opamp_dummy_magic_14_0.Vb2.t27 GNDA 0.031502f
C686 two_stage_opamp_dummy_magic_14_0.Vb2.n28 GNDA 0.094361f
C687 two_stage_opamp_dummy_magic_14_0.Vb2.n29 GNDA 0.154162f
C688 two_stage_opamp_dummy_magic_14_0.Vb2.n30 GNDA 0.287807f
C689 bgr_0.cap_res2.t6 GNDA 0.358376f
C690 bgr_0.cap_res2.t12 GNDA 0.359675f
C691 bgr_0.cap_res2.t14 GNDA 0.340442f
C692 bgr_0.cap_res2.t0 GNDA 0.358376f
C693 bgr_0.cap_res2.t5 GNDA 0.359675f
C694 bgr_0.cap_res2.t8 GNDA 0.340442f
C695 bgr_0.cap_res2.t4 GNDA 0.358376f
C696 bgr_0.cap_res2.t10 GNDA 0.359675f
C697 bgr_0.cap_res2.t13 GNDA 0.340442f
C698 bgr_0.cap_res2.t19 GNDA 0.358376f
C699 bgr_0.cap_res2.t3 GNDA 0.359675f
C700 bgr_0.cap_res2.t7 GNDA 0.340442f
C701 bgr_0.cap_res2.t15 GNDA 0.358376f
C702 bgr_0.cap_res2.t18 GNDA 0.359675f
C703 bgr_0.cap_res2.t1 GNDA 0.340442f
C704 bgr_0.cap_res2.n0 GNDA 0.24022f
C705 bgr_0.cap_res2.t2 GNDA 0.1913f
C706 bgr_0.cap_res2.n1 GNDA 0.260644f
C707 bgr_0.cap_res2.t9 GNDA 0.1913f
C708 bgr_0.cap_res2.n2 GNDA 0.260644f
C709 bgr_0.cap_res2.t16 GNDA 0.1913f
C710 bgr_0.cap_res2.n3 GNDA 0.260644f
C711 bgr_0.cap_res2.t11 GNDA 0.1913f
C712 bgr_0.cap_res2.n4 GNDA 0.260644f
C713 bgr_0.cap_res2.t17 GNDA 0.373116f
C714 bgr_0.cap_res2.t20 GNDA 0.086426f
C715 bgr_0.1st_Vout_2.n0 GNDA 0.723004f
C716 bgr_0.1st_Vout_2.n1 GNDA 0.237573f
C717 bgr_0.1st_Vout_2.n2 GNDA 1.43086f
C718 bgr_0.1st_Vout_2.n3 GNDA 0.104399f
C719 bgr_0.1st_Vout_2.n4 GNDA 1.45767f
C720 bgr_0.1st_Vout_2.n5 GNDA 0.010417f
C721 bgr_0.1st_Vout_2.t10 GNDA 0.015189f
C722 bgr_0.1st_Vout_2.n6 GNDA 0.157567f
C723 bgr_0.1st_Vout_2.t33 GNDA 0.017308f
C724 bgr_0.1st_Vout_2.n8 GNDA 0.018179f
C725 bgr_0.1st_Vout_2.t24 GNDA 0.010986f
C726 bgr_0.1st_Vout_2.t13 GNDA 0.010986f
C727 bgr_0.1st_Vout_2.n9 GNDA 0.024439f
C728 bgr_0.1st_Vout_2.t28 GNDA 0.288462f
C729 bgr_0.1st_Vout_2.t17 GNDA 0.293375f
C730 bgr_0.1st_Vout_2.t12 GNDA 0.288462f
C731 bgr_0.1st_Vout_2.t32 GNDA 0.288462f
C732 bgr_0.1st_Vout_2.t35 GNDA 0.293375f
C733 bgr_0.1st_Vout_2.t11 GNDA 0.293375f
C734 bgr_0.1st_Vout_2.t31 GNDA 0.288462f
C735 bgr_0.1st_Vout_2.t23 GNDA 0.288462f
C736 bgr_0.1st_Vout_2.t26 GNDA 0.293375f
C737 bgr_0.1st_Vout_2.t30 GNDA 0.293375f
C738 bgr_0.1st_Vout_2.t22 GNDA 0.288462f
C739 bgr_0.1st_Vout_2.t15 GNDA 0.288462f
C740 bgr_0.1st_Vout_2.t19 GNDA 0.293375f
C741 bgr_0.1st_Vout_2.t36 GNDA 0.293375f
C742 bgr_0.1st_Vout_2.t29 GNDA 0.288462f
C743 bgr_0.1st_Vout_2.t21 GNDA 0.288462f
C744 bgr_0.1st_Vout_2.t25 GNDA 0.293375f
C745 bgr_0.1st_Vout_2.t18 GNDA 0.293375f
C746 bgr_0.1st_Vout_2.t14 GNDA 0.288462f
C747 bgr_0.1st_Vout_2.t20 GNDA 0.288462f
C748 bgr_0.1st_Vout_2.t34 GNDA 0.018845f
C749 bgr_0.1st_Vout_2.n10 GNDA 0.018179f
C750 bgr_0.1st_Vout_2.t27 GNDA 0.010986f
C751 bgr_0.1st_Vout_2.t16 GNDA 0.010986f
C752 bgr_0.1st_Vout_2.n11 GNDA 0.024439f
C753 bgr_0.1st_Vout_2.n12 GNDA 0.017425f
C754 bgr_0.1st_Vout_1.n0 GNDA 0.538712f
C755 bgr_0.1st_Vout_1.n1 GNDA 0.236313f
C756 bgr_0.1st_Vout_1.n2 GNDA 0.973284f
C757 bgr_0.1st_Vout_1.n3 GNDA 0.907198f
C758 bgr_0.1st_Vout_1.n4 GNDA 0.891647f
C759 bgr_0.1st_Vout_1.t11 GNDA 0.358463f
C760 bgr_0.1st_Vout_1.t15 GNDA 0.35246f
C761 bgr_0.1st_Vout_1.t29 GNDA 0.358463f
C762 bgr_0.1st_Vout_1.t35 GNDA 0.35246f
C763 bgr_0.1st_Vout_1.t31 GNDA 0.358463f
C764 bgr_0.1st_Vout_1.t34 GNDA 0.35246f
C765 bgr_0.1st_Vout_1.t20 GNDA 0.358463f
C766 bgr_0.1st_Vout_1.t28 GNDA 0.35246f
C767 bgr_0.1st_Vout_1.t24 GNDA 0.358463f
C768 bgr_0.1st_Vout_1.t27 GNDA 0.35246f
C769 bgr_0.1st_Vout_1.t14 GNDA 0.358463f
C770 bgr_0.1st_Vout_1.t19 GNDA 0.35246f
C771 bgr_0.1st_Vout_1.t30 GNDA 0.358463f
C772 bgr_0.1st_Vout_1.t33 GNDA 0.35246f
C773 bgr_0.1st_Vout_1.t18 GNDA 0.358463f
C774 bgr_0.1st_Vout_1.t26 GNDA 0.35246f
C775 bgr_0.1st_Vout_1.t23 GNDA 0.358463f
C776 bgr_0.1st_Vout_1.t25 GNDA 0.35246f
C777 bgr_0.1st_Vout_1.t17 GNDA 0.35246f
C778 bgr_0.1st_Vout_1.t12 GNDA 0.35246f
C779 bgr_0.1st_Vout_1.t21 GNDA 0.023025f
C780 bgr_0.1st_Vout_1.n5 GNDA 0.715456f
C781 bgr_0.1st_Vout_1.n6 GNDA 0.022212f
C782 bgr_0.1st_Vout_1.n7 GNDA 0.104674f
C783 bgr_0.1st_Vout_1.t36 GNDA 0.013423f
C784 bgr_0.1st_Vout_1.t16 GNDA 0.013423f
C785 bgr_0.1st_Vout_1.n8 GNDA 0.029862f
C786 bgr_0.1st_Vout_1.n9 GNDA 0.082514f
C787 bgr_0.1st_Vout_1.t9 GNDA 0.018559f
C788 bgr_0.1st_Vout_1.n10 GNDA 0.012728f
C789 bgr_0.1st_Vout_1.n11 GNDA 0.192525f
C790 bgr_0.1st_Vout_1.n12 GNDA 0.011517f
C791 bgr_0.1st_Vout_1.n13 GNDA 0.048842f
C792 bgr_0.1st_Vout_1.n14 GNDA 0.021291f
C793 bgr_0.1st_Vout_1.n15 GNDA 0.078719f
C794 bgr_0.1st_Vout_1.n16 GNDA 0.038771f
C795 bgr_0.1st_Vout_1.t32 GNDA 0.013423f
C796 bgr_0.1st_Vout_1.t22 GNDA 0.013423f
C797 bgr_0.1st_Vout_1.n17 GNDA 0.029862f
C798 bgr_0.1st_Vout_1.n18 GNDA 0.082514f
C799 bgr_0.1st_Vout_1.n19 GNDA 0.022212f
C800 bgr_0.1st_Vout_1.n20 GNDA 0.104674f
C801 bgr_0.1st_Vout_1.t13 GNDA 0.021069f
C802 bgr_0.V_mir1.t10 GNDA 0.019293f
C803 bgr_0.V_mir1.t3 GNDA 0.02939f
C804 bgr_0.V_mir1.t7 GNDA 0.023151f
C805 bgr_0.V_mir1.t18 GNDA 0.023151f
C806 bgr_0.V_mir1.t20 GNDA 0.037369f
C807 bgr_0.V_mir1.n0 GNDA 0.041731f
C808 bgr_0.V_mir1.n1 GNDA 0.028507f
C809 bgr_0.V_mir1.n2 GNDA 0.044354f
C810 bgr_0.V_mir1.t4 GNDA 0.019293f
C811 bgr_0.V_mir1.t8 GNDA 0.019293f
C812 bgr_0.V_mir1.n3 GNDA 0.044166f
C813 bgr_0.V_mir1.n4 GNDA 0.109943f
C814 bgr_0.V_mir1.n5 GNDA 0.025223f
C815 bgr_0.V_mir1.t2 GNDA 0.041163f
C816 bgr_0.V_mir1.n6 GNDA 0.027381f
C817 bgr_0.V_mir1.n7 GNDA 0.451535f
C818 bgr_0.V_mir1.n8 GNDA 0.146338f
C819 bgr_0.V_mir1.t5 GNDA 0.02939f
C820 bgr_0.V_mir1.t11 GNDA 0.023151f
C821 bgr_0.V_mir1.t17 GNDA 0.023151f
C822 bgr_0.V_mir1.t21 GNDA 0.037369f
C823 bgr_0.V_mir1.n9 GNDA 0.041731f
C824 bgr_0.V_mir1.n10 GNDA 0.028507f
C825 bgr_0.V_mir1.n11 GNDA 0.044354f
C826 bgr_0.V_mir1.t6 GNDA 0.019293f
C827 bgr_0.V_mir1.t12 GNDA 0.019293f
C828 bgr_0.V_mir1.n12 GNDA 0.044166f
C829 bgr_0.V_mir1.n13 GNDA 0.085095f
C830 bgr_0.V_mir1.n14 GNDA 0.051125f
C831 bgr_0.V_mir1.n15 GNDA 0.381359f
C832 bgr_0.V_mir1.t9 GNDA 0.02939f
C833 bgr_0.V_mir1.t13 GNDA 0.023151f
C834 bgr_0.V_mir1.t22 GNDA 0.023151f
C835 bgr_0.V_mir1.t19 GNDA 0.037369f
C836 bgr_0.V_mir1.n16 GNDA 0.041731f
C837 bgr_0.V_mir1.n17 GNDA 0.028507f
C838 bgr_0.V_mir1.n18 GNDA 0.044354f
C839 bgr_0.V_mir1.n19 GNDA 0.111042f
C840 bgr_0.V_mir1.n20 GNDA 0.044166f
C841 bgr_0.V_mir1.t14 GNDA 0.019293f
C842 two_stage_opamp_dummy_magic_14_0.VD3.t30 GNDA 0.030951f
C843 two_stage_opamp_dummy_magic_14_0.VD3.t31 GNDA 0.030951f
C844 two_stage_opamp_dummy_magic_14_0.VD3.t25 GNDA 0.030951f
C845 two_stage_opamp_dummy_magic_14_0.VD3.n0 GNDA 0.108702f
C846 two_stage_opamp_dummy_magic_14_0.VD3.t23 GNDA 0.030951f
C847 two_stage_opamp_dummy_magic_14_0.VD3.t26 GNDA 0.030951f
C848 two_stage_opamp_dummy_magic_14_0.VD3.n1 GNDA 0.108329f
C849 two_stage_opamp_dummy_magic_14_0.VD3.n2 GNDA 0.202138f
C850 two_stage_opamp_dummy_magic_14_0.VD3.t28 GNDA 0.030951f
C851 two_stage_opamp_dummy_magic_14_0.VD3.t20 GNDA 0.030951f
C852 two_stage_opamp_dummy_magic_14_0.VD3.n3 GNDA 0.108329f
C853 two_stage_opamp_dummy_magic_14_0.VD3.n4 GNDA 0.104793f
C854 two_stage_opamp_dummy_magic_14_0.VD3.t21 GNDA 0.030951f
C855 two_stage_opamp_dummy_magic_14_0.VD3.t22 GNDA 0.030951f
C856 two_stage_opamp_dummy_magic_14_0.VD3.n5 GNDA 0.108329f
C857 two_stage_opamp_dummy_magic_14_0.VD3.n6 GNDA 0.104793f
C858 two_stage_opamp_dummy_magic_14_0.VD3.t24 GNDA 0.030951f
C859 two_stage_opamp_dummy_magic_14_0.VD3.t27 GNDA 0.030951f
C860 two_stage_opamp_dummy_magic_14_0.VD3.n7 GNDA 0.108329f
C861 two_stage_opamp_dummy_magic_14_0.VD3.n8 GNDA 0.104793f
C862 two_stage_opamp_dummy_magic_14_0.VD3.t3 GNDA 0.030951f
C863 two_stage_opamp_dummy_magic_14_0.VD3.t15 GNDA 0.030951f
C864 two_stage_opamp_dummy_magic_14_0.VD3.n9 GNDA 0.10726f
C865 two_stage_opamp_dummy_magic_14_0.VD3.n10 GNDA 0.104977f
C866 two_stage_opamp_dummy_magic_14_0.VD3.t11 GNDA 0.030951f
C867 two_stage_opamp_dummy_magic_14_0.VD3.n11 GNDA 0.092854f
C868 two_stage_opamp_dummy_magic_14_0.VD3.n12 GNDA 0.030951f
C869 two_stage_opamp_dummy_magic_14_0.VD3.n13 GNDA 0.017686f
C870 two_stage_opamp_dummy_magic_14_0.VD3.n15 GNDA 0.014321f
C871 two_stage_opamp_dummy_magic_14_0.VD3.n18 GNDA 0.014321f
C872 two_stage_opamp_dummy_magic_14_0.VD3.n19 GNDA 0.017686f
C873 two_stage_opamp_dummy_magic_14_0.VD3.t6 GNDA 0.054268f
C874 two_stage_opamp_dummy_magic_14_0.VD3.t13 GNDA 0.030951f
C875 two_stage_opamp_dummy_magic_14_0.VD3.t5 GNDA 0.030951f
C876 two_stage_opamp_dummy_magic_14_0.VD3.n20 GNDA 0.10726f
C877 two_stage_opamp_dummy_magic_14_0.VD3.n21 GNDA 0.104977f
C878 two_stage_opamp_dummy_magic_14_0.VD3.t35 GNDA 0.030951f
C879 two_stage_opamp_dummy_magic_14_0.VD3.t1 GNDA 0.030951f
C880 two_stage_opamp_dummy_magic_14_0.VD3.n22 GNDA 0.10726f
C881 two_stage_opamp_dummy_magic_14_0.VD3.n23 GNDA 0.104977f
C882 two_stage_opamp_dummy_magic_14_0.VD3.t33 GNDA 0.030951f
C883 two_stage_opamp_dummy_magic_14_0.VD3.t19 GNDA 0.030951f
C884 two_stage_opamp_dummy_magic_14_0.VD3.n24 GNDA 0.10726f
C885 two_stage_opamp_dummy_magic_14_0.VD3.n25 GNDA 0.104977f
C886 two_stage_opamp_dummy_magic_14_0.VD3.t37 GNDA 0.030951f
C887 two_stage_opamp_dummy_magic_14_0.VD3.t17 GNDA 0.030951f
C888 two_stage_opamp_dummy_magic_14_0.VD3.n26 GNDA 0.10726f
C889 two_stage_opamp_dummy_magic_14_0.VD3.n27 GNDA 0.134403f
C890 two_stage_opamp_dummy_magic_14_0.VD3.n28 GNDA 0.046089f
C891 two_stage_opamp_dummy_magic_14_0.VD3.t8 GNDA 0.030951f
C892 two_stage_opamp_dummy_magic_14_0.VD3.n29 GNDA 0.092854f
C893 two_stage_opamp_dummy_magic_14_0.VD3.n30 GNDA 0.031222f
C894 two_stage_opamp_dummy_magic_14_0.VD3.n31 GNDA 0.030951f
C895 two_stage_opamp_dummy_magic_14_0.VD3.n32 GNDA 0.017686f
C896 two_stage_opamp_dummy_magic_14_0.VD3.n33 GNDA 0.017686f
C897 two_stage_opamp_dummy_magic_14_0.VD3.n34 GNDA 0.030951f
C898 two_stage_opamp_dummy_magic_14_0.VD3.n36 GNDA 0.030951f
C899 two_stage_opamp_dummy_magic_14_0.VD3.n37 GNDA 0.017686f
C900 two_stage_opamp_dummy_magic_14_0.VD3.n38 GNDA 0.017686f
C901 two_stage_opamp_dummy_magic_14_0.VD3.n39 GNDA 0.030951f
C902 two_stage_opamp_dummy_magic_14_0.VD3.n41 GNDA 0.030951f
C903 two_stage_opamp_dummy_magic_14_0.VD3.n42 GNDA 0.029837f
C904 two_stage_opamp_dummy_magic_14_0.VD3.n43 GNDA 0.017686f
C905 two_stage_opamp_dummy_magic_14_0.VD3.n44 GNDA 0.258664f
C906 two_stage_opamp_dummy_magic_14_0.VD3.t7 GNDA 0.224175f
C907 two_stage_opamp_dummy_magic_14_0.VD3.t16 GNDA 0.206931f
C908 two_stage_opamp_dummy_magic_14_0.VD3.t36 GNDA 0.206931f
C909 two_stage_opamp_dummy_magic_14_0.VD3.t18 GNDA 0.206931f
C910 two_stage_opamp_dummy_magic_14_0.VD3.t32 GNDA 0.206931f
C911 two_stage_opamp_dummy_magic_14_0.VD3.t0 GNDA 0.206931f
C912 two_stage_opamp_dummy_magic_14_0.VD3.t34 GNDA 0.206931f
C913 two_stage_opamp_dummy_magic_14_0.VD3.t4 GNDA 0.206931f
C914 two_stage_opamp_dummy_magic_14_0.VD3.t12 GNDA 0.206931f
C915 two_stage_opamp_dummy_magic_14_0.VD3.t14 GNDA 0.206931f
C916 two_stage_opamp_dummy_magic_14_0.VD3.t2 GNDA 0.206931f
C917 two_stage_opamp_dummy_magic_14_0.VD3.t10 GNDA 0.224175f
C918 two_stage_opamp_dummy_magic_14_0.VD3.n45 GNDA 0.017686f
C919 two_stage_opamp_dummy_magic_14_0.VD3.n47 GNDA 0.031222f
C920 two_stage_opamp_dummy_magic_14_0.VD3.n48 GNDA 0.030951f
C921 two_stage_opamp_dummy_magic_14_0.VD3.n49 GNDA 0.017686f
C922 two_stage_opamp_dummy_magic_14_0.VD3.n50 GNDA 0.017686f
C923 two_stage_opamp_dummy_magic_14_0.VD3.n51 GNDA 0.030951f
C924 two_stage_opamp_dummy_magic_14_0.VD3.n53 GNDA 0.030951f
C925 two_stage_opamp_dummy_magic_14_0.VD3.n54 GNDA 0.030951f
C926 two_stage_opamp_dummy_magic_14_0.VD3.n55 GNDA 0.017686f
C927 two_stage_opamp_dummy_magic_14_0.VD3.n56 GNDA 0.258664f
C928 two_stage_opamp_dummy_magic_14_0.VD3.n57 GNDA 0.013727f
C929 two_stage_opamp_dummy_magic_14_0.VD3.n58 GNDA 0.033797f
C930 two_stage_opamp_dummy_magic_14_0.VD3.t9 GNDA 0.054268f
C931 two_stage_opamp_dummy_magic_14_0.VD3.n59 GNDA 0.044756f
C932 two_stage_opamp_dummy_magic_14_0.VD3.n60 GNDA 0.117031f
C933 two_stage_opamp_dummy_magic_14_0.VD3.n61 GNDA 0.19008f
C934 two_stage_opamp_dummy_magic_14_0.VD3.n62 GNDA 0.108328f
C935 two_stage_opamp_dummy_magic_14_0.VD3.t29 GNDA 0.030951f
C936 bgr_0.Vin+.t5 GNDA 0.173951f
C937 bgr_0.Vin+.t7 GNDA 0.010696f
C938 bgr_0.Vin+.t8 GNDA 0.025367f
C939 bgr_0.Vin+.t9 GNDA 0.01649f
C940 bgr_0.Vin+.n0 GNDA 0.054406f
C941 bgr_0.Vin+.t6 GNDA 0.01649f
C942 bgr_0.Vin+.n1 GNDA 0.042338f
C943 bgr_0.Vin+.t10 GNDA 0.01649f
C944 bgr_0.Vin+.n2 GNDA 0.042909f
C945 bgr_0.Vin+.n3 GNDA 0.130793f
C946 bgr_0.Vin+.t2 GNDA 0.05348f
C947 bgr_0.Vin+.t1 GNDA 0.05348f
C948 bgr_0.Vin+.n4 GNDA 0.176679f
C949 bgr_0.Vin+.n5 GNDA 1.27851f
C950 bgr_0.Vin+.t0 GNDA 0.05348f
C951 bgr_0.Vin+.t3 GNDA 0.05348f
C952 bgr_0.Vin+.n6 GNDA 0.176679f
C953 bgr_0.Vin+.n7 GNDA 1.06525f
C954 bgr_0.Vin+.n8 GNDA 1.7265f
C955 bgr_0.Vin+.t4 GNDA 0.232527f
C956 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t11 GNDA 0.010327f
C957 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t7 GNDA 0.010327f
C958 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n0 GNDA 0.02585f
C959 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t5 GNDA 0.010327f
C960 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t8 GNDA 0.010327f
C961 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n1 GNDA 0.02585f
C962 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t2 GNDA 0.010327f
C963 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t6 GNDA 0.010327f
C964 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n2 GNDA 0.025712f
C965 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n3 GNDA 0.174588f
C966 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n4 GNDA 0.146647f
C967 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t0 GNDA 0.010327f
C968 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t3 GNDA 0.010327f
C969 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n5 GNDA 0.020653f
C970 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n6 GNDA 0.036667f
C971 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t4 GNDA 0.01549f
C972 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t10 GNDA 0.01549f
C973 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n7 GNDA 0.052733f
C974 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t12 GNDA 0.027494f
C975 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t23 GNDA 0.027494f
C976 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t30 GNDA 0.027494f
C977 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t20 GNDA 0.027494f
C978 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t28 GNDA 0.027494f
C979 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t18 GNDA 0.027494f
C980 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t26 GNDA 0.027494f
C981 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t15 GNDA 0.027494f
C982 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t24 GNDA 0.027494f
C983 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t16 GNDA 0.03209f
C984 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n8 GNDA 0.030256f
C985 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n9 GNDA 0.018975f
C986 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n10 GNDA 0.018975f
C987 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n11 GNDA 0.018975f
C988 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n12 GNDA 0.018975f
C989 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n13 GNDA 0.018975f
C990 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n14 GNDA 0.018975f
C991 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n15 GNDA 0.018975f
C992 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n16 GNDA 0.016965f
C993 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t21 GNDA 0.027494f
C994 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t14 GNDA 0.027494f
C995 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t25 GNDA 0.027494f
C996 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t17 GNDA 0.027494f
C997 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t27 GNDA 0.027494f
C998 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t19 GNDA 0.027494f
C999 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t29 GNDA 0.027494f
C1000 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t22 GNDA 0.027494f
C1001 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t31 GNDA 0.027494f
C1002 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t13 GNDA 0.03209f
C1003 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n17 GNDA 0.030256f
C1004 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n18 GNDA 0.018975f
C1005 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n19 GNDA 0.018975f
C1006 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n20 GNDA 0.018975f
C1007 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n21 GNDA 0.018975f
C1008 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n22 GNDA 0.018975f
C1009 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n23 GNDA 0.018975f
C1010 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n24 GNDA 0.018975f
C1011 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n25 GNDA 0.016965f
C1012 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n26 GNDA 0.015749f
C1013 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n27 GNDA 0.237855f
C1014 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t9 GNDA 0.01549f
C1015 two_stage_opamp_dummy_magic_14_0.V_tail_gate.t1 GNDA 0.01549f
C1016 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n28 GNDA 0.030979f
C1017 two_stage_opamp_dummy_magic_14_0.V_tail_gate.n29 GNDA 0.052233f
C1018 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.t8 GNDA 0.042347f
C1019 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.t9 GNDA 0.041635f
C1020 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.n0 GNDA 0.301726f
C1021 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.t4 GNDA 0.19618f
C1022 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.t11 GNDA 0.030408f
C1023 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.t7 GNDA 0.01137f
C1024 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.n1 GNDA 0.035664f
C1025 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.t13 GNDA 0.01137f
C1026 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.n2 GNDA 0.029194f
C1027 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.t10 GNDA 0.01137f
C1028 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.n3 GNDA 0.029194f
C1029 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.t12 GNDA 0.01137f
C1030 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.n4 GNDA 0.050605f
C1031 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.n5 GNDA 1.02228f
C1032 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.t6 GNDA 0.036877f
C1033 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.t2 GNDA 0.036877f
C1034 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.n6 GNDA 0.12988f
C1035 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.t3 GNDA 0.036877f
C1036 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.t1 GNDA 0.036877f
C1037 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.n7 GNDA 0.123576f
C1038 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.n8 GNDA 0.577511f
C1039 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.t0 GNDA 0.036877f
C1040 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.t5 GNDA 0.036877f
C1041 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.n9 GNDA 0.123576f
C1042 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.n10 GNDA 0.412965f
C1043 two_stage_opamp_dummy_magic_14_0.V_err_amp_ref.n11 GNDA 0.850389f
C1044 two_stage_opamp_dummy_magic_14_0.V_b_2nd_stage.t1 GNDA 0.105964f
C1045 two_stage_opamp_dummy_magic_14_0.V_b_2nd_stage.t8 GNDA 0.265499f
C1046 two_stage_opamp_dummy_magic_14_0.V_b_2nd_stage.t5 GNDA 0.265499f
C1047 two_stage_opamp_dummy_magic_14_0.V_b_2nd_stage.t9 GNDA 0.315106f
C1048 two_stage_opamp_dummy_magic_14_0.V_b_2nd_stage.n0 GNDA 0.166436f
C1049 two_stage_opamp_dummy_magic_14_0.V_b_2nd_stage.n1 GNDA 0.105364f
C1050 two_stage_opamp_dummy_magic_14_0.V_b_2nd_stage.t2 GNDA 0.287618f
C1051 two_stage_opamp_dummy_magic_14_0.V_b_2nd_stage.n2 GNDA 0.102722f
C1052 two_stage_opamp_dummy_magic_14_0.V_b_2nd_stage.n3 GNDA 0.485792f
C1053 two_stage_opamp_dummy_magic_14_0.V_b_2nd_stage.t3 GNDA 0.287618f
C1054 two_stage_opamp_dummy_magic_14_0.V_b_2nd_stage.t6 GNDA 0.265499f
C1055 two_stage_opamp_dummy_magic_14_0.V_b_2nd_stage.t7 GNDA 0.265499f
C1056 two_stage_opamp_dummy_magic_14_0.V_b_2nd_stage.t4 GNDA 0.315106f
C1057 two_stage_opamp_dummy_magic_14_0.V_b_2nd_stage.n4 GNDA 0.166436f
C1058 two_stage_opamp_dummy_magic_14_0.V_b_2nd_stage.n5 GNDA 0.105364f
C1059 two_stage_opamp_dummy_magic_14_0.V_b_2nd_stage.n6 GNDA 0.102722f
C1060 two_stage_opamp_dummy_magic_14_0.V_b_2nd_stage.n7 GNDA 0.485792f
C1061 two_stage_opamp_dummy_magic_14_0.V_b_2nd_stage.t0 GNDA 0.105964f
C1062 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.t12 GNDA 0.019639f
C1063 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.t13 GNDA 0.019639f
C1064 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.n0 GNDA 0.071382f
C1065 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.t10 GNDA 0.019639f
C1066 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.t11 GNDA 0.019639f
C1067 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.n1 GNDA 0.059318f
C1068 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.n2 GNDA 1.15698f
C1069 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.t14 GNDA 0.241277f
C1070 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.t4 GNDA 0.058917f
C1071 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.t8 GNDA 0.058917f
C1072 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.n3 GNDA 0.245765f
C1073 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.t3 GNDA 0.058917f
C1074 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.t2 GNDA 0.058917f
C1075 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.n4 GNDA 0.244861f
C1076 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.n5 GNDA 0.336177f
C1077 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.t5 GNDA 0.058917f
C1078 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.t9 GNDA 0.058917f
C1079 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.n6 GNDA 0.244861f
C1080 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.n7 GNDA 0.175414f
C1081 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.t6 GNDA 0.058917f
C1082 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.t0 GNDA 0.058917f
C1083 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.n8 GNDA 0.244861f
C1084 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.n9 GNDA 0.175414f
C1085 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.t7 GNDA 0.058917f
C1086 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.t1 GNDA 0.058917f
C1087 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.n10 GNDA 0.244861f
C1088 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.n11 GNDA 0.243365f
C1089 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.n12 GNDA 1.30797f
C1090 two_stage_opamp_dummy_magic_14_0.V_CMFB_S2.n13 GNDA 1.92994f
C1091 two_stage_opamp_dummy_magic_14_0.X.t14 GNDA 0.030836f
C1092 two_stage_opamp_dummy_magic_14_0.X.t5 GNDA 0.030836f
C1093 two_stage_opamp_dummy_magic_14_0.X.n0 GNDA 0.108297f
C1094 two_stage_opamp_dummy_magic_14_0.X.t15 GNDA 0.030836f
C1095 two_stage_opamp_dummy_magic_14_0.X.t24 GNDA 0.030836f
C1096 two_stage_opamp_dummy_magic_14_0.X.n1 GNDA 0.107926f
C1097 two_stage_opamp_dummy_magic_14_0.X.n2 GNDA 0.201386f
C1098 two_stage_opamp_dummy_magic_14_0.X.t0 GNDA 0.030836f
C1099 two_stage_opamp_dummy_magic_14_0.X.t22 GNDA 0.030836f
C1100 two_stage_opamp_dummy_magic_14_0.X.n3 GNDA 0.107926f
C1101 two_stage_opamp_dummy_magic_14_0.X.n4 GNDA 0.104403f
C1102 two_stage_opamp_dummy_magic_14_0.X.t3 GNDA 0.030836f
C1103 two_stage_opamp_dummy_magic_14_0.X.t23 GNDA 0.030836f
C1104 two_stage_opamp_dummy_magic_14_0.X.n5 GNDA 0.107926f
C1105 two_stage_opamp_dummy_magic_14_0.X.n6 GNDA 0.104403f
C1106 two_stage_opamp_dummy_magic_14_0.X.t13 GNDA 0.030836f
C1107 two_stage_opamp_dummy_magic_14_0.X.t12 GNDA 0.030836f
C1108 two_stage_opamp_dummy_magic_14_0.X.n7 GNDA 0.107926f
C1109 two_stage_opamp_dummy_magic_14_0.X.n8 GNDA 0.122969f
C1110 two_stage_opamp_dummy_magic_14_0.X.t7 GNDA 0.030836f
C1111 two_stage_opamp_dummy_magic_14_0.X.t2 GNDA 0.030836f
C1112 two_stage_opamp_dummy_magic_14_0.X.n9 GNDA 0.105762f
C1113 two_stage_opamp_dummy_magic_14_0.X.n10 GNDA 0.180802f
C1114 two_stage_opamp_dummy_magic_14_0.X.t37 GNDA 0.018502f
C1115 two_stage_opamp_dummy_magic_14_0.X.t50 GNDA 0.018502f
C1116 two_stage_opamp_dummy_magic_14_0.X.t33 GNDA 0.018502f
C1117 two_stage_opamp_dummy_magic_14_0.X.t47 GNDA 0.018502f
C1118 two_stage_opamp_dummy_magic_14_0.X.t30 GNDA 0.018502f
C1119 two_stage_opamp_dummy_magic_14_0.X.t44 GNDA 0.022466f
C1120 two_stage_opamp_dummy_magic_14_0.X.n11 GNDA 0.022466f
C1121 two_stage_opamp_dummy_magic_14_0.X.n12 GNDA 0.014537f
C1122 two_stage_opamp_dummy_magic_14_0.X.n13 GNDA 0.014537f
C1123 two_stage_opamp_dummy_magic_14_0.X.n14 GNDA 0.014537f
C1124 two_stage_opamp_dummy_magic_14_0.X.n15 GNDA 0.012822f
C1125 two_stage_opamp_dummy_magic_14_0.X.t54 GNDA 0.018502f
C1126 two_stage_opamp_dummy_magic_14_0.X.t28 GNDA 0.018502f
C1127 two_stage_opamp_dummy_magic_14_0.X.t53 GNDA 0.018502f
C1128 two_stage_opamp_dummy_magic_14_0.X.t39 GNDA 0.022466f
C1129 two_stage_opamp_dummy_magic_14_0.X.n16 GNDA 0.022466f
C1130 two_stage_opamp_dummy_magic_14_0.X.n17 GNDA 0.014537f
C1131 two_stage_opamp_dummy_magic_14_0.X.n18 GNDA 0.012822f
C1132 two_stage_opamp_dummy_magic_14_0.X.n19 GNDA 0.013323f
C1133 two_stage_opamp_dummy_magic_14_0.X.t25 GNDA 0.028413f
C1134 two_stage_opamp_dummy_magic_14_0.X.t38 GNDA 0.028413f
C1135 two_stage_opamp_dummy_magic_14_0.X.t52 GNDA 0.028413f
C1136 two_stage_opamp_dummy_magic_14_0.X.t36 GNDA 0.028413f
C1137 two_stage_opamp_dummy_magic_14_0.X.t49 GNDA 0.028413f
C1138 two_stage_opamp_dummy_magic_14_0.X.t32 GNDA 0.032301f
C1139 two_stage_opamp_dummy_magic_14_0.X.n20 GNDA 0.029151f
C1140 two_stage_opamp_dummy_magic_14_0.X.n21 GNDA 0.017841f
C1141 two_stage_opamp_dummy_magic_14_0.X.n22 GNDA 0.017841f
C1142 two_stage_opamp_dummy_magic_14_0.X.n23 GNDA 0.017841f
C1143 two_stage_opamp_dummy_magic_14_0.X.n24 GNDA 0.016126f
C1144 two_stage_opamp_dummy_magic_14_0.X.t41 GNDA 0.028413f
C1145 two_stage_opamp_dummy_magic_14_0.X.t46 GNDA 0.028413f
C1146 two_stage_opamp_dummy_magic_14_0.X.t40 GNDA 0.028413f
C1147 two_stage_opamp_dummy_magic_14_0.X.t26 GNDA 0.032301f
C1148 two_stage_opamp_dummy_magic_14_0.X.n25 GNDA 0.029151f
C1149 two_stage_opamp_dummy_magic_14_0.X.n26 GNDA 0.017841f
C1150 two_stage_opamp_dummy_magic_14_0.X.n27 GNDA 0.016126f
C1151 two_stage_opamp_dummy_magic_14_0.X.n28 GNDA 0.013323f
C1152 two_stage_opamp_dummy_magic_14_0.X.n29 GNDA 0.108435f
C1153 two_stage_opamp_dummy_magic_14_0.X.t1 GNDA 0.013215f
C1154 two_stage_opamp_dummy_magic_14_0.X.t20 GNDA 0.013215f
C1155 two_stage_opamp_dummy_magic_14_0.X.n30 GNDA 0.048379f
C1156 two_stage_opamp_dummy_magic_14_0.X.t6 GNDA 0.013215f
C1157 two_stage_opamp_dummy_magic_14_0.X.t9 GNDA 0.013215f
C1158 two_stage_opamp_dummy_magic_14_0.X.n31 GNDA 0.047973f
C1159 two_stage_opamp_dummy_magic_14_0.X.n32 GNDA 0.175886f
C1160 two_stage_opamp_dummy_magic_14_0.X.t16 GNDA 0.013215f
C1161 two_stage_opamp_dummy_magic_14_0.X.t4 GNDA 0.013215f
C1162 two_stage_opamp_dummy_magic_14_0.X.n33 GNDA 0.047973f
C1163 two_stage_opamp_dummy_magic_14_0.X.n34 GNDA 0.091229f
C1164 two_stage_opamp_dummy_magic_14_0.X.t17 GNDA 0.013215f
C1165 two_stage_opamp_dummy_magic_14_0.X.t21 GNDA 0.013215f
C1166 two_stage_opamp_dummy_magic_14_0.X.n35 GNDA 0.047973f
C1167 two_stage_opamp_dummy_magic_14_0.X.n36 GNDA 0.091229f
C1168 two_stage_opamp_dummy_magic_14_0.X.t11 GNDA 0.013215f
C1169 two_stage_opamp_dummy_magic_14_0.X.t18 GNDA 0.013215f
C1170 two_stage_opamp_dummy_magic_14_0.X.n37 GNDA 0.047973f
C1171 two_stage_opamp_dummy_magic_14_0.X.n38 GNDA 0.091229f
C1172 two_stage_opamp_dummy_magic_14_0.X.t19 GNDA 0.013215f
C1173 two_stage_opamp_dummy_magic_14_0.X.t10 GNDA 0.013215f
C1174 two_stage_opamp_dummy_magic_14_0.X.n39 GNDA 0.047973f
C1175 two_stage_opamp_dummy_magic_14_0.X.n40 GNDA 0.137095f
C1176 two_stage_opamp_dummy_magic_14_0.X.n41 GNDA 0.114012f
C1177 two_stage_opamp_dummy_magic_14_0.X.n42 GNDA 0.217579f
C1178 two_stage_opamp_dummy_magic_14_0.X.t31 GNDA 0.058148f
C1179 two_stage_opamp_dummy_magic_14_0.X.t45 GNDA 0.058148f
C1180 two_stage_opamp_dummy_magic_14_0.X.t29 GNDA 0.058148f
C1181 two_stage_opamp_dummy_magic_14_0.X.t43 GNDA 0.058148f
C1182 two_stage_opamp_dummy_magic_14_0.X.t27 GNDA 0.061932f
C1183 two_stage_opamp_dummy_magic_14_0.X.n43 GNDA 0.049078f
C1184 two_stage_opamp_dummy_magic_14_0.X.n44 GNDA 0.027753f
C1185 two_stage_opamp_dummy_magic_14_0.X.n45 GNDA 0.027753f
C1186 two_stage_opamp_dummy_magic_14_0.X.n46 GNDA 0.026044f
C1187 two_stage_opamp_dummy_magic_14_0.X.t48 GNDA 0.058148f
C1188 two_stage_opamp_dummy_magic_14_0.X.t35 GNDA 0.058148f
C1189 two_stage_opamp_dummy_magic_14_0.X.t42 GNDA 0.058148f
C1190 two_stage_opamp_dummy_magic_14_0.X.t34 GNDA 0.058148f
C1191 two_stage_opamp_dummy_magic_14_0.X.t51 GNDA 0.061932f
C1192 two_stage_opamp_dummy_magic_14_0.X.n47 GNDA 0.049078f
C1193 two_stage_opamp_dummy_magic_14_0.X.n48 GNDA 0.027753f
C1194 two_stage_opamp_dummy_magic_14_0.X.n49 GNDA 0.027753f
C1195 two_stage_opamp_dummy_magic_14_0.X.n50 GNDA 0.026044f
C1196 two_stage_opamp_dummy_magic_14_0.X.n51 GNDA 0.015843f
C1197 two_stage_opamp_dummy_magic_14_0.X.n52 GNDA 0.500076f
C1198 two_stage_opamp_dummy_magic_14_0.X.t8 GNDA 0.428357f
C1199 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t2 GNDA 0.345142f
C1200 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t80 GNDA 0.346293f
C1201 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t38 GNDA 0.186001f
C1202 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n0 GNDA 0.198613f
C1203 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t37 GNDA 0.345142f
C1204 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t124 GNDA 0.346293f
C1205 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t79 GNDA 0.186001f
C1206 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n1 GNDA 0.217197f
C1207 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t22 GNDA 0.345142f
C1208 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t100 GNDA 0.346293f
C1209 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t60 GNDA 0.186001f
C1210 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n2 GNDA 0.217197f
C1211 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t54 GNDA 0.345142f
C1212 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t131 GNDA 0.346293f
C1213 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t96 GNDA 0.186001f
C1214 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n3 GNDA 0.217197f
C1215 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t94 GNDA 0.345142f
C1216 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t42 GNDA 0.346293f
C1217 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t136 GNDA 0.364878f
C1218 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t32 GNDA 0.364878f
C1219 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t130 GNDA 0.186001f
C1220 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n4 GNDA 0.217197f
C1221 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t74 GNDA 0.345142f
C1222 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t97 GNDA 0.346293f
C1223 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t120 GNDA 0.364878f
C1224 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t13 GNDA 0.364878f
C1225 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t116 GNDA 0.186001f
C1226 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n5 GNDA 0.217197f
C1227 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t137 GNDA 0.346293f
C1228 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t102 GNDA 0.347548f
C1229 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t101 GNDA 0.346293f
C1230 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t61 GNDA 0.349008f
C1231 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t25 GNDA 0.379597f
C1232 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t126 GNDA 0.328964f
C1233 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t36 GNDA 0.346293f
C1234 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t1 GNDA 0.347548f
C1235 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t90 GNDA 0.328964f
C1236 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t5 GNDA 0.346293f
C1237 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t110 GNDA 0.347548f
C1238 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t26 GNDA 0.346293f
C1239 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t63 GNDA 0.347548f
C1240 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t39 GNDA 0.346293f
C1241 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t11 GNDA 0.347548f
C1242 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t68 GNDA 0.346293f
C1243 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t104 GNDA 0.347548f
C1244 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t81 GNDA 0.346293f
C1245 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t45 GNDA 0.347548f
C1246 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t30 GNDA 0.346293f
C1247 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t69 GNDA 0.347548f
C1248 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t47 GNDA 0.346293f
C1249 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t17 GNDA 0.347548f
C1250 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t73 GNDA 0.346293f
C1251 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t111 GNDA 0.347548f
C1252 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t89 GNDA 0.346293f
C1253 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t53 GNDA 0.347548f
C1254 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t115 GNDA 0.346293f
C1255 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t8 GNDA 0.347548f
C1256 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t127 GNDA 0.346293f
C1257 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t92 GNDA 0.347548f
C1258 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t76 GNDA 0.346293f
C1259 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t117 GNDA 0.347548f
C1260 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t93 GNDA 0.346293f
C1261 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t59 GNDA 0.347548f
C1262 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t121 GNDA 0.346293f
C1263 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t14 GNDA 0.347548f
C1264 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t129 GNDA 0.346293f
C1265 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t99 GNDA 0.347548f
C1266 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t20 GNDA 0.346293f
C1267 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t51 GNDA 0.347548f
C1268 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t31 GNDA 0.346293f
C1269 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t135 GNDA 0.347548f
C1270 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t55 GNDA 0.346293f
C1271 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t91 GNDA 0.347548f
C1272 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t75 GNDA 0.346293f
C1273 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t34 GNDA 0.347548f
C1274 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t23 GNDA 0.346293f
C1275 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t57 GNDA 0.347548f
C1276 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t35 GNDA 0.346293f
C1277 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t4 GNDA 0.347548f
C1278 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t62 GNDA 0.346293f
C1279 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t98 GNDA 0.347548f
C1280 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t78 GNDA 0.346293f
C1281 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t40 GNDA 0.347548f
C1282 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t103 GNDA 0.346293f
C1283 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t133 GNDA 0.347548f
C1284 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t123 GNDA 0.346293f
C1285 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t83 GNDA 0.347548f
C1286 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t108 GNDA 0.345142f
C1287 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t6 GNDA 0.346293f
C1288 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t72 GNDA 0.186001f
C1289 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n6 GNDA 0.198613f
C1290 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t138 GNDA 0.345142f
C1291 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t95 GNDA 0.346293f
C1292 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t109 GNDA 0.186001f
C1293 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n7 GNDA 0.217197f
C1294 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t49 GNDA 0.345142f
C1295 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t134 GNDA 0.346293f
C1296 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t19 GNDA 0.186001f
C1297 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n8 GNDA 0.217197f
C1298 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t84 GNDA 0.345142f
C1299 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t87 GNDA 0.346293f
C1300 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t50 GNDA 0.186001f
C1301 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n9 GNDA 0.217197f
C1302 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t125 GNDA 0.345142f
C1303 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t33 GNDA 0.346293f
C1304 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t86 GNDA 0.186001f
C1305 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n10 GNDA 0.217197f
C1306 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t29 GNDA 0.345142f
C1307 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t77 GNDA 0.346293f
C1308 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t132 GNDA 0.186001f
C1309 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n11 GNDA 0.217197f
C1310 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t67 GNDA 0.345142f
C1311 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t27 GNDA 0.346293f
C1312 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t28 GNDA 0.186001f
C1313 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n12 GNDA 0.217197f
C1314 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t119 GNDA 0.346293f
C1315 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t70 GNDA 0.186001f
C1316 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n13 GNDA 0.197462f
C1317 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t66 GNDA 0.346293f
C1318 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t105 GNDA 0.186001f
C1319 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n14 GNDA 0.197462f
C1320 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t82 GNDA 0.346293f
C1321 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t46 GNDA 0.347548f
C1322 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t7 GNDA 0.346293f
C1323 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t56 GNDA 0.347548f
C1324 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t112 GNDA 0.167416f
C1325 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n15 GNDA 0.215942f
C1326 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t16 GNDA 0.18485f
C1327 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n16 GNDA 0.234527f
C1328 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t43 GNDA 0.18485f
C1329 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n17 GNDA 0.251856f
C1330 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t9 GNDA 0.18485f
C1331 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n18 GNDA 0.251856f
C1332 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t113 GNDA 0.18485f
C1333 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n19 GNDA 0.251856f
C1334 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t3 GNDA 0.18485f
C1335 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n20 GNDA 0.251856f
C1336 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t106 GNDA 0.18485f
C1337 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n21 GNDA 0.251856f
C1338 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t64 GNDA 0.18485f
C1339 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n22 GNDA 0.251856f
C1340 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t24 GNDA 0.18485f
C1341 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n23 GNDA 0.251856f
C1342 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t58 GNDA 0.18485f
C1343 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n24 GNDA 0.251856f
C1344 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t21 GNDA 0.18485f
C1345 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n25 GNDA 0.251856f
C1346 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t122 GNDA 0.18485f
C1347 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n26 GNDA 0.251856f
C1348 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t15 GNDA 0.18485f
C1349 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n27 GNDA 0.251856f
C1350 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t118 GNDA 0.18485f
C1351 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n28 GNDA 0.251856f
C1352 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t71 GNDA 0.18485f
C1353 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n29 GNDA 0.251856f
C1354 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t107 GNDA 0.18485f
C1355 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n30 GNDA 0.251856f
C1356 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t65 GNDA 0.18485f
C1357 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n31 GNDA 0.234527f
C1358 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t41 GNDA 0.345142f
C1359 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t85 GNDA 0.167416f
C1360 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n32 GNDA 0.217197f
C1361 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t10 GNDA 0.345142f
C1362 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t52 GNDA 0.346293f
C1363 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t88 GNDA 0.364878f
C1364 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t44 GNDA 0.186001f
C1365 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n33 GNDA 0.217197f
C1366 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t114 GNDA 0.345142f
C1367 two_stage_opamp_dummy_magic_14_0.cap_res_Y.n34 GNDA 0.217197f
C1368 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t12 GNDA 0.186001f
C1369 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t48 GNDA 0.364878f
C1370 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t18 GNDA 0.364878f
C1371 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t128 GNDA 0.730561f
C1372 two_stage_opamp_dummy_magic_14_0.cap_res_Y.t0 GNDA 0.29977f
C1373 VOUT+.t14 GNDA 0.048668f
C1374 VOUT+.t2 GNDA 0.048668f
C1375 VOUT+.n0 GNDA 0.225914f
C1376 VOUT+.t18 GNDA 0.048668f
C1377 VOUT+.t3 GNDA 0.048668f
C1378 VOUT+.n1 GNDA 0.225185f
C1379 VOUT+.n2 GNDA 0.138481f
C1380 VOUT+.t11 GNDA 0.048668f
C1381 VOUT+.t13 GNDA 0.048668f
C1382 VOUT+.n3 GNDA 0.225185f
C1383 VOUT+.n4 GNDA 0.077142f
C1384 VOUT+.t0 GNDA 0.081011f
C1385 VOUT+.n5 GNDA 0.091611f
C1386 VOUT+.t15 GNDA 0.041716f
C1387 VOUT+.t6 GNDA 0.041716f
C1388 VOUT+.n6 GNDA 0.168663f
C1389 VOUT+.t7 GNDA 0.041716f
C1390 VOUT+.t5 GNDA 0.041716f
C1391 VOUT+.n7 GNDA 0.168362f
C1392 VOUT+.n8 GNDA 0.164256f
C1393 VOUT+.t8 GNDA 0.041716f
C1394 VOUT+.t4 GNDA 0.041716f
C1395 VOUT+.n9 GNDA 0.168362f
C1396 VOUT+.n10 GNDA 0.084712f
C1397 VOUT+.t12 GNDA 0.041716f
C1398 VOUT+.t1 GNDA 0.041716f
C1399 VOUT+.n11 GNDA 0.168362f
C1400 VOUT+.n12 GNDA 0.084712f
C1401 VOUT+.t10 GNDA 0.041716f
C1402 VOUT+.t16 GNDA 0.041716f
C1403 VOUT+.n13 GNDA 0.168663f
C1404 VOUT+.n14 GNDA 0.100402f
C1405 VOUT+.t17 GNDA 0.041716f
C1406 VOUT+.t9 GNDA 0.041716f
C1407 VOUT+.n15 GNDA 0.166369f
C1408 VOUT+.n16 GNDA 0.14091f
C1409 VOUT+.t45 GNDA 0.278104f
C1410 VOUT+.t150 GNDA 0.282841f
C1411 VOUT+.t101 GNDA 0.278104f
C1412 VOUT+.n17 GNDA 0.186459f
C1413 VOUT+.n18 GNDA 0.12167f
C1414 VOUT+.t91 GNDA 0.282247f
C1415 VOUT+.t38 GNDA 0.282247f
C1416 VOUT+.t130 GNDA 0.282247f
C1417 VOUT+.t90 GNDA 0.282247f
C1418 VOUT+.t80 GNDA 0.282247f
C1419 VOUT+.t128 GNDA 0.282247f
C1420 VOUT+.t124 GNDA 0.282247f
C1421 VOUT+.t32 GNDA 0.282247f
C1422 VOUT+.t70 GNDA 0.282247f
C1423 VOUT+.t73 GNDA 0.282247f
C1424 VOUT+.t23 GNDA 0.282247f
C1425 VOUT+.t108 GNDA 0.282247f
C1426 VOUT+.t62 GNDA 0.282247f
C1427 VOUT+.t19 GNDA 0.282247f
C1428 VOUT+.t151 GNDA 0.282247f
C1429 VOUT+.t49 GNDA 0.282247f
C1430 VOUT+.t85 GNDA 0.278104f
C1431 VOUT+.n19 GNDA 0.304579f
C1432 VOUT+.t48 GNDA 0.278104f
C1433 VOUT+.n20 GNDA 0.356724f
C1434 VOUT+.t138 GNDA 0.278104f
C1435 VOUT+.n21 GNDA 0.356724f
C1436 VOUT+.t107 GNDA 0.278104f
C1437 VOUT+.n22 GNDA 0.356724f
C1438 VOUT+.t71 GNDA 0.278104f
C1439 VOUT+.n23 GNDA 0.356724f
C1440 VOUT+.t25 GNDA 0.278104f
C1441 VOUT+.n24 GNDA 0.356724f
C1442 VOUT+.t129 GNDA 0.278104f
C1443 VOUT+.n25 GNDA 0.356724f
C1444 VOUT+.t87 GNDA 0.278104f
C1445 VOUT+.n26 GNDA 0.239197f
C1446 VOUT+.t52 GNDA 0.278104f
C1447 VOUT+.n27 GNDA 0.239197f
C1448 VOUT+.t141 GNDA 0.278104f
C1449 VOUT+.t75 GNDA 0.282841f
C1450 VOUT+.t111 GNDA 0.278104f
C1451 VOUT+.n28 GNDA 0.186459f
C1452 VOUT+.n29 GNDA 0.225959f
C1453 VOUT+.t54 GNDA 0.282841f
C1454 VOUT+.t24 GNDA 0.278104f
C1455 VOUT+.n30 GNDA 0.186459f
C1456 VOUT+.t114 GNDA 0.278104f
C1457 VOUT+.t34 GNDA 0.282841f
C1458 VOUT+.t74 GNDA 0.278104f
C1459 VOUT+.n31 GNDA 0.186459f
C1460 VOUT+.n32 GNDA 0.225959f
C1461 VOUT+.t95 GNDA 0.282841f
C1462 VOUT+.t59 GNDA 0.278104f
C1463 VOUT+.n33 GNDA 0.186459f
C1464 VOUT+.t148 GNDA 0.278104f
C1465 VOUT+.t79 GNDA 0.282841f
C1466 VOUT+.t117 GNDA 0.278104f
C1467 VOUT+.n34 GNDA 0.186459f
C1468 VOUT+.n35 GNDA 0.225959f
C1469 VOUT+.t134 GNDA 0.282841f
C1470 VOUT+.t100 GNDA 0.278104f
C1471 VOUT+.n36 GNDA 0.186459f
C1472 VOUT+.t44 GNDA 0.278104f
C1473 VOUT+.t122 GNDA 0.282841f
C1474 VOUT+.t153 GNDA 0.278104f
C1475 VOUT+.n37 GNDA 0.186459f
C1476 VOUT+.n38 GNDA 0.225959f
C1477 VOUT+.t102 GNDA 0.282841f
C1478 VOUT+.t66 GNDA 0.278104f
C1479 VOUT+.n39 GNDA 0.186459f
C1480 VOUT+.t154 GNDA 0.278104f
C1481 VOUT+.t82 GNDA 0.282841f
C1482 VOUT+.t123 GNDA 0.278104f
C1483 VOUT+.n40 GNDA 0.186459f
C1484 VOUT+.n41 GNDA 0.225959f
C1485 VOUT+.t137 GNDA 0.282841f
C1486 VOUT+.t106 GNDA 0.278104f
C1487 VOUT+.n42 GNDA 0.186459f
C1488 VOUT+.t51 GNDA 0.278104f
C1489 VOUT+.t126 GNDA 0.282841f
C1490 VOUT+.t22 GNDA 0.278104f
C1491 VOUT+.n43 GNDA 0.186459f
C1492 VOUT+.n44 GNDA 0.225959f
C1493 VOUT+.t132 GNDA 0.278104f
C1494 VOUT+.t56 GNDA 0.282841f
C1495 VOUT+.t96 GNDA 0.278104f
C1496 VOUT+.n45 GNDA 0.186459f
C1497 VOUT+.n46 GNDA 0.12167f
C1498 VOUT+.t116 GNDA 0.282247f
C1499 VOUT+.t105 GNDA 0.282841f
C1500 VOUT+.t69 GNDA 0.278104f
C1501 VOUT+.n47 GNDA 0.182114f
C1502 VOUT+.t147 GNDA 0.282247f
C1503 VOUT+.t29 GNDA 0.282841f
C1504 VOUT+.t139 GNDA 0.278104f
C1505 VOUT+.n48 GNDA 0.186459f
C1506 VOUT+.t109 GNDA 0.278104f
C1507 VOUT+.n49 GNDA 0.117325f
C1508 VOUT+.t43 GNDA 0.282247f
C1509 VOUT+.t60 GNDA 0.282841f
C1510 VOUT+.t37 GNDA 0.278104f
C1511 VOUT+.n50 GNDA 0.186459f
C1512 VOUT+.t144 GNDA 0.278104f
C1513 VOUT+.n51 GNDA 0.117325f
C1514 VOUT+.t83 GNDA 0.282247f
C1515 VOUT+.t115 GNDA 0.282841f
C1516 VOUT+.t21 GNDA 0.278104f
C1517 VOUT+.n52 GNDA 0.186459f
C1518 VOUT+.t125 GNDA 0.278104f
C1519 VOUT+.n53 GNDA 0.117325f
C1520 VOUT+.t63 GNDA 0.282247f
C1521 VOUT+.t26 GNDA 0.282247f
C1522 VOUT+.t103 GNDA 0.282247f
C1523 VOUT+.t57 GNDA 0.28248f
C1524 VOUT+.t135 GNDA 0.282247f
C1525 VOUT+.t33 GNDA 0.28248f
C1526 VOUT+.t120 GNDA 0.282247f
C1527 VOUT+.t77 GNDA 0.28248f
C1528 VOUT+.t155 GNDA 0.282247f
C1529 VOUT+.t119 GNDA 0.278104f
C1530 VOUT+.n54 GNDA 0.307823f
C1531 VOUT+.t78 GNDA 0.278104f
C1532 VOUT+.n55 GNDA 0.359967f
C1533 VOUT+.t97 GNDA 0.278104f
C1534 VOUT+.n56 GNDA 0.359967f
C1535 VOUT+.t61 GNDA 0.278104f
C1536 VOUT+.n57 GNDA 0.356724f
C1537 VOUT+.t27 GNDA 0.278104f
C1538 VOUT+.n58 GNDA 0.295687f
C1539 VOUT+.t41 GNDA 0.278104f
C1540 VOUT+.n59 GNDA 0.295687f
C1541 VOUT+.t145 GNDA 0.278104f
C1542 VOUT+.n60 GNDA 0.295687f
C1543 VOUT+.t113 GNDA 0.278104f
C1544 VOUT+.n61 GNDA 0.295687f
C1545 VOUT+.t72 GNDA 0.278104f
C1546 VOUT+.n62 GNDA 0.239197f
C1547 VOUT+.t92 GNDA 0.278104f
C1548 VOUT+.t20 GNDA 0.282841f
C1549 VOUT+.t55 GNDA 0.278104f
C1550 VOUT+.n63 GNDA 0.186459f
C1551 VOUT+.n64 GNDA 0.225959f
C1552 VOUT+.t31 GNDA 0.282841f
C1553 VOUT+.t50 GNDA 0.278104f
C1554 VOUT+.t121 GNDA 0.282841f
C1555 VOUT+.t156 GNDA 0.278104f
C1556 VOUT+.n65 GNDA 0.186459f
C1557 VOUT+.n66 GNDA 0.290748f
C1558 VOUT+.t67 GNDA 0.282841f
C1559 VOUT+.t86 GNDA 0.278104f
C1560 VOUT+.t152 GNDA 0.282841f
C1561 VOUT+.t47 GNDA 0.278104f
C1562 VOUT+.n67 GNDA 0.186459f
C1563 VOUT+.n68 GNDA 0.290748f
C1564 VOUT+.t131 GNDA 0.282841f
C1565 VOUT+.t94 GNDA 0.278104f
C1566 VOUT+.n69 GNDA 0.186459f
C1567 VOUT+.t39 GNDA 0.278104f
C1568 VOUT+.t118 GNDA 0.282841f
C1569 VOUT+.t146 GNDA 0.278104f
C1570 VOUT+.n70 GNDA 0.186459f
C1571 VOUT+.n71 GNDA 0.225959f
C1572 VOUT+.t89 GNDA 0.282841f
C1573 VOUT+.t53 GNDA 0.278104f
C1574 VOUT+.n72 GNDA 0.186459f
C1575 VOUT+.t142 GNDA 0.278104f
C1576 VOUT+.t76 GNDA 0.282841f
C1577 VOUT+.t112 GNDA 0.278104f
C1578 VOUT+.n73 GNDA 0.186459f
C1579 VOUT+.n74 GNDA 0.225959f
C1580 VOUT+.t127 GNDA 0.282841f
C1581 VOUT+.t88 GNDA 0.278104f
C1582 VOUT+.n75 GNDA 0.186459f
C1583 VOUT+.t35 GNDA 0.278104f
C1584 VOUT+.t110 GNDA 0.282841f
C1585 VOUT+.t140 GNDA 0.278104f
C1586 VOUT+.n76 GNDA 0.186459f
C1587 VOUT+.n77 GNDA 0.225959f
C1588 VOUT+.t84 GNDA 0.282841f
C1589 VOUT+.t46 GNDA 0.278104f
C1590 VOUT+.n78 GNDA 0.186459f
C1591 VOUT+.t136 GNDA 0.278104f
C1592 VOUT+.t68 GNDA 0.282841f
C1593 VOUT+.t104 GNDA 0.278104f
C1594 VOUT+.n79 GNDA 0.186459f
C1595 VOUT+.n80 GNDA 0.225959f
C1596 VOUT+.t42 GNDA 0.282841f
C1597 VOUT+.t149 GNDA 0.278104f
C1598 VOUT+.n81 GNDA 0.186459f
C1599 VOUT+.t99 GNDA 0.278104f
C1600 VOUT+.t30 GNDA 0.282841f
C1601 VOUT+.t65 GNDA 0.278104f
C1602 VOUT+.n82 GNDA 0.186459f
C1603 VOUT+.n83 GNDA 0.225959f
C1604 VOUT+.t81 GNDA 0.282841f
C1605 VOUT+.t40 GNDA 0.278104f
C1606 VOUT+.n84 GNDA 0.186459f
C1607 VOUT+.t133 GNDA 0.278104f
C1608 VOUT+.t64 GNDA 0.282841f
C1609 VOUT+.t98 GNDA 0.278104f
C1610 VOUT+.n85 GNDA 0.186459f
C1611 VOUT+.n86 GNDA 0.225959f
C1612 VOUT+.t28 GNDA 0.282841f
C1613 VOUT+.t58 GNDA 0.278104f
C1614 VOUT+.n87 GNDA 0.186459f
C1615 VOUT+.t93 GNDA 0.278104f
C1616 VOUT+.n88 GNDA 0.225959f
C1617 VOUT+.t143 GNDA 0.278104f
C1618 VOUT+.n89 GNDA 0.12167f
C1619 VOUT+.t36 GNDA 0.278104f
C1620 VOUT+.n90 GNDA 0.177423f
C1621 VOUT+.n91 GNDA 0.210673f
C1622 two_stage_opamp_dummy_magic_14_0.cap_res_X.t128 GNDA 0.346251f
C1623 two_stage_opamp_dummy_magic_14_0.cap_res_X.t105 GNDA 0.347506f
C1624 two_stage_opamp_dummy_magic_14_0.cap_res_X.t89 GNDA 0.346251f
C1625 two_stage_opamp_dummy_magic_14_0.cap_res_X.t71 GNDA 0.348966f
C1626 two_stage_opamp_dummy_magic_14_0.cap_res_X.t103 GNDA 0.379551f
C1627 two_stage_opamp_dummy_magic_14_0.cap_res_X.t32 GNDA 0.346251f
C1628 two_stage_opamp_dummy_magic_14_0.cap_res_X.t5 GNDA 0.347506f
C1629 two_stage_opamp_dummy_magic_14_0.cap_res_X.t84 GNDA 0.328924f
C1630 two_stage_opamp_dummy_magic_14_0.cap_res_X.t134 GNDA 0.346251f
C1631 two_stage_opamp_dummy_magic_14_0.cap_res_X.t110 GNDA 0.347506f
C1632 two_stage_opamp_dummy_magic_14_0.cap_res_X.t48 GNDA 0.328924f
C1633 two_stage_opamp_dummy_magic_14_0.cap_res_X.t81 GNDA 0.346251f
C1634 two_stage_opamp_dummy_magic_14_0.cap_res_X.t130 GNDA 0.347506f
C1635 two_stage_opamp_dummy_magic_14_0.cap_res_X.t113 GNDA 0.346251f
C1636 two_stage_opamp_dummy_magic_14_0.cap_res_X.t60 GNDA 0.347506f
C1637 two_stage_opamp_dummy_magic_14_0.cap_res_X.t120 GNDA 0.346251f
C1638 two_stage_opamp_dummy_magic_14_0.cap_res_X.t34 GNDA 0.347506f
C1639 two_stage_opamp_dummy_magic_14_0.cap_res_X.t14 GNDA 0.346251f
C1640 two_stage_opamp_dummy_magic_14_0.cap_res_X.t100 GNDA 0.347506f
C1641 two_stage_opamp_dummy_magic_14_0.cap_res_X.t87 GNDA 0.346251f
C1642 two_stage_opamp_dummy_magic_14_0.cap_res_X.t137 GNDA 0.347506f
C1643 two_stage_opamp_dummy_magic_14_0.cap_res_X.t118 GNDA 0.346251f
C1644 two_stage_opamp_dummy_magic_14_0.cap_res_X.t70 GNDA 0.347506f
C1645 two_stage_opamp_dummy_magic_14_0.cap_res_X.t125 GNDA 0.346251f
C1646 two_stage_opamp_dummy_magic_14_0.cap_res_X.t39 GNDA 0.347506f
C1647 two_stage_opamp_dummy_magic_14_0.cap_res_X.t19 GNDA 0.346251f
C1648 two_stage_opamp_dummy_magic_14_0.cap_res_X.t104 GNDA 0.347506f
C1649 two_stage_opamp_dummy_magic_14_0.cap_res_X.t26 GNDA 0.346251f
C1650 two_stage_opamp_dummy_magic_14_0.cap_res_X.t78 GNDA 0.347506f
C1651 two_stage_opamp_dummy_magic_14_0.cap_res_X.t56 GNDA 0.346251f
C1652 two_stage_opamp_dummy_magic_14_0.cap_res_X.t4 GNDA 0.347506f
C1653 two_stage_opamp_dummy_magic_14_0.cap_res_X.t129 GNDA 0.346251f
C1654 two_stage_opamp_dummy_magic_14_0.cap_res_X.t40 GNDA 0.347506f
C1655 two_stage_opamp_dummy_magic_14_0.cap_res_X.t24 GNDA 0.346251f
C1656 two_stage_opamp_dummy_magic_14_0.cap_res_X.t111 GNDA 0.347506f
C1657 two_stage_opamp_dummy_magic_14_0.cap_res_X.t33 GNDA 0.346251f
C1658 two_stage_opamp_dummy_magic_14_0.cap_res_X.t82 GNDA 0.347506f
C1659 two_stage_opamp_dummy_magic_14_0.cap_res_X.t61 GNDA 0.346251f
C1660 two_stage_opamp_dummy_magic_14_0.cap_res_X.t12 GNDA 0.347506f
C1661 two_stage_opamp_dummy_magic_14_0.cap_res_X.t72 GNDA 0.346251f
C1662 two_stage_opamp_dummy_magic_14_0.cap_res_X.t123 GNDA 0.347506f
C1663 two_stage_opamp_dummy_magic_14_0.cap_res_X.t102 GNDA 0.346251f
C1664 two_stage_opamp_dummy_magic_14_0.cap_res_X.t51 GNDA 0.347506f
C1665 two_stage_opamp_dummy_magic_14_0.cap_res_X.t108 GNDA 0.346251f
C1666 two_stage_opamp_dummy_magic_14_0.cap_res_X.t22 GNDA 0.347506f
C1667 two_stage_opamp_dummy_magic_14_0.cap_res_X.t138 GNDA 0.346251f
C1668 two_stage_opamp_dummy_magic_14_0.cap_res_X.t90 GNDA 0.347506f
C1669 two_stage_opamp_dummy_magic_14_0.cap_res_X.t77 GNDA 0.346251f
C1670 two_stage_opamp_dummy_magic_14_0.cap_res_X.t127 GNDA 0.347506f
C1671 two_stage_opamp_dummy_magic_14_0.cap_res_X.t106 GNDA 0.346251f
C1672 two_stage_opamp_dummy_magic_14_0.cap_res_X.t54 GNDA 0.347506f
C1673 two_stage_opamp_dummy_magic_14_0.cap_res_X.t116 GNDA 0.346251f
C1674 two_stage_opamp_dummy_magic_14_0.cap_res_X.t28 GNDA 0.347506f
C1675 two_stage_opamp_dummy_magic_14_0.cap_res_X.t6 GNDA 0.346251f
C1676 two_stage_opamp_dummy_magic_14_0.cap_res_X.t94 GNDA 0.347506f
C1677 two_stage_opamp_dummy_magic_14_0.cap_res_X.t17 GNDA 0.346251f
C1678 two_stage_opamp_dummy_magic_14_0.cap_res_X.t68 GNDA 0.347506f
C1679 two_stage_opamp_dummy_magic_14_0.cap_res_X.t46 GNDA 0.346251f
C1680 two_stage_opamp_dummy_magic_14_0.cap_res_X.t136 GNDA 0.347506f
C1681 two_stage_opamp_dummy_magic_14_0.cap_res_X.t121 GNDA 0.346251f
C1682 two_stage_opamp_dummy_magic_14_0.cap_res_X.t35 GNDA 0.347506f
C1683 two_stage_opamp_dummy_magic_14_0.cap_res_X.t44 GNDA 0.3451f
C1684 two_stage_opamp_dummy_magic_14_0.cap_res_X.t86 GNDA 0.346251f
C1685 two_stage_opamp_dummy_magic_14_0.cap_res_X.t9 GNDA 0.185978f
C1686 two_stage_opamp_dummy_magic_14_0.cap_res_X.n0 GNDA 0.198589f
C1687 two_stage_opamp_dummy_magic_14_0.cap_res_X.t133 GNDA 0.3451f
C1688 two_stage_opamp_dummy_magic_14_0.cap_res_X.t43 GNDA 0.346251f
C1689 two_stage_opamp_dummy_magic_14_0.cap_res_X.t97 GNDA 0.185978f
C1690 two_stage_opamp_dummy_magic_14_0.cap_res_X.n1 GNDA 0.217171f
C1691 two_stage_opamp_dummy_magic_14_0.cap_res_X.t95 GNDA 0.3451f
C1692 two_stage_opamp_dummy_magic_14_0.cap_res_X.t92 GNDA 0.346251f
C1693 two_stage_opamp_dummy_magic_14_0.cap_res_X.t64 GNDA 0.185978f
C1694 two_stage_opamp_dummy_magic_14_0.cap_res_X.n2 GNDA 0.217171f
C1695 two_stage_opamp_dummy_magic_14_0.cap_res_X.t62 GNDA 0.3451f
C1696 two_stage_opamp_dummy_magic_14_0.cap_res_X.t3 GNDA 0.346251f
C1697 two_stage_opamp_dummy_magic_14_0.cap_res_X.t30 GNDA 0.185978f
C1698 two_stage_opamp_dummy_magic_14_0.cap_res_X.n3 GNDA 0.217171f
C1699 two_stage_opamp_dummy_magic_14_0.cap_res_X.t31 GNDA 0.3451f
C1700 two_stage_opamp_dummy_magic_14_0.cap_res_X.t52 GNDA 0.346251f
C1701 two_stage_opamp_dummy_magic_14_0.cap_res_X.t132 GNDA 0.185978f
C1702 two_stage_opamp_dummy_magic_14_0.cap_res_X.n4 GNDA 0.217171f
C1703 two_stage_opamp_dummy_magic_14_0.cap_res_X.t119 GNDA 0.3451f
C1704 two_stage_opamp_dummy_magic_14_0.cap_res_X.t16 GNDA 0.346251f
C1705 two_stage_opamp_dummy_magic_14_0.cap_res_X.t85 GNDA 0.185978f
C1706 two_stage_opamp_dummy_magic_14_0.cap_res_X.n5 GNDA 0.217171f
C1707 two_stage_opamp_dummy_magic_14_0.cap_res_X.t83 GNDA 0.3451f
C1708 two_stage_opamp_dummy_magic_14_0.cap_res_X.t65 GNDA 0.346251f
C1709 two_stage_opamp_dummy_magic_14_0.cap_res_X.t47 GNDA 0.185978f
C1710 two_stage_opamp_dummy_magic_14_0.cap_res_X.n6 GNDA 0.217171f
C1711 two_stage_opamp_dummy_magic_14_0.cap_res_X.t115 GNDA 0.346251f
C1712 two_stage_opamp_dummy_magic_14_0.cap_res_X.t15 GNDA 0.185978f
C1713 two_stage_opamp_dummy_magic_14_0.cap_res_X.n7 GNDA 0.197438f
C1714 two_stage_opamp_dummy_magic_14_0.cap_res_X.t75 GNDA 0.346251f
C1715 two_stage_opamp_dummy_magic_14_0.cap_res_X.t101 GNDA 0.185978f
C1716 two_stage_opamp_dummy_magic_14_0.cap_res_X.n8 GNDA 0.197438f
C1717 two_stage_opamp_dummy_magic_14_0.cap_res_X.t131 GNDA 0.346251f
C1718 two_stage_opamp_dummy_magic_14_0.cap_res_X.t38 GNDA 0.347506f
C1719 two_stage_opamp_dummy_magic_14_0.cap_res_X.t124 GNDA 0.167396f
C1720 two_stage_opamp_dummy_magic_14_0.cap_res_X.n9 GNDA 0.215916f
C1721 two_stage_opamp_dummy_magic_14_0.cap_res_X.t67 GNDA 0.184828f
C1722 two_stage_opamp_dummy_magic_14_0.cap_res_X.n10 GNDA 0.234498f
C1723 two_stage_opamp_dummy_magic_14_0.cap_res_X.t98 GNDA 0.184828f
C1724 two_stage_opamp_dummy_magic_14_0.cap_res_X.n11 GNDA 0.251826f
C1725 two_stage_opamp_dummy_magic_14_0.cap_res_X.t59 GNDA 0.184828f
C1726 two_stage_opamp_dummy_magic_14_0.cap_res_X.n12 GNDA 0.251826f
C1727 two_stage_opamp_dummy_magic_14_0.cap_res_X.t23 GNDA 0.184828f
C1728 two_stage_opamp_dummy_magic_14_0.cap_res_X.n13 GNDA 0.251826f
C1729 two_stage_opamp_dummy_magic_14_0.cap_res_X.t55 GNDA 0.184828f
C1730 two_stage_opamp_dummy_magic_14_0.cap_res_X.n14 GNDA 0.251826f
C1731 two_stage_opamp_dummy_magic_14_0.cap_res_X.t18 GNDA 0.184828f
C1732 two_stage_opamp_dummy_magic_14_0.cap_res_X.n15 GNDA 0.251826f
C1733 two_stage_opamp_dummy_magic_14_0.cap_res_X.t117 GNDA 0.184828f
C1734 two_stage_opamp_dummy_magic_14_0.cap_res_X.n16 GNDA 0.251826f
C1735 two_stage_opamp_dummy_magic_14_0.cap_res_X.t79 GNDA 0.184828f
C1736 two_stage_opamp_dummy_magic_14_0.cap_res_X.n17 GNDA 0.251826f
C1737 two_stage_opamp_dummy_magic_14_0.cap_res_X.t109 GNDA 0.184828f
C1738 two_stage_opamp_dummy_magic_14_0.cap_res_X.n18 GNDA 0.251826f
C1739 two_stage_opamp_dummy_magic_14_0.cap_res_X.t73 GNDA 0.184828f
C1740 two_stage_opamp_dummy_magic_14_0.cap_res_X.n19 GNDA 0.251826f
C1741 two_stage_opamp_dummy_magic_14_0.cap_res_X.t36 GNDA 0.184828f
C1742 two_stage_opamp_dummy_magic_14_0.cap_res_X.n20 GNDA 0.251826f
C1743 two_stage_opamp_dummy_magic_14_0.cap_res_X.t69 GNDA 0.184828f
C1744 two_stage_opamp_dummy_magic_14_0.cap_res_X.n21 GNDA 0.251826f
C1745 two_stage_opamp_dummy_magic_14_0.cap_res_X.t29 GNDA 0.184828f
C1746 two_stage_opamp_dummy_magic_14_0.cap_res_X.n22 GNDA 0.251826f
C1747 two_stage_opamp_dummy_magic_14_0.cap_res_X.t10 GNDA 0.184828f
C1748 two_stage_opamp_dummy_magic_14_0.cap_res_X.n23 GNDA 0.251826f
C1749 two_stage_opamp_dummy_magic_14_0.cap_res_X.t45 GNDA 0.184828f
C1750 two_stage_opamp_dummy_magic_14_0.cap_res_X.n24 GNDA 0.251826f
C1751 two_stage_opamp_dummy_magic_14_0.cap_res_X.t2 GNDA 0.184828f
C1752 two_stage_opamp_dummy_magic_14_0.cap_res_X.n25 GNDA 0.234498f
C1753 two_stage_opamp_dummy_magic_14_0.cap_res_X.t1 GNDA 0.3451f
C1754 two_stage_opamp_dummy_magic_14_0.cap_res_X.t41 GNDA 0.167396f
C1755 two_stage_opamp_dummy_magic_14_0.cap_res_X.n26 GNDA 0.217171f
C1756 two_stage_opamp_dummy_magic_14_0.cap_res_X.t122 GNDA 0.3451f
C1757 two_stage_opamp_dummy_magic_14_0.cap_res_X.t25 GNDA 0.346251f
C1758 two_stage_opamp_dummy_magic_14_0.cap_res_X.t58 GNDA 0.364834f
C1759 two_stage_opamp_dummy_magic_14_0.cap_res_X.t21 GNDA 0.185978f
C1760 two_stage_opamp_dummy_magic_14_0.cap_res_X.n27 GNDA 0.217171f
C1761 two_stage_opamp_dummy_magic_14_0.cap_res_X.t126 GNDA 0.3451f
C1762 two_stage_opamp_dummy_magic_14_0.cap_res_X.t66 GNDA 0.346251f
C1763 two_stage_opamp_dummy_magic_14_0.cap_res_X.t27 GNDA 0.185978f
C1764 two_stage_opamp_dummy_magic_14_0.cap_res_X.n28 GNDA 0.198589f
C1765 two_stage_opamp_dummy_magic_14_0.cap_res_X.t8 GNDA 0.3451f
C1766 two_stage_opamp_dummy_magic_14_0.cap_res_X.t88 GNDA 0.346251f
C1767 two_stage_opamp_dummy_magic_14_0.cap_res_X.t49 GNDA 0.185978f
C1768 two_stage_opamp_dummy_magic_14_0.cap_res_X.n29 GNDA 0.217171f
C1769 two_stage_opamp_dummy_magic_14_0.cap_res_X.t107 GNDA 0.3451f
C1770 two_stage_opamp_dummy_magic_14_0.cap_res_X.t50 GNDA 0.346251f
C1771 two_stage_opamp_dummy_magic_14_0.cap_res_X.t11 GNDA 0.185978f
C1772 two_stage_opamp_dummy_magic_14_0.cap_res_X.n30 GNDA 0.217171f
C1773 two_stage_opamp_dummy_magic_14_0.cap_res_X.t74 GNDA 0.3451f
C1774 two_stage_opamp_dummy_magic_14_0.cap_res_X.t13 GNDA 0.346251f
C1775 two_stage_opamp_dummy_magic_14_0.cap_res_X.t112 GNDA 0.185978f
C1776 two_stage_opamp_dummy_magic_14_0.cap_res_X.n31 GNDA 0.217171f
C1777 two_stage_opamp_dummy_magic_14_0.cap_res_X.t37 GNDA 0.3451f
C1778 two_stage_opamp_dummy_magic_14_0.cap_res_X.t91 GNDA 0.346251f
C1779 two_stage_opamp_dummy_magic_14_0.cap_res_X.t80 GNDA 0.364834f
C1780 two_stage_opamp_dummy_magic_14_0.cap_res_X.t114 GNDA 0.364834f
C1781 two_stage_opamp_dummy_magic_14_0.cap_res_X.t76 GNDA 0.185978f
C1782 two_stage_opamp_dummy_magic_14_0.cap_res_X.n32 GNDA 0.217171f
C1783 two_stage_opamp_dummy_magic_14_0.cap_res_X.t53 GNDA 0.3451f
C1784 two_stage_opamp_dummy_magic_14_0.cap_res_X.t42 GNDA 0.346251f
C1785 two_stage_opamp_dummy_magic_14_0.cap_res_X.t99 GNDA 0.364834f
C1786 two_stage_opamp_dummy_magic_14_0.cap_res_X.t135 GNDA 0.364834f
C1787 two_stage_opamp_dummy_magic_14_0.cap_res_X.t93 GNDA 0.185978f
C1788 two_stage_opamp_dummy_magic_14_0.cap_res_X.n33 GNDA 0.217171f
C1789 two_stage_opamp_dummy_magic_14_0.cap_res_X.t20 GNDA 0.3451f
C1790 two_stage_opamp_dummy_magic_14_0.cap_res_X.n34 GNDA 0.217171f
C1791 two_stage_opamp_dummy_magic_14_0.cap_res_X.t57 GNDA 0.185978f
C1792 two_stage_opamp_dummy_magic_14_0.cap_res_X.t96 GNDA 0.364834f
C1793 two_stage_opamp_dummy_magic_14_0.cap_res_X.t63 GNDA 0.364834f
C1794 two_stage_opamp_dummy_magic_14_0.cap_res_X.t7 GNDA 0.430822f
C1795 two_stage_opamp_dummy_magic_14_0.cap_res_X.t0 GNDA 0.292647f
C1796 VOUT-.t16 GNDA 0.041786f
C1797 VOUT-.t2 GNDA 0.041786f
C1798 VOUT-.n0 GNDA 0.16895f
C1799 VOUT-.t9 GNDA 0.041786f
C1800 VOUT-.t17 GNDA 0.041786f
C1801 VOUT-.n1 GNDA 0.168949f
C1802 VOUT-.t10 GNDA 0.041786f
C1803 VOUT-.t12 GNDA 0.041786f
C1804 VOUT-.n2 GNDA 0.168648f
C1805 VOUT-.n3 GNDA 0.164536f
C1806 VOUT-.t4 GNDA 0.041786f
C1807 VOUT-.t13 GNDA 0.041786f
C1808 VOUT-.n4 GNDA 0.168648f
C1809 VOUT-.n5 GNDA 0.084856f
C1810 VOUT-.t7 GNDA 0.041786f
C1811 VOUT-.t8 GNDA 0.041786f
C1812 VOUT-.n6 GNDA 0.168648f
C1813 VOUT-.n7 GNDA 0.084856f
C1814 VOUT-.n8 GNDA 0.100572f
C1815 VOUT-.t11 GNDA 0.041786f
C1816 VOUT-.t0 GNDA 0.041786f
C1817 VOUT-.n9 GNDA 0.166651f
C1818 VOUT-.n10 GNDA 0.141149f
C1819 VOUT-.t26 GNDA 0.283321f
C1820 VOUT-.t119 GNDA 0.278576f
C1821 VOUT-.n11 GNDA 0.186776f
C1822 VOUT-.t33 GNDA 0.278576f
C1823 VOUT-.n12 GNDA 0.121877f
C1824 VOUT-.t36 GNDA 0.283321f
C1825 VOUT-.t122 GNDA 0.278576f
C1826 VOUT-.n13 GNDA 0.186776f
C1827 VOUT-.t90 GNDA 0.278576f
C1828 VOUT-.t82 GNDA 0.282727f
C1829 VOUT-.t42 GNDA 0.282727f
C1830 VOUT-.t92 GNDA 0.282727f
C1831 VOUT-.t74 GNDA 0.282727f
C1832 VOUT-.t141 GNDA 0.282727f
C1833 VOUT-.t38 GNDA 0.282727f
C1834 VOUT-.t105 GNDA 0.282727f
C1835 VOUT-.t126 GNDA 0.282727f
C1836 VOUT-.t154 GNDA 0.282727f
C1837 VOUT-.t95 GNDA 0.282727f
C1838 VOUT-.t65 GNDA 0.282727f
C1839 VOUT-.t62 GNDA 0.282727f
C1840 VOUT-.t114 GNDA 0.282727f
C1841 VOUT-.t24 GNDA 0.282727f
C1842 VOUT-.t71 GNDA 0.282727f
C1843 VOUT-.t113 GNDA 0.282727f
C1844 VOUT-.t148 GNDA 0.278576f
C1845 VOUT-.n14 GNDA 0.305096f
C1846 VOUT-.t60 GNDA 0.278576f
C1847 VOUT-.n15 GNDA 0.357329f
C1848 VOUT-.t93 GNDA 0.278576f
C1849 VOUT-.n16 GNDA 0.357329f
C1850 VOUT-.t127 GNDA 0.278576f
C1851 VOUT-.n17 GNDA 0.357329f
C1852 VOUT-.t25 GNDA 0.278576f
C1853 VOUT-.n18 GNDA 0.357329f
C1854 VOUT-.t72 GNDA 0.278576f
C1855 VOUT-.n19 GNDA 0.357329f
C1856 VOUT-.t110 GNDA 0.278576f
C1857 VOUT-.n20 GNDA 0.357329f
C1858 VOUT-.t142 GNDA 0.278576f
C1859 VOUT-.n21 GNDA 0.239603f
C1860 VOUT-.t56 GNDA 0.278576f
C1861 VOUT-.n22 GNDA 0.239603f
C1862 VOUT-.n23 GNDA 0.226343f
C1863 VOUT-.t140 GNDA 0.283321f
C1864 VOUT-.t89 GNDA 0.278576f
C1865 VOUT-.n24 GNDA 0.186776f
C1866 VOUT-.t59 GNDA 0.278576f
C1867 VOUT-.t111 GNDA 0.283321f
C1868 VOUT-.t21 GNDA 0.278576f
C1869 VOUT-.n25 GNDA 0.186776f
C1870 VOUT-.n26 GNDA 0.226343f
C1871 VOUT-.t41 GNDA 0.283321f
C1872 VOUT-.t129 GNDA 0.278576f
C1873 VOUT-.n27 GNDA 0.186776f
C1874 VOUT-.t98 GNDA 0.278576f
C1875 VOUT-.t151 GNDA 0.283321f
C1876 VOUT-.t63 GNDA 0.278576f
C1877 VOUT-.n28 GNDA 0.186776f
C1878 VOUT-.n29 GNDA 0.226343f
C1879 VOUT-.t80 GNDA 0.283321f
C1880 VOUT-.t30 GNDA 0.278576f
C1881 VOUT-.n30 GNDA 0.186776f
C1882 VOUT-.t134 GNDA 0.278576f
C1883 VOUT-.t51 GNDA 0.283321f
C1884 VOUT-.t103 GNDA 0.278576f
C1885 VOUT-.n31 GNDA 0.186776f
C1886 VOUT-.n32 GNDA 0.226343f
C1887 VOUT-.t49 GNDA 0.283321f
C1888 VOUT-.t135 GNDA 0.278576f
C1889 VOUT-.n33 GNDA 0.186776f
C1890 VOUT-.t102 GNDA 0.278576f
C1891 VOUT-.t19 GNDA 0.283321f
C1892 VOUT-.t67 GNDA 0.278576f
C1893 VOUT-.n34 GNDA 0.186776f
C1894 VOUT-.n35 GNDA 0.226343f
C1895 VOUT-.t85 GNDA 0.283321f
C1896 VOUT-.t34 GNDA 0.278576f
C1897 VOUT-.n36 GNDA 0.186776f
C1898 VOUT-.t139 GNDA 0.278576f
C1899 VOUT-.t55 GNDA 0.283321f
C1900 VOUT-.t106 GNDA 0.278576f
C1901 VOUT-.n37 GNDA 0.186776f
C1902 VOUT-.n38 GNDA 0.226343f
C1903 VOUT-.t68 GNDA 0.283321f
C1904 VOUT-.t86 GNDA 0.278576f
C1905 VOUT-.n39 GNDA 0.186776f
C1906 VOUT-.t54 GNDA 0.278576f
C1907 VOUT-.n40 GNDA 0.121877f
C1908 VOUT-.t29 GNDA 0.283321f
C1909 VOUT-.t52 GNDA 0.278576f
C1910 VOUT-.n41 GNDA 0.186776f
C1911 VOUT-.t155 GNDA 0.278576f
C1912 VOUT-.t156 GNDA 0.282727f
C1913 VOUT-.t132 GNDA 0.283321f
C1914 VOUT-.t99 GNDA 0.278576f
C1915 VOUT-.n42 GNDA 0.182423f
C1916 VOUT-.t35 GNDA 0.282727f
C1917 VOUT-.t150 GNDA 0.283321f
C1918 VOUT-.t94 GNDA 0.278576f
C1919 VOUT-.n43 GNDA 0.186776f
C1920 VOUT-.t61 GNDA 0.278576f
C1921 VOUT-.n44 GNDA 0.117524f
C1922 VOUT-.t137 GNDA 0.282727f
C1923 VOUT-.t115 GNDA 0.283321f
C1924 VOUT-.t58 GNDA 0.278576f
C1925 VOUT-.n45 GNDA 0.186776f
C1926 VOUT-.t22 GNDA 0.278576f
C1927 VOUT-.n46 GNDA 0.117524f
C1928 VOUT-.t104 GNDA 0.282727f
C1929 VOUT-.t66 GNDA 0.283321f
C1930 VOUT-.t77 GNDA 0.278576f
C1931 VOUT-.n47 GNDA 0.186776f
C1932 VOUT-.t43 GNDA 0.278576f
C1933 VOUT-.n48 GNDA 0.117524f
C1934 VOUT-.t120 GNDA 0.282727f
C1935 VOUT-.t144 GNDA 0.282727f
C1936 VOUT-.t83 GNDA 0.282727f
C1937 VOUT-.t107 GNDA 0.28296f
C1938 VOUT-.t50 GNDA 0.282727f
C1939 VOUT-.t69 GNDA 0.28296f
C1940 VOUT-.t149 GNDA 0.282727f
C1941 VOUT-.t91 GNDA 0.28296f
C1942 VOUT-.t31 GNDA 0.282727f
C1943 VOUT-.t130 GNDA 0.278576f
C1944 VOUT-.n49 GNDA 0.308345f
C1945 VOUT-.t108 GNDA 0.278576f
C1946 VOUT-.n50 GNDA 0.360578f
C1947 VOUT-.t146 GNDA 0.278576f
C1948 VOUT-.n51 GNDA 0.360578f
C1949 VOUT-.t45 GNDA 0.278576f
C1950 VOUT-.n52 GNDA 0.357329f
C1951 VOUT-.t81 GNDA 0.278576f
C1952 VOUT-.n53 GNDA 0.296189f
C1953 VOUT-.t64 GNDA 0.278576f
C1954 VOUT-.n54 GNDA 0.296189f
C1955 VOUT-.t100 GNDA 0.278576f
C1956 VOUT-.n55 GNDA 0.296189f
C1957 VOUT-.t136 GNDA 0.278576f
C1958 VOUT-.n56 GNDA 0.296189f
C1959 VOUT-.t116 GNDA 0.278576f
C1960 VOUT-.n57 GNDA 0.239603f
C1961 VOUT-.n58 GNDA 0.226343f
C1962 VOUT-.t125 GNDA 0.283321f
C1963 VOUT-.t152 GNDA 0.278576f
C1964 VOUT-.n59 GNDA 0.186776f
C1965 VOUT-.t112 GNDA 0.278576f
C1966 VOUT-.t73 GNDA 0.283321f
C1967 VOUT-.n60 GNDA 0.291242f
C1968 VOUT-.t23 GNDA 0.283321f
C1969 VOUT-.t47 GNDA 0.278576f
C1970 VOUT-.n61 GNDA 0.186776f
C1971 VOUT-.t147 GNDA 0.278576f
C1972 VOUT-.t109 GNDA 0.283321f
C1973 VOUT-.n62 GNDA 0.291242f
C1974 VOUT-.t76 GNDA 0.283321f
C1975 VOUT-.t27 GNDA 0.278576f
C1976 VOUT-.n63 GNDA 0.186776f
C1977 VOUT-.t128 GNDA 0.278576f
C1978 VOUT-.t44 GNDA 0.283321f
C1979 VOUT-.t97 GNDA 0.278576f
C1980 VOUT-.n64 GNDA 0.186776f
C1981 VOUT-.n65 GNDA 0.226343f
C1982 VOUT-.t37 GNDA 0.283321f
C1983 VOUT-.t123 GNDA 0.278576f
C1984 VOUT-.n66 GNDA 0.186776f
C1985 VOUT-.t88 GNDA 0.278576f
C1986 VOUT-.t143 GNDA 0.283321f
C1987 VOUT-.t57 GNDA 0.278576f
C1988 VOUT-.n67 GNDA 0.186776f
C1989 VOUT-.n68 GNDA 0.226343f
C1990 VOUT-.t70 GNDA 0.283321f
C1991 VOUT-.t20 GNDA 0.278576f
C1992 VOUT-.n69 GNDA 0.186776f
C1993 VOUT-.t121 GNDA 0.278576f
C1994 VOUT-.t39 GNDA 0.283321f
C1995 VOUT-.t87 GNDA 0.278576f
C1996 VOUT-.n70 GNDA 0.186776f
C1997 VOUT-.n71 GNDA 0.226343f
C1998 VOUT-.t32 GNDA 0.283321f
C1999 VOUT-.t118 GNDA 0.278576f
C2000 VOUT-.n72 GNDA 0.186776f
C2001 VOUT-.t84 GNDA 0.278576f
C2002 VOUT-.t138 GNDA 0.283321f
C2003 VOUT-.t53 GNDA 0.278576f
C2004 VOUT-.n73 GNDA 0.186776f
C2005 VOUT-.n74 GNDA 0.226343f
C2006 VOUT-.t131 GNDA 0.283321f
C2007 VOUT-.t79 GNDA 0.278576f
C2008 VOUT-.n75 GNDA 0.186776f
C2009 VOUT-.t48 GNDA 0.278576f
C2010 VOUT-.t101 GNDA 0.283321f
C2011 VOUT-.t153 GNDA 0.278576f
C2012 VOUT-.n76 GNDA 0.186776f
C2013 VOUT-.n77 GNDA 0.226343f
C2014 VOUT-.t28 GNDA 0.283321f
C2015 VOUT-.t117 GNDA 0.278576f
C2016 VOUT-.n78 GNDA 0.186776f
C2017 VOUT-.t78 GNDA 0.278576f
C2018 VOUT-.t133 GNDA 0.283321f
C2019 VOUT-.t46 GNDA 0.278576f
C2020 VOUT-.n79 GNDA 0.186776f
C2021 VOUT-.n80 GNDA 0.226343f
C2022 VOUT-.t124 GNDA 0.283321f
C2023 VOUT-.t75 GNDA 0.278576f
C2024 VOUT-.n81 GNDA 0.186776f
C2025 VOUT-.t40 GNDA 0.278576f
C2026 VOUT-.n82 GNDA 0.226343f
C2027 VOUT-.t145 GNDA 0.278576f
C2028 VOUT-.n83 GNDA 0.121877f
C2029 VOUT-.t96 GNDA 0.278576f
C2030 VOUT-.n84 GNDA 0.177725f
C2031 VOUT-.n85 GNDA 0.212227f
C2032 VOUT-.t18 GNDA 0.048751f
C2033 VOUT-.t14 GNDA 0.048751f
C2034 VOUT-.n86 GNDA 0.226297f
C2035 VOUT-.t1 GNDA 0.048751f
C2036 VOUT-.t5 GNDA 0.048751f
C2037 VOUT-.n87 GNDA 0.225568f
C2038 VOUT-.n88 GNDA 0.138716f
C2039 VOUT-.t15 GNDA 0.048751f
C2040 VOUT-.t6 GNDA 0.048751f
C2041 VOUT-.n89 GNDA 0.225568f
C2042 VOUT-.n90 GNDA 0.077273f
C2043 VOUT-.t3 GNDA 0.081149f
C2044 VOUT-.n91 GNDA 0.089317f
C2045 bgr_0.V_TOP.t24 GNDA 0.095448f
C2046 bgr_0.V_TOP.t33 GNDA 0.095448f
C2047 bgr_0.V_TOP.t39 GNDA 0.095448f
C2048 bgr_0.V_TOP.t16 GNDA 0.095448f
C2049 bgr_0.V_TOP.t15 GNDA 0.095448f
C2050 bgr_0.V_TOP.t28 GNDA 0.095448f
C2051 bgr_0.V_TOP.t38 GNDA 0.095448f
C2052 bgr_0.V_TOP.t14 GNDA 0.095448f
C2053 bgr_0.V_TOP.t27 GNDA 0.095448f
C2054 bgr_0.V_TOP.t26 GNDA 0.095448f
C2055 bgr_0.V_TOP.t37 GNDA 0.095448f
C2056 bgr_0.V_TOP.t46 GNDA 0.095448f
C2057 bgr_0.V_TOP.t18 GNDA 0.095448f
C2058 bgr_0.V_TOP.t30 GNDA 0.095448f
C2059 bgr_0.V_TOP.t29 GNDA 0.124774f
C2060 bgr_0.V_TOP.n0 GNDA 0.069758f
C2061 bgr_0.V_TOP.n1 GNDA 0.050905f
C2062 bgr_0.V_TOP.n2 GNDA 0.050905f
C2063 bgr_0.V_TOP.n3 GNDA 0.050905f
C2064 bgr_0.V_TOP.n4 GNDA 0.050905f
C2065 bgr_0.V_TOP.n5 GNDA 0.04747f
C2066 bgr_0.V_TOP.t5 GNDA 0.122745f
C2067 bgr_0.V_TOP.t40 GNDA 0.36361f
C2068 bgr_0.V_TOP.t31 GNDA 0.369803f
C2069 bgr_0.V_TOP.t35 GNDA 0.36361f
C2070 bgr_0.V_TOP.n6 GNDA 0.243789f
C2071 bgr_0.V_TOP.t32 GNDA 0.36361f
C2072 bgr_0.V_TOP.t22 GNDA 0.369803f
C2073 bgr_0.V_TOP.n7 GNDA 0.311966f
C2074 bgr_0.V_TOP.t20 GNDA 0.369803f
C2075 bgr_0.V_TOP.t25 GNDA 0.36361f
C2076 bgr_0.V_TOP.n8 GNDA 0.243789f
C2077 bgr_0.V_TOP.t21 GNDA 0.36361f
C2078 bgr_0.V_TOP.t45 GNDA 0.369803f
C2079 bgr_0.V_TOP.n9 GNDA 0.380142f
C2080 bgr_0.V_TOP.t42 GNDA 0.369803f
C2081 bgr_0.V_TOP.t49 GNDA 0.36361f
C2082 bgr_0.V_TOP.n10 GNDA 0.243789f
C2083 bgr_0.V_TOP.t44 GNDA 0.36361f
C2084 bgr_0.V_TOP.t36 GNDA 0.369803f
C2085 bgr_0.V_TOP.n11 GNDA 0.380142f
C2086 bgr_0.V_TOP.t17 GNDA 0.369803f
C2087 bgr_0.V_TOP.t23 GNDA 0.36361f
C2088 bgr_0.V_TOP.n12 GNDA 0.243789f
C2089 bgr_0.V_TOP.t19 GNDA 0.36361f
C2090 bgr_0.V_TOP.t43 GNDA 0.369803f
C2091 bgr_0.V_TOP.n13 GNDA 0.380142f
C2092 bgr_0.V_TOP.t34 GNDA 0.369803f
C2093 bgr_0.V_TOP.t41 GNDA 0.36361f
C2094 bgr_0.V_TOP.n14 GNDA 0.311966f
C2095 bgr_0.V_TOP.t47 GNDA 0.36361f
C2096 bgr_0.V_TOP.n15 GNDA 0.159079f
C2097 bgr_0.V_TOP.n16 GNDA 0.544408f
C2098 bgr_0.V_TOP.t12 GNDA 0.102288f
C2099 bgr_0.V_TOP.n17 GNDA 0.724299f
C2100 bgr_0.V_TOP.n18 GNDA 0.022634f
C2101 bgr_0.V_TOP.n19 GNDA 0.414649f
C2102 bgr_0.V_TOP.n20 GNDA 0.021924f
C2103 bgr_0.V_TOP.n21 GNDA 0.022786f
C2104 bgr_0.V_TOP.n22 GNDA 0.022634f
C2105 bgr_0.V_TOP.n23 GNDA 0.209756f
C2106 bgr_0.V_TOP.n24 GNDA 0.127416f
C2107 bgr_0.V_TOP.n25 GNDA 0.072722f
C2108 bgr_0.V_TOP.n26 GNDA 0.022634f
C2109 bgr_0.V_TOP.n27 GNDA 0.125537f
C2110 bgr_0.V_TOP.n28 GNDA 0.022634f
C2111 bgr_0.V_TOP.n29 GNDA 0.124344f
C2112 bgr_0.V_TOP.n30 GNDA 0.273328f
C2113 bgr_0.V_TOP.n31 GNDA 0.019234f
C2114 bgr_0.V_TOP.n32 GNDA 0.04747f
C2115 bgr_0.V_TOP.n33 GNDA 0.050905f
C2116 bgr_0.V_TOP.n34 GNDA 0.050905f
C2117 bgr_0.V_TOP.n35 GNDA 0.050905f
C2118 bgr_0.V_TOP.n36 GNDA 0.050905f
C2119 bgr_0.V_TOP.n37 GNDA 0.050905f
C2120 bgr_0.V_TOP.n38 GNDA 0.050905f
C2121 bgr_0.V_TOP.n39 GNDA 0.04747f
C2122 bgr_0.V_TOP.t48 GNDA 0.109989f
C2123 VDDA.t253 GNDA 0.021244f
C2124 VDDA.t259 GNDA 0.021244f
C2125 VDDA.n0 GNDA 0.07362f
C2126 VDDA.n1 GNDA 0.072052f
C2127 VDDA.t274 GNDA 0.021244f
C2128 VDDA.n2 GNDA 0.063731f
C2129 VDDA.n3 GNDA 0.021244f
C2130 VDDA.n4 GNDA 0.012139f
C2131 VDDA.n8 GNDA 0.012139f
C2132 VDDA.t318 GNDA 0.037247f
C2133 VDDA.t245 GNDA 0.021244f
C2134 VDDA.t241 GNDA 0.021244f
C2135 VDDA.n9 GNDA 0.07362f
C2136 VDDA.n10 GNDA 0.092249f
C2137 VDDA.n11 GNDA 0.031634f
C2138 VDDA.n12 GNDA 0.021244f
C2139 VDDA.n14 GNDA 0.021244f
C2140 VDDA.n15 GNDA 0.012139f
C2141 VDDA.n16 GNDA 0.012139f
C2142 VDDA.n17 GNDA 0.021244f
C2143 VDDA.n19 GNDA 0.021244f
C2144 VDDA.n20 GNDA 0.012139f
C2145 VDDA.n21 GNDA 0.012139f
C2146 VDDA.n22 GNDA 0.021244f
C2147 VDDA.n23 GNDA 0.021429f
C2148 VDDA.t320 GNDA 0.021244f
C2149 VDDA.n24 GNDA 0.063731f
C2150 VDDA.n25 GNDA 0.020479f
C2151 VDDA.n26 GNDA 0.012139f
C2152 VDDA.n27 GNDA 0.177538f
C2153 VDDA.t319 GNDA 0.153866f
C2154 VDDA.t244 GNDA 0.14203f
C2155 VDDA.t240 GNDA 0.14203f
C2156 VDDA.t252 GNDA 0.14203f
C2157 VDDA.t258 GNDA 0.14203f
C2158 VDDA.t220 GNDA 0.14203f
C2159 VDDA.t222 GNDA 0.14203f
C2160 VDDA.t234 GNDA 0.14203f
C2161 VDDA.t242 GNDA 0.14203f
C2162 VDDA.t254 GNDA 0.14203f
C2163 VDDA.t260 GNDA 0.14203f
C2164 VDDA.t273 GNDA 0.153866f
C2165 VDDA.n30 GNDA 0.012139f
C2166 VDDA.n32 GNDA 0.021429f
C2167 VDDA.n33 GNDA 0.021244f
C2168 VDDA.n34 GNDA 0.012139f
C2169 VDDA.n35 GNDA 0.012139f
C2170 VDDA.n36 GNDA 0.021244f
C2171 VDDA.n38 GNDA 0.021244f
C2172 VDDA.n39 GNDA 0.021244f
C2173 VDDA.n40 GNDA 0.012139f
C2174 VDDA.n41 GNDA 0.177538f
C2175 VDDA.n43 GNDA 0.023197f
C2176 VDDA.t272 GNDA 0.037247f
C2177 VDDA.n44 GNDA 0.031634f
C2178 VDDA.t255 GNDA 0.021244f
C2179 VDDA.t261 GNDA 0.021244f
C2180 VDDA.n45 GNDA 0.07362f
C2181 VDDA.n46 GNDA 0.092249f
C2182 VDDA.t235 GNDA 0.021244f
C2183 VDDA.t243 GNDA 0.021244f
C2184 VDDA.n47 GNDA 0.07362f
C2185 VDDA.n48 GNDA 0.072052f
C2186 VDDA.n49 GNDA 0.019423f
C2187 VDDA.t221 GNDA 0.021244f
C2188 VDDA.t223 GNDA 0.021244f
C2189 VDDA.n50 GNDA 0.072095f
C2190 VDDA.n51 GNDA 0.083053f
C2191 VDDA.t264 GNDA 0.018209f
C2192 VDDA.t149 GNDA 0.018209f
C2193 VDDA.n52 GNDA 0.075302f
C2194 VDDA.t61 GNDA 0.018209f
C2195 VDDA.t79 GNDA 0.018209f
C2196 VDDA.n53 GNDA 0.075013f
C2197 VDDA.n54 GNDA 0.104005f
C2198 VDDA.t127 GNDA 0.018209f
C2199 VDDA.t147 GNDA 0.018209f
C2200 VDDA.n55 GNDA 0.075013f
C2201 VDDA.n56 GNDA 0.054271f
C2202 VDDA.t75 GNDA 0.018209f
C2203 VDDA.t140 GNDA 0.018209f
C2204 VDDA.n57 GNDA 0.075013f
C2205 VDDA.n58 GNDA 0.054271f
C2206 VDDA.t62 GNDA 0.018209f
C2207 VDDA.t139 GNDA 0.018209f
C2208 VDDA.n59 GNDA 0.075013f
C2209 VDDA.n60 GNDA 0.054271f
C2210 VDDA.t39 GNDA 0.018209f
C2211 VDDA.t265 GNDA 0.018209f
C2212 VDDA.n61 GNDA 0.075013f
C2213 VDDA.n62 GNDA 0.109478f
C2214 VDDA.t366 GNDA 0.018349f
C2215 VDDA.n64 GNDA 0.012139f
C2216 VDDA.n66 GNDA 0.012139f
C2217 VDDA.t351 GNDA 0.019177f
C2218 VDDA.n67 GNDA 0.021244f
C2219 VDDA.n68 GNDA 0.012139f
C2220 VDDA.n69 GNDA 0.021244f
C2221 VDDA.n70 GNDA 0.029557f
C2222 VDDA.t353 GNDA 0.032005f
C2223 VDDA.n72 GNDA 0.048593f
C2224 VDDA.n74 GNDA 0.107433f
C2225 VDDA.t352 GNDA 0.089224f
C2226 VDDA.t72 GNDA 0.08012f
C2227 VDDA.t76 GNDA 0.08012f
C2228 VDDA.t63 GNDA 0.08012f
C2229 VDDA.t150 GNDA 0.08012f
C2230 VDDA.t124 GNDA 0.08012f
C2231 VDDA.t80 GNDA 0.08012f
C2232 VDDA.t38 GNDA 0.08012f
C2233 VDDA.t10 GNDA 0.08012f
C2234 VDDA.t128 GNDA 0.08012f
C2235 VDDA.t148 GNDA 0.08012f
C2236 VDDA.t367 GNDA 0.089224f
C2237 VDDA.n76 GNDA 0.012139f
C2238 VDDA.n77 GNDA 0.021244f
C2239 VDDA.n78 GNDA 0.021244f
C2240 VDDA.t368 GNDA 0.032005f
C2241 VDDA.n79 GNDA 0.026759f
C2242 VDDA.n80 GNDA 0.012776f
C2243 VDDA.n81 GNDA 0.107433f
C2244 VDDA.n82 GNDA 0.012139f
C2245 VDDA.n83 GNDA 0.024075f
C2246 VDDA.n84 GNDA 0.038904f
C2247 VDDA.n85 GNDA 0.171f
C2248 VDDA.t142 GNDA 0.036418f
C2249 VDDA.t126 GNDA 0.036418f
C2250 VDDA.n86 GNDA 0.146104f
C2251 VDDA.n87 GNDA 0.074225f
C2252 VDDA.n89 GNDA 0.012139f
C2253 VDDA.n95 GNDA 0.012776f
C2254 VDDA.n96 GNDA 0.012139f
C2255 VDDA.t306 GNDA 0.044126f
C2256 VDDA.t144 GNDA 0.036418f
C2257 VDDA.t136 GNDA 0.036418f
C2258 VDDA.n97 GNDA 0.146104f
C2259 VDDA.n98 GNDA 0.074225f
C2260 VDDA.t78 GNDA 0.036418f
C2261 VDDA.t60 GNDA 0.036418f
C2262 VDDA.n99 GNDA 0.146104f
C2263 VDDA.n100 GNDA 0.074225f
C2264 VDDA.t12 GNDA 0.036418f
C2265 VDDA.t74 GNDA 0.036418f
C2266 VDDA.n101 GNDA 0.146104f
C2267 VDDA.n102 GNDA 0.074225f
C2268 VDDA.t41 GNDA 0.036418f
C2269 VDDA.t138 GNDA 0.036418f
C2270 VDDA.n103 GNDA 0.146104f
C2271 VDDA.n104 GNDA 0.093927f
C2272 VDDA.n105 GNDA 0.036327f
C2273 VDDA.n106 GNDA 0.024151f
C2274 VDDA.n107 GNDA 0.012139f
C2275 VDDA.n108 GNDA 0.012139f
C2276 VDDA.n109 GNDA 0.021244f
C2277 VDDA.n110 GNDA 0.012139f
C2278 VDDA.n111 GNDA 0.012139f
C2279 VDDA.n112 GNDA 0.012139f
C2280 VDDA.n113 GNDA 0.012139f
C2281 VDDA.n114 GNDA 0.021244f
C2282 VDDA.n115 GNDA 0.024151f
C2283 VDDA.n116 GNDA 0.012139f
C2284 VDDA.n117 GNDA 0.012139f
C2285 VDDA.n118 GNDA 0.012139f
C2286 VDDA.n119 GNDA 0.03075f
C2287 VDDA.n120 GNDA 0.021244f
C2288 VDDA.n121 GNDA 0.021244f
C2289 VDDA.n122 GNDA 0.021244f
C2290 VDDA.n123 GNDA 0.012139f
C2291 VDDA.n124 GNDA 0.012139f
C2292 VDDA.n126 GNDA 0.021244f
C2293 VDDA.n127 GNDA 0.021244f
C2294 VDDA.n129 GNDA 0.012139f
C2295 VDDA.n130 GNDA 0.012139f
C2296 VDDA.n131 GNDA 0.021244f
C2297 VDDA.n132 GNDA 0.021244f
C2298 VDDA.n133 GNDA 0.021244f
C2299 VDDA.n135 GNDA 0.024075f
C2300 VDDA.n136 GNDA 0.012139f
C2301 VDDA.n137 GNDA 0.286488f
C2302 VDDA.t307 GNDA 0.237931f
C2303 VDDA.t40 GNDA 0.213652f
C2304 VDDA.t137 GNDA 0.213652f
C2305 VDDA.t11 GNDA 0.213652f
C2306 VDDA.t73 GNDA 0.213652f
C2307 VDDA.t77 GNDA 0.213652f
C2308 VDDA.t59 GNDA 0.213652f
C2309 VDDA.t143 GNDA 0.213652f
C2310 VDDA.t135 GNDA 0.213652f
C2311 VDDA.t141 GNDA 0.213652f
C2312 VDDA.t125 GNDA 0.213652f
C2313 VDDA.t322 GNDA 0.237931f
C2314 VDDA.n142 GNDA 0.012776f
C2315 VDDA.n143 GNDA 0.012139f
C2316 VDDA.n144 GNDA 0.021244f
C2317 VDDA.n145 GNDA 0.024151f
C2318 VDDA.n146 GNDA 0.012139f
C2319 VDDA.n147 GNDA 0.012139f
C2320 VDDA.n150 GNDA 0.012139f
C2321 VDDA.n151 GNDA 0.012139f
C2322 VDDA.n152 GNDA 0.024151f
C2323 VDDA.n153 GNDA 0.03075f
C2324 VDDA.n154 GNDA 0.012139f
C2325 VDDA.n155 GNDA 0.021244f
C2326 VDDA.n156 GNDA 0.021244f
C2327 VDDA.n157 GNDA 0.012139f
C2328 VDDA.n158 GNDA 0.012139f
C2329 VDDA.n159 GNDA 0.021244f
C2330 VDDA.n160 GNDA 0.021244f
C2331 VDDA.n161 GNDA 0.012139f
C2332 VDDA.n162 GNDA 0.012139f
C2333 VDDA.n163 GNDA 0.021244f
C2334 VDDA.n164 GNDA 0.021244f
C2335 VDDA.n165 GNDA 0.012139f
C2336 VDDA.n166 GNDA 0.012139f
C2337 VDDA.n167 GNDA 0.021244f
C2338 VDDA.n168 GNDA 0.021244f
C2339 VDDA.n169 GNDA 0.021244f
C2340 VDDA.n170 GNDA 0.012139f
C2341 VDDA.n171 GNDA 0.286488f
C2342 VDDA.n173 GNDA 0.026793f
C2343 VDDA.t321 GNDA 0.044126f
C2344 VDDA.n174 GNDA 0.035525f
C2345 VDDA.n175 GNDA 0.049381f
C2346 VDDA.n176 GNDA 0.065204f
C2347 VDDA.t191 GNDA 0.015174f
C2348 VDDA.t189 GNDA 0.015174f
C2349 VDDA.n177 GNDA 0.052323f
C2350 VDDA.n178 GNDA 0.067661f
C2351 VDDA.t371 GNDA 0.015174f
C2352 VDDA.n179 GNDA 0.045522f
C2353 VDDA.n180 GNDA 0.021244f
C2354 VDDA.n181 GNDA 0.012139f
C2355 VDDA.t328 GNDA 0.107813f
C2356 VDDA.n184 GNDA 0.012139f
C2357 VDDA.n185 GNDA 0.012139f
C2358 VDDA.t284 GNDA 0.022803f
C2359 VDDA.n186 GNDA 0.031107f
C2360 VDDA.n187 GNDA 0.026369f
C2361 VDDA.t330 GNDA 0.022803f
C2362 VDDA.t332 GNDA 0.015174f
C2363 VDDA.n188 GNDA 0.045522f
C2364 VDDA.n189 GNDA 0.021244f
C2365 VDDA.n190 GNDA 0.012139f
C2366 VDDA.t375 GNDA 0.096811f
C2367 VDDA.t172 GNDA 0.096811f
C2368 VDDA.t162 GNDA 0.096811f
C2369 VDDA.t171 GNDA 0.096811f
C2370 VDDA.t331 GNDA 0.107813f
C2371 VDDA.n192 GNDA 0.012139f
C2372 VDDA.n194 GNDA 0.012139f
C2373 VDDA.n195 GNDA 0.021244f
C2374 VDDA.n196 GNDA 0.021244f
C2375 VDDA.n197 GNDA 0.021429f
C2376 VDDA.n199 GNDA 0.129815f
C2377 VDDA.n200 GNDA 0.012139f
C2378 VDDA.n201 GNDA 0.023274f
C2379 VDDA.n202 GNDA 0.033246f
C2380 VDDA.t173 GNDA 0.015174f
C2381 VDDA.t163 GNDA 0.015174f
C2382 VDDA.n203 GNDA 0.052323f
C2383 VDDA.n204 GNDA 0.090103f
C2384 VDDA.n205 GNDA 0.026369f
C2385 VDDA.t327 GNDA 0.022803f
C2386 VDDA.n206 GNDA 0.031107f
C2387 VDDA.n207 GNDA 0.016267f
C2388 VDDA.t286 GNDA 0.015174f
C2389 VDDA.n209 GNDA 0.033383f
C2390 VDDA.n211 GNDA 0.012139f
C2391 VDDA.n212 GNDA 0.033383f
C2392 VDDA.n213 GNDA 0.033383f
C2393 VDDA.t329 GNDA 0.015174f
C2394 VDDA.n215 GNDA 0.045522f
C2395 VDDA.n216 GNDA 0.032763f
C2396 VDDA.n218 GNDA 0.045522f
C2397 VDDA.n219 GNDA 0.026086f
C2398 VDDA.n221 GNDA 0.118814f
C2399 VDDA.t285 GNDA 0.107813f
C2400 VDDA.t376 GNDA 0.096811f
C2401 VDDA.t188 GNDA 0.096811f
C2402 VDDA.t190 GNDA 0.096811f
C2403 VDDA.t170 GNDA 0.096811f
C2404 VDDA.t370 GNDA 0.107813f
C2405 VDDA.n222 GNDA 0.012139f
C2406 VDDA.n224 GNDA 0.021429f
C2407 VDDA.n225 GNDA 0.021244f
C2408 VDDA.n226 GNDA 0.021244f
C2409 VDDA.n227 GNDA 0.012139f
C2410 VDDA.n228 GNDA 0.129815f
C2411 VDDA.n230 GNDA 0.025992f
C2412 VDDA.t369 GNDA 0.022803f
C2413 VDDA.n231 GNDA 0.031747f
C2414 VDDA.n232 GNDA 0.082891f
C2415 VDDA.n233 GNDA 0.093085f
C2416 VDDA.n234 GNDA 0.144098f
C2417 VDDA.t237 GNDA 0.021244f
C2418 VDDA.t247 GNDA 0.021244f
C2419 VDDA.n235 GNDA 0.07362f
C2420 VDDA.n236 GNDA 0.072052f
C2421 VDDA.t362 GNDA 0.021244f
C2422 VDDA.n237 GNDA 0.063731f
C2423 VDDA.n238 GNDA 0.021244f
C2424 VDDA.n239 GNDA 0.012139f
C2425 VDDA.n243 GNDA 0.012139f
C2426 VDDA.t287 GNDA 0.037247f
C2427 VDDA.t233 GNDA 0.021244f
C2428 VDDA.t229 GNDA 0.021244f
C2429 VDDA.n244 GNDA 0.07362f
C2430 VDDA.n245 GNDA 0.092249f
C2431 VDDA.n246 GNDA 0.031634f
C2432 VDDA.n247 GNDA 0.021244f
C2433 VDDA.n249 GNDA 0.021244f
C2434 VDDA.n250 GNDA 0.012139f
C2435 VDDA.n251 GNDA 0.012139f
C2436 VDDA.n252 GNDA 0.021244f
C2437 VDDA.n254 GNDA 0.021244f
C2438 VDDA.n255 GNDA 0.012139f
C2439 VDDA.n256 GNDA 0.012139f
C2440 VDDA.n257 GNDA 0.021244f
C2441 VDDA.n258 GNDA 0.021429f
C2442 VDDA.t289 GNDA 0.021244f
C2443 VDDA.n259 GNDA 0.063731f
C2444 VDDA.n260 GNDA 0.020479f
C2445 VDDA.n261 GNDA 0.012139f
C2446 VDDA.n262 GNDA 0.177538f
C2447 VDDA.t288 GNDA 0.153866f
C2448 VDDA.t232 GNDA 0.14203f
C2449 VDDA.t228 GNDA 0.14203f
C2450 VDDA.t236 GNDA 0.14203f
C2451 VDDA.t246 GNDA 0.14203f
C2452 VDDA.t256 GNDA 0.14203f
C2453 VDDA.t226 GNDA 0.14203f
C2454 VDDA.t224 GNDA 0.14203f
C2455 VDDA.t230 GNDA 0.14203f
C2456 VDDA.t238 GNDA 0.14203f
C2457 VDDA.t250 GNDA 0.14203f
C2458 VDDA.t361 GNDA 0.153866f
C2459 VDDA.n265 GNDA 0.012139f
C2460 VDDA.n267 GNDA 0.021429f
C2461 VDDA.n268 GNDA 0.021244f
C2462 VDDA.n269 GNDA 0.012139f
C2463 VDDA.n270 GNDA 0.012139f
C2464 VDDA.n271 GNDA 0.021244f
C2465 VDDA.n273 GNDA 0.021244f
C2466 VDDA.n274 GNDA 0.021244f
C2467 VDDA.n275 GNDA 0.012139f
C2468 VDDA.n276 GNDA 0.177538f
C2469 VDDA.n278 GNDA 0.023197f
C2470 VDDA.t360 GNDA 0.037247f
C2471 VDDA.n279 GNDA 0.031634f
C2472 VDDA.t239 GNDA 0.021244f
C2473 VDDA.t251 GNDA 0.021244f
C2474 VDDA.n280 GNDA 0.07362f
C2475 VDDA.n281 GNDA 0.092249f
C2476 VDDA.t225 GNDA 0.021244f
C2477 VDDA.t231 GNDA 0.021244f
C2478 VDDA.n282 GNDA 0.07362f
C2479 VDDA.n283 GNDA 0.072052f
C2480 VDDA.n284 GNDA 0.019423f
C2481 VDDA.t257 GNDA 0.021244f
C2482 VDDA.t227 GNDA 0.021244f
C2483 VDDA.n285 GNDA 0.072095f
C2484 VDDA.n286 GNDA 0.083053f
C2485 VDDA.t387 GNDA 0.018209f
C2486 VDDA.t263 GNDA 0.018209f
C2487 VDDA.n287 GNDA 0.075302f
C2488 VDDA.t66 GNDA 0.018209f
C2489 VDDA.t386 GNDA 0.018209f
C2490 VDDA.n288 GNDA 0.075013f
C2491 VDDA.n289 GNDA 0.104005f
C2492 VDDA.t193 GNDA 0.018209f
C2493 VDDA.t169 GNDA 0.018209f
C2494 VDDA.n290 GNDA 0.075013f
C2495 VDDA.n291 GNDA 0.054271f
C2496 VDDA.t71 GNDA 0.018209f
C2497 VDDA.t116 GNDA 0.018209f
C2498 VDDA.n292 GNDA 0.075013f
C2499 VDDA.n293 GNDA 0.054271f
C2500 VDDA.t198 GNDA 0.018209f
C2501 VDDA.t196 GNDA 0.018209f
C2502 VDDA.n294 GNDA 0.075013f
C2503 VDDA.n295 GNDA 0.054271f
C2504 VDDA.t262 GNDA 0.018209f
C2505 VDDA.t168 GNDA 0.018209f
C2506 VDDA.n296 GNDA 0.075013f
C2507 VDDA.n297 GNDA 0.109478f
C2508 VDDA.t333 GNDA 0.018349f
C2509 VDDA.n298 GNDA 0.012139f
C2510 VDDA.t335 GNDA 0.032005f
C2511 VDDA.n299 GNDA 0.012139f
C2512 VDDA.n300 GNDA 0.012139f
C2513 VDDA.n303 GNDA 0.012139f
C2514 VDDA.t345 GNDA 0.019177f
C2515 VDDA.n304 GNDA 0.021244f
C2516 VDDA.n305 GNDA 0.012139f
C2517 VDDA.n306 GNDA 0.021244f
C2518 VDDA.n307 GNDA 0.029557f
C2519 VDDA.t347 GNDA 0.032005f
C2520 VDDA.n309 GNDA 0.048593f
C2521 VDDA.n311 GNDA 0.107433f
C2522 VDDA.t346 GNDA 0.089224f
C2523 VDDA.t69 GNDA 0.08012f
C2524 VDDA.t70 GNDA 0.08012f
C2525 VDDA.t211 GNDA 0.08012f
C2526 VDDA.t35 GNDA 0.08012f
C2527 VDDA.t385 GNDA 0.08012f
C2528 VDDA.t197 GNDA 0.08012f
C2529 VDDA.t209 GNDA 0.08012f
C2530 VDDA.t113 GNDA 0.08012f
C2531 VDDA.t210 GNDA 0.08012f
C2532 VDDA.t192 GNDA 0.08012f
C2533 VDDA.t334 GNDA 0.089224f
C2534 VDDA.n312 GNDA 0.107433f
C2535 VDDA.n313 GNDA 0.012776f
C2536 VDDA.n314 GNDA 0.026759f
C2537 VDDA.n315 GNDA 0.021244f
C2538 VDDA.n316 GNDA 0.021244f
C2539 VDDA.n318 GNDA 0.024075f
C2540 VDDA.n319 GNDA 0.038904f
C2541 VDDA.n320 GNDA 0.171f
C2542 VDDA.t58 GNDA 0.036418f
C2543 VDDA.t68 GNDA 0.036418f
C2544 VDDA.n321 GNDA 0.146104f
C2545 VDDA.n322 GNDA 0.074225f
C2546 VDDA.n324 GNDA 0.012139f
C2547 VDDA.n329 GNDA 0.012776f
C2548 VDDA.n335 GNDA 0.012776f
C2549 VDDA.n336 GNDA 0.012139f
C2550 VDDA.t290 GNDA 0.044126f
C2551 VDDA.t56 GNDA 0.036418f
C2552 VDDA.t115 GNDA 0.036418f
C2553 VDDA.n337 GNDA 0.146104f
C2554 VDDA.n338 GNDA 0.074225f
C2555 VDDA.t54 GNDA 0.036418f
C2556 VDDA.t195 GNDA 0.036418f
C2557 VDDA.n339 GNDA 0.146104f
C2558 VDDA.n340 GNDA 0.074225f
C2559 VDDA.t20 GNDA 0.036418f
C2560 VDDA.t393 GNDA 0.036418f
C2561 VDDA.n341 GNDA 0.146104f
C2562 VDDA.n342 GNDA 0.074225f
C2563 VDDA.t118 GNDA 0.036418f
C2564 VDDA.t120 GNDA 0.036418f
C2565 VDDA.n343 GNDA 0.146104f
C2566 VDDA.n344 GNDA 0.093927f
C2567 VDDA.n345 GNDA 0.036327f
C2568 VDDA.n346 GNDA 0.021244f
C2569 VDDA.n347 GNDA 0.012139f
C2570 VDDA.n348 GNDA 0.012139f
C2571 VDDA.n351 GNDA 0.012139f
C2572 VDDA.n352 GNDA 0.012139f
C2573 VDDA.n353 GNDA 0.024151f
C2574 VDDA.n354 GNDA 0.03075f
C2575 VDDA.n355 GNDA 0.012139f
C2576 VDDA.n356 GNDA 0.021244f
C2577 VDDA.n357 GNDA 0.021244f
C2578 VDDA.n358 GNDA 0.012139f
C2579 VDDA.n359 GNDA 0.012139f
C2580 VDDA.n360 GNDA 0.021244f
C2581 VDDA.n361 GNDA 0.021244f
C2582 VDDA.n362 GNDA 0.012139f
C2583 VDDA.n363 GNDA 0.012139f
C2584 VDDA.n364 GNDA 0.021244f
C2585 VDDA.n365 GNDA 0.021244f
C2586 VDDA.n366 GNDA 0.012139f
C2587 VDDA.n367 GNDA 0.012139f
C2588 VDDA.n368 GNDA 0.021244f
C2589 VDDA.n369 GNDA 0.021244f
C2590 VDDA.n370 GNDA 0.012139f
C2591 VDDA.n371 GNDA 0.012139f
C2592 VDDA.n372 GNDA 0.021244f
C2593 VDDA.n373 GNDA 0.024151f
C2594 VDDA.n375 GNDA 0.024075f
C2595 VDDA.n376 GNDA 0.012139f
C2596 VDDA.n377 GNDA 0.286488f
C2597 VDDA.t291 GNDA 0.237931f
C2598 VDDA.t119 GNDA 0.213652f
C2599 VDDA.t117 GNDA 0.213652f
C2600 VDDA.t392 GNDA 0.213652f
C2601 VDDA.t19 GNDA 0.213652f
C2602 VDDA.t194 GNDA 0.213652f
C2603 VDDA.t53 GNDA 0.213652f
C2604 VDDA.t114 GNDA 0.213652f
C2605 VDDA.t55 GNDA 0.213652f
C2606 VDDA.t67 GNDA 0.213652f
C2607 VDDA.t57 GNDA 0.213652f
C2608 VDDA.t279 GNDA 0.237931f
C2609 VDDA.n378 GNDA 0.012139f
C2610 VDDA.n379 GNDA 0.021244f
C2611 VDDA.n380 GNDA 0.024151f
C2612 VDDA.n381 GNDA 0.012139f
C2613 VDDA.n382 GNDA 0.012139f
C2614 VDDA.n385 GNDA 0.012139f
C2615 VDDA.n386 GNDA 0.012139f
C2616 VDDA.n387 GNDA 0.024151f
C2617 VDDA.n388 GNDA 0.03075f
C2618 VDDA.n389 GNDA 0.012139f
C2619 VDDA.n390 GNDA 0.021244f
C2620 VDDA.n391 GNDA 0.021244f
C2621 VDDA.n392 GNDA 0.012139f
C2622 VDDA.n393 GNDA 0.012139f
C2623 VDDA.n394 GNDA 0.021244f
C2624 VDDA.n395 GNDA 0.021244f
C2625 VDDA.n396 GNDA 0.012139f
C2626 VDDA.n397 GNDA 0.012139f
C2627 VDDA.n398 GNDA 0.021244f
C2628 VDDA.n399 GNDA 0.021244f
C2629 VDDA.n400 GNDA 0.012139f
C2630 VDDA.n401 GNDA 0.012139f
C2631 VDDA.n402 GNDA 0.021244f
C2632 VDDA.n403 GNDA 0.021244f
C2633 VDDA.n404 GNDA 0.021244f
C2634 VDDA.n405 GNDA 0.012139f
C2635 VDDA.n406 GNDA 0.286488f
C2636 VDDA.n408 GNDA 0.026793f
C2637 VDDA.t278 GNDA 0.044126f
C2638 VDDA.n409 GNDA 0.035525f
C2639 VDDA.n410 GNDA 0.049381f
C2640 VDDA.n411 GNDA 0.128991f
C2641 VDDA.n412 GNDA 0.148584f
C2642 VDDA.n413 GNDA 0.132787f
C2643 VDDA.t208 GNDA 0.010925f
C2644 VDDA.t304 GNDA 0.010925f
C2645 VDDA.n414 GNDA 0.02535f
C2646 VDDA.n415 GNDA 0.082247f
C2647 VDDA.t295 GNDA 0.038764f
C2648 VDDA.t302 GNDA 0.022412f
C2649 VDDA.n416 GNDA 0.044333f
C2650 VDDA.t305 GNDA 0.038764f
C2651 VDDA.n417 GNDA 0.072776f
C2652 VDDA.t303 GNDA 0.12989f
C2653 VDDA.t207 GNDA 0.08012f
C2654 VDDA.t294 GNDA 0.12989f
C2655 VDDA.n418 GNDA 0.072776f
C2656 VDDA.t293 GNDA 0.022412f
C2657 VDDA.n419 GNDA 0.044023f
C2658 VDDA.n420 GNDA 0.04119f
C2659 VDDA.n421 GNDA 0.058359f
C2660 VDDA.n422 GNDA 0.08557f
C2661 VDDA.t356 GNDA 0.021244f
C2662 VDDA.n423 GNDA 0.063731f
C2663 VDDA.n424 GNDA 0.021244f
C2664 VDDA.n425 GNDA 0.012139f
C2665 VDDA.n429 GNDA 0.012139f
C2666 VDDA.t324 GNDA 0.037247f
C2667 VDDA.n430 GNDA 0.03103f
C2668 VDDA.n431 GNDA 0.021244f
C2669 VDDA.n433 GNDA 0.021244f
C2670 VDDA.n434 GNDA 0.012139f
C2671 VDDA.n435 GNDA 0.012139f
C2672 VDDA.n436 GNDA 0.021244f
C2673 VDDA.n438 GNDA 0.021244f
C2674 VDDA.n439 GNDA 0.012139f
C2675 VDDA.n440 GNDA 0.012139f
C2676 VDDA.n441 GNDA 0.021244f
C2677 VDDA.n442 GNDA 0.021429f
C2678 VDDA.t249 GNDA 0.021244f
C2679 VDDA.n443 GNDA 0.07362f
C2680 VDDA.t326 GNDA 0.042488f
C2681 VDDA.n444 GNDA 0.063731f
C2682 VDDA.n445 GNDA 0.020479f
C2683 VDDA.n446 GNDA 0.012139f
C2684 VDDA.n447 GNDA 0.177538f
C2685 VDDA.t325 GNDA 0.153866f
C2686 VDDA.t248 GNDA 0.14203f
C2687 VDDA.t355 GNDA 0.153866f
C2688 VDDA.n450 GNDA 0.012139f
C2689 VDDA.n452 GNDA 0.021429f
C2690 VDDA.n453 GNDA 0.021244f
C2691 VDDA.n454 GNDA 0.012139f
C2692 VDDA.n455 GNDA 0.012139f
C2693 VDDA.n456 GNDA 0.021244f
C2694 VDDA.n458 GNDA 0.021244f
C2695 VDDA.n459 GNDA 0.021244f
C2696 VDDA.n460 GNDA 0.012139f
C2697 VDDA.n461 GNDA 0.177538f
C2698 VDDA.n463 GNDA 0.023197f
C2699 VDDA.t354 GNDA 0.037247f
C2700 VDDA.n464 GNDA 0.030719f
C2701 VDDA.n465 GNDA 0.04119f
C2702 VDDA.n466 GNDA 0.17223f
C2703 VDDA.n467 GNDA 3.26143f
C2704 VDDA.t2 GNDA 0.339295f
C2705 VDDA.t95 GNDA 0.340524f
C2706 VDDA.t390 GNDA 0.322315f
C2707 VDDA.t100 GNDA 0.339295f
C2708 VDDA.t123 GNDA 0.340524f
C2709 VDDA.t51 GNDA 0.322315f
C2710 VDDA.t50 GNDA 0.339295f
C2711 VDDA.t83 GNDA 0.340524f
C2712 VDDA.t23 GNDA 0.322315f
C2713 VDDA.t104 GNDA 0.339295f
C2714 VDDA.t408 GNDA 0.340524f
C2715 VDDA.t92 GNDA 0.322315f
C2716 VDDA.t133 GNDA 0.339295f
C2717 VDDA.t391 GNDA 0.340524f
C2718 VDDA.t122 GNDA 0.322315f
C2719 VDDA.n468 GNDA 0.22743f
C2720 VDDA.t134 GNDA 0.181114f
C2721 VDDA.n469 GNDA 0.246766f
C2722 VDDA.t121 GNDA 0.181114f
C2723 VDDA.n470 GNDA 0.246766f
C2724 VDDA.t52 GNDA 0.181114f
C2725 VDDA.n471 GNDA 0.246766f
C2726 VDDA.t103 GNDA 0.181114f
C2727 VDDA.n472 GNDA 0.246766f
C2728 VDDA.t3 GNDA 0.317282f
C2729 VDDA.n473 GNDA 2.81776f
C2730 VDDA.t415 GNDA 0.671028f
C2731 VDDA.t417 GNDA 0.715187f
C2732 VDDA.t418 GNDA 0.714907f
C2733 VDDA.t416 GNDA 0.687995f
C2734 VDDA.n474 GNDA 0.478915f
C2735 VDDA.n475 GNDA 0.235185f
C2736 VDDA.n476 GNDA 0.341859f
C2737 VDDA.n477 GNDA 0.624023f
C2738 VDDA.n478 GNDA 0.015267f
C2739 VDDA.n479 GNDA 0.061818f
C2740 VDDA.n480 GNDA 0.02567f
C2741 VDDA.t317 GNDA 0.021113f
C2742 VDDA.n482 GNDA 0.02567f
C2743 VDDA.n483 GNDA 0.015267f
C2744 VDDA.n484 GNDA 0.061818f
C2745 VDDA.t301 GNDA 0.02126f
C2746 VDDA.n485 GNDA 0.02567f
C2747 VDDA.n486 GNDA 0.015267f
C2748 VDDA.n487 GNDA 0.061818f
C2749 VDDA.n488 GNDA 0.015267f
C2750 VDDA.n489 GNDA 0.061818f
C2751 VDDA.n490 GNDA 0.015267f
C2752 VDDA.n491 GNDA 0.061818f
C2753 VDDA.n492 GNDA 0.015267f
C2754 VDDA.n493 GNDA 0.061818f
C2755 VDDA.n494 GNDA 0.015267f
C2756 VDDA.n495 GNDA 0.061818f
C2757 VDDA.n496 GNDA 0.015267f
C2758 VDDA.n497 GNDA 0.061818f
C2759 VDDA.n498 GNDA 0.015267f
C2760 VDDA.n499 GNDA 0.061818f
C2761 VDDA.n500 GNDA 0.015267f
C2762 VDDA.n501 GNDA 0.088837f
C2763 VDDA.n502 GNDA 0.023536f
C2764 VDDA.t275 GNDA 0.022406f
C2765 VDDA.t277 GNDA 0.021113f
C2766 VDDA.n503 GNDA 0.040469f
C2767 VDDA.n504 GNDA 0.061517f
C2768 VDDA.t276 GNDA 0.076292f
C2769 VDDA.t396 GNDA 0.050985f
C2770 VDDA.t166 GNDA 0.050985f
C2771 VDDA.t42 GNDA 0.050985f
C2772 VDDA.t178 GNDA 0.050985f
C2773 VDDA.t160 GNDA 0.050985f
C2774 VDDA.t174 GNDA 0.050985f
C2775 VDDA.t154 GNDA 0.050985f
C2776 VDDA.t400 GNDA 0.050985f
C2777 VDDA.t205 GNDA 0.050985f
C2778 VDDA.t17 GNDA 0.050985f
C2779 VDDA.t186 GNDA 0.050985f
C2780 VDDA.t64 GNDA 0.050985f
C2781 VDDA.t411 GNDA 0.050985f
C2782 VDDA.t413 GNDA 0.050985f
C2783 VDDA.t383 GNDA 0.050985f
C2784 VDDA.t158 GNDA 0.050985f
C2785 VDDA.t184 GNDA 0.050985f
C2786 VDDA.t398 GNDA 0.050985f
C2787 VDDA.t300 GNDA 0.077771f
C2788 VDDA.n505 GNDA 0.110736f
C2789 VDDA.t299 GNDA 0.015025f
C2790 VDDA.n506 GNDA 0.024829f
C2791 VDDA.n507 GNDA 0.045214f
C2792 VDDA.n508 GNDA 0.015267f
C2793 VDDA.n509 GNDA 0.061818f
C2794 VDDA.n510 GNDA 0.015267f
C2795 VDDA.n511 GNDA 0.061818f
C2796 VDDA.n512 GNDA 0.015267f
C2797 VDDA.n513 GNDA 0.061818f
C2798 VDDA.n514 GNDA 0.015267f
C2799 VDDA.n515 GNDA 0.061818f
C2800 VDDA.n516 GNDA 0.015267f
C2801 VDDA.n517 GNDA 0.061818f
C2802 VDDA.n518 GNDA 0.015267f
C2803 VDDA.n519 GNDA 0.061818f
C2804 VDDA.n520 GNDA 0.015267f
C2805 VDDA.n521 GNDA 0.061818f
C2806 VDDA.n522 GNDA 0.015267f
C2807 VDDA.n523 GNDA 0.061818f
C2808 VDDA.n524 GNDA 0.045214f
C2809 VDDA.n525 GNDA 0.022336f
C2810 VDDA.t339 GNDA 0.022406f
C2811 VDDA.t341 GNDA 0.021113f
C2812 VDDA.n526 GNDA 0.040469f
C2813 VDDA.n527 GNDA 0.061517f
C2814 VDDA.t340 GNDA 0.076292f
C2815 VDDA.t15 GNDA 0.050985f
C2816 VDDA.t203 GNDA 0.050985f
C2817 VDDA.t394 GNDA 0.050985f
C2818 VDDA.t182 GNDA 0.050985f
C2819 VDDA.t201 GNDA 0.050985f
C2820 VDDA.t129 GNDA 0.050985f
C2821 VDDA.t404 GNDA 0.050985f
C2822 VDDA.t33 GNDA 0.050985f
C2823 VDDA.t36 GNDA 0.050985f
C2824 VDDA.t180 GNDA 0.050985f
C2825 VDDA.t86 GNDA 0.050985f
C2826 VDDA.t402 GNDA 0.050985f
C2827 VDDA.t156 GNDA 0.050985f
C2828 VDDA.t381 GNDA 0.050985f
C2829 VDDA.t44 GNDA 0.050985f
C2830 VDDA.t379 GNDA 0.050985f
C2831 VDDA.t84 GNDA 0.050985f
C2832 VDDA.t176 GNDA 0.050985f
C2833 VDDA.t316 GNDA 0.06299f
C2834 VDDA.n528 GNDA 0.074818f
C2835 VDDA.n529 GNDA 0.040632f
C2836 VDDA.t315 GNDA 0.022395f
C2837 VDDA.n530 GNDA 0.022336f
C2838 VDDA.n531 GNDA 0.104784f
C2839 VDDA.n532 GNDA 0.202032f
C2840 VDDA.t407 GNDA 0.018209f
C2841 VDDA.t82 GNDA 0.018209f
C2842 VDDA.n533 GNDA 0.060157f
C2843 VDDA.n534 GNDA 0.077625f
C2844 VDDA.n536 GNDA 0.012139f
C2845 VDDA.n539 GNDA 0.012139f
C2846 VDDA.n540 GNDA 0.012139f
C2847 VDDA.n541 GNDA 0.021117f
C2848 VDDA.n542 GNDA 0.012139f
C2849 VDDA.n543 GNDA 0.012139f
C2850 VDDA.n544 GNDA 0.012139f
C2851 VDDA.n545 GNDA 0.021244f
C2852 VDDA.t296 GNDA 0.086828f
C2853 VDDA.t336 GNDA 0.011507f
C2854 VDDA.n546 GNDA 0.029817f
C2855 VDDA.t374 GNDA 0.024234f
C2856 VDDA.t338 GNDA 0.02126f
C2857 VDDA.n547 GNDA 0.106358f
C2858 VDDA.t337 GNDA 0.073651f
C2859 VDDA.t153 GNDA 0.046736f
C2860 VDDA.t32 GNDA 0.046736f
C2861 VDDA.t373 GNDA 0.075272f
C2862 VDDA.n548 GNDA 0.111391f
C2863 VDDA.t372 GNDA 0.011507f
C2864 VDDA.n549 GNDA 0.02959f
C2865 VDDA.n550 GNDA 0.089011f
C2866 VDDA.t1 GNDA 0.018209f
C2867 VDDA.t389 GNDA 0.018209f
C2868 VDDA.n551 GNDA 0.060157f
C2869 VDDA.n552 GNDA 0.077625f
C2870 VDDA.t97 GNDA 0.018209f
C2871 VDDA.t99 GNDA 0.018209f
C2872 VDDA.n553 GNDA 0.060157f
C2873 VDDA.n554 GNDA 0.077625f
C2874 VDDA.t27 GNDA 0.018209f
C2875 VDDA.t108 GNDA 0.018209f
C2876 VDDA.n555 GNDA 0.060157f
C2877 VDDA.n556 GNDA 0.077625f
C2878 VDDA.t106 GNDA 0.018209f
C2879 VDDA.t29 GNDA 0.018209f
C2880 VDDA.n557 GNDA 0.060157f
C2881 VDDA.n558 GNDA 0.077625f
C2882 VDDA.t25 GNDA 0.018209f
C2883 VDDA.t410 GNDA 0.018209f
C2884 VDDA.n559 GNDA 0.060157f
C2885 VDDA.n560 GNDA 0.077625f
C2886 VDDA.t102 GNDA 0.018209f
C2887 VDDA.t94 GNDA 0.018209f
C2888 VDDA.n561 GNDA 0.060157f
C2889 VDDA.n562 GNDA 0.077625f
C2890 VDDA.t110 GNDA 0.018209f
C2891 VDDA.t132 GNDA 0.018209f
C2892 VDDA.n563 GNDA 0.060157f
C2893 VDDA.n564 GNDA 0.077625f
C2894 VDDA.n565 GNDA 0.041445f
C2895 VDDA.n566 GNDA 0.032427f
C2896 VDDA.n567 GNDA 0.024075f
C2897 VDDA.n569 GNDA 0.021117f
C2898 VDDA.n570 GNDA 0.021244f
C2899 VDDA.n571 GNDA 0.021244f
C2900 VDDA.n572 GNDA 0.021244f
C2901 VDDA.n573 GNDA 0.03075f
C2902 VDDA.n574 GNDA 0.012776f
C2903 VDDA.n575 GNDA 0.170254f
C2904 VDDA.t297 GNDA 0.180573f
C2905 VDDA.t109 GNDA 0.185732f
C2906 VDDA.t131 GNDA 0.185732f
C2907 VDDA.t101 GNDA 0.185732f
C2908 VDDA.t93 GNDA 0.185732f
C2909 VDDA.t24 GNDA 0.185732f
C2910 VDDA.t409 GNDA 0.185732f
C2911 VDDA.t105 GNDA 0.185732f
C2912 VDDA.t28 GNDA 0.185732f
C2913 VDDA.t26 GNDA 0.185732f
C2914 VDDA.t107 GNDA 0.185732f
C2915 VDDA.t96 GNDA 0.185732f
C2916 VDDA.t98 GNDA 0.185732f
C2917 VDDA.t0 GNDA 0.185732f
C2918 VDDA.t388 GNDA 0.185732f
C2919 VDDA.t406 GNDA 0.185732f
C2920 VDDA.t81 GNDA 0.185732f
C2921 VDDA.t267 GNDA 0.180573f
C2922 VDDA.n577 GNDA 0.012139f
C2923 VDDA.n578 GNDA 0.012139f
C2924 VDDA.n579 GNDA 0.021244f
C2925 VDDA.n580 GNDA 0.021117f
C2926 VDDA.n581 GNDA 0.021244f
C2927 VDDA.n582 GNDA 0.012139f
C2928 VDDA.n583 GNDA 0.021244f
C2929 VDDA.n584 GNDA 0.021244f
C2930 VDDA.n585 GNDA 0.021117f
C2931 VDDA.n586 GNDA 0.033547f
C2932 VDDA.n588 GNDA 0.170254f
C2933 VDDA.n589 GNDA 0.012139f
C2934 VDDA.n590 GNDA 0.024075f
C2935 VDDA.t266 GNDA 0.086828f
C2936 VDDA.n591 GNDA 0.032427f
C2937 VDDA.n592 GNDA 0.047819f
C2938 VDDA.t312 GNDA 0.011209f
C2939 VDDA.n593 GNDA 0.023952f
C2940 VDDA.t311 GNDA 0.02126f
C2941 VDDA.t314 GNDA 0.02126f
C2942 VDDA.n594 GNDA 0.105759f
C2943 VDDA.t313 GNDA 0.073651f
C2944 VDDA.t30 GNDA 0.046736f
C2945 VDDA.t218 GNDA 0.046736f
C2946 VDDA.t310 GNDA 0.073651f
C2947 VDDA.n595 GNDA 0.10576f
C2948 VDDA.t309 GNDA 0.011209f
C2949 VDDA.n596 GNDA 0.023952f
C2950 VDDA.n597 GNDA 0.057613f
C2951 VDDA.n598 GNDA 0.014639f
C2952 VDDA.n599 GNDA 0.051399f
C2953 VDDA.n600 GNDA 0.119345f
C2954 VDDA.n601 GNDA 0.164837f
C2955 VDDA.n602 GNDA 0.015141f
C2956 VDDA.n603 GNDA 0.053446f
C2957 VDDA.t359 GNDA 0.022129f
C2958 VDDA.t283 GNDA 0.022129f
C2959 VDDA.t281 GNDA 0.011953f
C2960 VDDA.n604 GNDA 0.015113f
C2961 VDDA.n605 GNDA 0.053475f
C2962 VDDA.t363 GNDA 0.011953f
C2963 VDDA.n606 GNDA 0.015147f
C2964 VDDA.n607 GNDA 0.05344f
C2965 VDDA.t271 GNDA 0.02214f
C2966 VDDA.t350 GNDA 0.02214f
C2967 VDDA.t348 GNDA 0.011953f
C2968 VDDA.n608 GNDA 0.015147f
C2969 VDDA.n609 GNDA 0.073142f
C2970 VDDA.n610 GNDA 0.025387f
C2971 VDDA.n611 GNDA 0.063181f
C2972 VDDA.t349 GNDA 0.066585f
C2973 VDDA.t21 GNDA 0.046736f
C2974 VDDA.t145 GNDA 0.046736f
C2975 VDDA.t214 GNDA 0.046736f
C2976 VDDA.t48 GNDA 0.046736f
C2977 VDDA.t270 GNDA 0.066585f
C2978 VDDA.n612 GNDA 0.063181f
C2979 VDDA.t269 GNDA 0.012332f
C2980 VDDA.n613 GNDA 0.024963f
C2981 VDDA.n614 GNDA 0.036893f
C2982 VDDA.n615 GNDA 0.015113f
C2983 VDDA.n616 GNDA 0.053475f
C2984 VDDA.n617 GNDA 0.015113f
C2985 VDDA.n618 GNDA 0.053475f
C2986 VDDA.n619 GNDA 0.015113f
C2987 VDDA.n620 GNDA 0.053475f
C2988 VDDA.n621 GNDA 0.015113f
C2989 VDDA.n622 GNDA 0.053475f
C2990 VDDA.n623 GNDA 0.036893f
C2991 VDDA.n624 GNDA 0.023615f
C2992 VDDA.t365 GNDA 0.021217f
C2993 VDDA.n625 GNDA 0.064903f
C2994 VDDA.t364 GNDA 0.066755f
C2995 VDDA.t90 GNDA 0.046736f
C2996 VDDA.t377 GNDA 0.046736f
C2997 VDDA.t199 GNDA 0.046736f
C2998 VDDA.t6 GNDA 0.046736f
C2999 VDDA.t88 GNDA 0.046736f
C3000 VDDA.t46 GNDA 0.046736f
C3001 VDDA.t164 GNDA 0.046736f
C3002 VDDA.t111 GNDA 0.046736f
C3003 VDDA.t212 GNDA 0.046736f
C3004 VDDA.t216 GNDA 0.046736f
C3005 VDDA.t343 GNDA 0.066755f
C3006 VDDA.t344 GNDA 0.021217f
C3007 VDDA.n626 GNDA 0.064903f
C3008 VDDA.t342 GNDA 0.011953f
C3009 VDDA.n627 GNDA 0.023615f
C3010 VDDA.n628 GNDA 0.036893f
C3011 VDDA.n629 GNDA 0.015141f
C3012 VDDA.n630 GNDA 0.053446f
C3013 VDDA.n631 GNDA 0.036893f
C3014 VDDA.n632 GNDA 0.024584f
C3015 VDDA.n633 GNDA 0.063193f
C3016 VDDA.t282 GNDA 0.066585f
C3017 VDDA.t8 GNDA 0.046736f
C3018 VDDA.t4 GNDA 0.046736f
C3019 VDDA.t151 GNDA 0.046736f
C3020 VDDA.t13 GNDA 0.046736f
C3021 VDDA.t358 GNDA 0.066585f
C3022 VDDA.n634 GNDA 0.063193f
C3023 VDDA.t357 GNDA 0.011953f
C3024 VDDA.n635 GNDA 0.024584f
C3025 VDDA.n636 GNDA 0.122741f
C3026 VDDA.n637 GNDA 0.143295f
C3027 VDDA.n638 GNDA 0.683128f
C3028 two_stage_opamp_dummy_magic_14_0.Vb3.t4 GNDA 0.014599f
C3029 two_stage_opamp_dummy_magic_14_0.Vb3.t6 GNDA 0.014599f
C3030 two_stage_opamp_dummy_magic_14_0.Vb3.n0 GNDA 0.047024f
C3031 two_stage_opamp_dummy_magic_14_0.Vb3.t3 GNDA 0.014599f
C3032 two_stage_opamp_dummy_magic_14_0.Vb3.t7 GNDA 0.014599f
C3033 two_stage_opamp_dummy_magic_14_0.Vb3.n1 GNDA 0.047024f
C3034 two_stage_opamp_dummy_magic_14_0.Vb3.n2 GNDA 0.25924f
C3035 two_stage_opamp_dummy_magic_14_0.Vb3.t2 GNDA 0.014599f
C3036 two_stage_opamp_dummy_magic_14_0.Vb3.t5 GNDA 0.014599f
C3037 two_stage_opamp_dummy_magic_14_0.Vb3.n3 GNDA 0.044094f
C3038 two_stage_opamp_dummy_magic_14_0.Vb3.n4 GNDA 0.785193f
C3039 two_stage_opamp_dummy_magic_14_0.Vb3.t1 GNDA 0.051095f
C3040 two_stage_opamp_dummy_magic_14_0.Vb3.t0 GNDA 0.051095f
C3041 two_stage_opamp_dummy_magic_14_0.Vb3.n5 GNDA 0.180135f
C3042 two_stage_opamp_dummy_magic_14_0.Vb3.t28 GNDA 0.072263f
C3043 two_stage_opamp_dummy_magic_14_0.Vb3.t9 GNDA 0.072263f
C3044 two_stage_opamp_dummy_magic_14_0.Vb3.t12 GNDA 0.072263f
C3045 two_stage_opamp_dummy_magic_14_0.Vb3.t18 GNDA 0.072263f
C3046 two_stage_opamp_dummy_magic_14_0.Vb3.t16 GNDA 0.083391f
C3047 two_stage_opamp_dummy_magic_14_0.Vb3.n6 GNDA 0.067705f
C3048 two_stage_opamp_dummy_magic_14_0.Vb3.n7 GNDA 0.041606f
C3049 two_stage_opamp_dummy_magic_14_0.Vb3.n8 GNDA 0.041606f
C3050 two_stage_opamp_dummy_magic_14_0.Vb3.n9 GNDA 0.038604f
C3051 two_stage_opamp_dummy_magic_14_0.Vb3.t27 GNDA 0.072263f
C3052 two_stage_opamp_dummy_magic_14_0.Vb3.t21 GNDA 0.072263f
C3053 two_stage_opamp_dummy_magic_14_0.Vb3.t17 GNDA 0.072263f
C3054 two_stage_opamp_dummy_magic_14_0.Vb3.t11 GNDA 0.072263f
C3055 two_stage_opamp_dummy_magic_14_0.Vb3.t8 GNDA 0.083391f
C3056 two_stage_opamp_dummy_magic_14_0.Vb3.n10 GNDA 0.067705f
C3057 two_stage_opamp_dummy_magic_14_0.Vb3.n11 GNDA 0.041606f
C3058 two_stage_opamp_dummy_magic_14_0.Vb3.n12 GNDA 0.041606f
C3059 two_stage_opamp_dummy_magic_14_0.Vb3.n13 GNDA 0.038604f
C3060 two_stage_opamp_dummy_magic_14_0.Vb3.n14 GNDA 0.040946f
C3061 two_stage_opamp_dummy_magic_14_0.Vb3.t10 GNDA 0.072263f
C3062 two_stage_opamp_dummy_magic_14_0.Vb3.t15 GNDA 0.072263f
C3063 two_stage_opamp_dummy_magic_14_0.Vb3.t20 GNDA 0.072263f
C3064 two_stage_opamp_dummy_magic_14_0.Vb3.t24 GNDA 0.072263f
C3065 two_stage_opamp_dummy_magic_14_0.Vb3.t22 GNDA 0.083391f
C3066 two_stage_opamp_dummy_magic_14_0.Vb3.n15 GNDA 0.067705f
C3067 two_stage_opamp_dummy_magic_14_0.Vb3.n16 GNDA 0.041606f
C3068 two_stage_opamp_dummy_magic_14_0.Vb3.n17 GNDA 0.041606f
C3069 two_stage_opamp_dummy_magic_14_0.Vb3.n18 GNDA 0.038604f
C3070 two_stage_opamp_dummy_magic_14_0.Vb3.t25 GNDA 0.072263f
C3071 two_stage_opamp_dummy_magic_14_0.Vb3.t26 GNDA 0.072263f
C3072 two_stage_opamp_dummy_magic_14_0.Vb3.t23 GNDA 0.072263f
C3073 two_stage_opamp_dummy_magic_14_0.Vb3.t19 GNDA 0.072263f
C3074 two_stage_opamp_dummy_magic_14_0.Vb3.t13 GNDA 0.083391f
C3075 two_stage_opamp_dummy_magic_14_0.Vb3.n19 GNDA 0.067705f
C3076 two_stage_opamp_dummy_magic_14_0.Vb3.n20 GNDA 0.041606f
C3077 two_stage_opamp_dummy_magic_14_0.Vb3.n21 GNDA 0.041606f
C3078 two_stage_opamp_dummy_magic_14_0.Vb3.n22 GNDA 0.038604f
C3079 two_stage_opamp_dummy_magic_14_0.Vb3.n23 GNDA 0.04262f
C3080 two_stage_opamp_dummy_magic_14_0.Vb3.n24 GNDA 1.17334f
C3081 two_stage_opamp_dummy_magic_14_0.Vb3.t14 GNDA 0.08858f
C3082 two_stage_opamp_dummy_magic_14_0.Vb3.n25 GNDA 0.307922f
C3083 two_stage_opamp_dummy_magic_14_0.Vb3.n26 GNDA 0.912484f
C3084 bgr_0.VB3_CUR_BIAS GNDA 1.63375f
C3085 bgr_0.NFET_GATE_10uA.t1 GNDA 0.01496f
C3086 bgr_0.NFET_GATE_10uA.t4 GNDA 0.01496f
C3087 bgr_0.NFET_GATE_10uA.n0 GNDA 0.042091f
C3088 bgr_0.NFET_GATE_10uA.t18 GNDA 0.014586f
C3089 bgr_0.NFET_GATE_10uA.t6 GNDA 0.014586f
C3090 bgr_0.NFET_GATE_10uA.t14 GNDA 0.014586f
C3091 bgr_0.NFET_GATE_10uA.t19 GNDA 0.014586f
C3092 bgr_0.NFET_GATE_10uA.t5 GNDA 0.014586f
C3093 bgr_0.NFET_GATE_10uA.t13 GNDA 0.014586f
C3094 bgr_0.NFET_GATE_10uA.t12 GNDA 0.021563f
C3095 bgr_0.NFET_GATE_10uA.n1 GNDA 0.026685f
C3096 bgr_0.NFET_GATE_10uA.n2 GNDA 0.019075f
C3097 bgr_0.NFET_GATE_10uA.n3 GNDA 0.016149f
C3098 bgr_0.NFET_GATE_10uA.t15 GNDA 0.014586f
C3099 bgr_0.NFET_GATE_10uA.t8 GNDA 0.014586f
C3100 bgr_0.NFET_GATE_10uA.t21 GNDA 0.014586f
C3101 bgr_0.NFET_GATE_10uA.t16 GNDA 0.021563f
C3102 bgr_0.NFET_GATE_10uA.n4 GNDA 0.026685f
C3103 bgr_0.NFET_GATE_10uA.n5 GNDA 0.019075f
C3104 bgr_0.NFET_GATE_10uA.n6 GNDA 0.016149f
C3105 bgr_0.NFET_GATE_10uA.t20 GNDA 0.014586f
C3106 bgr_0.NFET_GATE_10uA.t7 GNDA 0.021563f
C3107 bgr_0.NFET_GATE_10uA.n7 GNDA 0.02376f
C3108 bgr_0.NFET_GATE_10uA.n8 GNDA 0.026114f
C3109 bgr_0.NFET_GATE_10uA.t11 GNDA 0.014586f
C3110 bgr_0.NFET_GATE_10uA.t22 GNDA 0.021563f
C3111 bgr_0.NFET_GATE_10uA.n9 GNDA 0.02376f
C3112 bgr_0.NFET_GATE_10uA.t9 GNDA 0.014586f
C3113 bgr_0.NFET_GATE_10uA.t17 GNDA 0.014586f
C3114 bgr_0.NFET_GATE_10uA.t23 GNDA 0.014586f
C3115 bgr_0.NFET_GATE_10uA.t10 GNDA 0.021563f
C3116 bgr_0.NFET_GATE_10uA.n10 GNDA 0.026685f
C3117 bgr_0.NFET_GATE_10uA.n11 GNDA 0.019075f
C3118 bgr_0.NFET_GATE_10uA.n12 GNDA 0.016149f
C3119 bgr_0.NFET_GATE_10uA.n13 GNDA 0.026114f
C3120 bgr_0.NFET_GATE_10uA.n14 GNDA 0.605807f
C3121 bgr_0.NFET_GATE_10uA.n15 GNDA 0.022264f
C3122 bgr_0.NFET_GATE_10uA.n16 GNDA 0.016149f
C3123 bgr_0.NFET_GATE_10uA.n17 GNDA 0.019075f
C3124 bgr_0.NFET_GATE_10uA.n18 GNDA 0.026685f
C3125 bgr_0.NFET_GATE_10uA.t3 GNDA 0.034164f
C3126 bgr_0.NFET_GATE_10uA.n19 GNDA 0.327308f
C3127 bgr_0.NFET_GATE_10uA.t0 GNDA 0.01496f
C3128 bgr_0.NFET_GATE_10uA.t2 GNDA 0.01496f
C3129 bgr_0.NFET_GATE_10uA.n20 GNDA 0.088541f
.ends

