* PEX produced on Sat Feb  1 02:26:17 PM CET 2025 using /foss/tools/osic-multitool/iic-pex.sh with m=3 and s=1
* NGSPICE file created from TSPC_FF_ratioed_divide3_magic.ext - technology: sky130A

.subckt TSPC_FF_ratioed_divide3_magic VOUT VIN VDDA GNDA
X0 C.t3 A.t2 VDDA.t17 VDDA.t16 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X1 VDDA.t15 I.t2 VOUT.t2 VDDA.t14 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X2 VOUT.t0 I.t3 GNDA.t9 GNDA.t8 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X3 D.t0 CLK.t3 VDDA.t11 VDDA.t10 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X4 C.t2 CLK.t4 GNDA.t11 GNDA.t10 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X5 GNDA.t15 VIN.t0 CLK.t2 GNDA.t14 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X6 GNDA.t13 CLK.t5 H.t3 GNDA.t12 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X7 GNDA.t7 I.t4 G.t1 GNDA.t6 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X8 I.t0 CLK.t6 VDDA.t9 VDDA.t8 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X9 VDDA.t5 D.t2 E.t1 VDDA.t4 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X10 GNDA.t2 CLK.t7 C.t0 GNDA.t1 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X11 GNDA.t22 CLK.t8 H.t2 GNDA.t21 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X12 A.t1 CLK.t9 B.t0 GNDA.t20 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X13 F.t0 CLK.t10 E.t0 GNDA.t5 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X14 CLK.t0 VIN.t1 VDDA.t3 VDDA.t2 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X15 VDDA.t7 VOUT.t3 A.t0 VDDA.t6 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X16 VOUT.t1 I.t5 VDDA.t21 VDDA.t20 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X17 I.t1 H.t4 GNDA.t19 GNDA.t18 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X18 GNDA.t4 CLK.t11 C.t1 GNDA.t3 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X19 VDDA.t13 VIN.t2 CLK.t1 VDDA.t12 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X20 E.t2 I.t6 VDDA.t19 VDDA.t18 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X21 D.t1 C.t4 GNDA.t24 GNDA.t23 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X22 H.t1 CLK.t12 GNDA.t26 GNDA.t25 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X23 G.t0 D.t3 F.t1 GNDA.t0 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X24 VDDA.t1 E.t3 H.t0 VDDA.t0 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X25 B.t1 VOUT.t4 GNDA.t17 GNDA.t16 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
R0 A.n0 A.t0 713.933
R1 A.n0 A.t2 314.233
R2 A.t1 A.n0 308.2
R3 VDDA.t10 VDDA.t4 2307.14
R4 VDDA.t8 VDDA.t20 2126.19
R5 VDDA.t18 VDDA.t0 1492.86
R6 VDDA.t6 VDDA.t2 1130.95
R7 VDDA.n7 VDDA.t16 927.381
R8 VDDA.n0 VDDA.t15 673.375
R9 VDDA.n0 VDDA.t21 673.101
R10 VDDA.n6 VDDA.t11 663.801
R11 VDDA.n7 VDDA.t10 610.715
R12 VDDA.n13 VDDA.n12 594.301
R13 VDDA.n11 VDDA.n10 594.301
R14 VDDA.n4 VDDA.n3 594.301
R15 VDDA.n2 VDDA.n1 594.301
R16 VDDA.t20 VDDA.t14 497.62
R17 VDDA.t0 VDDA.t8 497.62
R18 VDDA.t4 VDDA.t18 497.62
R19 VDDA.t16 VDDA.t6 497.62
R20 VDDA.t2 VDDA.t12 497.62
R21 VDDA.n8 VDDA.n7 370
R22 VDDA.n12 VDDA.t3 78.8005
R23 VDDA.n12 VDDA.t13 78.8005
R24 VDDA.n10 VDDA.t17 78.8005
R25 VDDA.n10 VDDA.t7 78.8005
R26 VDDA.n3 VDDA.t19 78.8005
R27 VDDA.n3 VDDA.t5 78.8005
R28 VDDA.n1 VDDA.t9 78.8005
R29 VDDA.n1 VDDA.t1 78.8005
R30 VDDA.n8 VDDA.n6 12.8005
R31 VDDA.n6 VDDA.n5 9.3005
R32 VDDA.n9 VDDA.n8 9.3005
R33 VDDA.n5 VDDA.n4 0.7755
R34 VDDA.n2 VDDA.n0 0.588
R35 VDDA.n4 VDDA.n2 0.5505
R36 VDDA.n13 VDDA.n11 0.4505
R37 VDDA.n11 VDDA.n9 0.3255
R38 VDDA VDDA.n13 0.238
R39 VDDA.n9 VDDA.n5 0.1005
R40 C.n0 C.t3 721.4
R41 C.n1 C.t4 350.349
R42 C.n0 C.t1 276.733
R43 C.n2 C.n1 206.333
R44 C.n1 C.n0 48.0005
R45 C.t0 C.n2 48.0005
R46 C.n2 C.t2 48.0005
R47 I.n0 I.t0 663.801
R48 I.n0 I.t6 568.067
R49 I.t6 I.t4 514.134
R50 I.n3 I.n2 344.8
R51 I.n1 I.t2 289.2
R52 I.t1 I.n3 275.454
R53 I.n2 I.t3 241
R54 I.n1 I.t5 112.468
R55 I.n3 I.n0 97.9205
R56 I.n2 I.n1 64.2672
R57 VOUT.n2 VOUT.t4 4394.23
R58 VOUT.t4 VOUT.t3 819.4
R59 VOUT.n1 VOUT.n0 633
R60 VOUT.n1 VOUT.t0 261.8
R61 VOUT VOUT.n2 256.062
R62 VOUT.n2 VOUT.n1 152
R63 VOUT.n0 VOUT.t2 78.8005
R64 VOUT.n0 VOUT.t1 78.8005
R65 GNDA.t5 GNDA.t23 3723.08
R66 GNDA.t3 GNDA.t20 3723.08
R67 GNDA.t18 GNDA.t8 2820.51
R68 GNDA.n5 GNDA.t21 2200
R69 GNDA.n5 GNDA.t6 1523.08
R70 GNDA.t12 GNDA.t18 1241.03
R71 GNDA.t25 GNDA.t12 1241.03
R72 GNDA.t21 GNDA.t25 1241.03
R73 GNDA.t6 GNDA.t0 1241.03
R74 GNDA.t0 GNDA.t5 1241.03
R75 GNDA.t23 GNDA.t1 1241.03
R76 GNDA.t1 GNDA.t10 1241.03
R77 GNDA.t10 GNDA.t3 1241.03
R78 GNDA.t20 GNDA.t16 1241.03
R79 GNDA.t16 GNDA.t14 1241.03
R80 GNDA.n6 GNDA.n5 1170
R81 GNDA.n1 GNDA.t9 242.613
R82 GNDA.n7 GNDA.t7 233
R83 GNDA.n14 GNDA.n13 194.3
R84 GNDA.n12 GNDA.n11 194.3
R85 GNDA.n10 GNDA.n9 194.3
R86 GNDA.n3 GNDA.n2 194.3
R87 GNDA.n1 GNDA.n0 194.3
R88 GNDA.n13 GNDA.t17 48.0005
R89 GNDA.n13 GNDA.t15 48.0005
R90 GNDA.n11 GNDA.t11 48.0005
R91 GNDA.n11 GNDA.t4 48.0005
R92 GNDA.n9 GNDA.t24 48.0005
R93 GNDA.n9 GNDA.t2 48.0005
R94 GNDA.n2 GNDA.t26 48.0005
R95 GNDA.n2 GNDA.t22 48.0005
R96 GNDA.n0 GNDA.t19 48.0005
R97 GNDA.n0 GNDA.t13 48.0005
R98 GNDA.n7 GNDA.n6 12.8005
R99 GNDA.n6 GNDA.n4 9.3005
R100 GNDA.n8 GNDA.n7 9.3005
R101 GNDA.n10 GNDA.n8 0.8255
R102 GNDA.n14 GNDA.n12 0.688
R103 GNDA.n4 GNDA.n3 0.313
R104 GNDA.n3 GNDA.n1 0.2755
R105 GNDA.n12 GNDA.n10 0.2755
R106 GNDA GNDA.n14 0.238
R107 GNDA.n8 GNDA.n4 0.1005
R108 CLK.n3 CLK.n2 742.51
R109 CLK.n9 CLK.t1 723.534
R110 CLK.n8 CLK.t0 723.534
R111 CLK.n2 CLK.n1 684.806
R112 CLK.n7 CLK.n6 366.856
R113 CLK.n0 CLK.t6 337.401
R114 CLK.n0 CLK.t5 305.267
R115 CLK.t2 CLK.n9 254.333
R116 CLK.n4 CLK.n3 224.934
R117 CLK.n7 CLK.t9 190.123
R118 CLK.n8 CLK.n7 187.201
R119 CLK.n1 CLK.n0 176.733
R120 CLK.n5 CLK.n4 176.733
R121 CLK.n6 CLK.n5 176.733
R122 CLK.n3 CLK.t3 144.601
R123 CLK.n2 CLK.t10 131.976
R124 CLK.n0 CLK.t12 128.534
R125 CLK.n1 CLK.t8 128.534
R126 CLK.n4 CLK.t7 112.468
R127 CLK.n6 CLK.t11 112.468
R128 CLK.n5 CLK.t4 112.468
R129 CLK.n9 CLK.n8 70.4005
R130 D.n1 D.n0 701.467
R131 D.n1 D.t0 694.201
R132 D.n0 D.t3 321.334
R133 D.t1 D.n1 314.921
R134 D.n0 D.t2 144.601
R135 VIN.t2 VIN.t1 401.668
R136 VIN.n0 VIN.t2 257.067
R137 VIN VIN.n0 216.9
R138 VIN.n0 VIN.t0 208.868
R139 H.n0 H.t0 723.534
R140 H.n1 H.t4 553.534
R141 H.n0 H.t2 254.333
R142 H.n2 H.n1 206.333
R143 H.n1 H.n0 70.4005
R144 H.t3 H.n2 48.0005
R145 H.n2 H.t1 48.0005
R146 G.t0 G.t1 96.0005
R147 E.n0 E.t2 685.134
R148 E.n1 E.t1 663.801
R149 E.n0 E.t3 534.268
R150 E.t0 E.n1 362.921
R151 E.n1 E.n0 91.7338
R152 B.t0 B.t1 96.0005
R153 F.t0 F.t1 96.0005
C0 VIN VDDA 0.126677f
C1 VOUT VDDA 0.230937f
C2 VIN VOUT 0.055436f
C3 VOUT GNDA 2.12981f
C4 VIN GNDA 0.291288f
C5 VDDA GNDA 2.83767f
.ends

