magic
tech sky130A
magscale 1 2
timestamp 1756256667
<< nwell >>
rect 33830 840 35470 1120
rect 35730 840 37370 1120
rect 32750 40 33520 320
rect 33820 -160 37380 520
rect 32720 -1320 35450 -1040
rect 35750 -1320 38480 -1040
<< pwell >>
rect 35560 -8550 35640 -8240
<< nmos >>
rect 33760 -2120 33800 -2020
rect 33880 -2120 33920 -2020
rect 34000 -2120 34040 -2020
rect 34120 -2120 34160 -2020
rect 34240 -2120 34280 -2020
rect 34360 -2120 34400 -2020
rect 34480 -2120 34520 -2020
rect 34600 -2120 34640 -2020
rect 34720 -2120 34760 -2020
rect 34840 -2120 34880 -2020
rect 36320 -2120 36360 -2020
rect 36440 -2120 36480 -2020
rect 36560 -2120 36600 -2020
rect 36680 -2120 36720 -2020
rect 36800 -2120 36840 -2020
rect 36920 -2120 36960 -2020
rect 37040 -2120 37080 -2020
rect 37160 -2120 37200 -2020
rect 37280 -2120 37320 -2020
rect 37400 -2120 37440 -2020
rect 33140 -3130 34140 -2630
rect 34380 -3130 35380 -2630
rect 35820 -3130 36820 -2630
rect 37060 -3130 38060 -2630
rect 33560 -3740 35560 -3540
rect 35640 -3740 37640 -3540
<< pmos >>
rect 34030 880 34060 1080
rect 34140 880 34170 1080
rect 34250 880 34280 1080
rect 34360 880 34390 1080
rect 34470 880 34500 1080
rect 34580 880 34610 1080
rect 34690 880 34720 1080
rect 34800 880 34830 1080
rect 34910 880 34940 1080
rect 35020 880 35050 1080
rect 35130 880 35160 1080
rect 35240 880 35270 1080
rect 35930 880 35960 1080
rect 36040 880 36070 1080
rect 36150 880 36180 1080
rect 36260 880 36290 1080
rect 36370 880 36400 1080
rect 36480 880 36510 1080
rect 36590 880 36620 1080
rect 36700 880 36730 1080
rect 36810 880 36840 1080
rect 36920 880 36950 1080
rect 37030 880 37060 1080
rect 37140 880 37170 1080
rect 32950 80 32980 280
rect 33060 80 33090 280
rect 33170 80 33200 280
rect 33280 80 33310 280
rect 34020 -120 34120 480
rect 34200 -120 34300 480
rect 34380 -120 34480 480
rect 34560 -120 34660 480
rect 34740 -120 34840 480
rect 34920 -120 35020 480
rect 35100 -120 35200 480
rect 35280 -120 35380 480
rect 35460 -120 35560 480
rect 35640 -120 35740 480
rect 35820 -120 35920 480
rect 36000 -120 36100 480
rect 36180 -120 36280 480
rect 36360 -120 36460 480
rect 36540 -120 36640 480
rect 36720 -120 36820 480
rect 36900 -120 37000 480
rect 37080 -120 37180 480
rect 32920 -1280 32960 -1080
rect 33040 -1280 33080 -1080
rect 33160 -1280 33200 -1080
rect 33280 -1280 33320 -1080
rect 33400 -1280 33440 -1080
rect 33520 -1280 33560 -1080
rect 33640 -1280 33680 -1080
rect 33760 -1280 33800 -1080
rect 33880 -1280 33920 -1080
rect 34000 -1280 34040 -1080
rect 34120 -1280 34160 -1080
rect 34240 -1280 34280 -1080
rect 34360 -1280 34400 -1080
rect 34480 -1280 34520 -1080
rect 34600 -1280 34640 -1080
rect 34720 -1280 34760 -1080
rect 34840 -1280 34880 -1080
rect 34960 -1280 35000 -1080
rect 35080 -1280 35120 -1080
rect 35200 -1280 35240 -1080
rect 35960 -1280 36000 -1080
rect 36080 -1280 36120 -1080
rect 36200 -1280 36240 -1080
rect 36320 -1280 36360 -1080
rect 36440 -1280 36480 -1080
rect 36560 -1280 36600 -1080
rect 36680 -1280 36720 -1080
rect 36800 -1280 36840 -1080
rect 36920 -1280 36960 -1080
rect 37040 -1280 37080 -1080
rect 37160 -1280 37200 -1080
rect 37280 -1280 37320 -1080
rect 37400 -1280 37440 -1080
rect 37520 -1280 37560 -1080
rect 37640 -1280 37680 -1080
rect 37760 -1280 37800 -1080
rect 37880 -1280 37920 -1080
rect 38000 -1280 38040 -1080
rect 38120 -1280 38160 -1080
rect 38240 -1280 38280 -1080
<< ndiff >>
rect 33680 -2050 33760 -2020
rect 33680 -2090 33700 -2050
rect 33740 -2090 33760 -2050
rect 33680 -2120 33760 -2090
rect 33800 -2050 33880 -2020
rect 33800 -2090 33820 -2050
rect 33860 -2090 33880 -2050
rect 33800 -2120 33880 -2090
rect 33920 -2050 34000 -2020
rect 33920 -2090 33940 -2050
rect 33980 -2090 34000 -2050
rect 33920 -2120 34000 -2090
rect 34040 -2050 34120 -2020
rect 34040 -2090 34060 -2050
rect 34100 -2090 34120 -2050
rect 34040 -2120 34120 -2090
rect 34160 -2050 34240 -2020
rect 34160 -2090 34180 -2050
rect 34220 -2090 34240 -2050
rect 34160 -2120 34240 -2090
rect 34280 -2050 34360 -2020
rect 34280 -2090 34300 -2050
rect 34340 -2090 34360 -2050
rect 34280 -2120 34360 -2090
rect 34400 -2050 34480 -2020
rect 34400 -2090 34420 -2050
rect 34460 -2090 34480 -2050
rect 34400 -2120 34480 -2090
rect 34520 -2050 34600 -2020
rect 34520 -2090 34540 -2050
rect 34580 -2090 34600 -2050
rect 34520 -2120 34600 -2090
rect 34640 -2050 34720 -2020
rect 34640 -2090 34660 -2050
rect 34700 -2090 34720 -2050
rect 34640 -2120 34720 -2090
rect 34760 -2050 34840 -2020
rect 34760 -2090 34780 -2050
rect 34820 -2090 34840 -2050
rect 34760 -2120 34840 -2090
rect 34880 -2050 34960 -2020
rect 34880 -2090 34900 -2050
rect 34940 -2090 34960 -2050
rect 34880 -2120 34960 -2090
rect 36240 -2050 36320 -2020
rect 36240 -2090 36260 -2050
rect 36300 -2090 36320 -2050
rect 36240 -2120 36320 -2090
rect 36360 -2050 36440 -2020
rect 36360 -2090 36380 -2050
rect 36420 -2090 36440 -2050
rect 36360 -2120 36440 -2090
rect 36480 -2050 36560 -2020
rect 36480 -2090 36500 -2050
rect 36540 -2090 36560 -2050
rect 36480 -2120 36560 -2090
rect 36600 -2050 36680 -2020
rect 36600 -2090 36620 -2050
rect 36660 -2090 36680 -2050
rect 36600 -2120 36680 -2090
rect 36720 -2050 36800 -2020
rect 36720 -2090 36740 -2050
rect 36780 -2090 36800 -2050
rect 36720 -2120 36800 -2090
rect 36840 -2050 36920 -2020
rect 36840 -2090 36860 -2050
rect 36900 -2090 36920 -2050
rect 36840 -2120 36920 -2090
rect 36960 -2050 37040 -2020
rect 36960 -2090 36980 -2050
rect 37020 -2090 37040 -2050
rect 36960 -2120 37040 -2090
rect 37080 -2050 37160 -2020
rect 37080 -2090 37100 -2050
rect 37140 -2090 37160 -2050
rect 37080 -2120 37160 -2090
rect 37200 -2050 37280 -2020
rect 37200 -2090 37220 -2050
rect 37260 -2090 37280 -2050
rect 37200 -2120 37280 -2090
rect 37320 -2050 37400 -2020
rect 37320 -2090 37340 -2050
rect 37380 -2090 37400 -2050
rect 37320 -2120 37400 -2090
rect 37440 -2050 37520 -2020
rect 37440 -2090 37460 -2050
rect 37500 -2090 37520 -2050
rect 37440 -2120 37520 -2090
rect 33060 -2660 33140 -2630
rect 33060 -2700 33080 -2660
rect 33120 -2700 33140 -2660
rect 33060 -2760 33140 -2700
rect 33060 -2800 33080 -2760
rect 33120 -2800 33140 -2760
rect 33060 -2860 33140 -2800
rect 33060 -2900 33080 -2860
rect 33120 -2900 33140 -2860
rect 33060 -2960 33140 -2900
rect 33060 -3000 33080 -2960
rect 33120 -3000 33140 -2960
rect 33060 -3060 33140 -3000
rect 33060 -3100 33080 -3060
rect 33120 -3100 33140 -3060
rect 33060 -3130 33140 -3100
rect 34140 -2660 34220 -2630
rect 34300 -2660 34380 -2630
rect 34140 -2700 34160 -2660
rect 34200 -2700 34220 -2660
rect 34300 -2700 34320 -2660
rect 34360 -2700 34380 -2660
rect 34140 -2760 34220 -2700
rect 34300 -2760 34380 -2700
rect 34140 -2800 34160 -2760
rect 34200 -2800 34220 -2760
rect 34300 -2800 34320 -2760
rect 34360 -2800 34380 -2760
rect 34140 -2860 34220 -2800
rect 34300 -2860 34380 -2800
rect 34140 -2900 34160 -2860
rect 34200 -2900 34220 -2860
rect 34300 -2900 34320 -2860
rect 34360 -2900 34380 -2860
rect 34140 -2960 34220 -2900
rect 34300 -2960 34380 -2900
rect 34140 -3000 34160 -2960
rect 34200 -3000 34220 -2960
rect 34300 -3000 34320 -2960
rect 34360 -3000 34380 -2960
rect 34140 -3060 34220 -3000
rect 34300 -3060 34380 -3000
rect 34140 -3100 34160 -3060
rect 34200 -3100 34220 -3060
rect 34300 -3100 34320 -3060
rect 34360 -3100 34380 -3060
rect 34140 -3120 34220 -3100
rect 34300 -3120 34380 -3100
rect 34140 -3130 34380 -3120
rect 35380 -2660 35460 -2630
rect 35380 -2700 35400 -2660
rect 35440 -2700 35460 -2660
rect 35380 -2760 35460 -2700
rect 35380 -2800 35400 -2760
rect 35440 -2800 35460 -2760
rect 35380 -2860 35460 -2800
rect 35380 -2900 35400 -2860
rect 35440 -2900 35460 -2860
rect 35380 -2960 35460 -2900
rect 35380 -3000 35400 -2960
rect 35440 -3000 35460 -2960
rect 35380 -3060 35460 -3000
rect 35380 -3100 35400 -3060
rect 35440 -3100 35460 -3060
rect 35380 -3130 35460 -3100
rect 35740 -2660 35820 -2630
rect 35740 -2700 35760 -2660
rect 35800 -2700 35820 -2660
rect 35740 -2760 35820 -2700
rect 35740 -2800 35760 -2760
rect 35800 -2800 35820 -2760
rect 35740 -2860 35820 -2800
rect 35740 -2900 35760 -2860
rect 35800 -2900 35820 -2860
rect 35740 -2960 35820 -2900
rect 35740 -3000 35760 -2960
rect 35800 -3000 35820 -2960
rect 35740 -3060 35820 -3000
rect 35740 -3100 35760 -3060
rect 35800 -3100 35820 -3060
rect 35740 -3130 35820 -3100
rect 36820 -2660 36900 -2630
rect 36980 -2660 37060 -2630
rect 36820 -2700 36840 -2660
rect 36880 -2700 36900 -2660
rect 36980 -2700 37000 -2660
rect 37040 -2700 37060 -2660
rect 36820 -2760 36900 -2700
rect 36980 -2760 37060 -2700
rect 36820 -2800 36840 -2760
rect 36880 -2800 36900 -2760
rect 36980 -2800 37000 -2760
rect 37040 -2800 37060 -2760
rect 36820 -2860 36900 -2800
rect 36980 -2860 37060 -2800
rect 36820 -2900 36840 -2860
rect 36880 -2900 36900 -2860
rect 36980 -2900 37000 -2860
rect 37040 -2900 37060 -2860
rect 36820 -2960 36900 -2900
rect 36980 -2960 37060 -2900
rect 36820 -3000 36840 -2960
rect 36880 -3000 36900 -2960
rect 36980 -3000 37000 -2960
rect 37040 -3000 37060 -2960
rect 36820 -3060 36900 -3000
rect 36980 -3060 37060 -3000
rect 36820 -3100 36840 -3060
rect 36880 -3100 36900 -3060
rect 36980 -3100 37000 -3060
rect 37040 -3100 37060 -3060
rect 36820 -3130 36900 -3100
rect 36980 -3130 37060 -3100
rect 38060 -2660 38140 -2630
rect 38060 -2700 38080 -2660
rect 38120 -2700 38140 -2660
rect 38060 -2760 38140 -2700
rect 38060 -2800 38080 -2760
rect 38120 -2800 38140 -2760
rect 38060 -2860 38140 -2800
rect 38060 -2900 38080 -2860
rect 38120 -2900 38140 -2860
rect 38060 -2960 38140 -2900
rect 38060 -3000 38080 -2960
rect 38120 -3000 38140 -2960
rect 38060 -3060 38140 -3000
rect 38060 -3100 38080 -3060
rect 38120 -3100 38140 -3060
rect 38060 -3130 38140 -3100
rect 33480 -3570 33560 -3540
rect 33480 -3610 33500 -3570
rect 33540 -3610 33560 -3570
rect 33480 -3670 33560 -3610
rect 33480 -3710 33500 -3670
rect 33540 -3710 33560 -3670
rect 33480 -3740 33560 -3710
rect 35560 -3570 35640 -3540
rect 35560 -3610 35580 -3570
rect 35620 -3610 35640 -3570
rect 35560 -3670 35640 -3610
rect 35560 -3710 35580 -3670
rect 35620 -3710 35640 -3670
rect 35560 -3740 35640 -3710
rect 37640 -3570 37720 -3540
rect 37640 -3610 37660 -3570
rect 37700 -3610 37720 -3570
rect 37640 -3670 37720 -3610
rect 37640 -3710 37660 -3670
rect 37700 -3710 37720 -3670
rect 37640 -3740 37720 -3710
<< pdiff >>
rect 33950 1050 34030 1080
rect 33950 1010 33970 1050
rect 34010 1010 34030 1050
rect 33950 950 34030 1010
rect 33950 910 33970 950
rect 34010 910 34030 950
rect 33950 880 34030 910
rect 34060 1050 34140 1080
rect 34060 1010 34080 1050
rect 34120 1010 34140 1050
rect 34060 950 34140 1010
rect 34060 910 34080 950
rect 34120 910 34140 950
rect 34060 880 34140 910
rect 34170 1050 34250 1080
rect 34170 1010 34190 1050
rect 34230 1010 34250 1050
rect 34170 950 34250 1010
rect 34170 910 34190 950
rect 34230 910 34250 950
rect 34170 880 34250 910
rect 34280 1050 34360 1080
rect 34280 1010 34300 1050
rect 34340 1010 34360 1050
rect 34280 950 34360 1010
rect 34280 910 34300 950
rect 34340 910 34360 950
rect 34280 880 34360 910
rect 34390 1050 34470 1080
rect 34390 1010 34410 1050
rect 34450 1010 34470 1050
rect 34390 950 34470 1010
rect 34390 910 34410 950
rect 34450 910 34470 950
rect 34390 880 34470 910
rect 34500 1050 34580 1080
rect 34500 1010 34520 1050
rect 34560 1010 34580 1050
rect 34500 950 34580 1010
rect 34500 910 34520 950
rect 34560 910 34580 950
rect 34500 880 34580 910
rect 34610 1050 34690 1080
rect 34610 1010 34630 1050
rect 34670 1010 34690 1050
rect 34610 950 34690 1010
rect 34610 910 34630 950
rect 34670 910 34690 950
rect 34610 880 34690 910
rect 34720 1050 34800 1080
rect 34720 1010 34740 1050
rect 34780 1010 34800 1050
rect 34720 950 34800 1010
rect 34720 910 34740 950
rect 34780 910 34800 950
rect 34720 880 34800 910
rect 34830 1050 34910 1080
rect 34830 1010 34850 1050
rect 34890 1010 34910 1050
rect 34830 950 34910 1010
rect 34830 910 34850 950
rect 34890 910 34910 950
rect 34830 880 34910 910
rect 34940 1050 35020 1080
rect 34940 1010 34960 1050
rect 35000 1010 35020 1050
rect 34940 950 35020 1010
rect 34940 910 34960 950
rect 35000 910 35020 950
rect 34940 880 35020 910
rect 35050 1050 35130 1080
rect 35050 1010 35070 1050
rect 35110 1010 35130 1050
rect 35050 950 35130 1010
rect 35050 910 35070 950
rect 35110 910 35130 950
rect 35050 880 35130 910
rect 35160 1050 35240 1080
rect 35160 1010 35180 1050
rect 35220 1010 35240 1050
rect 35160 950 35240 1010
rect 35160 910 35180 950
rect 35220 910 35240 950
rect 35160 880 35240 910
rect 35270 1050 35350 1080
rect 35270 1010 35290 1050
rect 35330 1010 35350 1050
rect 35270 950 35350 1010
rect 35270 910 35290 950
rect 35330 910 35350 950
rect 35270 880 35350 910
rect 35850 1050 35930 1080
rect 35850 1010 35870 1050
rect 35910 1010 35930 1050
rect 35850 950 35930 1010
rect 35850 910 35870 950
rect 35910 910 35930 950
rect 35850 880 35930 910
rect 35960 1050 36040 1080
rect 35960 1010 35980 1050
rect 36020 1010 36040 1050
rect 35960 950 36040 1010
rect 35960 910 35980 950
rect 36020 910 36040 950
rect 35960 880 36040 910
rect 36070 1050 36150 1080
rect 36070 1010 36090 1050
rect 36130 1010 36150 1050
rect 36070 950 36150 1010
rect 36070 910 36090 950
rect 36130 910 36150 950
rect 36070 880 36150 910
rect 36180 1050 36260 1080
rect 36180 1010 36200 1050
rect 36240 1010 36260 1050
rect 36180 950 36260 1010
rect 36180 910 36200 950
rect 36240 910 36260 950
rect 36180 880 36260 910
rect 36290 1050 36370 1080
rect 36290 1010 36310 1050
rect 36350 1010 36370 1050
rect 36290 950 36370 1010
rect 36290 910 36310 950
rect 36350 910 36370 950
rect 36290 880 36370 910
rect 36400 1050 36480 1080
rect 36400 1010 36420 1050
rect 36460 1010 36480 1050
rect 36400 950 36480 1010
rect 36400 910 36420 950
rect 36460 910 36480 950
rect 36400 880 36480 910
rect 36510 1050 36590 1080
rect 36510 1010 36530 1050
rect 36570 1010 36590 1050
rect 36510 950 36590 1010
rect 36510 910 36530 950
rect 36570 910 36590 950
rect 36510 880 36590 910
rect 36620 1050 36700 1080
rect 36620 1010 36640 1050
rect 36680 1010 36700 1050
rect 36620 950 36700 1010
rect 36620 910 36640 950
rect 36680 910 36700 950
rect 36620 880 36700 910
rect 36730 1050 36810 1080
rect 36730 1010 36750 1050
rect 36790 1010 36810 1050
rect 36730 950 36810 1010
rect 36730 910 36750 950
rect 36790 910 36810 950
rect 36730 880 36810 910
rect 36840 1050 36920 1080
rect 36840 1010 36860 1050
rect 36900 1010 36920 1050
rect 36840 950 36920 1010
rect 36840 910 36860 950
rect 36900 910 36920 950
rect 36840 880 36920 910
rect 36950 1050 37030 1080
rect 36950 1010 36970 1050
rect 37010 1010 37030 1050
rect 36950 950 37030 1010
rect 36950 910 36970 950
rect 37010 910 37030 950
rect 36950 880 37030 910
rect 37060 1050 37140 1080
rect 37060 1010 37080 1050
rect 37120 1010 37140 1050
rect 37060 950 37140 1010
rect 37060 910 37080 950
rect 37120 910 37140 950
rect 37060 880 37140 910
rect 37170 1050 37250 1080
rect 37170 1010 37190 1050
rect 37230 1010 37250 1050
rect 37170 950 37250 1010
rect 37170 910 37190 950
rect 37230 910 37250 950
rect 37170 880 37250 910
rect 33940 450 34020 480
rect 33940 410 33960 450
rect 34000 410 34020 450
rect 33940 350 34020 410
rect 33940 310 33960 350
rect 34000 310 34020 350
rect 32870 250 32950 280
rect 32870 210 32890 250
rect 32930 210 32950 250
rect 32870 150 32950 210
rect 32870 110 32890 150
rect 32930 110 32950 150
rect 32870 80 32950 110
rect 32980 250 33060 280
rect 32980 210 33000 250
rect 33040 210 33060 250
rect 32980 150 33060 210
rect 32980 110 33000 150
rect 33040 110 33060 150
rect 32980 80 33060 110
rect 33090 250 33170 280
rect 33090 210 33110 250
rect 33150 210 33170 250
rect 33090 150 33170 210
rect 33090 110 33110 150
rect 33150 110 33170 150
rect 33090 80 33170 110
rect 33200 250 33280 280
rect 33200 210 33220 250
rect 33260 210 33280 250
rect 33200 150 33280 210
rect 33200 110 33220 150
rect 33260 110 33280 150
rect 33200 80 33280 110
rect 33310 250 33400 280
rect 33310 210 33330 250
rect 33370 210 33400 250
rect 33310 150 33400 210
rect 33310 110 33330 150
rect 33370 110 33400 150
rect 33310 80 33400 110
rect 33940 250 34020 310
rect 33940 210 33960 250
rect 34000 210 34020 250
rect 33940 150 34020 210
rect 33940 110 33960 150
rect 34000 110 34020 150
rect 33940 50 34020 110
rect 33940 10 33960 50
rect 34000 10 34020 50
rect 33940 -50 34020 10
rect 33940 -90 33960 -50
rect 34000 -90 34020 -50
rect 33940 -120 34020 -90
rect 34120 450 34200 480
rect 34120 410 34140 450
rect 34180 410 34200 450
rect 34120 350 34200 410
rect 34120 310 34140 350
rect 34180 310 34200 350
rect 34120 250 34200 310
rect 34120 210 34140 250
rect 34180 210 34200 250
rect 34120 150 34200 210
rect 34120 110 34140 150
rect 34180 110 34200 150
rect 34120 50 34200 110
rect 34120 10 34140 50
rect 34180 10 34200 50
rect 34120 -50 34200 10
rect 34120 -90 34140 -50
rect 34180 -90 34200 -50
rect 34120 -120 34200 -90
rect 34300 450 34380 480
rect 34300 410 34320 450
rect 34360 410 34380 450
rect 34300 350 34380 410
rect 34300 310 34320 350
rect 34360 310 34380 350
rect 34300 250 34380 310
rect 34300 210 34320 250
rect 34360 210 34380 250
rect 34300 150 34380 210
rect 34300 110 34320 150
rect 34360 110 34380 150
rect 34300 50 34380 110
rect 34300 10 34320 50
rect 34360 10 34380 50
rect 34300 -50 34380 10
rect 34300 -90 34320 -50
rect 34360 -90 34380 -50
rect 34300 -120 34380 -90
rect 34480 450 34560 480
rect 34480 410 34500 450
rect 34540 410 34560 450
rect 34480 350 34560 410
rect 34480 310 34500 350
rect 34540 310 34560 350
rect 34480 250 34560 310
rect 34480 210 34500 250
rect 34540 210 34560 250
rect 34480 150 34560 210
rect 34480 110 34500 150
rect 34540 110 34560 150
rect 34480 50 34560 110
rect 34480 10 34500 50
rect 34540 10 34560 50
rect 34480 -50 34560 10
rect 34480 -90 34500 -50
rect 34540 -90 34560 -50
rect 34480 -120 34560 -90
rect 34660 450 34740 480
rect 34660 410 34680 450
rect 34720 410 34740 450
rect 34660 350 34740 410
rect 34660 310 34680 350
rect 34720 310 34740 350
rect 34660 250 34740 310
rect 34660 210 34680 250
rect 34720 210 34740 250
rect 34660 150 34740 210
rect 34660 110 34680 150
rect 34720 110 34740 150
rect 34660 50 34740 110
rect 34660 10 34680 50
rect 34720 10 34740 50
rect 34660 -50 34740 10
rect 34660 -90 34680 -50
rect 34720 -90 34740 -50
rect 34660 -120 34740 -90
rect 34840 450 34920 480
rect 34840 410 34860 450
rect 34900 410 34920 450
rect 34840 350 34920 410
rect 34840 310 34860 350
rect 34900 310 34920 350
rect 34840 250 34920 310
rect 34840 210 34860 250
rect 34900 210 34920 250
rect 34840 150 34920 210
rect 34840 110 34860 150
rect 34900 110 34920 150
rect 34840 50 34920 110
rect 34840 10 34860 50
rect 34900 10 34920 50
rect 34840 -50 34920 10
rect 34840 -90 34860 -50
rect 34900 -90 34920 -50
rect 34840 -120 34920 -90
rect 35020 450 35100 480
rect 35020 410 35040 450
rect 35080 410 35100 450
rect 35020 350 35100 410
rect 35020 310 35040 350
rect 35080 310 35100 350
rect 35020 250 35100 310
rect 35020 210 35040 250
rect 35080 210 35100 250
rect 35020 150 35100 210
rect 35020 110 35040 150
rect 35080 110 35100 150
rect 35020 50 35100 110
rect 35020 10 35040 50
rect 35080 10 35100 50
rect 35020 -50 35100 10
rect 35020 -90 35040 -50
rect 35080 -90 35100 -50
rect 35020 -120 35100 -90
rect 35200 450 35280 480
rect 35200 410 35220 450
rect 35260 410 35280 450
rect 35200 350 35280 410
rect 35200 310 35220 350
rect 35260 310 35280 350
rect 35200 250 35280 310
rect 35200 210 35220 250
rect 35260 210 35280 250
rect 35200 150 35280 210
rect 35200 110 35220 150
rect 35260 110 35280 150
rect 35200 50 35280 110
rect 35200 10 35220 50
rect 35260 10 35280 50
rect 35200 -50 35280 10
rect 35200 -90 35220 -50
rect 35260 -90 35280 -50
rect 35200 -120 35280 -90
rect 35380 450 35460 480
rect 35380 410 35400 450
rect 35440 410 35460 450
rect 35380 350 35460 410
rect 35380 310 35400 350
rect 35440 310 35460 350
rect 35380 250 35460 310
rect 35380 210 35400 250
rect 35440 210 35460 250
rect 35380 150 35460 210
rect 35380 110 35400 150
rect 35440 110 35460 150
rect 35380 50 35460 110
rect 35380 10 35400 50
rect 35440 10 35460 50
rect 35380 -50 35460 10
rect 35380 -90 35400 -50
rect 35440 -90 35460 -50
rect 35380 -120 35460 -90
rect 35560 450 35640 480
rect 35560 410 35580 450
rect 35620 410 35640 450
rect 35560 350 35640 410
rect 35560 310 35580 350
rect 35620 310 35640 350
rect 35560 250 35640 310
rect 35560 210 35580 250
rect 35620 210 35640 250
rect 35560 150 35640 210
rect 35560 110 35580 150
rect 35620 110 35640 150
rect 35560 50 35640 110
rect 35560 10 35580 50
rect 35620 10 35640 50
rect 35560 -50 35640 10
rect 35560 -90 35580 -50
rect 35620 -90 35640 -50
rect 35560 -120 35640 -90
rect 35740 450 35820 480
rect 35740 410 35760 450
rect 35800 410 35820 450
rect 35740 350 35820 410
rect 35740 310 35760 350
rect 35800 310 35820 350
rect 35740 250 35820 310
rect 35740 210 35760 250
rect 35800 210 35820 250
rect 35740 150 35820 210
rect 35740 110 35760 150
rect 35800 110 35820 150
rect 35740 50 35820 110
rect 35740 10 35760 50
rect 35800 10 35820 50
rect 35740 -50 35820 10
rect 35740 -90 35760 -50
rect 35800 -90 35820 -50
rect 35740 -120 35820 -90
rect 35920 450 36000 480
rect 35920 410 35940 450
rect 35980 410 36000 450
rect 35920 350 36000 410
rect 35920 310 35940 350
rect 35980 310 36000 350
rect 35920 250 36000 310
rect 35920 210 35940 250
rect 35980 210 36000 250
rect 35920 150 36000 210
rect 35920 110 35940 150
rect 35980 110 36000 150
rect 35920 50 36000 110
rect 35920 10 35940 50
rect 35980 10 36000 50
rect 35920 -50 36000 10
rect 35920 -90 35940 -50
rect 35980 -90 36000 -50
rect 35920 -120 36000 -90
rect 36100 450 36180 480
rect 36100 410 36120 450
rect 36160 410 36180 450
rect 36100 350 36180 410
rect 36100 310 36120 350
rect 36160 310 36180 350
rect 36100 250 36180 310
rect 36100 210 36120 250
rect 36160 210 36180 250
rect 36100 150 36180 210
rect 36100 110 36120 150
rect 36160 110 36180 150
rect 36100 50 36180 110
rect 36100 10 36120 50
rect 36160 10 36180 50
rect 36100 -50 36180 10
rect 36100 -90 36120 -50
rect 36160 -90 36180 -50
rect 36100 -120 36180 -90
rect 36280 450 36360 480
rect 36280 410 36300 450
rect 36340 410 36360 450
rect 36280 350 36360 410
rect 36280 310 36300 350
rect 36340 310 36360 350
rect 36280 250 36360 310
rect 36280 210 36300 250
rect 36340 210 36360 250
rect 36280 150 36360 210
rect 36280 110 36300 150
rect 36340 110 36360 150
rect 36280 50 36360 110
rect 36280 10 36300 50
rect 36340 10 36360 50
rect 36280 -50 36360 10
rect 36280 -90 36300 -50
rect 36340 -90 36360 -50
rect 36280 -120 36360 -90
rect 36460 450 36540 480
rect 36460 410 36480 450
rect 36520 410 36540 450
rect 36460 350 36540 410
rect 36460 310 36480 350
rect 36520 310 36540 350
rect 36460 250 36540 310
rect 36460 210 36480 250
rect 36520 210 36540 250
rect 36460 150 36540 210
rect 36460 110 36480 150
rect 36520 110 36540 150
rect 36460 50 36540 110
rect 36460 10 36480 50
rect 36520 10 36540 50
rect 36460 -50 36540 10
rect 36460 -90 36480 -50
rect 36520 -90 36540 -50
rect 36460 -120 36540 -90
rect 36640 450 36720 480
rect 36640 410 36660 450
rect 36700 410 36720 450
rect 36640 350 36720 410
rect 36640 310 36660 350
rect 36700 310 36720 350
rect 36640 250 36720 310
rect 36640 210 36660 250
rect 36700 210 36720 250
rect 36640 150 36720 210
rect 36640 110 36660 150
rect 36700 110 36720 150
rect 36640 50 36720 110
rect 36640 10 36660 50
rect 36700 10 36720 50
rect 36640 -50 36720 10
rect 36640 -90 36660 -50
rect 36700 -90 36720 -50
rect 36640 -120 36720 -90
rect 36820 450 36900 480
rect 36820 410 36840 450
rect 36880 410 36900 450
rect 36820 350 36900 410
rect 36820 310 36840 350
rect 36880 310 36900 350
rect 36820 250 36900 310
rect 36820 210 36840 250
rect 36880 210 36900 250
rect 36820 150 36900 210
rect 36820 110 36840 150
rect 36880 110 36900 150
rect 36820 50 36900 110
rect 36820 10 36840 50
rect 36880 10 36900 50
rect 36820 -50 36900 10
rect 36820 -90 36840 -50
rect 36880 -90 36900 -50
rect 36820 -120 36900 -90
rect 37000 450 37080 480
rect 37000 410 37020 450
rect 37060 410 37080 450
rect 37000 350 37080 410
rect 37000 310 37020 350
rect 37060 310 37080 350
rect 37000 250 37080 310
rect 37000 210 37020 250
rect 37060 210 37080 250
rect 37000 150 37080 210
rect 37000 110 37020 150
rect 37060 110 37080 150
rect 37000 50 37080 110
rect 37000 10 37020 50
rect 37060 10 37080 50
rect 37000 -50 37080 10
rect 37000 -90 37020 -50
rect 37060 -90 37080 -50
rect 37000 -120 37080 -90
rect 37180 450 37260 480
rect 37180 410 37200 450
rect 37240 410 37260 450
rect 37180 350 37260 410
rect 37180 310 37200 350
rect 37240 310 37260 350
rect 37180 250 37260 310
rect 37180 210 37200 250
rect 37240 210 37260 250
rect 37180 150 37260 210
rect 37180 110 37200 150
rect 37240 110 37260 150
rect 37180 50 37260 110
rect 37180 10 37200 50
rect 37240 10 37260 50
rect 37180 -50 37260 10
rect 37180 -90 37200 -50
rect 37240 -90 37260 -50
rect 37180 -120 37260 -90
rect 32840 -1110 32920 -1080
rect 32840 -1150 32860 -1110
rect 32900 -1150 32920 -1110
rect 32840 -1210 32920 -1150
rect 32840 -1250 32860 -1210
rect 32900 -1250 32920 -1210
rect 32840 -1280 32920 -1250
rect 32960 -1110 33040 -1080
rect 32960 -1150 32980 -1110
rect 33020 -1150 33040 -1110
rect 32960 -1210 33040 -1150
rect 32960 -1250 32980 -1210
rect 33020 -1250 33040 -1210
rect 32960 -1280 33040 -1250
rect 33080 -1110 33160 -1080
rect 33080 -1150 33100 -1110
rect 33140 -1150 33160 -1110
rect 33080 -1210 33160 -1150
rect 33080 -1250 33100 -1210
rect 33140 -1250 33160 -1210
rect 33080 -1280 33160 -1250
rect 33200 -1110 33280 -1080
rect 33200 -1150 33220 -1110
rect 33260 -1150 33280 -1110
rect 33200 -1210 33280 -1150
rect 33200 -1250 33220 -1210
rect 33260 -1250 33280 -1210
rect 33200 -1280 33280 -1250
rect 33320 -1110 33400 -1080
rect 33320 -1150 33340 -1110
rect 33380 -1150 33400 -1110
rect 33320 -1210 33400 -1150
rect 33320 -1250 33340 -1210
rect 33380 -1250 33400 -1210
rect 33320 -1280 33400 -1250
rect 33440 -1110 33520 -1080
rect 33440 -1150 33460 -1110
rect 33500 -1150 33520 -1110
rect 33440 -1210 33520 -1150
rect 33440 -1250 33460 -1210
rect 33500 -1250 33520 -1210
rect 33440 -1280 33520 -1250
rect 33560 -1110 33640 -1080
rect 33560 -1150 33580 -1110
rect 33620 -1150 33640 -1110
rect 33560 -1210 33640 -1150
rect 33560 -1250 33580 -1210
rect 33620 -1250 33640 -1210
rect 33560 -1280 33640 -1250
rect 33680 -1110 33760 -1080
rect 33680 -1150 33700 -1110
rect 33740 -1150 33760 -1110
rect 33680 -1210 33760 -1150
rect 33680 -1250 33700 -1210
rect 33740 -1250 33760 -1210
rect 33680 -1280 33760 -1250
rect 33800 -1110 33880 -1080
rect 33800 -1150 33820 -1110
rect 33860 -1150 33880 -1110
rect 33800 -1210 33880 -1150
rect 33800 -1250 33820 -1210
rect 33860 -1250 33880 -1210
rect 33800 -1280 33880 -1250
rect 33920 -1110 34000 -1080
rect 33920 -1150 33940 -1110
rect 33980 -1150 34000 -1110
rect 33920 -1210 34000 -1150
rect 33920 -1250 33940 -1210
rect 33980 -1250 34000 -1210
rect 33920 -1280 34000 -1250
rect 34040 -1110 34120 -1080
rect 34040 -1150 34060 -1110
rect 34100 -1150 34120 -1110
rect 34040 -1210 34120 -1150
rect 34040 -1250 34060 -1210
rect 34100 -1250 34120 -1210
rect 34040 -1280 34120 -1250
rect 34160 -1110 34240 -1080
rect 34160 -1150 34180 -1110
rect 34220 -1150 34240 -1110
rect 34160 -1210 34240 -1150
rect 34160 -1250 34180 -1210
rect 34220 -1250 34240 -1210
rect 34160 -1280 34240 -1250
rect 34280 -1110 34360 -1080
rect 34280 -1150 34300 -1110
rect 34340 -1150 34360 -1110
rect 34280 -1210 34360 -1150
rect 34280 -1250 34300 -1210
rect 34340 -1250 34360 -1210
rect 34280 -1280 34360 -1250
rect 34400 -1110 34480 -1080
rect 34400 -1150 34420 -1110
rect 34460 -1150 34480 -1110
rect 34400 -1210 34480 -1150
rect 34400 -1250 34420 -1210
rect 34460 -1250 34480 -1210
rect 34400 -1280 34480 -1250
rect 34520 -1110 34600 -1080
rect 34520 -1150 34540 -1110
rect 34580 -1150 34600 -1110
rect 34520 -1210 34600 -1150
rect 34520 -1250 34540 -1210
rect 34580 -1250 34600 -1210
rect 34520 -1280 34600 -1250
rect 34640 -1110 34720 -1080
rect 34640 -1150 34660 -1110
rect 34700 -1150 34720 -1110
rect 34640 -1210 34720 -1150
rect 34640 -1250 34660 -1210
rect 34700 -1250 34720 -1210
rect 34640 -1280 34720 -1250
rect 34760 -1110 34840 -1080
rect 34760 -1150 34780 -1110
rect 34820 -1150 34840 -1110
rect 34760 -1210 34840 -1150
rect 34760 -1250 34780 -1210
rect 34820 -1250 34840 -1210
rect 34760 -1280 34840 -1250
rect 34880 -1110 34960 -1080
rect 34880 -1150 34900 -1110
rect 34940 -1150 34960 -1110
rect 34880 -1210 34960 -1150
rect 34880 -1250 34900 -1210
rect 34940 -1250 34960 -1210
rect 34880 -1280 34960 -1250
rect 35000 -1110 35080 -1080
rect 35000 -1150 35020 -1110
rect 35060 -1150 35080 -1110
rect 35000 -1210 35080 -1150
rect 35000 -1250 35020 -1210
rect 35060 -1250 35080 -1210
rect 35000 -1280 35080 -1250
rect 35120 -1110 35200 -1080
rect 35120 -1150 35140 -1110
rect 35180 -1150 35200 -1110
rect 35120 -1210 35200 -1150
rect 35120 -1250 35140 -1210
rect 35180 -1250 35200 -1210
rect 35120 -1280 35200 -1250
rect 35240 -1110 35320 -1080
rect 35240 -1150 35260 -1110
rect 35300 -1150 35320 -1110
rect 35240 -1210 35320 -1150
rect 35240 -1250 35260 -1210
rect 35300 -1250 35320 -1210
rect 35240 -1280 35320 -1250
rect 35880 -1110 35960 -1080
rect 35880 -1150 35900 -1110
rect 35940 -1150 35960 -1110
rect 35880 -1210 35960 -1150
rect 35880 -1250 35900 -1210
rect 35940 -1250 35960 -1210
rect 35880 -1280 35960 -1250
rect 36000 -1110 36080 -1080
rect 36000 -1150 36020 -1110
rect 36060 -1150 36080 -1110
rect 36000 -1210 36080 -1150
rect 36000 -1250 36020 -1210
rect 36060 -1250 36080 -1210
rect 36000 -1280 36080 -1250
rect 36120 -1110 36200 -1080
rect 36120 -1150 36140 -1110
rect 36180 -1150 36200 -1110
rect 36120 -1210 36200 -1150
rect 36120 -1250 36140 -1210
rect 36180 -1250 36200 -1210
rect 36120 -1280 36200 -1250
rect 36240 -1110 36320 -1080
rect 36240 -1150 36260 -1110
rect 36300 -1150 36320 -1110
rect 36240 -1210 36320 -1150
rect 36240 -1250 36260 -1210
rect 36300 -1250 36320 -1210
rect 36240 -1280 36320 -1250
rect 36360 -1110 36440 -1080
rect 36360 -1150 36380 -1110
rect 36420 -1150 36440 -1110
rect 36360 -1210 36440 -1150
rect 36360 -1250 36380 -1210
rect 36420 -1250 36440 -1210
rect 36360 -1280 36440 -1250
rect 36480 -1110 36560 -1080
rect 36480 -1150 36500 -1110
rect 36540 -1150 36560 -1110
rect 36480 -1210 36560 -1150
rect 36480 -1250 36500 -1210
rect 36540 -1250 36560 -1210
rect 36480 -1280 36560 -1250
rect 36600 -1110 36680 -1080
rect 36600 -1150 36620 -1110
rect 36660 -1150 36680 -1110
rect 36600 -1210 36680 -1150
rect 36600 -1250 36620 -1210
rect 36660 -1250 36680 -1210
rect 36600 -1280 36680 -1250
rect 36720 -1110 36800 -1080
rect 36720 -1150 36740 -1110
rect 36780 -1150 36800 -1110
rect 36720 -1210 36800 -1150
rect 36720 -1250 36740 -1210
rect 36780 -1250 36800 -1210
rect 36720 -1280 36800 -1250
rect 36840 -1110 36920 -1080
rect 36840 -1150 36860 -1110
rect 36900 -1150 36920 -1110
rect 36840 -1210 36920 -1150
rect 36840 -1250 36860 -1210
rect 36900 -1250 36920 -1210
rect 36840 -1280 36920 -1250
rect 36960 -1110 37040 -1080
rect 36960 -1150 36980 -1110
rect 37020 -1150 37040 -1110
rect 36960 -1210 37040 -1150
rect 36960 -1250 36980 -1210
rect 37020 -1250 37040 -1210
rect 36960 -1280 37040 -1250
rect 37080 -1110 37160 -1080
rect 37080 -1150 37100 -1110
rect 37140 -1150 37160 -1110
rect 37080 -1210 37160 -1150
rect 37080 -1250 37100 -1210
rect 37140 -1250 37160 -1210
rect 37080 -1280 37160 -1250
rect 37200 -1110 37280 -1080
rect 37200 -1150 37220 -1110
rect 37260 -1150 37280 -1110
rect 37200 -1210 37280 -1150
rect 37200 -1250 37220 -1210
rect 37260 -1250 37280 -1210
rect 37200 -1280 37280 -1250
rect 37320 -1110 37400 -1080
rect 37320 -1150 37340 -1110
rect 37380 -1150 37400 -1110
rect 37320 -1210 37400 -1150
rect 37320 -1250 37340 -1210
rect 37380 -1250 37400 -1210
rect 37320 -1280 37400 -1250
rect 37440 -1110 37520 -1080
rect 37440 -1150 37460 -1110
rect 37500 -1150 37520 -1110
rect 37440 -1210 37520 -1150
rect 37440 -1250 37460 -1210
rect 37500 -1250 37520 -1210
rect 37440 -1280 37520 -1250
rect 37560 -1110 37640 -1080
rect 37560 -1150 37580 -1110
rect 37620 -1150 37640 -1110
rect 37560 -1210 37640 -1150
rect 37560 -1250 37580 -1210
rect 37620 -1250 37640 -1210
rect 37560 -1280 37640 -1250
rect 37680 -1110 37760 -1080
rect 37680 -1150 37700 -1110
rect 37740 -1150 37760 -1110
rect 37680 -1210 37760 -1150
rect 37680 -1250 37700 -1210
rect 37740 -1250 37760 -1210
rect 37680 -1280 37760 -1250
rect 37800 -1110 37880 -1080
rect 37800 -1150 37820 -1110
rect 37860 -1150 37880 -1110
rect 37800 -1210 37880 -1150
rect 37800 -1250 37820 -1210
rect 37860 -1250 37880 -1210
rect 37800 -1280 37880 -1250
rect 37920 -1110 38000 -1080
rect 37920 -1150 37940 -1110
rect 37980 -1150 38000 -1110
rect 37920 -1210 38000 -1150
rect 37920 -1250 37940 -1210
rect 37980 -1250 38000 -1210
rect 37920 -1280 38000 -1250
rect 38040 -1110 38120 -1080
rect 38040 -1150 38060 -1110
rect 38100 -1150 38120 -1110
rect 38040 -1210 38120 -1150
rect 38040 -1250 38060 -1210
rect 38100 -1250 38120 -1210
rect 38040 -1280 38120 -1250
rect 38160 -1110 38240 -1080
rect 38160 -1150 38180 -1110
rect 38220 -1150 38240 -1110
rect 38160 -1210 38240 -1150
rect 38160 -1250 38180 -1210
rect 38220 -1250 38240 -1210
rect 38160 -1280 38240 -1250
rect 38280 -1110 38360 -1080
rect 38280 -1150 38300 -1110
rect 38340 -1150 38360 -1110
rect 38280 -1210 38360 -1150
rect 38280 -1250 38300 -1210
rect 38340 -1250 38360 -1210
rect 38280 -1280 38360 -1250
<< ndiffc >>
rect 33700 -2090 33740 -2050
rect 33820 -2090 33860 -2050
rect 33940 -2090 33980 -2050
rect 34060 -2090 34100 -2050
rect 34180 -2090 34220 -2050
rect 34300 -2090 34340 -2050
rect 34420 -2090 34460 -2050
rect 34540 -2090 34580 -2050
rect 34660 -2090 34700 -2050
rect 34780 -2090 34820 -2050
rect 34900 -2090 34940 -2050
rect 36260 -2090 36300 -2050
rect 36380 -2090 36420 -2050
rect 36500 -2090 36540 -2050
rect 36620 -2090 36660 -2050
rect 36740 -2090 36780 -2050
rect 36860 -2090 36900 -2050
rect 36980 -2090 37020 -2050
rect 37100 -2090 37140 -2050
rect 37220 -2090 37260 -2050
rect 37340 -2090 37380 -2050
rect 37460 -2090 37500 -2050
rect 33080 -2700 33120 -2660
rect 33080 -2800 33120 -2760
rect 33080 -2900 33120 -2860
rect 33080 -3000 33120 -2960
rect 33080 -3100 33120 -3060
rect 34160 -2700 34200 -2660
rect 34320 -2700 34360 -2660
rect 34160 -2800 34200 -2760
rect 34320 -2800 34360 -2760
rect 34160 -2900 34200 -2860
rect 34320 -2900 34360 -2860
rect 34160 -3000 34200 -2960
rect 34320 -3000 34360 -2960
rect 34160 -3100 34200 -3060
rect 34320 -3100 34360 -3060
rect 35400 -2700 35440 -2660
rect 35400 -2800 35440 -2760
rect 35400 -2900 35440 -2860
rect 35400 -3000 35440 -2960
rect 35400 -3100 35440 -3060
rect 35760 -2700 35800 -2660
rect 35760 -2800 35800 -2760
rect 35760 -2900 35800 -2860
rect 35760 -3000 35800 -2960
rect 35760 -3100 35800 -3060
rect 36840 -2700 36880 -2660
rect 37000 -2700 37040 -2660
rect 36840 -2800 36880 -2760
rect 37000 -2800 37040 -2760
rect 36840 -2900 36880 -2860
rect 37000 -2900 37040 -2860
rect 36840 -3000 36880 -2960
rect 37000 -3000 37040 -2960
rect 36840 -3100 36880 -3060
rect 37000 -3100 37040 -3060
rect 38080 -2700 38120 -2660
rect 38080 -2800 38120 -2760
rect 38080 -2900 38120 -2860
rect 38080 -3000 38120 -2960
rect 38080 -3100 38120 -3060
rect 33500 -3610 33540 -3570
rect 33500 -3710 33540 -3670
rect 35580 -3610 35620 -3570
rect 35580 -3710 35620 -3670
rect 37660 -3610 37700 -3570
rect 37660 -3710 37700 -3670
<< pdiffc >>
rect 33970 1010 34010 1050
rect 33970 910 34010 950
rect 34080 1010 34120 1050
rect 34080 910 34120 950
rect 34190 1010 34230 1050
rect 34190 910 34230 950
rect 34300 1010 34340 1050
rect 34300 910 34340 950
rect 34410 1010 34450 1050
rect 34410 910 34450 950
rect 34520 1010 34560 1050
rect 34520 910 34560 950
rect 34630 1010 34670 1050
rect 34630 910 34670 950
rect 34740 1010 34780 1050
rect 34740 910 34780 950
rect 34850 1010 34890 1050
rect 34850 910 34890 950
rect 34960 1010 35000 1050
rect 34960 910 35000 950
rect 35070 1010 35110 1050
rect 35070 910 35110 950
rect 35180 1010 35220 1050
rect 35180 910 35220 950
rect 35290 1010 35330 1050
rect 35290 910 35330 950
rect 35870 1010 35910 1050
rect 35870 910 35910 950
rect 35980 1010 36020 1050
rect 35980 910 36020 950
rect 36090 1010 36130 1050
rect 36090 910 36130 950
rect 36200 1010 36240 1050
rect 36200 910 36240 950
rect 36310 1010 36350 1050
rect 36310 910 36350 950
rect 36420 1010 36460 1050
rect 36420 910 36460 950
rect 36530 1010 36570 1050
rect 36530 910 36570 950
rect 36640 1010 36680 1050
rect 36640 910 36680 950
rect 36750 1010 36790 1050
rect 36750 910 36790 950
rect 36860 1010 36900 1050
rect 36860 910 36900 950
rect 36970 1010 37010 1050
rect 36970 910 37010 950
rect 37080 1010 37120 1050
rect 37080 910 37120 950
rect 37190 1010 37230 1050
rect 37190 910 37230 950
rect 33960 410 34000 450
rect 33960 310 34000 350
rect 32890 210 32930 250
rect 32890 110 32930 150
rect 33000 210 33040 250
rect 33000 110 33040 150
rect 33110 210 33150 250
rect 33110 110 33150 150
rect 33220 210 33260 250
rect 33220 110 33260 150
rect 33330 210 33370 250
rect 33330 110 33370 150
rect 33960 210 34000 250
rect 33960 110 34000 150
rect 33960 10 34000 50
rect 33960 -90 34000 -50
rect 34140 410 34180 450
rect 34140 310 34180 350
rect 34140 210 34180 250
rect 34140 110 34180 150
rect 34140 10 34180 50
rect 34140 -90 34180 -50
rect 34320 410 34360 450
rect 34320 310 34360 350
rect 34320 210 34360 250
rect 34320 110 34360 150
rect 34320 10 34360 50
rect 34320 -90 34360 -50
rect 34500 410 34540 450
rect 34500 310 34540 350
rect 34500 210 34540 250
rect 34500 110 34540 150
rect 34500 10 34540 50
rect 34500 -90 34540 -50
rect 34680 410 34720 450
rect 34680 310 34720 350
rect 34680 210 34720 250
rect 34680 110 34720 150
rect 34680 10 34720 50
rect 34680 -90 34720 -50
rect 34860 410 34900 450
rect 34860 310 34900 350
rect 34860 210 34900 250
rect 34860 110 34900 150
rect 34860 10 34900 50
rect 34860 -90 34900 -50
rect 35040 410 35080 450
rect 35040 310 35080 350
rect 35040 210 35080 250
rect 35040 110 35080 150
rect 35040 10 35080 50
rect 35040 -90 35080 -50
rect 35220 410 35260 450
rect 35220 310 35260 350
rect 35220 210 35260 250
rect 35220 110 35260 150
rect 35220 10 35260 50
rect 35220 -90 35260 -50
rect 35400 410 35440 450
rect 35400 310 35440 350
rect 35400 210 35440 250
rect 35400 110 35440 150
rect 35400 10 35440 50
rect 35400 -90 35440 -50
rect 35580 410 35620 450
rect 35580 310 35620 350
rect 35580 210 35620 250
rect 35580 110 35620 150
rect 35580 10 35620 50
rect 35580 -90 35620 -50
rect 35760 410 35800 450
rect 35760 310 35800 350
rect 35760 210 35800 250
rect 35760 110 35800 150
rect 35760 10 35800 50
rect 35760 -90 35800 -50
rect 35940 410 35980 450
rect 35940 310 35980 350
rect 35940 210 35980 250
rect 35940 110 35980 150
rect 35940 10 35980 50
rect 35940 -90 35980 -50
rect 36120 410 36160 450
rect 36120 310 36160 350
rect 36120 210 36160 250
rect 36120 110 36160 150
rect 36120 10 36160 50
rect 36120 -90 36160 -50
rect 36300 410 36340 450
rect 36300 310 36340 350
rect 36300 210 36340 250
rect 36300 110 36340 150
rect 36300 10 36340 50
rect 36300 -90 36340 -50
rect 36480 410 36520 450
rect 36480 310 36520 350
rect 36480 210 36520 250
rect 36480 110 36520 150
rect 36480 10 36520 50
rect 36480 -90 36520 -50
rect 36660 410 36700 450
rect 36660 310 36700 350
rect 36660 210 36700 250
rect 36660 110 36700 150
rect 36660 10 36700 50
rect 36660 -90 36700 -50
rect 36840 410 36880 450
rect 36840 310 36880 350
rect 36840 210 36880 250
rect 36840 110 36880 150
rect 36840 10 36880 50
rect 36840 -90 36880 -50
rect 37020 410 37060 450
rect 37020 310 37060 350
rect 37020 210 37060 250
rect 37020 110 37060 150
rect 37020 10 37060 50
rect 37020 -90 37060 -50
rect 37200 410 37240 450
rect 37200 310 37240 350
rect 37200 210 37240 250
rect 37200 110 37240 150
rect 37200 10 37240 50
rect 37200 -90 37240 -50
rect 32860 -1150 32900 -1110
rect 32860 -1250 32900 -1210
rect 32980 -1150 33020 -1110
rect 32980 -1250 33020 -1210
rect 33100 -1150 33140 -1110
rect 33100 -1250 33140 -1210
rect 33220 -1150 33260 -1110
rect 33220 -1250 33260 -1210
rect 33340 -1150 33380 -1110
rect 33340 -1250 33380 -1210
rect 33460 -1150 33500 -1110
rect 33460 -1250 33500 -1210
rect 33580 -1150 33620 -1110
rect 33580 -1250 33620 -1210
rect 33700 -1150 33740 -1110
rect 33700 -1250 33740 -1210
rect 33820 -1150 33860 -1110
rect 33820 -1250 33860 -1210
rect 33940 -1150 33980 -1110
rect 33940 -1250 33980 -1210
rect 34060 -1150 34100 -1110
rect 34060 -1250 34100 -1210
rect 34180 -1150 34220 -1110
rect 34180 -1250 34220 -1210
rect 34300 -1150 34340 -1110
rect 34300 -1250 34340 -1210
rect 34420 -1150 34460 -1110
rect 34420 -1250 34460 -1210
rect 34540 -1150 34580 -1110
rect 34540 -1250 34580 -1210
rect 34660 -1150 34700 -1110
rect 34660 -1250 34700 -1210
rect 34780 -1150 34820 -1110
rect 34780 -1250 34820 -1210
rect 34900 -1150 34940 -1110
rect 34900 -1250 34940 -1210
rect 35020 -1150 35060 -1110
rect 35020 -1250 35060 -1210
rect 35140 -1150 35180 -1110
rect 35140 -1250 35180 -1210
rect 35260 -1150 35300 -1110
rect 35260 -1250 35300 -1210
rect 35900 -1150 35940 -1110
rect 35900 -1250 35940 -1210
rect 36020 -1150 36060 -1110
rect 36020 -1250 36060 -1210
rect 36140 -1150 36180 -1110
rect 36140 -1250 36180 -1210
rect 36260 -1150 36300 -1110
rect 36260 -1250 36300 -1210
rect 36380 -1150 36420 -1110
rect 36380 -1250 36420 -1210
rect 36500 -1150 36540 -1110
rect 36500 -1250 36540 -1210
rect 36620 -1150 36660 -1110
rect 36620 -1250 36660 -1210
rect 36740 -1150 36780 -1110
rect 36740 -1250 36780 -1210
rect 36860 -1150 36900 -1110
rect 36860 -1250 36900 -1210
rect 36980 -1150 37020 -1110
rect 36980 -1250 37020 -1210
rect 37100 -1150 37140 -1110
rect 37100 -1250 37140 -1210
rect 37220 -1150 37260 -1110
rect 37220 -1250 37260 -1210
rect 37340 -1150 37380 -1110
rect 37340 -1250 37380 -1210
rect 37460 -1150 37500 -1110
rect 37460 -1250 37500 -1210
rect 37580 -1150 37620 -1110
rect 37580 -1250 37620 -1210
rect 37700 -1150 37740 -1110
rect 37700 -1250 37740 -1210
rect 37820 -1150 37860 -1110
rect 37820 -1250 37860 -1210
rect 37940 -1150 37980 -1110
rect 37940 -1250 37980 -1210
rect 38060 -1150 38100 -1110
rect 38060 -1250 38100 -1210
rect 38180 -1150 38220 -1110
rect 38180 -1250 38220 -1210
rect 38300 -1150 38340 -1110
rect 38300 -1250 38340 -1210
<< psubdiff >>
rect 35120 -1980 35200 -1950
rect 35120 -2020 35140 -1980
rect 35180 -2020 35200 -1980
rect 35120 -2060 35200 -2020
rect 35120 -2100 35140 -2060
rect 35180 -2100 35200 -2060
rect 35120 -2140 35200 -2100
rect 35120 -2180 35140 -2140
rect 35180 -2180 35200 -2140
rect 35120 -2210 35200 -2180
rect 36000 -1980 36080 -1950
rect 36000 -2020 36020 -1980
rect 36060 -2020 36080 -1980
rect 36000 -2060 36080 -2020
rect 36000 -2100 36020 -2060
rect 36060 -2100 36080 -2060
rect 36000 -2140 36080 -2100
rect 36000 -2180 36020 -2140
rect 36060 -2180 36080 -2140
rect 36000 -2210 36080 -2180
rect 34220 -2660 34300 -2630
rect 34220 -2700 34240 -2660
rect 34280 -2700 34300 -2660
rect 34220 -2760 34300 -2700
rect 34220 -2800 34240 -2760
rect 34280 -2800 34300 -2760
rect 34220 -2860 34300 -2800
rect 34220 -2900 34240 -2860
rect 34280 -2900 34300 -2860
rect 34220 -2960 34300 -2900
rect 34220 -3000 34240 -2960
rect 34280 -3000 34300 -2960
rect 34220 -3060 34300 -3000
rect 34220 -3100 34240 -3060
rect 34280 -3100 34300 -3060
rect 34220 -3120 34300 -3100
rect 36900 -2660 36980 -2630
rect 36900 -2700 36920 -2660
rect 36960 -2700 36980 -2660
rect 36900 -2760 36980 -2700
rect 36900 -2800 36920 -2760
rect 36960 -2800 36980 -2760
rect 36900 -2860 36980 -2800
rect 36900 -2900 36920 -2860
rect 36960 -2900 36980 -2860
rect 36900 -2960 36980 -2900
rect 36900 -3000 36920 -2960
rect 36960 -3000 36980 -2960
rect 36900 -3060 36980 -3000
rect 36900 -3100 36920 -3060
rect 36960 -3100 36980 -3060
rect 36900 -3130 36980 -3100
rect 33400 -3570 33480 -3540
rect 33400 -3610 33420 -3570
rect 33460 -3610 33480 -3570
rect 33400 -3670 33480 -3610
rect 33400 -3710 33420 -3670
rect 33460 -3710 33480 -3670
rect 33400 -3740 33480 -3710
rect 35550 -8330 35650 -8300
rect 35550 -8370 35580 -8330
rect 35620 -8370 35650 -8330
rect 35550 -8410 35650 -8370
rect 35550 -8450 35580 -8410
rect 35620 -8450 35650 -8410
rect 35550 -8490 35650 -8450
rect 35550 -8530 35580 -8490
rect 35620 -8530 35650 -8490
rect 35550 -8560 35650 -8530
<< nsubdiff >>
rect 33870 1050 33950 1080
rect 33870 1010 33890 1050
rect 33930 1010 33950 1050
rect 33870 950 33950 1010
rect 33870 910 33890 950
rect 33930 910 33950 950
rect 33870 880 33950 910
rect 35350 1050 35430 1080
rect 35350 1010 35370 1050
rect 35410 1010 35430 1050
rect 35350 950 35430 1010
rect 35350 910 35370 950
rect 35410 910 35430 950
rect 35350 880 35430 910
rect 35770 1050 35850 1080
rect 35770 1010 35790 1050
rect 35830 1010 35850 1050
rect 35770 950 35850 1010
rect 35770 910 35790 950
rect 35830 910 35850 950
rect 35770 880 35850 910
rect 37250 1050 37330 1080
rect 37250 1010 37270 1050
rect 37310 1010 37330 1050
rect 37250 950 37330 1010
rect 37250 910 37270 950
rect 37310 910 37330 950
rect 37250 880 37330 910
rect 33860 450 33940 480
rect 33860 410 33880 450
rect 33920 410 33940 450
rect 33860 350 33940 410
rect 33860 310 33880 350
rect 33920 310 33940 350
rect 32790 250 32870 280
rect 32790 210 32810 250
rect 32850 210 32870 250
rect 32790 150 32870 210
rect 32790 110 32810 150
rect 32850 110 32870 150
rect 32790 80 32870 110
rect 33400 250 33480 280
rect 33400 210 33420 250
rect 33460 210 33480 250
rect 33400 150 33480 210
rect 33400 110 33420 150
rect 33460 110 33480 150
rect 33400 80 33480 110
rect 33860 250 33940 310
rect 33860 210 33880 250
rect 33920 210 33940 250
rect 33860 150 33940 210
rect 33860 110 33880 150
rect 33920 110 33940 150
rect 33860 50 33940 110
rect 33860 10 33880 50
rect 33920 10 33940 50
rect 33860 -50 33940 10
rect 33860 -90 33880 -50
rect 33920 -90 33940 -50
rect 33860 -120 33940 -90
rect 37260 450 37340 480
rect 37260 410 37280 450
rect 37320 410 37340 450
rect 37260 350 37340 410
rect 37260 310 37280 350
rect 37320 310 37340 350
rect 37260 250 37340 310
rect 37260 210 37280 250
rect 37320 210 37340 250
rect 37260 150 37340 210
rect 37260 110 37280 150
rect 37320 110 37340 150
rect 37260 50 37340 110
rect 37260 10 37280 50
rect 37320 10 37340 50
rect 37260 -50 37340 10
rect 37260 -90 37280 -50
rect 37320 -90 37340 -50
rect 37260 -120 37340 -90
rect 32760 -1110 32840 -1080
rect 32760 -1150 32780 -1110
rect 32820 -1150 32840 -1110
rect 32760 -1210 32840 -1150
rect 32760 -1250 32780 -1210
rect 32820 -1250 32840 -1210
rect 32760 -1280 32840 -1250
rect 35320 -1110 35400 -1080
rect 35320 -1150 35340 -1110
rect 35380 -1150 35400 -1110
rect 35320 -1210 35400 -1150
rect 35320 -1250 35340 -1210
rect 35380 -1250 35400 -1210
rect 35320 -1280 35400 -1250
rect 35800 -1110 35880 -1080
rect 35800 -1150 35820 -1110
rect 35860 -1150 35880 -1110
rect 35800 -1210 35880 -1150
rect 35800 -1250 35820 -1210
rect 35860 -1250 35880 -1210
rect 35800 -1280 35880 -1250
rect 38360 -1110 38440 -1080
rect 38360 -1150 38380 -1110
rect 38420 -1150 38440 -1110
rect 38360 -1210 38440 -1150
rect 38360 -1250 38380 -1210
rect 38420 -1250 38440 -1210
rect 38360 -1280 38440 -1250
<< psubdiffcont >>
rect 35140 -2020 35180 -1980
rect 35140 -2100 35180 -2060
rect 35140 -2180 35180 -2140
rect 36020 -2020 36060 -1980
rect 36020 -2100 36060 -2060
rect 36020 -2180 36060 -2140
rect 34240 -2700 34280 -2660
rect 34240 -2800 34280 -2760
rect 34240 -2900 34280 -2860
rect 34240 -3000 34280 -2960
rect 34240 -3100 34280 -3060
rect 36920 -2700 36960 -2660
rect 36920 -2800 36960 -2760
rect 36920 -2900 36960 -2860
rect 36920 -3000 36960 -2960
rect 36920 -3100 36960 -3060
rect 33420 -3610 33460 -3570
rect 33420 -3710 33460 -3670
rect 35580 -8370 35620 -8330
rect 35580 -8450 35620 -8410
rect 35580 -8530 35620 -8490
<< nsubdiffcont >>
rect 33890 1010 33930 1050
rect 33890 910 33930 950
rect 35370 1010 35410 1050
rect 35370 910 35410 950
rect 35790 1010 35830 1050
rect 35790 910 35830 950
rect 37270 1010 37310 1050
rect 37270 910 37310 950
rect 33880 410 33920 450
rect 33880 310 33920 350
rect 32810 210 32850 250
rect 32810 110 32850 150
rect 33420 210 33460 250
rect 33420 110 33460 150
rect 33880 210 33920 250
rect 33880 110 33920 150
rect 33880 10 33920 50
rect 33880 -90 33920 -50
rect 37280 410 37320 450
rect 37280 310 37320 350
rect 37280 210 37320 250
rect 37280 110 37320 150
rect 37280 10 37320 50
rect 37280 -90 37320 -50
rect 32780 -1150 32820 -1110
rect 32780 -1250 32820 -1210
rect 35340 -1150 35380 -1110
rect 35340 -1250 35380 -1210
rect 35820 -1150 35860 -1110
rect 35820 -1250 35860 -1210
rect 38380 -1150 38420 -1110
rect 38380 -1250 38420 -1210
<< poly >>
rect 33950 1170 34030 1190
rect 33950 1130 33970 1170
rect 34010 1140 34030 1170
rect 35270 1170 35350 1190
rect 35270 1140 35290 1170
rect 34010 1130 34060 1140
rect 33950 1110 34060 1130
rect 35240 1130 35290 1140
rect 35330 1130 35350 1170
rect 35240 1110 35350 1130
rect 35850 1170 35930 1190
rect 35850 1130 35870 1170
rect 35910 1140 35930 1170
rect 37170 1170 37250 1190
rect 37170 1140 37190 1170
rect 35910 1130 35960 1140
rect 35850 1110 35960 1130
rect 37140 1130 37190 1140
rect 37230 1130 37250 1170
rect 37140 1110 37250 1130
rect 34030 1080 34060 1110
rect 34140 1080 34170 1110
rect 34250 1080 34280 1110
rect 34360 1080 34390 1110
rect 34470 1080 34500 1110
rect 34580 1080 34610 1110
rect 34690 1080 34720 1110
rect 34800 1080 34830 1110
rect 34910 1080 34940 1110
rect 35020 1080 35050 1110
rect 35130 1080 35160 1110
rect 35240 1080 35270 1110
rect 35930 1080 35960 1110
rect 36040 1080 36070 1110
rect 36150 1080 36180 1110
rect 36260 1080 36290 1110
rect 36370 1080 36400 1110
rect 36480 1080 36510 1110
rect 36590 1080 36620 1110
rect 36700 1080 36730 1110
rect 36810 1080 36840 1110
rect 36920 1080 36950 1110
rect 37030 1080 37060 1110
rect 37140 1080 37170 1110
rect 34030 850 34060 880
rect 34140 850 34170 880
rect 34250 850 34280 880
rect 34360 850 34390 880
rect 34470 850 34500 880
rect 34580 850 34610 880
rect 34690 850 34720 880
rect 34800 850 34830 880
rect 34910 850 34940 880
rect 35020 850 35050 880
rect 35130 850 35160 880
rect 35240 850 35270 880
rect 35930 850 35960 880
rect 36040 850 36070 880
rect 36150 850 36180 880
rect 36260 850 36290 880
rect 36370 850 36400 880
rect 36480 850 36510 880
rect 36590 850 36620 880
rect 36700 850 36730 880
rect 36810 850 36840 880
rect 36920 850 36950 880
rect 37030 850 37060 880
rect 37140 850 37170 880
rect 34126 832 34184 850
rect 34126 798 34138 832
rect 34172 798 34184 832
rect 34126 780 34184 798
rect 34236 832 34294 850
rect 34236 798 34248 832
rect 34282 798 34294 832
rect 34236 780 34294 798
rect 34346 832 34404 850
rect 34346 798 34358 832
rect 34392 798 34404 832
rect 34346 780 34404 798
rect 34456 832 34514 850
rect 34456 798 34468 832
rect 34502 798 34514 832
rect 34456 780 34514 798
rect 34566 832 34624 850
rect 34566 798 34578 832
rect 34612 798 34624 832
rect 34566 780 34624 798
rect 34676 832 34734 850
rect 34676 798 34688 832
rect 34722 798 34734 832
rect 34676 780 34734 798
rect 34786 832 34844 850
rect 34786 798 34798 832
rect 34832 798 34844 832
rect 34786 780 34844 798
rect 34896 832 34954 850
rect 34896 798 34908 832
rect 34942 798 34954 832
rect 34896 780 34954 798
rect 35006 832 35064 850
rect 35006 798 35018 832
rect 35052 798 35064 832
rect 35006 780 35064 798
rect 35116 832 35174 850
rect 35116 798 35128 832
rect 35162 798 35174 832
rect 35116 780 35174 798
rect 36026 832 36084 850
rect 36026 798 36038 832
rect 36072 798 36084 832
rect 36026 780 36084 798
rect 36136 832 36194 850
rect 36136 798 36148 832
rect 36182 798 36194 832
rect 36136 780 36194 798
rect 36246 832 36304 850
rect 36246 798 36258 832
rect 36292 798 36304 832
rect 36246 780 36304 798
rect 36356 832 36414 850
rect 36356 798 36368 832
rect 36402 798 36414 832
rect 36356 780 36414 798
rect 36466 832 36524 850
rect 36466 798 36478 832
rect 36512 798 36524 832
rect 36466 780 36524 798
rect 36576 832 36634 850
rect 36576 798 36588 832
rect 36622 798 36634 832
rect 36576 780 36634 798
rect 36686 832 36744 850
rect 36686 798 36698 832
rect 36732 798 36744 832
rect 36686 780 36744 798
rect 36796 832 36854 850
rect 36796 798 36808 832
rect 36842 798 36854 832
rect 36796 780 36854 798
rect 36906 832 36964 850
rect 36906 798 36918 832
rect 36952 798 36964 832
rect 36906 780 36964 798
rect 37016 832 37074 850
rect 37016 798 37028 832
rect 37062 798 37074 832
rect 37016 780 37074 798
rect 33940 570 34020 590
rect 33940 530 33960 570
rect 34000 540 34020 570
rect 37180 570 37260 590
rect 37180 540 37200 570
rect 34000 530 34120 540
rect 33940 510 34120 530
rect 37080 530 37200 540
rect 37240 530 37260 570
rect 37080 510 37260 530
rect 34020 480 34120 510
rect 34200 480 34300 510
rect 34380 480 34480 510
rect 34560 480 34660 510
rect 34740 480 34840 510
rect 34920 480 35020 510
rect 35100 480 35200 510
rect 35280 480 35380 510
rect 35460 480 35560 510
rect 35640 480 35740 510
rect 35820 480 35920 510
rect 36000 480 36100 510
rect 36180 480 36280 510
rect 36360 480 36460 510
rect 36540 480 36640 510
rect 36720 480 36820 510
rect 36900 480 37000 510
rect 37080 480 37180 510
rect 32880 370 32940 390
rect 32880 330 32890 370
rect 32930 330 32940 370
rect 33320 370 33380 390
rect 33320 330 33330 370
rect 33370 330 33380 370
rect 32880 300 32980 330
rect 32950 280 32980 300
rect 33060 280 33090 310
rect 33170 280 33200 310
rect 33280 300 33380 330
rect 33280 280 33310 300
rect 32950 50 32980 80
rect 33060 60 33090 80
rect 33170 60 33200 80
rect 33060 30 33200 60
rect 33280 50 33310 80
rect 33090 -10 33110 30
rect 33150 -10 33170 30
rect 33090 -30 33170 -10
rect 34020 -150 34120 -120
rect 34200 -160 34300 -120
rect 34380 -150 34480 -120
rect 34560 -150 34660 -120
rect 34740 -150 34840 -120
rect 34920 -150 35020 -120
rect 35100 -150 35200 -120
rect 35280 -150 35380 -120
rect 35460 -150 35560 -120
rect 35640 -150 35740 -120
rect 35820 -150 35920 -120
rect 36000 -150 36100 -120
rect 36180 -150 36280 -120
rect 36360 -150 36460 -120
rect 36540 -150 36640 -120
rect 36720 -150 36820 -120
rect 36900 -150 37000 -120
rect 37080 -150 37180 -120
rect 34220 -170 34290 -160
rect 34220 -210 34230 -170
rect 34270 -210 34290 -170
rect 34220 -230 34290 -210
rect 34390 -170 34470 -150
rect 34390 -210 34410 -170
rect 34450 -210 34470 -170
rect 34390 -230 34470 -210
rect 34570 -170 34650 -150
rect 34570 -210 34590 -170
rect 34630 -210 34650 -170
rect 34570 -230 34650 -210
rect 34750 -170 34830 -150
rect 34750 -210 34770 -170
rect 34810 -210 34830 -170
rect 34750 -230 34830 -210
rect 34930 -170 35010 -150
rect 34930 -210 34950 -170
rect 34990 -210 35010 -170
rect 34930 -230 35010 -210
rect 35110 -170 35190 -150
rect 35110 -210 35130 -170
rect 35170 -210 35190 -170
rect 35110 -230 35190 -210
rect 35290 -170 35370 -150
rect 35290 -210 35310 -170
rect 35350 -210 35370 -170
rect 35290 -230 35370 -210
rect 35470 -170 35540 -150
rect 35470 -210 35490 -170
rect 35530 -210 35540 -170
rect 35470 -230 35540 -210
rect 35660 -170 35730 -150
rect 35660 -210 35670 -170
rect 35710 -210 35730 -170
rect 35660 -230 35730 -210
rect 35830 -170 35910 -150
rect 35830 -210 35850 -170
rect 35890 -210 35910 -170
rect 35830 -230 35910 -210
rect 36010 -170 36090 -150
rect 36010 -210 36030 -170
rect 36070 -210 36090 -170
rect 36010 -230 36090 -210
rect 36190 -170 36270 -150
rect 36190 -210 36210 -170
rect 36250 -210 36270 -170
rect 36190 -230 36270 -210
rect 36370 -170 36450 -150
rect 36370 -210 36390 -170
rect 36430 -210 36450 -170
rect 36370 -230 36450 -210
rect 36550 -170 36630 -150
rect 36550 -210 36570 -170
rect 36610 -210 36630 -170
rect 36550 -230 36630 -210
rect 36730 -170 36810 -150
rect 36730 -210 36750 -170
rect 36790 -210 36810 -170
rect 36730 -230 36810 -210
rect 36910 -170 36980 -150
rect 36910 -210 36930 -170
rect 36970 -210 36980 -170
rect 36910 -230 36980 -210
rect 32850 -990 32910 -970
rect 32850 -1030 32860 -990
rect 32900 -1020 32910 -990
rect 35250 -990 35310 -970
rect 35250 -1020 35260 -990
rect 32900 -1030 32960 -1020
rect 32850 -1050 32960 -1030
rect 35200 -1030 35260 -1020
rect 35300 -1030 35310 -990
rect 35200 -1050 35310 -1030
rect 35890 -990 35950 -970
rect 35890 -1030 35900 -990
rect 35940 -1020 35950 -990
rect 38290 -990 38350 -970
rect 38290 -1020 38300 -990
rect 35940 -1030 36000 -1020
rect 35890 -1050 36000 -1030
rect 38240 -1030 38300 -1020
rect 38340 -1030 38350 -990
rect 38240 -1050 38350 -1030
rect 32920 -1080 32960 -1050
rect 33040 -1080 33080 -1050
rect 33160 -1080 33200 -1050
rect 33280 -1080 33320 -1050
rect 33400 -1080 33440 -1050
rect 33520 -1080 33560 -1050
rect 33640 -1080 33680 -1050
rect 33760 -1080 33800 -1050
rect 33880 -1080 33920 -1050
rect 34000 -1080 34040 -1050
rect 34120 -1080 34160 -1050
rect 34240 -1080 34280 -1050
rect 34360 -1080 34400 -1050
rect 34480 -1080 34520 -1050
rect 34600 -1080 34640 -1050
rect 34720 -1080 34760 -1050
rect 34840 -1080 34880 -1050
rect 34960 -1080 35000 -1050
rect 35080 -1080 35120 -1050
rect 35200 -1080 35240 -1050
rect 35960 -1080 36000 -1050
rect 36080 -1080 36120 -1050
rect 36200 -1080 36240 -1050
rect 36320 -1080 36360 -1050
rect 36440 -1080 36480 -1050
rect 36560 -1080 36600 -1050
rect 36680 -1080 36720 -1050
rect 36800 -1080 36840 -1050
rect 36920 -1080 36960 -1050
rect 37040 -1080 37080 -1050
rect 37160 -1080 37200 -1050
rect 37280 -1080 37320 -1050
rect 37400 -1080 37440 -1050
rect 37520 -1080 37560 -1050
rect 37640 -1080 37680 -1050
rect 37760 -1080 37800 -1050
rect 37880 -1080 37920 -1050
rect 38000 -1080 38040 -1050
rect 38120 -1080 38160 -1050
rect 38240 -1080 38280 -1050
rect 32920 -1310 32960 -1280
rect 33040 -1320 33080 -1280
rect 33160 -1300 33200 -1280
rect 33280 -1300 33320 -1280
rect 33400 -1300 33440 -1280
rect 33520 -1300 33560 -1280
rect 33030 -1340 33090 -1320
rect 33160 -1330 33560 -1300
rect 33640 -1300 33680 -1280
rect 33760 -1300 33800 -1280
rect 33640 -1330 33800 -1300
rect 33880 -1300 33920 -1280
rect 34000 -1300 34040 -1280
rect 34120 -1300 34160 -1280
rect 34240 -1300 34280 -1280
rect 33880 -1330 34280 -1300
rect 34360 -1300 34400 -1280
rect 34480 -1300 34520 -1280
rect 34360 -1330 34520 -1300
rect 34600 -1300 34640 -1280
rect 34720 -1300 34760 -1280
rect 34840 -1300 34880 -1280
rect 34960 -1300 35000 -1280
rect 34600 -1330 35000 -1300
rect 35080 -1310 35120 -1280
rect 35200 -1310 35240 -1280
rect 35960 -1310 36000 -1280
rect 36080 -1310 36120 -1280
rect 36200 -1300 36240 -1280
rect 36320 -1300 36360 -1280
rect 36440 -1300 36480 -1280
rect 36560 -1300 36600 -1280
rect 35070 -1330 35130 -1310
rect 33030 -1380 33040 -1340
rect 33080 -1380 33090 -1340
rect 33030 -1400 33090 -1380
rect 33200 -1370 33220 -1330
rect 33260 -1370 33280 -1330
rect 33200 -1390 33280 -1370
rect 33690 -1370 33700 -1330
rect 33740 -1370 33750 -1330
rect 33690 -1390 33750 -1370
rect 33920 -1370 33940 -1330
rect 33980 -1370 34000 -1330
rect 33920 -1390 34000 -1370
rect 34410 -1370 34420 -1330
rect 34460 -1370 34470 -1330
rect 34410 -1390 34470 -1370
rect 34640 -1370 34660 -1330
rect 34700 -1370 34720 -1330
rect 34640 -1390 34720 -1370
rect 35070 -1370 35080 -1330
rect 35120 -1370 35130 -1330
rect 35070 -1390 35130 -1370
rect 36070 -1330 36130 -1310
rect 36200 -1330 36600 -1300
rect 36680 -1300 36720 -1280
rect 36800 -1300 36840 -1280
rect 36680 -1330 36840 -1300
rect 36920 -1300 36960 -1280
rect 37040 -1300 37080 -1280
rect 37160 -1300 37200 -1280
rect 37280 -1300 37320 -1280
rect 36920 -1330 37320 -1300
rect 37400 -1300 37440 -1280
rect 37520 -1300 37560 -1280
rect 37400 -1330 37560 -1300
rect 37640 -1300 37680 -1280
rect 37760 -1300 37800 -1280
rect 37880 -1300 37920 -1280
rect 38000 -1300 38040 -1280
rect 37640 -1330 38040 -1300
rect 38120 -1320 38160 -1280
rect 38240 -1310 38280 -1280
rect 36070 -1370 36080 -1330
rect 36120 -1370 36130 -1330
rect 36070 -1390 36130 -1370
rect 36480 -1370 36500 -1330
rect 36540 -1370 36560 -1330
rect 36480 -1390 36560 -1370
rect 36730 -1370 36740 -1330
rect 36780 -1370 36790 -1330
rect 36730 -1390 36790 -1370
rect 37200 -1370 37220 -1330
rect 37260 -1370 37280 -1330
rect 37200 -1390 37280 -1370
rect 37450 -1370 37460 -1330
rect 37500 -1370 37510 -1330
rect 37450 -1390 37510 -1370
rect 37920 -1370 37940 -1330
rect 37980 -1370 38000 -1330
rect 37920 -1390 38000 -1370
rect 38110 -1340 38170 -1320
rect 38110 -1380 38120 -1340
rect 38160 -1380 38170 -1340
rect 38110 -1400 38170 -1380
rect 33852 -1938 33920 -1920
rect 33852 -1972 33864 -1938
rect 33898 -1972 33920 -1938
rect 33852 -1990 33920 -1972
rect 33760 -2020 33800 -1990
rect 33880 -2020 33920 -1990
rect 34000 -1938 34068 -1920
rect 34000 -1972 34022 -1938
rect 34056 -1972 34068 -1938
rect 34000 -1990 34068 -1972
rect 34334 -1938 34400 -1920
rect 34334 -1972 34346 -1938
rect 34380 -1972 34400 -1938
rect 34334 -1990 34400 -1972
rect 34000 -2020 34040 -1990
rect 34120 -2020 34160 -1990
rect 34240 -2020 34280 -1990
rect 34360 -2020 34400 -1990
rect 34480 -1938 34546 -1920
rect 34480 -1972 34500 -1938
rect 34534 -1972 34546 -1938
rect 34480 -1990 34546 -1972
rect 34812 -1938 34880 -1920
rect 34812 -1972 34824 -1938
rect 34858 -1972 34880 -1938
rect 36320 -1938 36388 -1920
rect 34812 -1990 34880 -1972
rect 34480 -2020 34520 -1990
rect 34600 -2020 34640 -1990
rect 34720 -2020 34760 -1990
rect 34840 -2020 34880 -1990
rect 33760 -2150 33800 -2120
rect 33880 -2150 33920 -2120
rect 34000 -2150 34040 -2120
rect 34120 -2150 34160 -2120
rect 34240 -2150 34280 -2120
rect 34360 -2150 34400 -2120
rect 34480 -2150 34520 -2120
rect 34600 -2150 34640 -2120
rect 34720 -2150 34760 -2120
rect 34840 -2150 34880 -2120
rect 33751 -2168 33809 -2150
rect 33751 -2202 33763 -2168
rect 33797 -2202 33809 -2168
rect 33751 -2220 33809 -2202
rect 34111 -2168 34169 -2150
rect 34111 -2202 34123 -2168
rect 34157 -2202 34169 -2168
rect 34111 -2220 34169 -2202
rect 34231 -2168 34289 -2150
rect 34231 -2202 34243 -2168
rect 34277 -2202 34289 -2168
rect 34231 -2220 34289 -2202
rect 34591 -2168 34649 -2150
rect 34591 -2202 34603 -2168
rect 34637 -2202 34649 -2168
rect 34591 -2220 34649 -2202
rect 34711 -2168 34769 -2150
rect 34711 -2202 34723 -2168
rect 34757 -2202 34769 -2168
rect 34711 -2220 34769 -2202
rect 36320 -1972 36342 -1938
rect 36376 -1972 36388 -1938
rect 36320 -1990 36388 -1972
rect 36654 -1938 36720 -1920
rect 36654 -1972 36666 -1938
rect 36700 -1972 36720 -1938
rect 36654 -1990 36720 -1972
rect 36320 -2020 36360 -1990
rect 36440 -2020 36480 -1990
rect 36560 -2020 36600 -1990
rect 36680 -2020 36720 -1990
rect 36800 -1938 36866 -1920
rect 36800 -1972 36820 -1938
rect 36854 -1972 36866 -1938
rect 36800 -1990 36866 -1972
rect 37132 -1938 37200 -1920
rect 37132 -1972 37144 -1938
rect 37178 -1972 37200 -1938
rect 37132 -1990 37200 -1972
rect 36800 -2020 36840 -1990
rect 36920 -2020 36960 -1990
rect 37040 -2020 37080 -1990
rect 37160 -2020 37200 -1990
rect 37280 -1938 37348 -1920
rect 37280 -1972 37302 -1938
rect 37336 -1972 37348 -1938
rect 37280 -1990 37348 -1972
rect 37280 -2020 37320 -1990
rect 37400 -2020 37440 -1990
rect 36320 -2150 36360 -2120
rect 36440 -2150 36480 -2120
rect 36560 -2150 36600 -2120
rect 36680 -2150 36720 -2120
rect 36800 -2150 36840 -2120
rect 36920 -2150 36960 -2120
rect 37040 -2150 37080 -2120
rect 37160 -2150 37200 -2120
rect 37280 -2150 37320 -2120
rect 37400 -2150 37440 -2120
rect 36431 -2168 36489 -2150
rect 36431 -2202 36443 -2168
rect 36477 -2202 36489 -2168
rect 36431 -2220 36489 -2202
rect 36551 -2168 36609 -2150
rect 36551 -2202 36563 -2168
rect 36597 -2202 36609 -2168
rect 36551 -2220 36609 -2202
rect 36911 -2168 36969 -2150
rect 36911 -2202 36923 -2168
rect 36957 -2202 36969 -2168
rect 36911 -2220 36969 -2202
rect 37031 -2168 37089 -2150
rect 37031 -2202 37043 -2168
rect 37077 -2202 37089 -2168
rect 37031 -2220 37089 -2202
rect 37391 -2168 37449 -2150
rect 37391 -2202 37403 -2168
rect 37437 -2202 37449 -2168
rect 37391 -2220 37449 -2202
rect 33240 -2540 33320 -2520
rect 33240 -2580 33260 -2540
rect 33300 -2580 33320 -2540
rect 33240 -2600 33320 -2580
rect 33480 -2540 33560 -2520
rect 33480 -2580 33500 -2540
rect 33540 -2580 33560 -2540
rect 33480 -2600 33560 -2580
rect 33720 -2540 33800 -2520
rect 33720 -2580 33740 -2540
rect 33780 -2580 33800 -2540
rect 33720 -2600 33800 -2580
rect 33960 -2540 34040 -2520
rect 33960 -2580 33980 -2540
rect 34020 -2580 34040 -2540
rect 33960 -2600 34040 -2580
rect 34600 -2540 34680 -2520
rect 34600 -2580 34620 -2540
rect 34660 -2580 34680 -2540
rect 34600 -2600 34680 -2580
rect 34840 -2540 34920 -2520
rect 34840 -2580 34860 -2540
rect 34900 -2580 34920 -2540
rect 34840 -2600 34920 -2580
rect 35080 -2540 35160 -2520
rect 35080 -2580 35100 -2540
rect 35140 -2580 35160 -2540
rect 35080 -2600 35160 -2580
rect 36040 -2540 36120 -2520
rect 36040 -2580 36060 -2540
rect 36100 -2580 36120 -2540
rect 36040 -2600 36120 -2580
rect 36280 -2540 36360 -2520
rect 36280 -2580 36300 -2540
rect 36340 -2580 36360 -2540
rect 36280 -2600 36360 -2580
rect 36520 -2540 36600 -2520
rect 36520 -2580 36540 -2540
rect 36580 -2580 36600 -2540
rect 36520 -2600 36600 -2580
rect 37160 -2540 37240 -2520
rect 37160 -2580 37180 -2540
rect 37220 -2580 37240 -2540
rect 37160 -2600 37240 -2580
rect 37400 -2540 37480 -2520
rect 37400 -2580 37420 -2540
rect 37460 -2580 37480 -2540
rect 37400 -2600 37480 -2580
rect 37640 -2540 37720 -2520
rect 37640 -2580 37660 -2540
rect 37700 -2580 37720 -2540
rect 37640 -2600 37720 -2580
rect 37880 -2540 37960 -2520
rect 37880 -2580 37900 -2540
rect 37940 -2580 37960 -2540
rect 37880 -2600 37960 -2580
rect 33140 -2630 34140 -2600
rect 34380 -2630 35380 -2600
rect 35820 -2630 36820 -2600
rect 37060 -2630 38060 -2600
rect 33140 -3160 34140 -3130
rect 34380 -3160 35380 -3130
rect 35820 -3160 36820 -3130
rect 37060 -3160 38060 -3130
rect 33640 -3450 33720 -3430
rect 33640 -3490 33660 -3450
rect 33700 -3490 33720 -3450
rect 33640 -3510 33720 -3490
rect 33800 -3450 33880 -3430
rect 33800 -3490 33820 -3450
rect 33860 -3490 33880 -3450
rect 33800 -3510 33880 -3490
rect 33960 -3450 34040 -3430
rect 33960 -3490 33980 -3450
rect 34020 -3490 34040 -3450
rect 33960 -3510 34040 -3490
rect 34120 -3450 34200 -3430
rect 34120 -3490 34140 -3450
rect 34180 -3490 34200 -3450
rect 34120 -3510 34200 -3490
rect 34280 -3450 34360 -3430
rect 34280 -3490 34300 -3450
rect 34340 -3490 34360 -3450
rect 34280 -3510 34360 -3490
rect 34440 -3450 34520 -3430
rect 34440 -3490 34460 -3450
rect 34500 -3490 34520 -3450
rect 34440 -3510 34520 -3490
rect 34600 -3450 34680 -3430
rect 34600 -3490 34620 -3450
rect 34660 -3490 34680 -3450
rect 34600 -3510 34680 -3490
rect 34760 -3450 34840 -3430
rect 34760 -3490 34780 -3450
rect 34820 -3490 34840 -3450
rect 34760 -3510 34840 -3490
rect 34920 -3450 35000 -3430
rect 34920 -3490 34940 -3450
rect 34980 -3490 35000 -3450
rect 34920 -3510 35000 -3490
rect 35080 -3450 35160 -3430
rect 35080 -3490 35100 -3450
rect 35140 -3490 35160 -3450
rect 35080 -3510 35160 -3490
rect 35240 -3450 35320 -3430
rect 35240 -3490 35260 -3450
rect 35300 -3490 35320 -3450
rect 35240 -3510 35320 -3490
rect 35400 -3450 35480 -3430
rect 35400 -3490 35420 -3450
rect 35460 -3490 35480 -3450
rect 35400 -3510 35480 -3490
rect 35720 -3450 35800 -3430
rect 35720 -3490 35740 -3450
rect 35780 -3490 35800 -3450
rect 35720 -3510 35800 -3490
rect 35880 -3450 35960 -3430
rect 35880 -3490 35900 -3450
rect 35940 -3490 35960 -3450
rect 35880 -3510 35960 -3490
rect 36040 -3450 36120 -3430
rect 36040 -3490 36060 -3450
rect 36100 -3490 36120 -3450
rect 36040 -3510 36120 -3490
rect 36200 -3450 36280 -3430
rect 36200 -3490 36220 -3450
rect 36260 -3490 36280 -3450
rect 36200 -3510 36280 -3490
rect 36360 -3450 36440 -3430
rect 36360 -3490 36380 -3450
rect 36420 -3490 36440 -3450
rect 36360 -3510 36440 -3490
rect 36520 -3450 36600 -3430
rect 36520 -3490 36540 -3450
rect 36580 -3490 36600 -3450
rect 36520 -3510 36600 -3490
rect 36680 -3450 36760 -3430
rect 36680 -3490 36700 -3450
rect 36740 -3490 36760 -3450
rect 36680 -3510 36760 -3490
rect 36840 -3450 36920 -3430
rect 36840 -3490 36860 -3450
rect 36900 -3490 36920 -3450
rect 36840 -3510 36920 -3490
rect 37000 -3450 37080 -3430
rect 37000 -3490 37020 -3450
rect 37060 -3490 37080 -3450
rect 37000 -3510 37080 -3490
rect 37160 -3450 37240 -3430
rect 37160 -3490 37180 -3450
rect 37220 -3490 37240 -3450
rect 37160 -3510 37240 -3490
rect 37320 -3450 37400 -3430
rect 37320 -3490 37340 -3450
rect 37380 -3490 37400 -3450
rect 37320 -3510 37400 -3490
rect 37480 -3450 37560 -3430
rect 37480 -3490 37500 -3450
rect 37540 -3490 37560 -3450
rect 37480 -3510 37560 -3490
rect 33560 -3540 35560 -3510
rect 35640 -3540 37640 -3510
rect 33560 -3770 35560 -3740
rect 35640 -3770 37640 -3740
<< polycont >>
rect 33970 1130 34010 1170
rect 35290 1130 35330 1170
rect 35870 1130 35910 1170
rect 37190 1130 37230 1170
rect 34138 798 34172 832
rect 34248 798 34282 832
rect 34358 798 34392 832
rect 34468 798 34502 832
rect 34578 798 34612 832
rect 34688 798 34722 832
rect 34798 798 34832 832
rect 34908 798 34942 832
rect 35018 798 35052 832
rect 35128 798 35162 832
rect 36038 798 36072 832
rect 36148 798 36182 832
rect 36258 798 36292 832
rect 36368 798 36402 832
rect 36478 798 36512 832
rect 36588 798 36622 832
rect 36698 798 36732 832
rect 36808 798 36842 832
rect 36918 798 36952 832
rect 37028 798 37062 832
rect 33960 530 34000 570
rect 37200 530 37240 570
rect 32890 330 32930 370
rect 33330 330 33370 370
rect 33110 -10 33150 30
rect 34230 -210 34270 -170
rect 34410 -210 34450 -170
rect 34590 -210 34630 -170
rect 34770 -210 34810 -170
rect 34950 -210 34990 -170
rect 35130 -210 35170 -170
rect 35310 -210 35350 -170
rect 35490 -210 35530 -170
rect 35670 -210 35710 -170
rect 35850 -210 35890 -170
rect 36030 -210 36070 -170
rect 36210 -210 36250 -170
rect 36390 -210 36430 -170
rect 36570 -210 36610 -170
rect 36750 -210 36790 -170
rect 36930 -210 36970 -170
rect 32860 -1030 32900 -990
rect 35260 -1030 35300 -990
rect 35900 -1030 35940 -990
rect 38300 -1030 38340 -990
rect 33040 -1380 33080 -1340
rect 33220 -1370 33260 -1330
rect 33700 -1370 33740 -1330
rect 33940 -1370 33980 -1330
rect 34420 -1370 34460 -1330
rect 34660 -1370 34700 -1330
rect 35080 -1370 35120 -1330
rect 36080 -1370 36120 -1330
rect 36500 -1370 36540 -1330
rect 36740 -1370 36780 -1330
rect 37220 -1370 37260 -1330
rect 37460 -1370 37500 -1330
rect 37940 -1370 37980 -1330
rect 38120 -1380 38160 -1340
rect 33864 -1972 33898 -1938
rect 34022 -1972 34056 -1938
rect 34346 -1972 34380 -1938
rect 34500 -1972 34534 -1938
rect 34824 -1972 34858 -1938
rect 33763 -2202 33797 -2168
rect 34123 -2202 34157 -2168
rect 34243 -2202 34277 -2168
rect 34603 -2202 34637 -2168
rect 34723 -2202 34757 -2168
rect 36342 -1972 36376 -1938
rect 36666 -1972 36700 -1938
rect 36820 -1972 36854 -1938
rect 37144 -1972 37178 -1938
rect 37302 -1972 37336 -1938
rect 36443 -2202 36477 -2168
rect 36563 -2202 36597 -2168
rect 36923 -2202 36957 -2168
rect 37043 -2202 37077 -2168
rect 37403 -2202 37437 -2168
rect 33260 -2580 33300 -2540
rect 33500 -2580 33540 -2540
rect 33740 -2580 33780 -2540
rect 33980 -2580 34020 -2540
rect 34620 -2580 34660 -2540
rect 34860 -2580 34900 -2540
rect 35100 -2580 35140 -2540
rect 36060 -2580 36100 -2540
rect 36300 -2580 36340 -2540
rect 36540 -2580 36580 -2540
rect 37180 -2580 37220 -2540
rect 37420 -2580 37460 -2540
rect 37660 -2580 37700 -2540
rect 37900 -2580 37940 -2540
rect 33660 -3490 33700 -3450
rect 33820 -3490 33860 -3450
rect 33980 -3490 34020 -3450
rect 34140 -3490 34180 -3450
rect 34300 -3490 34340 -3450
rect 34460 -3490 34500 -3450
rect 34620 -3490 34660 -3450
rect 34780 -3490 34820 -3450
rect 34940 -3490 34980 -3450
rect 35100 -3490 35140 -3450
rect 35260 -3490 35300 -3450
rect 35420 -3490 35460 -3450
rect 35740 -3490 35780 -3450
rect 35900 -3490 35940 -3450
rect 36060 -3490 36100 -3450
rect 36220 -3490 36260 -3450
rect 36380 -3490 36420 -3450
rect 36540 -3490 36580 -3450
rect 36700 -3490 36740 -3450
rect 36860 -3490 36900 -3450
rect 37020 -3490 37060 -3450
rect 37180 -3490 37220 -3450
rect 37340 -3490 37380 -3450
rect 37500 -3490 37540 -3450
<< xpolycontact >>
rect 34940 -4070 35380 -4000
rect 35808 -4070 36248 -4000
rect 33120 -6320 33190 -5880
rect 32340 -6962 32410 -6522
rect 32340 -7778 32410 -7340
rect 33000 -7170 33070 -6730
rect 33000 -7778 33070 -7338
rect 33120 -7928 33190 -7488
rect 33240 -6320 33310 -5880
rect 33240 -7928 33310 -7488
rect 33360 -6320 33430 -5880
rect 33360 -7928 33430 -7488
rect 37890 -6320 37960 -5880
rect 37890 -7928 37960 -7488
rect 38010 -6320 38080 -5880
rect 38010 -7928 38080 -7488
rect 38130 -6320 38200 -5880
rect 38130 -7928 38200 -7488
rect 38320 -6700 38390 -6260
rect 38320 -7778 38390 -7338
rect 38440 -6700 38510 -6260
rect 38440 -7778 38510 -7338
rect 38560 -6700 38630 -6260
rect 38560 -7778 38630 -7338
rect 38680 -6752 38750 -6312
rect 38680 -7568 38750 -7130
<< ppolyres >>
rect 32340 -7340 32410 -6962
rect 38680 -7130 38750 -6752
<< xpolyres >>
rect 35380 -4070 35808 -4000
rect 33000 -7338 33070 -7170
rect 33120 -7488 33190 -6320
rect 33240 -7488 33310 -6320
rect 33360 -7488 33430 -6320
rect 37890 -7488 37960 -6320
rect 38010 -7488 38080 -6320
rect 38130 -7488 38200 -6320
rect 38320 -7338 38390 -6700
rect 38440 -7338 38510 -6700
rect 38560 -7338 38630 -6700
<< locali >>
rect 33950 1170 34030 1190
rect 33950 1130 33970 1170
rect 34010 1130 34030 1170
rect 33950 1110 34030 1130
rect 35270 1170 35350 1190
rect 35270 1130 35290 1170
rect 35330 1130 35350 1170
rect 35270 1110 35350 1130
rect 35850 1170 35930 1190
rect 35850 1130 35870 1170
rect 35910 1130 35930 1170
rect 35850 1110 35930 1130
rect 37170 1170 37250 1190
rect 37170 1130 37190 1170
rect 37230 1130 37250 1170
rect 37170 1110 37250 1130
rect 33880 1050 34020 1070
rect 33880 1010 33890 1050
rect 33930 1010 33970 1050
rect 34010 1010 34020 1050
rect 33880 950 34020 1010
rect 33880 910 33890 950
rect 33930 910 33970 950
rect 34010 910 34020 950
rect 33880 890 34020 910
rect 34070 1050 34130 1070
rect 34070 1010 34080 1050
rect 34120 1010 34130 1050
rect 34070 950 34130 1010
rect 34070 910 34080 950
rect 34120 910 34130 950
rect 34070 890 34130 910
rect 34180 1050 34240 1070
rect 34180 1010 34190 1050
rect 34230 1010 34240 1050
rect 34180 950 34240 1010
rect 34180 910 34190 950
rect 34230 910 34240 950
rect 34180 890 34240 910
rect 34290 1050 34350 1070
rect 34290 1010 34300 1050
rect 34340 1010 34350 1050
rect 34290 950 34350 1010
rect 34290 910 34300 950
rect 34340 910 34350 950
rect 34290 890 34350 910
rect 34400 1050 34460 1070
rect 34400 1010 34410 1050
rect 34450 1010 34460 1050
rect 34400 950 34460 1010
rect 34400 910 34410 950
rect 34450 910 34460 950
rect 34400 890 34460 910
rect 34510 1050 34570 1070
rect 34510 1010 34520 1050
rect 34560 1010 34570 1050
rect 34510 950 34570 1010
rect 34510 910 34520 950
rect 34560 910 34570 950
rect 34510 890 34570 910
rect 34620 1050 34680 1070
rect 34620 1010 34630 1050
rect 34670 1010 34680 1050
rect 34620 950 34680 1010
rect 34620 910 34630 950
rect 34670 910 34680 950
rect 34620 890 34680 910
rect 34730 1050 34790 1070
rect 34730 1010 34740 1050
rect 34780 1010 34790 1050
rect 34730 950 34790 1010
rect 34730 910 34740 950
rect 34780 910 34790 950
rect 34730 890 34790 910
rect 34840 1050 34900 1070
rect 34840 1010 34850 1050
rect 34890 1010 34900 1050
rect 34840 950 34900 1010
rect 34840 910 34850 950
rect 34890 910 34900 950
rect 34840 890 34900 910
rect 34950 1050 35010 1070
rect 34950 1010 34960 1050
rect 35000 1010 35010 1050
rect 34950 950 35010 1010
rect 34950 910 34960 950
rect 35000 910 35010 950
rect 34950 890 35010 910
rect 35060 1050 35120 1070
rect 35060 1010 35070 1050
rect 35110 1010 35120 1050
rect 35060 950 35120 1010
rect 35060 910 35070 950
rect 35110 910 35120 950
rect 35060 890 35120 910
rect 35170 1050 35230 1070
rect 35170 1010 35180 1050
rect 35220 1010 35230 1050
rect 35170 950 35230 1010
rect 35170 910 35180 950
rect 35220 910 35230 950
rect 35170 890 35230 910
rect 35280 1050 35420 1070
rect 35280 1010 35290 1050
rect 35330 1010 35370 1050
rect 35410 1010 35420 1050
rect 35280 950 35420 1010
rect 35280 910 35290 950
rect 35330 910 35370 950
rect 35410 910 35420 950
rect 35280 890 35420 910
rect 35780 1050 35920 1070
rect 35780 1010 35790 1050
rect 35830 1010 35870 1050
rect 35910 1010 35920 1050
rect 35780 950 35920 1010
rect 35780 910 35790 950
rect 35830 910 35870 950
rect 35910 910 35920 950
rect 35780 890 35920 910
rect 35970 1050 36030 1070
rect 35970 1010 35980 1050
rect 36020 1010 36030 1050
rect 35970 950 36030 1010
rect 35970 910 35980 950
rect 36020 910 36030 950
rect 35970 890 36030 910
rect 36080 1050 36140 1070
rect 36080 1010 36090 1050
rect 36130 1010 36140 1050
rect 36080 950 36140 1010
rect 36080 910 36090 950
rect 36130 910 36140 950
rect 36080 890 36140 910
rect 36190 1050 36250 1070
rect 36190 1010 36200 1050
rect 36240 1010 36250 1050
rect 36190 950 36250 1010
rect 36190 910 36200 950
rect 36240 910 36250 950
rect 36190 890 36250 910
rect 36300 1050 36360 1070
rect 36300 1010 36310 1050
rect 36350 1010 36360 1050
rect 36300 950 36360 1010
rect 36300 910 36310 950
rect 36350 910 36360 950
rect 36300 890 36360 910
rect 36410 1050 36470 1070
rect 36410 1010 36420 1050
rect 36460 1010 36470 1050
rect 36410 950 36470 1010
rect 36410 910 36420 950
rect 36460 910 36470 950
rect 36410 890 36470 910
rect 36520 1050 36580 1070
rect 36520 1010 36530 1050
rect 36570 1010 36580 1050
rect 36520 950 36580 1010
rect 36520 910 36530 950
rect 36570 910 36580 950
rect 36520 890 36580 910
rect 36630 1050 36690 1070
rect 36630 1010 36640 1050
rect 36680 1010 36690 1050
rect 36630 950 36690 1010
rect 36630 910 36640 950
rect 36680 910 36690 950
rect 36630 890 36690 910
rect 36740 1050 36800 1070
rect 36740 1010 36750 1050
rect 36790 1010 36800 1050
rect 36740 950 36800 1010
rect 36740 910 36750 950
rect 36790 910 36800 950
rect 36740 890 36800 910
rect 36850 1050 36910 1070
rect 36850 1010 36860 1050
rect 36900 1010 36910 1050
rect 36850 950 36910 1010
rect 36850 910 36860 950
rect 36900 910 36910 950
rect 36850 890 36910 910
rect 36960 1050 37020 1070
rect 36960 1010 36970 1050
rect 37010 1010 37020 1050
rect 36960 950 37020 1010
rect 36960 910 36970 950
rect 37010 910 37020 950
rect 36960 890 37020 910
rect 37070 1050 37130 1070
rect 37070 1010 37080 1050
rect 37120 1010 37130 1050
rect 37070 950 37130 1010
rect 37070 910 37080 950
rect 37120 910 37130 950
rect 37070 890 37130 910
rect 37180 1050 37320 1070
rect 37180 1010 37190 1050
rect 37230 1010 37270 1050
rect 37310 1010 37320 1050
rect 37180 950 37320 1010
rect 37180 910 37190 950
rect 37230 910 37270 950
rect 37310 910 37320 950
rect 37180 890 37320 910
rect 34126 832 34184 850
rect 34126 798 34138 832
rect 34172 798 34184 832
rect 34126 780 34184 798
rect 34236 832 34294 850
rect 34236 798 34248 832
rect 34282 798 34294 832
rect 34236 780 34294 798
rect 34346 832 34404 850
rect 34346 798 34358 832
rect 34392 798 34404 832
rect 34346 780 34404 798
rect 34456 832 34514 850
rect 34456 798 34468 832
rect 34502 798 34514 832
rect 34456 780 34514 798
rect 34566 832 34624 850
rect 34566 798 34578 832
rect 34612 798 34624 832
rect 34566 780 34624 798
rect 34676 832 34734 850
rect 34676 798 34688 832
rect 34722 798 34734 832
rect 34676 780 34734 798
rect 34786 832 34844 850
rect 34786 798 34798 832
rect 34832 798 34844 832
rect 34786 780 34844 798
rect 34896 832 34954 850
rect 34896 798 34908 832
rect 34942 798 34954 832
rect 34896 780 34954 798
rect 35006 832 35064 850
rect 35006 798 35018 832
rect 35052 798 35064 832
rect 35006 780 35064 798
rect 35116 832 35174 850
rect 35116 798 35128 832
rect 35162 798 35174 832
rect 35116 780 35174 798
rect 36026 832 36084 850
rect 36026 798 36038 832
rect 36072 798 36084 832
rect 36026 780 36084 798
rect 36136 832 36194 850
rect 36136 798 36148 832
rect 36182 798 36194 832
rect 36136 780 36194 798
rect 36246 832 36304 850
rect 36246 798 36258 832
rect 36292 798 36304 832
rect 36246 780 36304 798
rect 36356 832 36414 850
rect 36356 798 36368 832
rect 36402 798 36414 832
rect 36356 780 36414 798
rect 36466 832 36524 850
rect 36466 798 36478 832
rect 36512 798 36524 832
rect 36466 780 36524 798
rect 36576 832 36634 850
rect 36576 798 36588 832
rect 36622 798 36634 832
rect 36576 780 36634 798
rect 36686 832 36744 850
rect 36686 798 36698 832
rect 36732 798 36744 832
rect 36686 780 36744 798
rect 36796 832 36854 850
rect 36796 798 36808 832
rect 36842 798 36854 832
rect 36796 780 36854 798
rect 36906 832 36964 850
rect 36906 798 36918 832
rect 36952 798 36964 832
rect 36906 780 36964 798
rect 37016 832 37074 850
rect 37016 798 37028 832
rect 37062 798 37074 832
rect 37016 780 37074 798
rect 33940 570 34020 590
rect 33940 530 33960 570
rect 34000 530 34020 570
rect 33940 510 34020 530
rect 34300 570 34380 590
rect 34300 530 34320 570
rect 34360 530 34380 570
rect 34300 510 34380 530
rect 34660 570 34740 590
rect 34660 530 34680 570
rect 34720 530 34740 570
rect 34660 510 34740 530
rect 35020 570 35100 590
rect 35020 530 35040 570
rect 35080 530 35100 570
rect 35020 510 35100 530
rect 35380 570 35460 590
rect 35380 530 35400 570
rect 35440 530 35460 570
rect 35380 510 35460 530
rect 35740 570 35820 590
rect 35740 530 35760 570
rect 35800 530 35820 570
rect 35740 510 35820 530
rect 36100 570 36180 590
rect 36100 530 36120 570
rect 36160 530 36180 570
rect 36100 510 36180 530
rect 36460 570 36540 590
rect 36460 530 36480 570
rect 36520 530 36540 570
rect 36460 510 36540 530
rect 36820 570 36900 590
rect 36820 530 36840 570
rect 36880 530 36900 570
rect 36820 510 36900 530
rect 37180 570 37260 590
rect 37180 530 37200 570
rect 37240 530 37260 570
rect 37180 510 37260 530
rect 33960 470 34000 510
rect 34320 470 34360 510
rect 34680 470 34720 510
rect 35040 470 35080 510
rect 35400 470 35440 510
rect 35760 470 35800 510
rect 36120 470 36160 510
rect 36480 470 36520 510
rect 36840 470 36880 510
rect 37200 470 37240 510
rect 33870 450 34010 470
rect 33870 410 33880 450
rect 33920 410 33960 450
rect 34000 410 34010 450
rect 32880 370 32940 390
rect 32880 330 32890 370
rect 32930 330 32940 370
rect 32880 310 32940 330
rect 33090 370 33170 390
rect 33090 330 33110 370
rect 33150 330 33170 370
rect 33090 310 33170 330
rect 33310 370 33390 390
rect 33310 330 33330 370
rect 33370 330 33390 370
rect 33310 310 33390 330
rect 33870 350 34010 410
rect 33870 310 33880 350
rect 33920 310 33960 350
rect 34000 310 34010 350
rect 32800 250 32940 270
rect 32800 210 32810 250
rect 32850 210 32890 250
rect 32930 210 32940 250
rect 32800 150 32940 210
rect 32800 110 32810 150
rect 32850 110 32890 150
rect 32930 110 32940 150
rect 32800 90 32940 110
rect 32990 250 33050 270
rect 32990 210 33000 250
rect 33040 210 33050 250
rect 32990 150 33050 210
rect 32990 110 33000 150
rect 33040 110 33050 150
rect 32990 90 33050 110
rect 33100 250 33160 270
rect 33100 210 33110 250
rect 33150 210 33160 250
rect 33100 150 33160 210
rect 33100 110 33110 150
rect 33150 110 33160 150
rect 33100 90 33160 110
rect 33210 250 33270 270
rect 33210 210 33220 250
rect 33260 210 33270 250
rect 33210 150 33270 210
rect 33210 110 33220 150
rect 33260 110 33270 150
rect 33210 90 33270 110
rect 33320 250 33470 270
rect 33320 210 33330 250
rect 33370 210 33420 250
rect 33460 210 33470 250
rect 33320 150 33470 210
rect 33320 110 33330 150
rect 33370 110 33420 150
rect 33460 110 33470 150
rect 33320 90 33470 110
rect 33870 250 34010 310
rect 33870 210 33880 250
rect 33920 210 33960 250
rect 34000 210 34010 250
rect 33870 150 34010 210
rect 33870 110 33880 150
rect 33920 110 33960 150
rect 34000 110 34010 150
rect 33870 50 34010 110
rect 32970 30 33050 50
rect 32970 -10 32990 30
rect 33030 -10 33050 30
rect 32970 -30 33050 -10
rect 33090 30 33170 50
rect 33090 -10 33110 30
rect 33150 -10 33170 30
rect 33090 -30 33170 -10
rect 33210 30 33290 50
rect 33210 -10 33230 30
rect 33270 -10 33290 30
rect 33210 -30 33290 -10
rect 33870 10 33880 50
rect 33920 10 33960 50
rect 34000 10 34010 50
rect 33870 -50 34010 10
rect 33870 -90 33880 -50
rect 33920 -90 33960 -50
rect 34000 -90 34010 -50
rect 33870 -110 34010 -90
rect 34130 450 34190 470
rect 34130 410 34140 450
rect 34180 410 34190 450
rect 34130 350 34190 410
rect 34130 310 34140 350
rect 34180 310 34190 350
rect 34130 250 34190 310
rect 34130 210 34140 250
rect 34180 210 34190 250
rect 34130 150 34190 210
rect 34130 110 34140 150
rect 34180 110 34190 150
rect 34130 50 34190 110
rect 34130 10 34140 50
rect 34180 10 34190 50
rect 34130 -50 34190 10
rect 34130 -90 34140 -50
rect 34180 -90 34190 -50
rect 34130 -110 34190 -90
rect 34310 450 34370 470
rect 34310 410 34320 450
rect 34360 410 34370 450
rect 34310 350 34370 410
rect 34310 310 34320 350
rect 34360 310 34370 350
rect 34310 250 34370 310
rect 34310 210 34320 250
rect 34360 210 34370 250
rect 34310 150 34370 210
rect 34310 110 34320 150
rect 34360 110 34370 150
rect 34310 50 34370 110
rect 34310 10 34320 50
rect 34360 10 34370 50
rect 34310 -50 34370 10
rect 34310 -90 34320 -50
rect 34360 -90 34370 -50
rect 34310 -110 34370 -90
rect 34490 450 34550 470
rect 34490 410 34500 450
rect 34540 410 34550 450
rect 34490 350 34550 410
rect 34490 310 34500 350
rect 34540 310 34550 350
rect 34490 250 34550 310
rect 34490 210 34500 250
rect 34540 210 34550 250
rect 34490 150 34550 210
rect 34490 110 34500 150
rect 34540 110 34550 150
rect 34490 50 34550 110
rect 34490 10 34500 50
rect 34540 10 34550 50
rect 34490 -50 34550 10
rect 34490 -90 34500 -50
rect 34540 -90 34550 -50
rect 34490 -110 34550 -90
rect 34670 450 34730 470
rect 34670 410 34680 450
rect 34720 410 34730 450
rect 34670 350 34730 410
rect 34670 310 34680 350
rect 34720 310 34730 350
rect 34670 250 34730 310
rect 34670 210 34680 250
rect 34720 210 34730 250
rect 34670 150 34730 210
rect 34670 110 34680 150
rect 34720 110 34730 150
rect 34670 50 34730 110
rect 34670 10 34680 50
rect 34720 10 34730 50
rect 34670 -50 34730 10
rect 34670 -90 34680 -50
rect 34720 -90 34730 -50
rect 34670 -110 34730 -90
rect 34850 450 34910 470
rect 34850 410 34860 450
rect 34900 410 34910 450
rect 34850 350 34910 410
rect 34850 310 34860 350
rect 34900 310 34910 350
rect 34850 250 34910 310
rect 34850 210 34860 250
rect 34900 210 34910 250
rect 34850 150 34910 210
rect 34850 110 34860 150
rect 34900 110 34910 150
rect 34850 50 34910 110
rect 34850 10 34860 50
rect 34900 10 34910 50
rect 34850 -50 34910 10
rect 34850 -90 34860 -50
rect 34900 -90 34910 -50
rect 34850 -110 34910 -90
rect 35030 450 35090 470
rect 35030 410 35040 450
rect 35080 410 35090 450
rect 35030 350 35090 410
rect 35030 310 35040 350
rect 35080 310 35090 350
rect 35030 250 35090 310
rect 35030 210 35040 250
rect 35080 210 35090 250
rect 35030 150 35090 210
rect 35030 110 35040 150
rect 35080 110 35090 150
rect 35030 50 35090 110
rect 35030 10 35040 50
rect 35080 10 35090 50
rect 35030 -50 35090 10
rect 35030 -90 35040 -50
rect 35080 -90 35090 -50
rect 35030 -110 35090 -90
rect 35210 450 35270 470
rect 35210 410 35220 450
rect 35260 410 35270 450
rect 35210 350 35270 410
rect 35210 310 35220 350
rect 35260 310 35270 350
rect 35210 250 35270 310
rect 35210 210 35220 250
rect 35260 210 35270 250
rect 35210 150 35270 210
rect 35210 110 35220 150
rect 35260 110 35270 150
rect 35210 50 35270 110
rect 35210 10 35220 50
rect 35260 10 35270 50
rect 35210 -50 35270 10
rect 35210 -90 35220 -50
rect 35260 -90 35270 -50
rect 35210 -110 35270 -90
rect 35390 450 35450 470
rect 35390 410 35400 450
rect 35440 410 35450 450
rect 35390 350 35450 410
rect 35390 310 35400 350
rect 35440 310 35450 350
rect 35390 250 35450 310
rect 35390 210 35400 250
rect 35440 210 35450 250
rect 35390 150 35450 210
rect 35390 110 35400 150
rect 35440 110 35450 150
rect 35390 50 35450 110
rect 35390 10 35400 50
rect 35440 10 35450 50
rect 35390 -50 35450 10
rect 35390 -90 35400 -50
rect 35440 -90 35450 -50
rect 35390 -110 35450 -90
rect 35570 450 35630 470
rect 35570 410 35580 450
rect 35620 410 35630 450
rect 35570 350 35630 410
rect 35570 310 35580 350
rect 35620 310 35630 350
rect 35570 250 35630 310
rect 35570 210 35580 250
rect 35620 210 35630 250
rect 35570 150 35630 210
rect 35570 110 35580 150
rect 35620 110 35630 150
rect 35570 50 35630 110
rect 35570 10 35580 50
rect 35620 10 35630 50
rect 35570 -50 35630 10
rect 35570 -90 35580 -50
rect 35620 -90 35630 -50
rect 35570 -110 35630 -90
rect 35750 450 35810 470
rect 35750 410 35760 450
rect 35800 410 35810 450
rect 35750 350 35810 410
rect 35750 310 35760 350
rect 35800 310 35810 350
rect 35750 250 35810 310
rect 35750 210 35760 250
rect 35800 210 35810 250
rect 35750 150 35810 210
rect 35750 110 35760 150
rect 35800 110 35810 150
rect 35750 50 35810 110
rect 35750 10 35760 50
rect 35800 10 35810 50
rect 35750 -50 35810 10
rect 35750 -90 35760 -50
rect 35800 -90 35810 -50
rect 35750 -110 35810 -90
rect 35930 450 35990 470
rect 35930 410 35940 450
rect 35980 410 35990 450
rect 35930 350 35990 410
rect 35930 310 35940 350
rect 35980 310 35990 350
rect 35930 250 35990 310
rect 35930 210 35940 250
rect 35980 210 35990 250
rect 35930 150 35990 210
rect 35930 110 35940 150
rect 35980 110 35990 150
rect 35930 50 35990 110
rect 35930 10 35940 50
rect 35980 10 35990 50
rect 35930 -50 35990 10
rect 35930 -90 35940 -50
rect 35980 -90 35990 -50
rect 35930 -110 35990 -90
rect 36110 450 36170 470
rect 36110 410 36120 450
rect 36160 410 36170 450
rect 36110 350 36170 410
rect 36110 310 36120 350
rect 36160 310 36170 350
rect 36110 250 36170 310
rect 36110 210 36120 250
rect 36160 210 36170 250
rect 36110 150 36170 210
rect 36110 110 36120 150
rect 36160 110 36170 150
rect 36110 50 36170 110
rect 36110 10 36120 50
rect 36160 10 36170 50
rect 36110 -50 36170 10
rect 36110 -90 36120 -50
rect 36160 -90 36170 -50
rect 36110 -110 36170 -90
rect 36290 450 36350 470
rect 36290 410 36300 450
rect 36340 410 36350 450
rect 36290 350 36350 410
rect 36290 310 36300 350
rect 36340 310 36350 350
rect 36290 250 36350 310
rect 36290 210 36300 250
rect 36340 210 36350 250
rect 36290 150 36350 210
rect 36290 110 36300 150
rect 36340 110 36350 150
rect 36290 50 36350 110
rect 36290 10 36300 50
rect 36340 10 36350 50
rect 36290 -50 36350 10
rect 36290 -90 36300 -50
rect 36340 -90 36350 -50
rect 36290 -110 36350 -90
rect 36470 450 36530 470
rect 36470 410 36480 450
rect 36520 410 36530 450
rect 36470 350 36530 410
rect 36470 310 36480 350
rect 36520 310 36530 350
rect 36470 250 36530 310
rect 36470 210 36480 250
rect 36520 210 36530 250
rect 36470 150 36530 210
rect 36470 110 36480 150
rect 36520 110 36530 150
rect 36470 50 36530 110
rect 36470 10 36480 50
rect 36520 10 36530 50
rect 36470 -50 36530 10
rect 36470 -90 36480 -50
rect 36520 -90 36530 -50
rect 36470 -110 36530 -90
rect 36650 450 36710 470
rect 36650 410 36660 450
rect 36700 410 36710 450
rect 36650 350 36710 410
rect 36650 310 36660 350
rect 36700 310 36710 350
rect 36650 250 36710 310
rect 36650 210 36660 250
rect 36700 210 36710 250
rect 36650 150 36710 210
rect 36650 110 36660 150
rect 36700 110 36710 150
rect 36650 50 36710 110
rect 36650 10 36660 50
rect 36700 10 36710 50
rect 36650 -50 36710 10
rect 36650 -90 36660 -50
rect 36700 -90 36710 -50
rect 36650 -110 36710 -90
rect 36830 450 36890 470
rect 36830 410 36840 450
rect 36880 410 36890 450
rect 36830 350 36890 410
rect 36830 310 36840 350
rect 36880 310 36890 350
rect 36830 250 36890 310
rect 36830 210 36840 250
rect 36880 210 36890 250
rect 36830 150 36890 210
rect 36830 110 36840 150
rect 36880 110 36890 150
rect 36830 50 36890 110
rect 36830 10 36840 50
rect 36880 10 36890 50
rect 36830 -50 36890 10
rect 36830 -90 36840 -50
rect 36880 -90 36890 -50
rect 36830 -110 36890 -90
rect 37010 450 37070 470
rect 37010 410 37020 450
rect 37060 410 37070 450
rect 37010 350 37070 410
rect 37010 310 37020 350
rect 37060 310 37070 350
rect 37010 250 37070 310
rect 37010 210 37020 250
rect 37060 210 37070 250
rect 37010 150 37070 210
rect 37010 110 37020 150
rect 37060 110 37070 150
rect 37010 50 37070 110
rect 37010 10 37020 50
rect 37060 10 37070 50
rect 37010 -50 37070 10
rect 37010 -90 37020 -50
rect 37060 -90 37070 -50
rect 37010 -110 37070 -90
rect 37190 450 37330 470
rect 37190 410 37200 450
rect 37240 410 37280 450
rect 37320 410 37330 450
rect 37190 350 37330 410
rect 37190 310 37200 350
rect 37240 310 37280 350
rect 37320 310 37330 350
rect 37190 250 37330 310
rect 37190 210 37200 250
rect 37240 210 37280 250
rect 37320 210 37330 250
rect 37190 150 37330 210
rect 37190 110 37200 150
rect 37240 110 37280 150
rect 37320 110 37330 150
rect 37190 50 37330 110
rect 37190 10 37200 50
rect 37240 10 37280 50
rect 37320 10 37330 50
rect 37190 -50 37330 10
rect 37190 -90 37200 -50
rect 37240 -90 37280 -50
rect 37320 -90 37330 -50
rect 37190 -110 37330 -90
rect 34220 -170 34290 -150
rect 34220 -210 34230 -170
rect 34270 -210 34290 -170
rect 34220 -230 34290 -210
rect 34390 -170 34470 -150
rect 34390 -210 34410 -170
rect 34450 -210 34470 -170
rect 34390 -230 34470 -210
rect 34570 -170 34650 -150
rect 34570 -210 34590 -170
rect 34630 -210 34650 -170
rect 34570 -230 34650 -210
rect 34750 -170 34830 -150
rect 34750 -210 34770 -170
rect 34810 -210 34830 -170
rect 34750 -230 34830 -210
rect 34930 -170 35010 -150
rect 34930 -210 34950 -170
rect 34990 -210 35010 -170
rect 34930 -230 35010 -210
rect 35110 -170 35190 -150
rect 35110 -210 35130 -170
rect 35170 -210 35190 -170
rect 35110 -230 35190 -210
rect 35290 -170 35370 -150
rect 35290 -210 35310 -170
rect 35350 -210 35370 -170
rect 35290 -230 35370 -210
rect 35470 -170 35540 -150
rect 35470 -210 35490 -170
rect 35530 -210 35540 -170
rect 35470 -230 35540 -210
rect 35660 -170 35730 -150
rect 35660 -210 35670 -170
rect 35710 -210 35730 -170
rect 35660 -230 35730 -210
rect 35830 -170 35910 -150
rect 35830 -210 35850 -170
rect 35890 -210 35910 -170
rect 35830 -230 35910 -210
rect 36010 -170 36090 -150
rect 36010 -210 36030 -170
rect 36070 -210 36090 -170
rect 36010 -230 36090 -210
rect 36190 -170 36270 -150
rect 36190 -210 36210 -170
rect 36250 -210 36270 -170
rect 36190 -230 36270 -210
rect 36370 -170 36450 -150
rect 36370 -210 36390 -170
rect 36430 -210 36450 -170
rect 36370 -230 36450 -210
rect 36550 -170 36630 -150
rect 36550 -210 36570 -170
rect 36610 -210 36630 -170
rect 36550 -230 36630 -210
rect 36730 -170 36810 -150
rect 36730 -210 36750 -170
rect 36790 -210 36810 -170
rect 36730 -230 36810 -210
rect 36910 -170 36980 -150
rect 36910 -210 36930 -170
rect 36970 -210 36980 -170
rect 36910 -230 36980 -210
rect 32850 -990 32910 -970
rect 32850 -1030 32860 -990
rect 32900 -1030 32910 -990
rect 32850 -1050 32910 -1030
rect 35250 -990 35310 -970
rect 35250 -1030 35260 -990
rect 35300 -1030 35310 -990
rect 35250 -1050 35310 -1030
rect 35890 -990 35950 -970
rect 35890 -1030 35900 -990
rect 35940 -1030 35950 -990
rect 35890 -1050 35950 -1030
rect 38290 -990 38350 -970
rect 38290 -1030 38300 -990
rect 38340 -1030 38350 -990
rect 38290 -1050 38350 -1030
rect 32770 -1110 32910 -1090
rect 32770 -1150 32780 -1110
rect 32820 -1150 32860 -1110
rect 32900 -1150 32910 -1110
rect 32770 -1210 32910 -1150
rect 32770 -1250 32780 -1210
rect 32820 -1250 32860 -1210
rect 32900 -1250 32910 -1210
rect 32770 -1270 32910 -1250
rect 32970 -1110 33030 -1090
rect 32970 -1150 32980 -1110
rect 33020 -1150 33030 -1110
rect 32970 -1210 33030 -1150
rect 32970 -1250 32980 -1210
rect 33020 -1250 33030 -1210
rect 32970 -1270 33030 -1250
rect 33090 -1110 33150 -1090
rect 33090 -1150 33100 -1110
rect 33140 -1150 33150 -1110
rect 33090 -1210 33150 -1150
rect 33090 -1250 33100 -1210
rect 33140 -1250 33150 -1210
rect 33090 -1270 33150 -1250
rect 33210 -1110 33270 -1090
rect 33210 -1150 33220 -1110
rect 33260 -1150 33270 -1110
rect 33210 -1210 33270 -1150
rect 33210 -1250 33220 -1210
rect 33260 -1250 33270 -1210
rect 33210 -1270 33270 -1250
rect 33330 -1110 33390 -1090
rect 33330 -1150 33340 -1110
rect 33380 -1150 33390 -1110
rect 33330 -1210 33390 -1150
rect 33330 -1250 33340 -1210
rect 33380 -1250 33390 -1210
rect 33330 -1270 33390 -1250
rect 33450 -1110 33510 -1090
rect 33450 -1150 33460 -1110
rect 33500 -1150 33510 -1110
rect 33450 -1210 33510 -1150
rect 33450 -1250 33460 -1210
rect 33500 -1250 33510 -1210
rect 33450 -1270 33510 -1250
rect 33570 -1110 33630 -1090
rect 33570 -1150 33580 -1110
rect 33620 -1150 33630 -1110
rect 33570 -1210 33630 -1150
rect 33570 -1250 33580 -1210
rect 33620 -1250 33630 -1210
rect 33570 -1270 33630 -1250
rect 33690 -1110 33750 -1090
rect 33690 -1150 33700 -1110
rect 33740 -1150 33750 -1110
rect 33690 -1210 33750 -1150
rect 33690 -1250 33700 -1210
rect 33740 -1250 33750 -1210
rect 33690 -1270 33750 -1250
rect 33810 -1110 33870 -1090
rect 33810 -1150 33820 -1110
rect 33860 -1150 33870 -1110
rect 33810 -1210 33870 -1150
rect 33810 -1250 33820 -1210
rect 33860 -1250 33870 -1210
rect 33810 -1270 33870 -1250
rect 33930 -1110 33990 -1090
rect 33930 -1150 33940 -1110
rect 33980 -1150 33990 -1110
rect 33930 -1210 33990 -1150
rect 33930 -1250 33940 -1210
rect 33980 -1250 33990 -1210
rect 33930 -1270 33990 -1250
rect 34050 -1110 34110 -1090
rect 34050 -1150 34060 -1110
rect 34100 -1150 34110 -1110
rect 34050 -1210 34110 -1150
rect 34050 -1250 34060 -1210
rect 34100 -1250 34110 -1210
rect 34050 -1270 34110 -1250
rect 34170 -1110 34230 -1090
rect 34170 -1150 34180 -1110
rect 34220 -1150 34230 -1110
rect 34170 -1210 34230 -1150
rect 34170 -1250 34180 -1210
rect 34220 -1250 34230 -1210
rect 34170 -1270 34230 -1250
rect 34290 -1110 34350 -1090
rect 34290 -1150 34300 -1110
rect 34340 -1150 34350 -1110
rect 34290 -1210 34350 -1150
rect 34290 -1250 34300 -1210
rect 34340 -1250 34350 -1210
rect 34290 -1270 34350 -1250
rect 34410 -1110 34470 -1090
rect 34410 -1150 34420 -1110
rect 34460 -1150 34470 -1110
rect 34410 -1210 34470 -1150
rect 34410 -1250 34420 -1210
rect 34460 -1250 34470 -1210
rect 34410 -1270 34470 -1250
rect 34530 -1110 34590 -1090
rect 34530 -1150 34540 -1110
rect 34580 -1150 34590 -1110
rect 34530 -1210 34590 -1150
rect 34530 -1250 34540 -1210
rect 34580 -1250 34590 -1210
rect 34530 -1270 34590 -1250
rect 34650 -1110 34710 -1090
rect 34650 -1150 34660 -1110
rect 34700 -1150 34710 -1110
rect 34650 -1210 34710 -1150
rect 34650 -1250 34660 -1210
rect 34700 -1250 34710 -1210
rect 34650 -1270 34710 -1250
rect 34770 -1110 34830 -1090
rect 34770 -1150 34780 -1110
rect 34820 -1150 34830 -1110
rect 34770 -1210 34830 -1150
rect 34770 -1250 34780 -1210
rect 34820 -1250 34830 -1210
rect 34770 -1270 34830 -1250
rect 34890 -1110 34950 -1090
rect 34890 -1150 34900 -1110
rect 34940 -1150 34950 -1110
rect 34890 -1210 34950 -1150
rect 34890 -1250 34900 -1210
rect 34940 -1250 34950 -1210
rect 34890 -1270 34950 -1250
rect 35010 -1110 35070 -1090
rect 35010 -1150 35020 -1110
rect 35060 -1150 35070 -1110
rect 35010 -1210 35070 -1150
rect 35010 -1250 35020 -1210
rect 35060 -1250 35070 -1210
rect 35010 -1270 35070 -1250
rect 35130 -1110 35190 -1090
rect 35130 -1150 35140 -1110
rect 35180 -1150 35190 -1110
rect 35130 -1210 35190 -1150
rect 35130 -1250 35140 -1210
rect 35180 -1250 35190 -1210
rect 35130 -1270 35190 -1250
rect 35250 -1110 35390 -1090
rect 35250 -1150 35260 -1110
rect 35300 -1150 35340 -1110
rect 35380 -1150 35390 -1110
rect 35250 -1210 35390 -1150
rect 35250 -1250 35260 -1210
rect 35300 -1250 35340 -1210
rect 35380 -1250 35390 -1210
rect 35250 -1270 35390 -1250
rect 35810 -1110 35950 -1090
rect 35810 -1150 35820 -1110
rect 35860 -1150 35900 -1110
rect 35940 -1150 35950 -1110
rect 35810 -1210 35950 -1150
rect 35810 -1250 35820 -1210
rect 35860 -1250 35900 -1210
rect 35940 -1250 35950 -1210
rect 35810 -1270 35950 -1250
rect 36010 -1110 36070 -1090
rect 36010 -1150 36020 -1110
rect 36060 -1150 36070 -1110
rect 36010 -1210 36070 -1150
rect 36010 -1250 36020 -1210
rect 36060 -1250 36070 -1210
rect 36010 -1270 36070 -1250
rect 36130 -1110 36190 -1090
rect 36130 -1150 36140 -1110
rect 36180 -1150 36190 -1110
rect 36130 -1210 36190 -1150
rect 36130 -1250 36140 -1210
rect 36180 -1250 36190 -1210
rect 36130 -1270 36190 -1250
rect 36250 -1110 36310 -1090
rect 36250 -1150 36260 -1110
rect 36300 -1150 36310 -1110
rect 36250 -1210 36310 -1150
rect 36250 -1250 36260 -1210
rect 36300 -1250 36310 -1210
rect 36250 -1270 36310 -1250
rect 36370 -1110 36430 -1090
rect 36370 -1150 36380 -1110
rect 36420 -1150 36430 -1110
rect 36370 -1210 36430 -1150
rect 36370 -1250 36380 -1210
rect 36420 -1250 36430 -1210
rect 36370 -1270 36430 -1250
rect 36490 -1110 36550 -1090
rect 36490 -1150 36500 -1110
rect 36540 -1150 36550 -1110
rect 36490 -1210 36550 -1150
rect 36490 -1250 36500 -1210
rect 36540 -1250 36550 -1210
rect 36490 -1270 36550 -1250
rect 36610 -1110 36670 -1090
rect 36610 -1150 36620 -1110
rect 36660 -1150 36670 -1110
rect 36610 -1210 36670 -1150
rect 36610 -1250 36620 -1210
rect 36660 -1250 36670 -1210
rect 36610 -1270 36670 -1250
rect 36730 -1110 36790 -1090
rect 36730 -1150 36740 -1110
rect 36780 -1150 36790 -1110
rect 36730 -1210 36790 -1150
rect 36730 -1250 36740 -1210
rect 36780 -1250 36790 -1210
rect 36730 -1270 36790 -1250
rect 36850 -1110 36910 -1090
rect 36850 -1150 36860 -1110
rect 36900 -1150 36910 -1110
rect 36850 -1210 36910 -1150
rect 36850 -1250 36860 -1210
rect 36900 -1250 36910 -1210
rect 36850 -1270 36910 -1250
rect 36970 -1110 37030 -1090
rect 36970 -1150 36980 -1110
rect 37020 -1150 37030 -1110
rect 36970 -1210 37030 -1150
rect 36970 -1250 36980 -1210
rect 37020 -1250 37030 -1210
rect 36970 -1270 37030 -1250
rect 37090 -1110 37150 -1090
rect 37090 -1150 37100 -1110
rect 37140 -1150 37150 -1110
rect 37090 -1210 37150 -1150
rect 37090 -1250 37100 -1210
rect 37140 -1250 37150 -1210
rect 37090 -1270 37150 -1250
rect 37210 -1110 37270 -1090
rect 37210 -1150 37220 -1110
rect 37260 -1150 37270 -1110
rect 37210 -1210 37270 -1150
rect 37210 -1250 37220 -1210
rect 37260 -1250 37270 -1210
rect 37210 -1270 37270 -1250
rect 37330 -1110 37390 -1090
rect 37330 -1150 37340 -1110
rect 37380 -1150 37390 -1110
rect 37330 -1210 37390 -1150
rect 37330 -1250 37340 -1210
rect 37380 -1250 37390 -1210
rect 37330 -1270 37390 -1250
rect 37450 -1110 37510 -1090
rect 37450 -1150 37460 -1110
rect 37500 -1150 37510 -1110
rect 37450 -1210 37510 -1150
rect 37450 -1250 37460 -1210
rect 37500 -1250 37510 -1210
rect 37450 -1270 37510 -1250
rect 37570 -1110 37630 -1090
rect 37570 -1150 37580 -1110
rect 37620 -1150 37630 -1110
rect 37570 -1210 37630 -1150
rect 37570 -1250 37580 -1210
rect 37620 -1250 37630 -1210
rect 37570 -1270 37630 -1250
rect 37690 -1110 37750 -1090
rect 37690 -1150 37700 -1110
rect 37740 -1150 37750 -1110
rect 37690 -1210 37750 -1150
rect 37690 -1250 37700 -1210
rect 37740 -1250 37750 -1210
rect 37690 -1270 37750 -1250
rect 37810 -1110 37870 -1090
rect 37810 -1150 37820 -1110
rect 37860 -1150 37870 -1110
rect 37810 -1210 37870 -1150
rect 37810 -1250 37820 -1210
rect 37860 -1250 37870 -1210
rect 37810 -1270 37870 -1250
rect 37930 -1110 37990 -1090
rect 37930 -1150 37940 -1110
rect 37980 -1150 37990 -1110
rect 37930 -1210 37990 -1150
rect 37930 -1250 37940 -1210
rect 37980 -1250 37990 -1210
rect 37930 -1270 37990 -1250
rect 38050 -1110 38110 -1090
rect 38050 -1150 38060 -1110
rect 38100 -1150 38110 -1110
rect 38050 -1210 38110 -1150
rect 38050 -1250 38060 -1210
rect 38100 -1250 38110 -1210
rect 38050 -1270 38110 -1250
rect 38170 -1110 38230 -1090
rect 38170 -1150 38180 -1110
rect 38220 -1150 38230 -1110
rect 38170 -1210 38230 -1150
rect 38170 -1250 38180 -1210
rect 38220 -1250 38230 -1210
rect 38170 -1270 38230 -1250
rect 38290 -1110 38430 -1090
rect 38290 -1150 38300 -1110
rect 38340 -1150 38380 -1110
rect 38420 -1150 38430 -1110
rect 38290 -1210 38430 -1150
rect 38290 -1250 38300 -1210
rect 38340 -1250 38380 -1210
rect 38420 -1250 38430 -1210
rect 38290 -1270 38430 -1250
rect 33030 -1340 33090 -1320
rect 33030 -1380 33040 -1340
rect 33080 -1380 33090 -1340
rect 33030 -1400 33090 -1380
rect 33200 -1330 33280 -1310
rect 33200 -1370 33220 -1330
rect 33260 -1370 33280 -1330
rect 33200 -1390 33280 -1370
rect 33690 -1330 33750 -1310
rect 33690 -1370 33700 -1330
rect 33740 -1370 33750 -1330
rect 33690 -1390 33750 -1370
rect 33920 -1330 34000 -1310
rect 33920 -1370 33940 -1330
rect 33980 -1370 34000 -1330
rect 33920 -1390 34000 -1370
rect 34410 -1330 34470 -1310
rect 34410 -1370 34420 -1330
rect 34460 -1370 34470 -1330
rect 34410 -1390 34470 -1370
rect 34640 -1330 34720 -1310
rect 34640 -1370 34660 -1330
rect 34700 -1370 34720 -1330
rect 34640 -1390 34720 -1370
rect 35070 -1330 35130 -1310
rect 35070 -1370 35080 -1330
rect 35120 -1370 35130 -1330
rect 35070 -1390 35130 -1370
rect 36070 -1330 36130 -1310
rect 36070 -1370 36080 -1330
rect 36120 -1370 36130 -1330
rect 36070 -1390 36130 -1370
rect 36480 -1330 36560 -1310
rect 36480 -1370 36500 -1330
rect 36540 -1370 36560 -1330
rect 36480 -1390 36560 -1370
rect 36730 -1330 36790 -1310
rect 36730 -1370 36740 -1330
rect 36780 -1370 36790 -1330
rect 36730 -1390 36790 -1370
rect 37200 -1330 37280 -1310
rect 37200 -1370 37220 -1330
rect 37260 -1370 37280 -1330
rect 37200 -1390 37280 -1370
rect 37450 -1330 37510 -1310
rect 37450 -1370 37460 -1330
rect 37500 -1370 37510 -1330
rect 37450 -1390 37510 -1370
rect 37920 -1330 38000 -1310
rect 37920 -1370 37940 -1330
rect 37980 -1370 38000 -1330
rect 37920 -1390 38000 -1370
rect 38110 -1340 38170 -1320
rect 38110 -1380 38120 -1340
rect 38160 -1380 38170 -1340
rect 38110 -1400 38170 -1380
rect 33852 -1938 33910 -1920
rect 33852 -1972 33864 -1938
rect 33898 -1972 33910 -1938
rect 33852 -1990 33910 -1972
rect 34010 -1938 34068 -1920
rect 34010 -1972 34022 -1938
rect 34056 -1972 34068 -1938
rect 34010 -1990 34068 -1972
rect 34334 -1938 34392 -1920
rect 34334 -1972 34346 -1938
rect 34380 -1972 34392 -1938
rect 34334 -1990 34392 -1972
rect 34488 -1938 34546 -1920
rect 34488 -1972 34500 -1938
rect 34534 -1972 34546 -1938
rect 34488 -1990 34546 -1972
rect 34812 -1938 34870 -1920
rect 34812 -1972 34824 -1938
rect 34858 -1972 34870 -1938
rect 36330 -1938 36388 -1920
rect 34812 -1990 34870 -1972
rect 35120 -1980 35200 -1960
rect 35120 -2020 35140 -1980
rect 35180 -2020 35200 -1980
rect 33690 -2050 33750 -2030
rect 33690 -2090 33700 -2050
rect 33740 -2090 33750 -2050
rect 33690 -2110 33750 -2090
rect 33810 -2050 33870 -2030
rect 33810 -2090 33820 -2050
rect 33860 -2090 33870 -2050
rect 33810 -2110 33870 -2090
rect 33930 -2050 33990 -2030
rect 33930 -2090 33940 -2050
rect 33980 -2090 33990 -2050
rect 33930 -2110 33990 -2090
rect 34050 -2050 34110 -2030
rect 34050 -2090 34060 -2050
rect 34100 -2090 34110 -2050
rect 34050 -2110 34110 -2090
rect 34170 -2050 34230 -2030
rect 34170 -2090 34180 -2050
rect 34220 -2090 34230 -2050
rect 34170 -2110 34230 -2090
rect 34290 -2050 34350 -2030
rect 34290 -2090 34300 -2050
rect 34340 -2090 34350 -2050
rect 34290 -2110 34350 -2090
rect 34410 -2050 34470 -2030
rect 34410 -2090 34420 -2050
rect 34460 -2090 34470 -2050
rect 34410 -2110 34470 -2090
rect 34530 -2050 34590 -2030
rect 34530 -2090 34540 -2050
rect 34580 -2090 34590 -2050
rect 34530 -2110 34590 -2090
rect 34650 -2050 34710 -2030
rect 34650 -2090 34660 -2050
rect 34700 -2090 34710 -2050
rect 34650 -2110 34710 -2090
rect 34770 -2050 34830 -2030
rect 34770 -2090 34780 -2050
rect 34820 -2090 34830 -2050
rect 34770 -2110 34830 -2090
rect 34890 -2050 34950 -2030
rect 34890 -2090 34900 -2050
rect 34940 -2090 34950 -2050
rect 34890 -2110 34950 -2090
rect 35120 -2060 35200 -2020
rect 35120 -2100 35140 -2060
rect 35180 -2100 35200 -2060
rect 35120 -2140 35200 -2100
rect 33751 -2168 33809 -2150
rect 33751 -2202 33763 -2168
rect 33797 -2202 33809 -2168
rect 33751 -2220 33809 -2202
rect 34111 -2168 34169 -2150
rect 34111 -2202 34123 -2168
rect 34157 -2202 34169 -2168
rect 34111 -2220 34169 -2202
rect 34231 -2168 34289 -2150
rect 34231 -2202 34243 -2168
rect 34277 -2202 34289 -2168
rect 34231 -2220 34289 -2202
rect 34591 -2168 34649 -2150
rect 34591 -2202 34603 -2168
rect 34637 -2202 34649 -2168
rect 34591 -2220 34649 -2202
rect 34711 -2168 34769 -2150
rect 34711 -2202 34723 -2168
rect 34757 -2202 34769 -2168
rect 35120 -2180 35140 -2140
rect 35180 -2180 35200 -2140
rect 35120 -2200 35200 -2180
rect 36000 -1980 36080 -1960
rect 36000 -2020 36020 -1980
rect 36060 -2020 36080 -1980
rect 36330 -1972 36342 -1938
rect 36376 -1972 36388 -1938
rect 36330 -1990 36388 -1972
rect 36654 -1938 36712 -1920
rect 36654 -1972 36666 -1938
rect 36700 -1972 36712 -1938
rect 36654 -1990 36712 -1972
rect 36808 -1938 36866 -1920
rect 36808 -1972 36820 -1938
rect 36854 -1972 36866 -1938
rect 36808 -1990 36866 -1972
rect 37132 -1938 37190 -1920
rect 37132 -1972 37144 -1938
rect 37178 -1972 37190 -1938
rect 37132 -1990 37190 -1972
rect 37290 -1938 37348 -1920
rect 37290 -1972 37302 -1938
rect 37336 -1972 37348 -1938
rect 37290 -1990 37348 -1972
rect 36000 -2060 36080 -2020
rect 36000 -2100 36020 -2060
rect 36060 -2100 36080 -2060
rect 36000 -2140 36080 -2100
rect 36250 -2050 36310 -2030
rect 36250 -2090 36260 -2050
rect 36300 -2090 36310 -2050
rect 36250 -2110 36310 -2090
rect 36370 -2050 36430 -2030
rect 36370 -2090 36380 -2050
rect 36420 -2090 36430 -2050
rect 36370 -2110 36430 -2090
rect 36490 -2050 36550 -2030
rect 36490 -2090 36500 -2050
rect 36540 -2090 36550 -2050
rect 36490 -2110 36550 -2090
rect 36610 -2050 36670 -2030
rect 36610 -2090 36620 -2050
rect 36660 -2090 36670 -2050
rect 36610 -2110 36670 -2090
rect 36730 -2050 36790 -2030
rect 36730 -2090 36740 -2050
rect 36780 -2090 36790 -2050
rect 36730 -2110 36790 -2090
rect 36850 -2050 36910 -2030
rect 36850 -2090 36860 -2050
rect 36900 -2090 36910 -2050
rect 36850 -2110 36910 -2090
rect 36970 -2050 37030 -2030
rect 36970 -2090 36980 -2050
rect 37020 -2090 37030 -2050
rect 36970 -2110 37030 -2090
rect 37090 -2050 37150 -2030
rect 37090 -2090 37100 -2050
rect 37140 -2090 37150 -2050
rect 37090 -2110 37150 -2090
rect 37210 -2050 37270 -2030
rect 37210 -2090 37220 -2050
rect 37260 -2090 37270 -2050
rect 37210 -2110 37270 -2090
rect 37330 -2050 37390 -2030
rect 37330 -2090 37340 -2050
rect 37380 -2090 37390 -2050
rect 37330 -2110 37390 -2090
rect 37450 -2050 37510 -2030
rect 37450 -2090 37460 -2050
rect 37500 -2090 37510 -2050
rect 37450 -2110 37510 -2090
rect 36000 -2180 36020 -2140
rect 36060 -2180 36080 -2140
rect 36000 -2200 36080 -2180
rect 36431 -2168 36489 -2150
rect 34711 -2220 34769 -2202
rect 36431 -2202 36443 -2168
rect 36477 -2202 36489 -2168
rect 36431 -2220 36489 -2202
rect 36551 -2168 36609 -2150
rect 36551 -2202 36563 -2168
rect 36597 -2202 36609 -2168
rect 36551 -2220 36609 -2202
rect 36911 -2168 36969 -2150
rect 36911 -2202 36923 -2168
rect 36957 -2202 36969 -2168
rect 36911 -2220 36969 -2202
rect 37031 -2168 37089 -2150
rect 37031 -2202 37043 -2168
rect 37077 -2202 37089 -2168
rect 37031 -2220 37089 -2202
rect 37391 -2168 37449 -2150
rect 37391 -2202 37403 -2168
rect 37437 -2202 37449 -2168
rect 37391 -2220 37449 -2202
rect 33240 -2540 33320 -2520
rect 33240 -2580 33260 -2540
rect 33300 -2580 33320 -2540
rect 33240 -2600 33320 -2580
rect 33480 -2540 33560 -2520
rect 33480 -2580 33500 -2540
rect 33540 -2580 33560 -2540
rect 33480 -2600 33560 -2580
rect 33720 -2540 33800 -2520
rect 33720 -2580 33740 -2540
rect 33780 -2580 33800 -2540
rect 33720 -2600 33800 -2580
rect 33960 -2540 34040 -2520
rect 33960 -2580 33980 -2540
rect 34020 -2580 34040 -2540
rect 33960 -2600 34040 -2580
rect 34600 -2540 34680 -2520
rect 34600 -2580 34620 -2540
rect 34660 -2580 34680 -2540
rect 34600 -2600 34680 -2580
rect 34840 -2540 34920 -2520
rect 34840 -2580 34860 -2540
rect 34900 -2580 34920 -2540
rect 34840 -2600 34920 -2580
rect 35080 -2540 35160 -2520
rect 35080 -2580 35100 -2540
rect 35140 -2580 35160 -2540
rect 36040 -2540 36120 -2520
rect 35080 -2600 35160 -2580
rect 35390 -2570 35450 -2550
rect 35390 -2610 35400 -2570
rect 35440 -2610 35450 -2570
rect 33070 -2660 33130 -2640
rect 33070 -2700 33080 -2660
rect 33120 -2700 33130 -2660
rect 33070 -2760 33130 -2700
rect 33070 -2800 33080 -2760
rect 33120 -2800 33130 -2760
rect 33070 -2860 33130 -2800
rect 33070 -2900 33080 -2860
rect 33120 -2900 33130 -2860
rect 33070 -2960 33130 -2900
rect 33070 -3000 33080 -2960
rect 33120 -3000 33130 -2960
rect 33070 -3060 33130 -3000
rect 33070 -3100 33080 -3060
rect 33120 -3100 33130 -3060
rect 33070 -3120 33130 -3100
rect 34150 -2660 34370 -2640
rect 34150 -2700 34160 -2660
rect 34200 -2700 34240 -2660
rect 34280 -2700 34320 -2660
rect 34360 -2700 34370 -2660
rect 34150 -2760 34370 -2700
rect 34150 -2800 34160 -2760
rect 34200 -2800 34240 -2760
rect 34280 -2800 34320 -2760
rect 34360 -2800 34370 -2760
rect 34150 -2860 34370 -2800
rect 34150 -2900 34160 -2860
rect 34200 -2900 34240 -2860
rect 34280 -2900 34320 -2860
rect 34360 -2900 34370 -2860
rect 34150 -2960 34370 -2900
rect 34150 -3000 34160 -2960
rect 34200 -3000 34240 -2960
rect 34280 -3000 34320 -2960
rect 34360 -3000 34370 -2960
rect 34150 -3060 34370 -3000
rect 34150 -3100 34160 -3060
rect 34200 -3100 34240 -3060
rect 34280 -3100 34320 -3060
rect 34360 -3100 34370 -3060
rect 34150 -3120 34370 -3100
rect 35390 -2660 35450 -2610
rect 35390 -2700 35400 -2660
rect 35440 -2700 35450 -2660
rect 35390 -2760 35450 -2700
rect 35390 -2800 35400 -2760
rect 35440 -2800 35450 -2760
rect 35390 -2860 35450 -2800
rect 35390 -2900 35400 -2860
rect 35440 -2900 35450 -2860
rect 35390 -2960 35450 -2900
rect 35390 -3000 35400 -2960
rect 35440 -3000 35450 -2960
rect 35390 -3060 35450 -3000
rect 35390 -3100 35400 -3060
rect 35440 -3100 35450 -3060
rect 35390 -3120 35450 -3100
rect 35750 -2570 35810 -2550
rect 35750 -2610 35760 -2570
rect 35800 -2610 35810 -2570
rect 36040 -2580 36060 -2540
rect 36100 -2580 36120 -2540
rect 36040 -2600 36120 -2580
rect 36280 -2540 36360 -2520
rect 36280 -2580 36300 -2540
rect 36340 -2580 36360 -2540
rect 36280 -2600 36360 -2580
rect 36520 -2540 36600 -2520
rect 36520 -2580 36540 -2540
rect 36580 -2580 36600 -2540
rect 36520 -2600 36600 -2580
rect 37160 -2540 37240 -2520
rect 37160 -2580 37180 -2540
rect 37220 -2580 37240 -2540
rect 37160 -2600 37240 -2580
rect 37400 -2540 37480 -2520
rect 37400 -2580 37420 -2540
rect 37460 -2580 37480 -2540
rect 37400 -2600 37480 -2580
rect 37640 -2540 37720 -2520
rect 37640 -2580 37660 -2540
rect 37700 -2580 37720 -2540
rect 37640 -2600 37720 -2580
rect 37880 -2540 37960 -2520
rect 37880 -2580 37900 -2540
rect 37940 -2580 37960 -2540
rect 37880 -2600 37960 -2580
rect 38060 -2580 38140 -2560
rect 35750 -2660 35810 -2610
rect 38060 -2620 38080 -2580
rect 38120 -2620 38140 -2580
rect 38060 -2640 38140 -2620
rect 35750 -2700 35760 -2660
rect 35800 -2700 35810 -2660
rect 35750 -2760 35810 -2700
rect 35750 -2800 35760 -2760
rect 35800 -2800 35810 -2760
rect 35750 -2860 35810 -2800
rect 35750 -2900 35760 -2860
rect 35800 -2900 35810 -2860
rect 35750 -2960 35810 -2900
rect 35750 -3000 35760 -2960
rect 35800 -3000 35810 -2960
rect 35750 -3060 35810 -3000
rect 35750 -3100 35760 -3060
rect 35800 -3100 35810 -3060
rect 35750 -3120 35810 -3100
rect 36830 -2660 37050 -2640
rect 36830 -2700 36840 -2660
rect 36880 -2700 36920 -2660
rect 36960 -2700 37000 -2660
rect 37040 -2700 37050 -2660
rect 36830 -2760 37050 -2700
rect 36830 -2800 36840 -2760
rect 36880 -2800 36920 -2760
rect 36960 -2800 37000 -2760
rect 37040 -2800 37050 -2760
rect 36830 -2860 37050 -2800
rect 36830 -2900 36840 -2860
rect 36880 -2900 36920 -2860
rect 36960 -2900 37000 -2860
rect 37040 -2900 37050 -2860
rect 36830 -2960 37050 -2900
rect 36830 -3000 36840 -2960
rect 36880 -3000 36920 -2960
rect 36960 -3000 37000 -2960
rect 37040 -3000 37050 -2960
rect 36830 -3060 37050 -3000
rect 36830 -3100 36840 -3060
rect 36880 -3100 36920 -3060
rect 36960 -3100 37000 -3060
rect 37040 -3100 37050 -3060
rect 36830 -3120 37050 -3100
rect 38070 -2660 38130 -2640
rect 38070 -2700 38080 -2660
rect 38120 -2700 38130 -2660
rect 38070 -2760 38130 -2700
rect 38070 -2800 38080 -2760
rect 38120 -2800 38130 -2760
rect 38070 -2860 38130 -2800
rect 38070 -2900 38080 -2860
rect 38120 -2900 38130 -2860
rect 38070 -2960 38130 -2900
rect 38070 -3000 38080 -2960
rect 38120 -3000 38130 -2960
rect 38070 -3060 38130 -3000
rect 38070 -3100 38080 -3060
rect 38120 -3100 38130 -3060
rect 38070 -3120 38130 -3100
rect 34240 -3160 34280 -3120
rect 36920 -3160 36960 -3120
rect 34220 -3180 34300 -3160
rect 34220 -3220 34240 -3180
rect 34280 -3220 34300 -3180
rect 34220 -3240 34300 -3220
rect 36900 -3180 36980 -3160
rect 36900 -3220 36920 -3180
rect 36960 -3220 36980 -3180
rect 36900 -3240 36980 -3220
rect 33640 -3450 33720 -3430
rect 33640 -3490 33660 -3450
rect 33700 -3490 33720 -3450
rect 33640 -3510 33720 -3490
rect 33800 -3450 33880 -3430
rect 33800 -3490 33820 -3450
rect 33860 -3490 33880 -3450
rect 33800 -3510 33880 -3490
rect 33960 -3450 34040 -3430
rect 33960 -3490 33980 -3450
rect 34020 -3490 34040 -3450
rect 33960 -3510 34040 -3490
rect 34120 -3450 34200 -3430
rect 34120 -3490 34140 -3450
rect 34180 -3490 34200 -3450
rect 34120 -3510 34200 -3490
rect 34280 -3450 34360 -3430
rect 34280 -3490 34300 -3450
rect 34340 -3490 34360 -3450
rect 34280 -3510 34360 -3490
rect 34440 -3450 34520 -3430
rect 34440 -3490 34460 -3450
rect 34500 -3490 34520 -3450
rect 34440 -3510 34520 -3490
rect 34600 -3450 34680 -3430
rect 34600 -3490 34620 -3450
rect 34660 -3490 34680 -3450
rect 34600 -3510 34680 -3490
rect 34760 -3450 34840 -3430
rect 34760 -3490 34780 -3450
rect 34820 -3490 34840 -3450
rect 34760 -3510 34840 -3490
rect 34920 -3450 35000 -3430
rect 34920 -3490 34940 -3450
rect 34980 -3490 35000 -3450
rect 34920 -3510 35000 -3490
rect 35080 -3450 35160 -3430
rect 35080 -3490 35100 -3450
rect 35140 -3490 35160 -3450
rect 35080 -3510 35160 -3490
rect 35240 -3450 35320 -3430
rect 35240 -3490 35260 -3450
rect 35300 -3490 35320 -3450
rect 35240 -3510 35320 -3490
rect 35400 -3450 35480 -3430
rect 35400 -3490 35420 -3450
rect 35460 -3490 35480 -3450
rect 35400 -3510 35480 -3490
rect 35560 -3450 35640 -3430
rect 35560 -3490 35580 -3450
rect 35620 -3490 35640 -3450
rect 35560 -3510 35640 -3490
rect 35720 -3450 35800 -3430
rect 35720 -3490 35740 -3450
rect 35780 -3490 35800 -3450
rect 35720 -3510 35800 -3490
rect 35880 -3450 35960 -3430
rect 35880 -3490 35900 -3450
rect 35940 -3490 35960 -3450
rect 35880 -3510 35960 -3490
rect 36040 -3450 36120 -3430
rect 36040 -3490 36060 -3450
rect 36100 -3490 36120 -3450
rect 36040 -3510 36120 -3490
rect 36200 -3450 36280 -3430
rect 36200 -3490 36220 -3450
rect 36260 -3490 36280 -3450
rect 36200 -3510 36280 -3490
rect 36360 -3450 36440 -3430
rect 36360 -3490 36380 -3450
rect 36420 -3490 36440 -3450
rect 36360 -3510 36440 -3490
rect 36520 -3450 36600 -3430
rect 36520 -3490 36540 -3450
rect 36580 -3490 36600 -3450
rect 36520 -3510 36600 -3490
rect 36680 -3450 36760 -3430
rect 36680 -3490 36700 -3450
rect 36740 -3490 36760 -3450
rect 36680 -3510 36760 -3490
rect 36840 -3450 36920 -3430
rect 36840 -3490 36860 -3450
rect 36900 -3490 36920 -3450
rect 36840 -3510 36920 -3490
rect 37000 -3450 37080 -3430
rect 37000 -3490 37020 -3450
rect 37060 -3490 37080 -3450
rect 37000 -3510 37080 -3490
rect 37160 -3450 37240 -3430
rect 37160 -3490 37180 -3450
rect 37220 -3490 37240 -3450
rect 37160 -3510 37240 -3490
rect 37320 -3450 37400 -3430
rect 37320 -3490 37340 -3450
rect 37380 -3490 37400 -3450
rect 37320 -3510 37400 -3490
rect 37480 -3450 37560 -3430
rect 37480 -3490 37500 -3450
rect 37540 -3490 37560 -3450
rect 37480 -3510 37560 -3490
rect 37640 -3450 37720 -3430
rect 37640 -3490 37660 -3450
rect 37700 -3490 37720 -3450
rect 37640 -3510 37720 -3490
rect 35580 -3550 35620 -3510
rect 37660 -3550 37700 -3510
rect 33410 -3560 33550 -3550
rect 33330 -3570 33550 -3560
rect 33330 -3580 33420 -3570
rect 33330 -3620 33350 -3580
rect 33390 -3610 33420 -3580
rect 33460 -3610 33500 -3570
rect 33540 -3610 33550 -3570
rect 33390 -3620 33550 -3610
rect 33330 -3660 33550 -3620
rect 33330 -3700 33350 -3660
rect 33390 -3670 33550 -3660
rect 33390 -3700 33420 -3670
rect 33330 -3710 33420 -3700
rect 33460 -3710 33500 -3670
rect 33540 -3710 33550 -3670
rect 33330 -3720 33550 -3710
rect 33410 -3730 33550 -3720
rect 35570 -3570 35630 -3550
rect 35570 -3610 35580 -3570
rect 35620 -3610 35630 -3570
rect 35570 -3670 35630 -3610
rect 35570 -3710 35580 -3670
rect 35620 -3710 35630 -3670
rect 35570 -3730 35630 -3710
rect 37650 -3570 37710 -3550
rect 37650 -3610 37660 -3570
rect 37700 -3600 37710 -3570
rect 37700 -3610 37800 -3600
rect 37650 -3620 37800 -3610
rect 37650 -3660 37740 -3620
rect 37780 -3660 37800 -3620
rect 37650 -3670 37800 -3660
rect 37650 -3710 37660 -3670
rect 37700 -3680 37800 -3670
rect 37700 -3710 37710 -3680
rect 37650 -3730 37710 -3710
rect 34850 -4010 34940 -4000
rect 34850 -4060 34870 -4010
rect 34920 -4060 34940 -4010
rect 34850 -4070 34940 -4060
rect 36248 -4010 36338 -4000
rect 36248 -4060 36268 -4010
rect 36318 -4060 36338 -4010
rect 36248 -4070 36338 -4060
rect 33590 -4480 37610 -4230
rect 34880 -5590 34960 -4480
rect 36240 -5590 36320 -4480
rect 33120 -5810 33190 -5790
rect 33120 -5860 33130 -5810
rect 33180 -5860 33190 -5810
rect 33590 -5840 37610 -5590
rect 38130 -5810 38200 -5790
rect 33120 -5880 33190 -5860
rect 33310 -5950 33360 -5880
rect 32340 -6452 32410 -6430
rect 32340 -6502 32350 -6452
rect 32400 -6502 32410 -6452
rect 32340 -6522 32410 -6502
rect 33000 -6660 33070 -6640
rect 33000 -6710 33010 -6660
rect 33060 -6710 33070 -6660
rect 33000 -6730 33070 -6710
rect 34880 -6950 34960 -5840
rect 36240 -6950 36320 -5840
rect 38130 -5860 38140 -5810
rect 38190 -5860 38200 -5810
rect 38130 -5880 38200 -5860
rect 37960 -5950 38010 -5880
rect 38560 -6190 38630 -6170
rect 38560 -6240 38570 -6190
rect 38620 -6240 38630 -6190
rect 38560 -6260 38630 -6240
rect 38390 -6330 38440 -6260
rect 38680 -6240 38750 -6220
rect 38680 -6290 38690 -6240
rect 38740 -6290 38750 -6240
rect 38680 -6312 38750 -6290
rect 33590 -7200 37610 -6950
rect 32340 -7798 32410 -7778
rect 32340 -7848 32350 -7798
rect 32400 -7848 32410 -7798
rect 32340 -7868 32410 -7848
rect 33000 -7798 33070 -7778
rect 33000 -7848 33010 -7798
rect 33060 -7848 33070 -7798
rect 33000 -7868 33070 -7848
rect 33190 -7928 33240 -7858
rect 33360 -7948 33430 -7928
rect 33360 -7998 33370 -7948
rect 33420 -7998 33430 -7948
rect 33360 -8018 33430 -7998
rect 34880 -8250 34960 -7200
rect 35560 -8330 35640 -8240
rect 36240 -8250 36320 -7200
rect 38080 -7928 38130 -7858
rect 38510 -7778 38560 -7708
rect 38680 -7588 38750 -7568
rect 38680 -7638 38690 -7588
rect 38740 -7638 38750 -7588
rect 38680 -7658 38750 -7638
rect 38320 -7798 38390 -7778
rect 38320 -7848 38330 -7798
rect 38380 -7848 38390 -7798
rect 38320 -7868 38390 -7848
rect 37890 -7948 37960 -7928
rect 37890 -7998 37900 -7948
rect 37950 -7998 37960 -7948
rect 37890 -8018 37960 -7998
rect 35560 -8370 35580 -8330
rect 35620 -8370 35640 -8330
rect 35560 -8410 35640 -8370
rect 35560 -8450 35580 -8410
rect 35620 -8450 35640 -8410
rect 35560 -8490 35640 -8450
rect 35560 -8530 35580 -8490
rect 35620 -8530 35640 -8490
rect 35560 -8550 35640 -8530
<< viali >>
rect 33970 1130 34010 1170
rect 35290 1130 35330 1170
rect 35870 1130 35910 1170
rect 37190 1130 37230 1170
rect 33890 1010 33930 1050
rect 33970 1010 34010 1050
rect 33890 910 33930 950
rect 33970 910 34010 950
rect 34080 1010 34120 1050
rect 34080 910 34120 950
rect 34190 1010 34230 1050
rect 34190 910 34230 950
rect 34300 1010 34340 1050
rect 34300 910 34340 950
rect 34410 1010 34450 1050
rect 34410 910 34450 950
rect 34520 1010 34560 1050
rect 34520 910 34560 950
rect 34630 1010 34670 1050
rect 34630 910 34670 950
rect 34740 1010 34780 1050
rect 34740 910 34780 950
rect 34850 1010 34890 1050
rect 34850 910 34890 950
rect 34960 1010 35000 1050
rect 34960 910 35000 950
rect 35070 1010 35110 1050
rect 35070 910 35110 950
rect 35180 1010 35220 1050
rect 35180 910 35220 950
rect 35290 1010 35330 1050
rect 35370 1010 35410 1050
rect 35290 910 35330 950
rect 35370 910 35410 950
rect 35790 1010 35830 1050
rect 35870 1010 35910 1050
rect 35790 910 35830 950
rect 35870 910 35910 950
rect 35980 1010 36020 1050
rect 35980 910 36020 950
rect 36090 1010 36130 1050
rect 36090 910 36130 950
rect 36200 1010 36240 1050
rect 36200 910 36240 950
rect 36310 1010 36350 1050
rect 36310 910 36350 950
rect 36420 1010 36460 1050
rect 36420 910 36460 950
rect 36530 1010 36570 1050
rect 36530 910 36570 950
rect 36640 1010 36680 1050
rect 36640 910 36680 950
rect 36750 1010 36790 1050
rect 36750 910 36790 950
rect 36860 1010 36900 1050
rect 36860 910 36900 950
rect 36970 1010 37010 1050
rect 36970 910 37010 950
rect 37080 1010 37120 1050
rect 37080 910 37120 950
rect 37190 1010 37230 1050
rect 37270 1010 37310 1050
rect 37190 910 37230 950
rect 37270 910 37310 950
rect 34138 798 34172 832
rect 34248 798 34282 832
rect 34358 798 34392 832
rect 34468 798 34502 832
rect 34578 798 34612 832
rect 34688 798 34722 832
rect 34798 798 34832 832
rect 34908 798 34942 832
rect 35018 798 35052 832
rect 35128 798 35162 832
rect 36038 798 36072 832
rect 36148 798 36182 832
rect 36258 798 36292 832
rect 36368 798 36402 832
rect 36478 798 36512 832
rect 36588 798 36622 832
rect 36698 798 36732 832
rect 36808 798 36842 832
rect 36918 798 36952 832
rect 37028 798 37062 832
rect 33960 530 34000 570
rect 34320 530 34360 570
rect 34680 530 34720 570
rect 35040 530 35080 570
rect 35400 530 35440 570
rect 35760 530 35800 570
rect 36120 530 36160 570
rect 36480 530 36520 570
rect 36840 530 36880 570
rect 37200 530 37240 570
rect 33960 410 34000 450
rect 32890 330 32930 370
rect 33110 330 33150 370
rect 33330 330 33370 370
rect 33960 310 34000 350
rect 32890 210 32930 250
rect 32890 110 32930 150
rect 33000 210 33040 250
rect 33000 110 33040 150
rect 33110 210 33150 250
rect 33110 110 33150 150
rect 33220 210 33260 250
rect 33220 110 33260 150
rect 33330 210 33370 250
rect 33330 110 33370 150
rect 33960 210 34000 250
rect 33960 110 34000 150
rect 32990 -10 33030 30
rect 33110 -10 33150 30
rect 33230 -10 33270 30
rect 33960 10 34000 50
rect 33960 -90 34000 -50
rect 34140 410 34180 450
rect 34140 310 34180 350
rect 34140 210 34180 250
rect 34140 110 34180 150
rect 34140 10 34180 50
rect 34140 -90 34180 -50
rect 34320 410 34360 450
rect 34320 310 34360 350
rect 34320 210 34360 250
rect 34320 110 34360 150
rect 34320 10 34360 50
rect 34320 -90 34360 -50
rect 34500 410 34540 450
rect 34500 310 34540 350
rect 34500 210 34540 250
rect 34500 110 34540 150
rect 34500 10 34540 50
rect 34500 -90 34540 -50
rect 34680 410 34720 450
rect 34680 310 34720 350
rect 34680 210 34720 250
rect 34680 110 34720 150
rect 34680 10 34720 50
rect 34680 -90 34720 -50
rect 34860 410 34900 450
rect 34860 310 34900 350
rect 34860 210 34900 250
rect 34860 110 34900 150
rect 34860 10 34900 50
rect 34860 -90 34900 -50
rect 35040 410 35080 450
rect 35040 310 35080 350
rect 35040 210 35080 250
rect 35040 110 35080 150
rect 35040 10 35080 50
rect 35040 -90 35080 -50
rect 35220 410 35260 450
rect 35220 310 35260 350
rect 35220 210 35260 250
rect 35220 110 35260 150
rect 35220 10 35260 50
rect 35220 -90 35260 -50
rect 35400 410 35440 450
rect 35400 310 35440 350
rect 35400 210 35440 250
rect 35400 110 35440 150
rect 35400 10 35440 50
rect 35400 -90 35440 -50
rect 35580 410 35620 450
rect 35580 310 35620 350
rect 35580 210 35620 250
rect 35580 110 35620 150
rect 35580 10 35620 50
rect 35580 -90 35620 -50
rect 35760 410 35800 450
rect 35760 310 35800 350
rect 35760 210 35800 250
rect 35760 110 35800 150
rect 35760 10 35800 50
rect 35760 -90 35800 -50
rect 35940 410 35980 450
rect 35940 310 35980 350
rect 35940 210 35980 250
rect 35940 110 35980 150
rect 35940 10 35980 50
rect 35940 -90 35980 -50
rect 36120 410 36160 450
rect 36120 310 36160 350
rect 36120 210 36160 250
rect 36120 110 36160 150
rect 36120 10 36160 50
rect 36120 -90 36160 -50
rect 36300 410 36340 450
rect 36300 310 36340 350
rect 36300 210 36340 250
rect 36300 110 36340 150
rect 36300 10 36340 50
rect 36300 -90 36340 -50
rect 36480 410 36520 450
rect 36480 310 36520 350
rect 36480 210 36520 250
rect 36480 110 36520 150
rect 36480 10 36520 50
rect 36480 -90 36520 -50
rect 36660 410 36700 450
rect 36660 310 36700 350
rect 36660 210 36700 250
rect 36660 110 36700 150
rect 36660 10 36700 50
rect 36660 -90 36700 -50
rect 36840 410 36880 450
rect 36840 310 36880 350
rect 36840 210 36880 250
rect 36840 110 36880 150
rect 36840 10 36880 50
rect 36840 -90 36880 -50
rect 37020 410 37060 450
rect 37020 310 37060 350
rect 37020 210 37060 250
rect 37020 110 37060 150
rect 37020 10 37060 50
rect 37020 -90 37060 -50
rect 37200 410 37240 450
rect 37200 310 37240 350
rect 37200 210 37240 250
rect 37200 110 37240 150
rect 37200 10 37240 50
rect 37200 -90 37240 -50
rect 34230 -210 34270 -170
rect 34410 -210 34450 -170
rect 34590 -210 34630 -170
rect 34770 -210 34810 -170
rect 34950 -210 34990 -170
rect 35130 -210 35170 -170
rect 35310 -210 35350 -170
rect 35490 -210 35530 -170
rect 35670 -210 35710 -170
rect 35850 -210 35890 -170
rect 36030 -210 36070 -170
rect 36210 -210 36250 -170
rect 36390 -210 36430 -170
rect 36570 -210 36610 -170
rect 36750 -210 36790 -170
rect 36930 -210 36970 -170
rect 32860 -1030 32900 -990
rect 35260 -1030 35300 -990
rect 35900 -1030 35940 -990
rect 38300 -1030 38340 -990
rect 32860 -1150 32900 -1110
rect 32860 -1250 32900 -1210
rect 32980 -1150 33020 -1110
rect 32980 -1250 33020 -1210
rect 33100 -1150 33140 -1110
rect 33100 -1250 33140 -1210
rect 33220 -1150 33260 -1110
rect 33220 -1250 33260 -1210
rect 33340 -1150 33380 -1110
rect 33340 -1250 33380 -1210
rect 33460 -1150 33500 -1110
rect 33460 -1250 33500 -1210
rect 33580 -1150 33620 -1110
rect 33580 -1250 33620 -1210
rect 33700 -1150 33740 -1110
rect 33700 -1250 33740 -1210
rect 33820 -1150 33860 -1110
rect 33820 -1250 33860 -1210
rect 33940 -1150 33980 -1110
rect 33940 -1250 33980 -1210
rect 34060 -1150 34100 -1110
rect 34060 -1250 34100 -1210
rect 34180 -1150 34220 -1110
rect 34180 -1250 34220 -1210
rect 34300 -1150 34340 -1110
rect 34300 -1250 34340 -1210
rect 34420 -1150 34460 -1110
rect 34420 -1250 34460 -1210
rect 34540 -1150 34580 -1110
rect 34540 -1250 34580 -1210
rect 34660 -1150 34700 -1110
rect 34660 -1250 34700 -1210
rect 34780 -1150 34820 -1110
rect 34780 -1250 34820 -1210
rect 34900 -1150 34940 -1110
rect 34900 -1250 34940 -1210
rect 35020 -1150 35060 -1110
rect 35020 -1250 35060 -1210
rect 35140 -1150 35180 -1110
rect 35140 -1250 35180 -1210
rect 35260 -1150 35300 -1110
rect 35260 -1250 35300 -1210
rect 35900 -1150 35940 -1110
rect 35900 -1250 35940 -1210
rect 36020 -1150 36060 -1110
rect 36020 -1250 36060 -1210
rect 36140 -1150 36180 -1110
rect 36140 -1250 36180 -1210
rect 36260 -1150 36300 -1110
rect 36260 -1250 36300 -1210
rect 36380 -1150 36420 -1110
rect 36380 -1250 36420 -1210
rect 36500 -1150 36540 -1110
rect 36500 -1250 36540 -1210
rect 36620 -1150 36660 -1110
rect 36620 -1250 36660 -1210
rect 36740 -1150 36780 -1110
rect 36740 -1250 36780 -1210
rect 36860 -1150 36900 -1110
rect 36860 -1250 36900 -1210
rect 36980 -1150 37020 -1110
rect 36980 -1250 37020 -1210
rect 37100 -1150 37140 -1110
rect 37100 -1250 37140 -1210
rect 37220 -1150 37260 -1110
rect 37220 -1250 37260 -1210
rect 37340 -1150 37380 -1110
rect 37340 -1250 37380 -1210
rect 37460 -1150 37500 -1110
rect 37460 -1250 37500 -1210
rect 37580 -1150 37620 -1110
rect 37580 -1250 37620 -1210
rect 37700 -1150 37740 -1110
rect 37700 -1250 37740 -1210
rect 37820 -1150 37860 -1110
rect 37820 -1250 37860 -1210
rect 37940 -1150 37980 -1110
rect 37940 -1250 37980 -1210
rect 38060 -1150 38100 -1110
rect 38060 -1250 38100 -1210
rect 38180 -1150 38220 -1110
rect 38180 -1250 38220 -1210
rect 38300 -1150 38340 -1110
rect 38300 -1250 38340 -1210
rect 33040 -1380 33080 -1340
rect 33220 -1370 33260 -1330
rect 33700 -1370 33740 -1330
rect 33940 -1370 33980 -1330
rect 34420 -1370 34460 -1330
rect 34660 -1370 34700 -1330
rect 35080 -1370 35120 -1330
rect 36080 -1370 36120 -1330
rect 36500 -1370 36540 -1330
rect 36740 -1370 36780 -1330
rect 37220 -1370 37260 -1330
rect 37460 -1370 37500 -1330
rect 37940 -1370 37980 -1330
rect 38120 -1380 38160 -1340
rect 33864 -1972 33898 -1938
rect 34022 -1972 34056 -1938
rect 34346 -1972 34380 -1938
rect 34500 -1972 34534 -1938
rect 34824 -1972 34858 -1938
rect 35140 -2020 35180 -1980
rect 33700 -2090 33740 -2050
rect 33820 -2090 33860 -2050
rect 33940 -2090 33980 -2050
rect 34060 -2090 34100 -2050
rect 34180 -2090 34220 -2050
rect 34300 -2090 34340 -2050
rect 34420 -2090 34460 -2050
rect 34540 -2090 34580 -2050
rect 34660 -2090 34700 -2050
rect 34780 -2090 34820 -2050
rect 34900 -2090 34940 -2050
rect 35140 -2100 35180 -2060
rect 33763 -2202 33797 -2168
rect 34123 -2202 34157 -2168
rect 34243 -2202 34277 -2168
rect 34603 -2202 34637 -2168
rect 34723 -2202 34757 -2168
rect 35140 -2180 35180 -2140
rect 36020 -2020 36060 -1980
rect 36342 -1972 36376 -1938
rect 36666 -1972 36700 -1938
rect 36820 -1972 36854 -1938
rect 37144 -1972 37178 -1938
rect 37302 -1972 37336 -1938
rect 36020 -2100 36060 -2060
rect 36260 -2090 36300 -2050
rect 36380 -2090 36420 -2050
rect 36500 -2090 36540 -2050
rect 36620 -2090 36660 -2050
rect 36740 -2090 36780 -2050
rect 36860 -2090 36900 -2050
rect 36980 -2090 37020 -2050
rect 37100 -2090 37140 -2050
rect 37220 -2090 37260 -2050
rect 37340 -2090 37380 -2050
rect 37460 -2090 37500 -2050
rect 36020 -2180 36060 -2140
rect 36443 -2202 36477 -2168
rect 36563 -2202 36597 -2168
rect 36923 -2202 36957 -2168
rect 37043 -2202 37077 -2168
rect 37403 -2202 37437 -2168
rect 33260 -2580 33300 -2540
rect 33500 -2580 33540 -2540
rect 33740 -2580 33780 -2540
rect 33980 -2580 34020 -2540
rect 34620 -2580 34660 -2540
rect 34860 -2580 34900 -2540
rect 35100 -2580 35140 -2540
rect 35400 -2610 35440 -2570
rect 33080 -2700 33120 -2660
rect 33080 -2800 33120 -2760
rect 33080 -2900 33120 -2860
rect 33080 -3000 33120 -2960
rect 33080 -3100 33120 -3060
rect 35760 -2610 35800 -2570
rect 36060 -2580 36100 -2540
rect 36300 -2580 36340 -2540
rect 36540 -2580 36580 -2540
rect 37180 -2580 37220 -2540
rect 37420 -2580 37460 -2540
rect 37660 -2580 37700 -2540
rect 37900 -2580 37940 -2540
rect 38080 -2620 38120 -2580
rect 34240 -3220 34280 -3180
rect 36920 -3220 36960 -3180
rect 33660 -3490 33700 -3450
rect 33820 -3490 33860 -3450
rect 33980 -3490 34020 -3450
rect 34140 -3490 34180 -3450
rect 34300 -3490 34340 -3450
rect 34460 -3490 34500 -3450
rect 34620 -3490 34660 -3450
rect 34780 -3490 34820 -3450
rect 34940 -3490 34980 -3450
rect 35100 -3490 35140 -3450
rect 35260 -3490 35300 -3450
rect 35420 -3490 35460 -3450
rect 35580 -3490 35620 -3450
rect 35740 -3490 35780 -3450
rect 35900 -3490 35940 -3450
rect 36060 -3490 36100 -3450
rect 36220 -3490 36260 -3450
rect 36380 -3490 36420 -3450
rect 36540 -3490 36580 -3450
rect 36700 -3490 36740 -3450
rect 36860 -3490 36900 -3450
rect 37020 -3490 37060 -3450
rect 37180 -3490 37220 -3450
rect 37340 -3490 37380 -3450
rect 37500 -3490 37540 -3450
rect 37660 -3490 37700 -3450
rect 33350 -3620 33390 -3580
rect 33350 -3700 33390 -3660
rect 37740 -3660 37780 -3620
rect 34870 -4060 34920 -4010
rect 36268 -4060 36318 -4010
rect 33130 -5860 33180 -5810
rect 32350 -6502 32400 -6452
rect 33010 -6710 33060 -6660
rect 38140 -5860 38190 -5810
rect 38570 -6240 38620 -6190
rect 38690 -6290 38740 -6240
rect 32350 -7848 32400 -7798
rect 33010 -7848 33060 -7798
rect 33370 -7998 33420 -7948
rect 38690 -7638 38740 -7588
rect 38330 -7848 38380 -7798
rect 37900 -7998 37950 -7948
rect 35580 -8370 35620 -8330
rect 35580 -8450 35620 -8410
rect 35580 -8530 35620 -8490
<< metal1 >>
rect 34060 1290 34140 1300
rect 34060 1230 34070 1290
rect 34130 1230 34140 1290
rect 34060 1220 34140 1230
rect 34280 1290 34360 1300
rect 34280 1230 34290 1290
rect 34350 1230 34360 1290
rect 34280 1220 34360 1230
rect 34500 1290 34580 1300
rect 34500 1230 34510 1290
rect 34570 1230 34580 1290
rect 34500 1220 34580 1230
rect 34720 1290 34800 1300
rect 34720 1230 34730 1290
rect 34790 1230 34800 1290
rect 34720 1220 34800 1230
rect 34940 1290 35020 1300
rect 34940 1230 34950 1290
rect 35010 1230 35020 1290
rect 34940 1220 35020 1230
rect 35160 1290 35240 1300
rect 35160 1230 35170 1290
rect 35230 1230 35240 1290
rect 35160 1220 35240 1230
rect 35960 1290 36040 1300
rect 35960 1230 35970 1290
rect 36030 1230 36040 1290
rect 35960 1220 36040 1230
rect 36180 1290 36260 1300
rect 36180 1230 36190 1290
rect 36250 1230 36260 1290
rect 36180 1220 36260 1230
rect 36400 1290 36480 1300
rect 36400 1230 36410 1290
rect 36470 1230 36480 1290
rect 36400 1220 36480 1230
rect 36620 1290 36700 1300
rect 36620 1230 36630 1290
rect 36690 1230 36700 1290
rect 36620 1220 36700 1230
rect 36840 1290 36920 1300
rect 36840 1230 36850 1290
rect 36910 1230 36920 1290
rect 36840 1220 36920 1230
rect 37060 1290 37140 1300
rect 37060 1230 37070 1290
rect 37130 1230 37140 1290
rect 37060 1220 37140 1230
rect 38450 1290 38530 1300
rect 38450 1230 38460 1290
rect 38520 1230 38530 1290
rect 33950 1180 34030 1190
rect 33950 1120 33960 1180
rect 34020 1120 34030 1180
rect 33950 1110 34030 1120
rect 33960 1070 34020 1110
rect 33880 1050 34020 1070
rect 33880 1010 33890 1050
rect 33930 1010 33970 1050
rect 34010 1010 34020 1050
rect 33880 950 34020 1010
rect 33880 910 33890 950
rect 33930 910 33970 950
rect 34010 910 34020 950
rect 33880 890 34020 910
rect 34070 1050 34130 1220
rect 34170 1180 34250 1190
rect 34170 1120 34180 1180
rect 34240 1120 34250 1180
rect 34170 1110 34250 1120
rect 34070 1010 34080 1050
rect 34120 1010 34130 1050
rect 34070 950 34130 1010
rect 34070 910 34080 950
rect 34120 910 34130 950
rect 34070 890 34130 910
rect 34180 1050 34240 1110
rect 34180 1010 34190 1050
rect 34230 1010 34240 1050
rect 34180 950 34240 1010
rect 34180 910 34190 950
rect 34230 910 34240 950
rect 34180 890 34240 910
rect 34290 1050 34350 1220
rect 34390 1180 34470 1190
rect 34390 1120 34400 1180
rect 34460 1120 34470 1180
rect 34390 1110 34470 1120
rect 34290 1010 34300 1050
rect 34340 1010 34350 1050
rect 34290 950 34350 1010
rect 34290 910 34300 950
rect 34340 910 34350 950
rect 34290 890 34350 910
rect 34400 1050 34460 1110
rect 34400 1010 34410 1050
rect 34450 1010 34460 1050
rect 34400 950 34460 1010
rect 34400 910 34410 950
rect 34450 910 34460 950
rect 34400 890 34460 910
rect 34510 1050 34570 1220
rect 34610 1180 34690 1190
rect 34610 1120 34620 1180
rect 34680 1120 34690 1180
rect 34610 1110 34690 1120
rect 34510 1010 34520 1050
rect 34560 1010 34570 1050
rect 34510 950 34570 1010
rect 34510 910 34520 950
rect 34560 910 34570 950
rect 34510 890 34570 910
rect 34620 1050 34680 1110
rect 34620 1010 34630 1050
rect 34670 1010 34680 1050
rect 34620 950 34680 1010
rect 34620 910 34630 950
rect 34670 910 34680 950
rect 34620 890 34680 910
rect 34730 1050 34790 1220
rect 34830 1180 34910 1190
rect 34830 1120 34840 1180
rect 34900 1120 34910 1180
rect 34830 1110 34910 1120
rect 34730 1010 34740 1050
rect 34780 1010 34790 1050
rect 34730 950 34790 1010
rect 34730 910 34740 950
rect 34780 910 34790 950
rect 34730 890 34790 910
rect 34840 1050 34900 1110
rect 34840 1010 34850 1050
rect 34890 1010 34900 1050
rect 34840 950 34900 1010
rect 34840 910 34850 950
rect 34890 910 34900 950
rect 34840 890 34900 910
rect 34950 1050 35010 1220
rect 35050 1180 35130 1190
rect 35050 1120 35060 1180
rect 35120 1120 35130 1180
rect 35050 1110 35130 1120
rect 34950 1010 34960 1050
rect 35000 1010 35010 1050
rect 34950 950 35010 1010
rect 34950 910 34960 950
rect 35000 910 35010 950
rect 34950 890 35010 910
rect 35060 1050 35120 1110
rect 35060 1010 35070 1050
rect 35110 1010 35120 1050
rect 35060 950 35120 1010
rect 35060 910 35070 950
rect 35110 910 35120 950
rect 35060 890 35120 910
rect 35170 1050 35230 1220
rect 35270 1180 35350 1190
rect 35270 1120 35280 1180
rect 35340 1120 35350 1180
rect 35270 1110 35350 1120
rect 35850 1180 35930 1190
rect 35850 1120 35860 1180
rect 35920 1120 35930 1180
rect 35850 1110 35930 1120
rect 35170 1010 35180 1050
rect 35220 1010 35230 1050
rect 35170 950 35230 1010
rect 35170 910 35180 950
rect 35220 910 35230 950
rect 35170 890 35230 910
rect 35280 1070 35340 1110
rect 35860 1070 35920 1110
rect 35280 1050 35420 1070
rect 35280 1010 35290 1050
rect 35330 1010 35370 1050
rect 35410 1010 35420 1050
rect 35280 950 35420 1010
rect 35280 910 35290 950
rect 35330 910 35370 950
rect 35410 910 35420 950
rect 35280 890 35420 910
rect 35780 1050 35920 1070
rect 35780 1010 35790 1050
rect 35830 1010 35870 1050
rect 35910 1010 35920 1050
rect 35780 950 35920 1010
rect 35780 910 35790 950
rect 35830 910 35870 950
rect 35910 910 35920 950
rect 35780 890 35920 910
rect 35970 1050 36030 1220
rect 36070 1180 36150 1190
rect 36070 1120 36080 1180
rect 36140 1120 36150 1180
rect 36070 1110 36150 1120
rect 35970 1010 35980 1050
rect 36020 1010 36030 1050
rect 35970 950 36030 1010
rect 35970 910 35980 950
rect 36020 910 36030 950
rect 35970 890 36030 910
rect 36080 1050 36140 1110
rect 36080 1010 36090 1050
rect 36130 1010 36140 1050
rect 36080 950 36140 1010
rect 36080 910 36090 950
rect 36130 910 36140 950
rect 36080 890 36140 910
rect 36190 1050 36250 1220
rect 36290 1180 36370 1190
rect 36290 1120 36300 1180
rect 36360 1120 36370 1180
rect 36290 1110 36370 1120
rect 36190 1010 36200 1050
rect 36240 1010 36250 1050
rect 36190 950 36250 1010
rect 36190 910 36200 950
rect 36240 910 36250 950
rect 36190 890 36250 910
rect 36300 1050 36360 1110
rect 36300 1010 36310 1050
rect 36350 1010 36360 1050
rect 36300 950 36360 1010
rect 36300 910 36310 950
rect 36350 910 36360 950
rect 36300 890 36360 910
rect 36410 1050 36470 1220
rect 36510 1180 36590 1190
rect 36510 1120 36520 1180
rect 36580 1120 36590 1180
rect 36510 1110 36590 1120
rect 36410 1010 36420 1050
rect 36460 1010 36470 1050
rect 36410 950 36470 1010
rect 36410 910 36420 950
rect 36460 910 36470 950
rect 36410 890 36470 910
rect 36520 1050 36580 1110
rect 36520 1010 36530 1050
rect 36570 1010 36580 1050
rect 36520 950 36580 1010
rect 36520 910 36530 950
rect 36570 910 36580 950
rect 36520 890 36580 910
rect 36630 1050 36690 1220
rect 36730 1180 36810 1190
rect 36730 1120 36740 1180
rect 36800 1120 36810 1180
rect 36730 1110 36810 1120
rect 36630 1010 36640 1050
rect 36680 1010 36690 1050
rect 36630 950 36690 1010
rect 36630 910 36640 950
rect 36680 910 36690 950
rect 36630 890 36690 910
rect 36740 1050 36800 1110
rect 36740 1010 36750 1050
rect 36790 1010 36800 1050
rect 36740 950 36800 1010
rect 36740 910 36750 950
rect 36790 910 36800 950
rect 36740 890 36800 910
rect 36850 1050 36910 1220
rect 36950 1180 37030 1190
rect 36950 1120 36960 1180
rect 37020 1120 37030 1180
rect 36950 1110 37030 1120
rect 36850 1010 36860 1050
rect 36900 1010 36910 1050
rect 36850 950 36910 1010
rect 36850 910 36860 950
rect 36900 910 36910 950
rect 36850 890 36910 910
rect 36960 1050 37020 1110
rect 36960 1010 36970 1050
rect 37010 1010 37020 1050
rect 36960 950 37020 1010
rect 36960 910 36970 950
rect 37010 910 37020 950
rect 36960 890 37020 910
rect 37070 1050 37130 1220
rect 37170 1180 37250 1190
rect 37170 1120 37180 1180
rect 37240 1120 37250 1180
rect 37170 1110 37250 1120
rect 37070 1010 37080 1050
rect 37120 1010 37130 1050
rect 37070 950 37130 1010
rect 37070 910 37080 950
rect 37120 910 37130 950
rect 37070 890 37130 910
rect 37180 1070 37240 1110
rect 37180 1050 37320 1070
rect 37180 1010 37190 1050
rect 37230 1010 37270 1050
rect 37310 1010 37320 1050
rect 37180 950 37320 1010
rect 37180 910 37190 950
rect 37230 910 37270 950
rect 37310 910 37320 950
rect 37180 890 37320 910
rect 34126 842 34184 850
rect 34126 790 34130 842
rect 34182 790 34184 842
rect 34126 780 34184 790
rect 34236 842 34294 850
rect 34236 790 34240 842
rect 34292 790 34294 842
rect 34236 780 34294 790
rect 34346 842 34404 850
rect 34346 790 34350 842
rect 34402 790 34404 842
rect 34346 780 34404 790
rect 34456 842 34514 850
rect 34456 790 34460 842
rect 34512 790 34514 842
rect 34456 780 34514 790
rect 34566 842 34624 850
rect 34566 790 34570 842
rect 34622 790 34624 842
rect 34566 780 34624 790
rect 34676 842 34734 850
rect 34676 790 34680 842
rect 34732 790 34734 842
rect 34676 780 34734 790
rect 34786 842 34844 850
rect 34786 790 34790 842
rect 34842 790 34844 842
rect 34786 780 34844 790
rect 34896 842 34954 850
rect 34896 790 34900 842
rect 34952 790 34954 842
rect 34896 780 34954 790
rect 35006 842 35064 850
rect 35006 790 35010 842
rect 35062 790 35064 842
rect 35006 780 35064 790
rect 35116 842 35174 850
rect 35116 790 35120 842
rect 35172 790 35174 842
rect 35116 780 35174 790
rect 36026 842 36084 850
rect 36026 790 36030 842
rect 36082 790 36084 842
rect 36026 780 36084 790
rect 36136 842 36194 850
rect 36136 790 36140 842
rect 36192 790 36194 842
rect 36136 780 36194 790
rect 36246 842 36304 850
rect 36246 790 36250 842
rect 36302 790 36304 842
rect 36246 780 36304 790
rect 36356 842 36414 850
rect 36356 790 36360 842
rect 36412 790 36414 842
rect 36356 780 36414 790
rect 36466 842 36524 850
rect 36466 790 36470 842
rect 36522 790 36524 842
rect 36466 780 36524 790
rect 36576 842 36634 850
rect 36576 790 36580 842
rect 36632 790 36634 842
rect 36576 780 36634 790
rect 36686 842 36744 850
rect 36686 790 36690 842
rect 36742 790 36744 842
rect 36686 780 36744 790
rect 36796 842 36854 850
rect 36796 790 36800 842
rect 36852 790 36854 842
rect 36796 780 36854 790
rect 36906 842 36964 850
rect 36906 790 36910 842
rect 36962 790 36964 842
rect 36906 780 36964 790
rect 37016 842 37074 850
rect 37016 790 37020 842
rect 37072 790 37074 842
rect 37016 780 37074 790
rect 32870 740 32950 750
rect 32870 680 32880 740
rect 32940 680 32950 740
rect 32870 660 32950 680
rect 32870 600 32880 660
rect 32940 600 32950 660
rect 32870 580 32950 600
rect 32870 520 32880 580
rect 32940 520 32950 580
rect 32870 510 32950 520
rect 33310 740 33390 750
rect 33310 680 33320 740
rect 33380 680 33390 740
rect 33310 660 33390 680
rect 33310 600 33320 660
rect 33380 600 33390 660
rect 33310 580 33390 600
rect 33310 520 33320 580
rect 33380 520 33390 580
rect 33310 510 33390 520
rect 33940 740 34020 750
rect 33940 680 33950 740
rect 34010 680 34020 740
rect 33940 660 34020 680
rect 33940 600 33950 660
rect 34010 600 34020 660
rect 33940 580 34020 600
rect 33940 520 33950 580
rect 34010 520 34020 580
rect 33940 510 34020 520
rect 34300 740 34380 750
rect 34300 680 34310 740
rect 34370 680 34380 740
rect 34300 660 34380 680
rect 34300 600 34310 660
rect 34370 600 34380 660
rect 34300 580 34380 600
rect 34300 520 34310 580
rect 34370 520 34380 580
rect 34300 510 34380 520
rect 34660 740 34740 750
rect 34660 680 34670 740
rect 34730 680 34740 740
rect 34660 660 34740 680
rect 34660 600 34670 660
rect 34730 600 34740 660
rect 34660 580 34740 600
rect 34660 520 34670 580
rect 34730 520 34740 580
rect 34660 510 34740 520
rect 35020 740 35100 750
rect 35020 680 35030 740
rect 35090 680 35100 740
rect 35020 660 35100 680
rect 35020 600 35030 660
rect 35090 600 35100 660
rect 35020 580 35100 600
rect 35020 520 35030 580
rect 35090 520 35100 580
rect 35020 510 35100 520
rect 35380 740 35460 750
rect 35380 680 35390 740
rect 35450 680 35460 740
rect 35380 660 35460 680
rect 35380 600 35390 660
rect 35450 600 35460 660
rect 35380 580 35460 600
rect 35380 520 35390 580
rect 35450 520 35460 580
rect 35380 510 35460 520
rect 35740 740 35820 750
rect 35740 680 35750 740
rect 35810 680 35820 740
rect 35740 660 35820 680
rect 35740 600 35750 660
rect 35810 600 35820 660
rect 35740 580 35820 600
rect 35740 520 35750 580
rect 35810 520 35820 580
rect 35740 510 35820 520
rect 36100 740 36180 750
rect 36100 680 36110 740
rect 36170 680 36180 740
rect 36100 660 36180 680
rect 36100 600 36110 660
rect 36170 600 36180 660
rect 36100 580 36180 600
rect 36100 520 36110 580
rect 36170 520 36180 580
rect 36100 510 36180 520
rect 36460 740 36540 750
rect 36460 680 36470 740
rect 36530 680 36540 740
rect 36460 660 36540 680
rect 36460 600 36470 660
rect 36530 600 36540 660
rect 36460 580 36540 600
rect 36460 520 36470 580
rect 36530 520 36540 580
rect 36460 510 36540 520
rect 36820 740 36900 750
rect 36820 680 36830 740
rect 36890 680 36900 740
rect 36820 660 36900 680
rect 36820 600 36830 660
rect 36890 600 36900 660
rect 36820 580 36900 600
rect 36820 520 36830 580
rect 36890 520 36900 580
rect 36820 510 36900 520
rect 37180 740 37260 750
rect 37180 680 37190 740
rect 37250 680 37260 740
rect 37180 660 37260 680
rect 37180 600 37190 660
rect 37250 600 37260 660
rect 37180 580 37260 600
rect 37180 520 37190 580
rect 37250 520 37260 580
rect 37180 510 37260 520
rect 32880 390 32940 510
rect 33320 390 33380 510
rect 33950 450 34010 470
rect 33950 410 33960 450
rect 34000 410 34010 450
rect 32870 370 32950 390
rect 32870 330 32890 370
rect 32930 330 32950 370
rect 32870 310 32950 330
rect 33090 380 33170 390
rect 33090 320 33100 380
rect 33160 320 33170 380
rect 33090 310 33170 320
rect 33310 370 33390 390
rect 33310 330 33330 370
rect 33370 330 33390 370
rect 33310 310 33390 330
rect 33560 380 33640 390
rect 33560 320 33570 380
rect 33630 320 33640 380
rect 33560 310 33640 320
rect 33950 350 34010 410
rect 33950 310 33960 350
rect 34000 310 34010 350
rect 32880 250 32940 310
rect 32880 210 32890 250
rect 32930 210 32940 250
rect 32880 150 32940 210
rect 32880 110 32890 150
rect 32930 110 32940 150
rect 32880 90 32940 110
rect 32990 250 33050 270
rect 32990 210 33000 250
rect 33040 210 33050 250
rect 32990 150 33050 210
rect 32990 110 33000 150
rect 33040 110 33050 150
rect 32990 50 33050 110
rect 33100 250 33160 310
rect 33100 210 33110 250
rect 33150 210 33160 250
rect 33100 150 33160 210
rect 33100 110 33110 150
rect 33150 110 33160 150
rect 33100 90 33160 110
rect 33210 250 33270 270
rect 33210 210 33220 250
rect 33260 210 33270 250
rect 33210 150 33270 210
rect 33210 110 33220 150
rect 33260 110 33270 150
rect 33210 50 33270 110
rect 33320 250 33380 310
rect 33320 210 33330 250
rect 33370 210 33380 250
rect 33320 150 33380 210
rect 33320 110 33330 150
rect 33370 110 33380 150
rect 33320 90 33380 110
rect 32970 40 33050 50
rect 32970 -20 32980 40
rect 33040 -20 33050 40
rect 32970 -30 33050 -20
rect 33090 30 33170 50
rect 33090 -10 33110 30
rect 33150 -10 33170 30
rect 32650 -270 32730 -260
rect 32650 -330 32660 -270
rect 32720 -330 32730 -270
rect 32650 -340 32730 -330
rect 32560 -380 32640 -370
rect 32560 -440 32570 -380
rect 32630 -440 32640 -380
rect 32560 -450 32640 -440
rect 32330 -980 32410 -970
rect 32330 -1040 32340 -980
rect 32400 -1040 32410 -980
rect 32060 -1440 32300 -1430
rect 32060 -1500 32070 -1440
rect 32130 -1500 32150 -1440
rect 32210 -1500 32230 -1440
rect 32290 -1500 32300 -1440
rect 32060 -1520 32300 -1500
rect 32060 -1580 32070 -1520
rect 32130 -1580 32150 -1520
rect 32210 -1580 32230 -1520
rect 32290 -1580 32300 -1520
rect 32060 -1600 32300 -1580
rect 32060 -1660 32070 -1600
rect 32130 -1660 32150 -1600
rect 32210 -1660 32230 -1600
rect 32290 -1660 32300 -1600
rect 31830 -3780 31910 -3770
rect 31830 -3840 31840 -3780
rect 31900 -3840 31910 -3780
rect 31700 -4750 31800 -4730
rect 31700 -4810 31720 -4750
rect 31780 -4810 31800 -4750
rect 31700 -4830 31800 -4810
rect 31700 -6150 31800 -6130
rect 31700 -6210 31720 -6150
rect 31780 -6210 31800 -6150
rect 31700 -6230 31800 -6210
rect 31580 -6850 31660 -6840
rect 31580 -6910 31590 -6850
rect 31650 -6910 31660 -6850
rect 31580 -6920 31660 -6910
rect 31830 -7530 31910 -3840
rect 32060 -4750 32300 -1660
rect 32060 -4810 32070 -4750
rect 32130 -4810 32150 -4750
rect 32210 -4810 32230 -4750
rect 32290 -4810 32300 -4750
rect 32060 -4830 32300 -4810
rect 31950 -5450 32030 -5440
rect 31950 -5510 31960 -5450
rect 32020 -5510 32030 -5450
rect 31820 -7550 31920 -7530
rect 31820 -7610 31840 -7550
rect 31900 -7610 31920 -7550
rect 31820 -7630 31920 -7610
rect 31950 -7780 32030 -5510
rect 32330 -6150 32410 -1040
rect 32580 -1910 32620 -450
rect 32560 -1920 32640 -1910
rect 32560 -1980 32570 -1920
rect 32630 -1980 32640 -1920
rect 32560 -1990 32640 -1980
rect 32580 -4190 32620 -1990
rect 32670 -2140 32710 -340
rect 32840 -710 32920 -700
rect 32840 -770 32850 -710
rect 32910 -770 32920 -710
rect 32840 -790 32920 -770
rect 32840 -850 32850 -790
rect 32910 -850 32920 -790
rect 32840 -870 32920 -850
rect 32840 -930 32850 -870
rect 32910 -930 32920 -870
rect 32840 -940 32920 -930
rect 32850 -990 32910 -940
rect 32850 -1030 32860 -990
rect 32900 -1030 32910 -990
rect 32850 -1110 32910 -1030
rect 32960 -980 33040 -30
rect 33090 -490 33170 -10
rect 33210 40 33290 50
rect 33210 -20 33220 40
rect 33280 -20 33290 40
rect 33210 -30 33290 -20
rect 33580 -370 33620 310
rect 33950 250 34010 310
rect 33950 210 33960 250
rect 34000 210 34010 250
rect 33950 150 34010 210
rect 33950 110 33960 150
rect 34000 110 34010 150
rect 33950 50 34010 110
rect 33950 10 33960 50
rect 34000 10 34010 50
rect 33950 -50 34010 10
rect 33950 -90 33960 -50
rect 34000 -90 34010 -50
rect 33950 -110 34010 -90
rect 34130 450 34190 470
rect 34130 410 34140 450
rect 34180 410 34190 450
rect 34130 350 34190 410
rect 34130 310 34140 350
rect 34180 310 34190 350
rect 34130 250 34190 310
rect 34130 210 34140 250
rect 34180 210 34190 250
rect 34130 150 34190 210
rect 34130 110 34140 150
rect 34180 110 34190 150
rect 34130 50 34190 110
rect 34130 10 34140 50
rect 34180 10 34190 50
rect 34130 -50 34190 10
rect 34130 -90 34140 -50
rect 34180 -90 34190 -50
rect 33560 -380 33640 -370
rect 33560 -440 33570 -380
rect 33630 -440 33640 -380
rect 33560 -450 33640 -440
rect 33090 -550 33100 -490
rect 33160 -550 33170 -490
rect 33090 -560 33170 -550
rect 34130 -590 34190 -90
rect 34310 450 34370 470
rect 34310 410 34320 450
rect 34360 410 34370 450
rect 34310 350 34370 410
rect 34310 310 34320 350
rect 34360 310 34370 350
rect 34310 250 34370 310
rect 34310 210 34320 250
rect 34360 210 34370 250
rect 34310 150 34370 210
rect 34310 110 34320 150
rect 34360 110 34370 150
rect 34310 50 34370 110
rect 34310 10 34320 50
rect 34360 10 34370 50
rect 34310 -50 34370 10
rect 34310 -90 34320 -50
rect 34360 -90 34370 -50
rect 34310 -110 34370 -90
rect 34490 450 34550 470
rect 34490 410 34500 450
rect 34540 410 34550 450
rect 34490 350 34550 410
rect 34490 310 34500 350
rect 34540 310 34550 350
rect 34490 250 34550 310
rect 34490 210 34500 250
rect 34540 210 34550 250
rect 34490 150 34550 210
rect 34490 110 34500 150
rect 34540 110 34550 150
rect 34490 50 34550 110
rect 34490 10 34500 50
rect 34540 10 34550 50
rect 34490 -50 34550 10
rect 34490 -90 34500 -50
rect 34540 -90 34550 -50
rect 34490 -110 34550 -90
rect 34670 450 34730 470
rect 34670 410 34680 450
rect 34720 410 34730 450
rect 34670 350 34730 410
rect 34670 310 34680 350
rect 34720 310 34730 350
rect 34670 250 34730 310
rect 34670 210 34680 250
rect 34720 210 34730 250
rect 34670 150 34730 210
rect 34670 110 34680 150
rect 34720 110 34730 150
rect 34670 50 34730 110
rect 34670 10 34680 50
rect 34720 10 34730 50
rect 34670 -50 34730 10
rect 34670 -90 34680 -50
rect 34720 -90 34730 -50
rect 34670 -110 34730 -90
rect 34850 450 34910 470
rect 34850 410 34860 450
rect 34900 410 34910 450
rect 34850 350 34910 410
rect 34850 310 34860 350
rect 34900 310 34910 350
rect 34850 250 34910 310
rect 34850 210 34860 250
rect 34900 210 34910 250
rect 34850 150 34910 210
rect 34850 110 34860 150
rect 34900 110 34910 150
rect 34850 50 34910 110
rect 34850 10 34860 50
rect 34900 10 34910 50
rect 34850 -50 34910 10
rect 34850 -90 34860 -50
rect 34900 -90 34910 -50
rect 34850 -110 34910 -90
rect 35030 450 35090 470
rect 35030 410 35040 450
rect 35080 410 35090 450
rect 35030 350 35090 410
rect 35030 310 35040 350
rect 35080 310 35090 350
rect 35030 250 35090 310
rect 35030 210 35040 250
rect 35080 210 35090 250
rect 35030 150 35090 210
rect 35030 110 35040 150
rect 35080 110 35090 150
rect 35030 50 35090 110
rect 35030 10 35040 50
rect 35080 10 35090 50
rect 35030 -50 35090 10
rect 35030 -90 35040 -50
rect 35080 -90 35090 -50
rect 35030 -110 35090 -90
rect 35210 450 35270 470
rect 35210 410 35220 450
rect 35260 410 35270 450
rect 35210 350 35270 410
rect 35210 310 35220 350
rect 35260 310 35270 350
rect 35210 250 35270 310
rect 35210 210 35220 250
rect 35260 210 35270 250
rect 35210 150 35270 210
rect 35210 110 35220 150
rect 35260 110 35270 150
rect 35210 50 35270 110
rect 35210 10 35220 50
rect 35260 10 35270 50
rect 35210 -50 35270 10
rect 35210 -90 35220 -50
rect 35260 -90 35270 -50
rect 35210 -110 35270 -90
rect 35390 450 35450 470
rect 35390 410 35400 450
rect 35440 410 35450 450
rect 35390 350 35450 410
rect 35390 310 35400 350
rect 35440 310 35450 350
rect 35390 250 35450 310
rect 35390 210 35400 250
rect 35440 210 35450 250
rect 35390 150 35450 210
rect 35390 110 35400 150
rect 35440 110 35450 150
rect 35390 50 35450 110
rect 35390 10 35400 50
rect 35440 10 35450 50
rect 35390 -50 35450 10
rect 35390 -90 35400 -50
rect 35440 -90 35450 -50
rect 35390 -110 35450 -90
rect 35570 450 35630 470
rect 35570 410 35580 450
rect 35620 410 35630 450
rect 35570 350 35630 410
rect 35570 310 35580 350
rect 35620 310 35630 350
rect 35570 250 35630 310
rect 35570 210 35580 250
rect 35620 210 35630 250
rect 35570 150 35630 210
rect 35570 110 35580 150
rect 35620 110 35630 150
rect 35570 50 35630 110
rect 35570 10 35580 50
rect 35620 10 35630 50
rect 35570 -50 35630 10
rect 35570 -90 35580 -50
rect 35620 -90 35630 -50
rect 34220 -160 34290 -150
rect 34280 -220 34290 -160
rect 34220 -230 34290 -220
rect 34390 -160 34470 -150
rect 34390 -220 34400 -160
rect 34460 -220 34470 -160
rect 34390 -230 34470 -220
rect 34500 -480 34540 -110
rect 34570 -160 34650 -150
rect 34570 -220 34580 -160
rect 34640 -220 34650 -160
rect 34570 -230 34650 -220
rect 34750 -160 34830 -150
rect 34750 -220 34760 -160
rect 34820 -220 34830 -160
rect 34750 -230 34830 -220
rect 34860 -370 34900 -110
rect 34930 -160 35010 -150
rect 34930 -220 34940 -160
rect 35000 -220 35010 -160
rect 34930 -230 35010 -220
rect 35110 -160 35190 -150
rect 35110 -220 35120 -160
rect 35180 -220 35190 -160
rect 35110 -230 35190 -220
rect 35220 -260 35260 -110
rect 35290 -160 35540 -150
rect 35290 -220 35300 -160
rect 35360 -220 35390 -160
rect 35450 -220 35480 -160
rect 35290 -230 35540 -220
rect 35200 -270 35280 -260
rect 35200 -330 35210 -270
rect 35270 -330 35280 -270
rect 35200 -340 35280 -330
rect 34840 -380 34920 -370
rect 34840 -440 34850 -380
rect 34910 -440 34920 -380
rect 34840 -450 34920 -440
rect 34480 -490 34560 -480
rect 34480 -550 34490 -490
rect 34550 -550 34560 -490
rect 34480 -560 34560 -550
rect 34120 -600 34200 -590
rect 34120 -660 34130 -600
rect 34190 -660 34200 -600
rect 34120 -670 34200 -660
rect 33080 -710 33160 -700
rect 33080 -770 33090 -710
rect 33150 -770 33160 -710
rect 33080 -790 33160 -770
rect 33080 -850 33090 -790
rect 33150 -850 33160 -790
rect 33080 -870 33160 -850
rect 33080 -930 33090 -870
rect 33150 -930 33160 -870
rect 33080 -940 33160 -930
rect 33320 -710 33400 -700
rect 33320 -770 33330 -710
rect 33390 -770 33400 -710
rect 33320 -790 33400 -770
rect 33320 -850 33330 -790
rect 33390 -850 33400 -790
rect 33320 -870 33400 -850
rect 33320 -930 33330 -870
rect 33390 -930 33400 -870
rect 33320 -940 33400 -930
rect 33560 -710 33640 -700
rect 33560 -770 33570 -710
rect 33630 -770 33640 -710
rect 33560 -790 33640 -770
rect 33560 -850 33570 -790
rect 33630 -850 33640 -790
rect 33560 -870 33640 -850
rect 33560 -930 33570 -870
rect 33630 -930 33640 -870
rect 33560 -940 33640 -930
rect 33800 -710 33880 -700
rect 33800 -770 33810 -710
rect 33870 -770 33880 -710
rect 33800 -790 33880 -770
rect 33800 -850 33810 -790
rect 33870 -850 33880 -790
rect 33800 -870 33880 -850
rect 33800 -930 33810 -870
rect 33870 -930 33880 -870
rect 33800 -940 33880 -930
rect 34040 -710 34120 -700
rect 34040 -770 34050 -710
rect 34110 -770 34120 -710
rect 34040 -790 34120 -770
rect 34040 -850 34050 -790
rect 34110 -850 34120 -790
rect 34040 -870 34120 -850
rect 34040 -930 34050 -870
rect 34110 -930 34120 -870
rect 34040 -940 34120 -930
rect 34280 -710 34360 -700
rect 34280 -770 34290 -710
rect 34350 -770 34360 -710
rect 34280 -790 34360 -770
rect 34280 -850 34290 -790
rect 34350 -850 34360 -790
rect 34280 -870 34360 -850
rect 34280 -930 34290 -870
rect 34350 -930 34360 -870
rect 34280 -940 34360 -930
rect 34520 -710 34600 -700
rect 34520 -770 34530 -710
rect 34590 -770 34600 -710
rect 34520 -790 34600 -770
rect 34520 -850 34530 -790
rect 34590 -850 34600 -790
rect 34520 -870 34600 -850
rect 34520 -930 34530 -870
rect 34590 -930 34600 -870
rect 34520 -940 34600 -930
rect 34760 -710 34840 -700
rect 34760 -770 34770 -710
rect 34830 -770 34840 -710
rect 34760 -790 34840 -770
rect 34760 -850 34770 -790
rect 34830 -850 34840 -790
rect 34760 -870 34840 -850
rect 34760 -930 34770 -870
rect 34830 -930 34840 -870
rect 34760 -940 34840 -930
rect 35000 -710 35080 -700
rect 35000 -770 35010 -710
rect 35070 -770 35080 -710
rect 35000 -790 35080 -770
rect 35000 -850 35010 -790
rect 35070 -850 35080 -790
rect 35000 -870 35080 -850
rect 35000 -930 35010 -870
rect 35070 -930 35080 -870
rect 35000 -940 35080 -930
rect 35240 -710 35320 -700
rect 35240 -770 35250 -710
rect 35310 -770 35320 -710
rect 35240 -790 35320 -770
rect 35240 -850 35250 -790
rect 35310 -850 35320 -790
rect 35240 -870 35320 -850
rect 35240 -930 35250 -870
rect 35310 -930 35320 -870
rect 35240 -940 35320 -930
rect 32960 -1040 32970 -980
rect 33030 -1040 33040 -980
rect 32960 -1050 33040 -1040
rect 32850 -1150 32860 -1110
rect 32900 -1150 32910 -1110
rect 32850 -1210 32910 -1150
rect 32850 -1250 32860 -1210
rect 32900 -1250 32910 -1210
rect 32850 -1270 32910 -1250
rect 32970 -1110 33030 -1050
rect 32970 -1150 32980 -1110
rect 33020 -1150 33030 -1110
rect 32970 -1210 33030 -1150
rect 32970 -1250 32980 -1210
rect 33020 -1250 33030 -1210
rect 32970 -1270 33030 -1250
rect 33090 -1110 33150 -940
rect 33090 -1150 33100 -1110
rect 33140 -1150 33150 -1110
rect 33090 -1210 33150 -1150
rect 33090 -1250 33100 -1210
rect 33140 -1250 33150 -1210
rect 33090 -1270 33150 -1250
rect 33210 -1110 33270 -1090
rect 33210 -1150 33220 -1110
rect 33260 -1150 33270 -1110
rect 33210 -1210 33270 -1150
rect 33210 -1250 33220 -1210
rect 33260 -1250 33270 -1210
rect 33210 -1310 33270 -1250
rect 33330 -1110 33390 -940
rect 33330 -1150 33340 -1110
rect 33380 -1150 33390 -1110
rect 33330 -1210 33390 -1150
rect 33330 -1250 33340 -1210
rect 33380 -1250 33390 -1210
rect 33330 -1270 33390 -1250
rect 33450 -1110 33510 -1090
rect 33450 -1150 33460 -1110
rect 33500 -1150 33510 -1110
rect 33450 -1210 33510 -1150
rect 33450 -1250 33460 -1210
rect 33500 -1250 33510 -1210
rect 33200 -1320 33280 -1310
rect 33030 -1340 33090 -1320
rect 33030 -1380 33040 -1340
rect 33080 -1380 33090 -1340
rect 33030 -1430 33090 -1380
rect 33200 -1380 33210 -1320
rect 33270 -1380 33280 -1320
rect 33200 -1390 33280 -1380
rect 33450 -1430 33510 -1250
rect 33570 -1110 33630 -940
rect 33680 -980 33760 -970
rect 33680 -1040 33690 -980
rect 33750 -1040 33760 -980
rect 33680 -1050 33760 -1040
rect 33570 -1150 33580 -1110
rect 33620 -1150 33630 -1110
rect 33570 -1210 33630 -1150
rect 33570 -1250 33580 -1210
rect 33620 -1250 33630 -1210
rect 33570 -1270 33630 -1250
rect 33690 -1110 33750 -1050
rect 33690 -1150 33700 -1110
rect 33740 -1150 33750 -1110
rect 33690 -1210 33750 -1150
rect 33690 -1250 33700 -1210
rect 33740 -1250 33750 -1210
rect 33690 -1270 33750 -1250
rect 33810 -1110 33870 -940
rect 33810 -1150 33820 -1110
rect 33860 -1150 33870 -1110
rect 33810 -1210 33870 -1150
rect 33810 -1250 33820 -1210
rect 33860 -1250 33870 -1210
rect 33810 -1270 33870 -1250
rect 33930 -1110 33990 -1090
rect 33930 -1150 33940 -1110
rect 33980 -1150 33990 -1110
rect 33930 -1210 33990 -1150
rect 33930 -1250 33940 -1210
rect 33980 -1250 33990 -1210
rect 33930 -1310 33990 -1250
rect 34050 -1110 34110 -940
rect 34050 -1150 34060 -1110
rect 34100 -1150 34110 -1110
rect 34050 -1210 34110 -1150
rect 34050 -1250 34060 -1210
rect 34100 -1250 34110 -1210
rect 34050 -1270 34110 -1250
rect 34170 -1110 34230 -1090
rect 34170 -1150 34180 -1110
rect 34220 -1150 34230 -1110
rect 34170 -1210 34230 -1150
rect 34170 -1250 34180 -1210
rect 34220 -1250 34230 -1210
rect 33690 -1330 33750 -1310
rect 33690 -1370 33700 -1330
rect 33740 -1370 33750 -1330
rect 33690 -1430 33750 -1370
rect 33920 -1320 34000 -1310
rect 33920 -1380 33930 -1320
rect 33990 -1380 34000 -1320
rect 33020 -1440 33100 -1430
rect 33020 -1500 33030 -1440
rect 33090 -1500 33100 -1440
rect 33020 -1520 33100 -1500
rect 33020 -1580 33030 -1520
rect 33090 -1580 33100 -1520
rect 33020 -1600 33100 -1580
rect 33020 -1660 33030 -1600
rect 33090 -1660 33100 -1600
rect 33020 -1670 33100 -1660
rect 33440 -1440 33520 -1430
rect 33440 -1500 33450 -1440
rect 33510 -1500 33520 -1440
rect 33440 -1520 33520 -1500
rect 33440 -1580 33450 -1520
rect 33510 -1580 33520 -1520
rect 33440 -1600 33520 -1580
rect 33440 -1660 33450 -1600
rect 33510 -1660 33520 -1600
rect 33440 -1670 33520 -1660
rect 33680 -1440 33760 -1430
rect 33680 -1500 33690 -1440
rect 33750 -1500 33760 -1440
rect 33680 -1520 33760 -1500
rect 33680 -1580 33690 -1520
rect 33750 -1580 33760 -1520
rect 33680 -1600 33760 -1580
rect 33680 -1660 33690 -1600
rect 33750 -1660 33760 -1600
rect 33680 -1710 33760 -1660
rect 33680 -1770 33690 -1710
rect 33750 -1770 33760 -1710
rect 33680 -1780 33760 -1770
rect 33690 -2050 33750 -1780
rect 33920 -1820 34000 -1380
rect 34170 -1430 34230 -1250
rect 34290 -1110 34350 -940
rect 34400 -980 34480 -970
rect 34400 -1040 34410 -980
rect 34470 -1040 34480 -980
rect 34400 -1050 34480 -1040
rect 34290 -1150 34300 -1110
rect 34340 -1150 34350 -1110
rect 34290 -1210 34350 -1150
rect 34290 -1250 34300 -1210
rect 34340 -1250 34350 -1210
rect 34290 -1270 34350 -1250
rect 34410 -1110 34470 -1050
rect 34410 -1150 34420 -1110
rect 34460 -1150 34470 -1110
rect 34410 -1210 34470 -1150
rect 34410 -1250 34420 -1210
rect 34460 -1250 34470 -1210
rect 34410 -1270 34470 -1250
rect 34530 -1110 34590 -940
rect 34530 -1150 34540 -1110
rect 34580 -1150 34590 -1110
rect 34530 -1210 34590 -1150
rect 34530 -1250 34540 -1210
rect 34580 -1250 34590 -1210
rect 34530 -1270 34590 -1250
rect 34650 -1110 34710 -1090
rect 34650 -1150 34660 -1110
rect 34700 -1150 34710 -1110
rect 34650 -1210 34710 -1150
rect 34650 -1250 34660 -1210
rect 34700 -1250 34710 -1210
rect 34650 -1310 34710 -1250
rect 34770 -1110 34830 -940
rect 34770 -1150 34780 -1110
rect 34820 -1150 34830 -1110
rect 34770 -1210 34830 -1150
rect 34770 -1250 34780 -1210
rect 34820 -1250 34830 -1210
rect 34770 -1270 34830 -1250
rect 34890 -1110 34950 -1090
rect 34890 -1150 34900 -1110
rect 34940 -1150 34950 -1110
rect 34890 -1210 34950 -1150
rect 34890 -1250 34900 -1210
rect 34940 -1250 34950 -1210
rect 34410 -1330 34470 -1310
rect 34410 -1370 34420 -1330
rect 34460 -1370 34470 -1330
rect 34410 -1430 34470 -1370
rect 34640 -1320 34720 -1310
rect 34640 -1380 34650 -1320
rect 34710 -1380 34720 -1320
rect 34640 -1390 34720 -1380
rect 34890 -1430 34950 -1250
rect 35010 -1110 35070 -940
rect 35120 -980 35200 -970
rect 35120 -1040 35130 -980
rect 35190 -1040 35200 -980
rect 35120 -1050 35200 -1040
rect 35250 -990 35310 -940
rect 35250 -1030 35260 -990
rect 35300 -1030 35310 -990
rect 35010 -1150 35020 -1110
rect 35060 -1150 35070 -1110
rect 35010 -1210 35070 -1150
rect 35010 -1250 35020 -1210
rect 35060 -1250 35070 -1210
rect 35010 -1270 35070 -1250
rect 35130 -1110 35190 -1050
rect 35130 -1150 35140 -1110
rect 35180 -1150 35190 -1110
rect 35130 -1210 35190 -1150
rect 35130 -1250 35140 -1210
rect 35180 -1250 35190 -1210
rect 35130 -1270 35190 -1250
rect 35250 -1110 35310 -1030
rect 35380 -980 35460 -230
rect 35570 -590 35630 -90
rect 35750 450 35810 470
rect 35750 410 35760 450
rect 35800 410 35810 450
rect 35750 350 35810 410
rect 35750 310 35760 350
rect 35800 310 35810 350
rect 35750 250 35810 310
rect 35750 210 35760 250
rect 35800 210 35810 250
rect 35750 150 35810 210
rect 35750 110 35760 150
rect 35800 110 35810 150
rect 35750 50 35810 110
rect 35750 10 35760 50
rect 35800 10 35810 50
rect 35750 -50 35810 10
rect 35750 -90 35760 -50
rect 35800 -90 35810 -50
rect 35750 -110 35810 -90
rect 35930 450 35990 470
rect 35930 410 35940 450
rect 35980 410 35990 450
rect 35930 350 35990 410
rect 35930 310 35940 350
rect 35980 310 35990 350
rect 35930 250 35990 310
rect 35930 210 35940 250
rect 35980 210 35990 250
rect 35930 150 35990 210
rect 35930 110 35940 150
rect 35980 110 35990 150
rect 35930 50 35990 110
rect 35930 10 35940 50
rect 35980 10 35990 50
rect 35930 -50 35990 10
rect 35930 -90 35940 -50
rect 35980 -90 35990 -50
rect 35930 -110 35990 -90
rect 36110 450 36170 470
rect 36110 410 36120 450
rect 36160 410 36170 450
rect 36110 350 36170 410
rect 36110 310 36120 350
rect 36160 310 36170 350
rect 36110 250 36170 310
rect 36110 210 36120 250
rect 36160 210 36170 250
rect 36110 150 36170 210
rect 36110 110 36120 150
rect 36160 110 36170 150
rect 36110 50 36170 110
rect 36110 10 36120 50
rect 36160 10 36170 50
rect 36110 -50 36170 10
rect 36110 -90 36120 -50
rect 36160 -90 36170 -50
rect 36110 -110 36170 -90
rect 36290 450 36350 470
rect 36290 410 36300 450
rect 36340 410 36350 450
rect 36290 350 36350 410
rect 36290 310 36300 350
rect 36340 310 36350 350
rect 36290 250 36350 310
rect 36290 210 36300 250
rect 36340 210 36350 250
rect 36290 150 36350 210
rect 36290 110 36300 150
rect 36340 110 36350 150
rect 36290 50 36350 110
rect 36290 10 36300 50
rect 36340 10 36350 50
rect 36290 -50 36350 10
rect 36290 -90 36300 -50
rect 36340 -90 36350 -50
rect 36290 -110 36350 -90
rect 36470 450 36530 470
rect 36470 410 36480 450
rect 36520 410 36530 450
rect 36470 350 36530 410
rect 36470 310 36480 350
rect 36520 310 36530 350
rect 36470 250 36530 310
rect 36470 210 36480 250
rect 36520 210 36530 250
rect 36470 150 36530 210
rect 36470 110 36480 150
rect 36520 110 36530 150
rect 36470 50 36530 110
rect 36470 10 36480 50
rect 36520 10 36530 50
rect 36470 -50 36530 10
rect 36470 -90 36480 -50
rect 36520 -90 36530 -50
rect 36470 -110 36530 -90
rect 36650 450 36710 470
rect 36650 410 36660 450
rect 36700 410 36710 450
rect 36650 350 36710 410
rect 36650 310 36660 350
rect 36700 310 36710 350
rect 36650 250 36710 310
rect 36650 210 36660 250
rect 36700 210 36710 250
rect 36650 150 36710 210
rect 36650 110 36660 150
rect 36700 110 36710 150
rect 36650 50 36710 110
rect 36650 10 36660 50
rect 36700 10 36710 50
rect 36650 -50 36710 10
rect 36650 -90 36660 -50
rect 36700 -90 36710 -50
rect 36650 -110 36710 -90
rect 36830 450 36890 470
rect 36830 410 36840 450
rect 36880 410 36890 450
rect 36830 350 36890 410
rect 36830 310 36840 350
rect 36880 310 36890 350
rect 36830 250 36890 310
rect 36830 210 36840 250
rect 36880 210 36890 250
rect 36830 150 36890 210
rect 36830 110 36840 150
rect 36880 110 36890 150
rect 36830 50 36890 110
rect 36830 10 36840 50
rect 36880 10 36890 50
rect 36830 -50 36890 10
rect 36830 -90 36840 -50
rect 36880 -90 36890 -50
rect 36830 -110 36890 -90
rect 37010 450 37070 470
rect 37010 410 37020 450
rect 37060 410 37070 450
rect 37010 350 37070 410
rect 37010 310 37020 350
rect 37060 310 37070 350
rect 37010 250 37070 310
rect 37010 210 37020 250
rect 37060 210 37070 250
rect 37010 150 37070 210
rect 37010 110 37020 150
rect 37060 110 37070 150
rect 37010 50 37070 110
rect 37010 10 37020 50
rect 37060 10 37070 50
rect 37010 -50 37070 10
rect 37010 -90 37020 -50
rect 37060 -90 37070 -50
rect 35660 -160 35730 -150
rect 35720 -220 35730 -160
rect 35660 -230 35730 -220
rect 35830 -160 35910 -150
rect 35830 -220 35840 -160
rect 35900 -220 35910 -160
rect 35830 -230 35910 -220
rect 35940 -260 35980 -110
rect 36010 -160 36090 -150
rect 36010 -220 36020 -160
rect 36080 -220 36090 -160
rect 36010 -230 36090 -220
rect 36190 -160 36270 -150
rect 36190 -220 36200 -160
rect 36260 -220 36270 -160
rect 36190 -230 36270 -220
rect 35920 -270 36000 -260
rect 35920 -330 35930 -270
rect 35990 -330 36000 -270
rect 35920 -340 36000 -330
rect 36300 -370 36340 -110
rect 36370 -160 36450 -150
rect 36370 -220 36380 -160
rect 36440 -220 36450 -160
rect 36370 -230 36450 -220
rect 36550 -160 36630 -150
rect 36550 -220 36560 -160
rect 36620 -220 36630 -160
rect 36550 -230 36630 -220
rect 36280 -380 36360 -370
rect 36280 -440 36290 -380
rect 36350 -440 36360 -380
rect 36280 -450 36360 -440
rect 36660 -480 36700 -110
rect 36730 -160 36810 -150
rect 36730 -220 36740 -160
rect 36800 -220 36810 -160
rect 36730 -230 36810 -220
rect 36910 -160 36980 -150
rect 36910 -220 36920 -160
rect 36910 -230 36980 -220
rect 36640 -490 36720 -480
rect 36640 -550 36650 -490
rect 36710 -550 36720 -490
rect 36640 -560 36720 -550
rect 37010 -590 37070 -90
rect 37190 450 37250 470
rect 37190 410 37200 450
rect 37240 410 37250 450
rect 37190 350 37250 410
rect 37190 310 37200 350
rect 37240 310 37250 350
rect 37190 250 37250 310
rect 37190 210 37200 250
rect 37240 210 37250 250
rect 37190 150 37250 210
rect 37190 110 37200 150
rect 37240 110 37250 150
rect 37190 50 37250 110
rect 37190 10 37200 50
rect 37240 10 37250 50
rect 37190 -50 37250 10
rect 37190 -90 37200 -50
rect 37240 -90 37250 -50
rect 37190 -110 37250 -90
rect 35560 -600 35640 -590
rect 35560 -660 35570 -600
rect 35630 -660 35640 -600
rect 35560 -670 35640 -660
rect 37000 -600 37080 -590
rect 37000 -660 37010 -600
rect 37070 -660 37080 -600
rect 37000 -670 37080 -660
rect 35880 -710 35960 -700
rect 35880 -770 35890 -710
rect 35950 -770 35960 -710
rect 35880 -790 35960 -770
rect 35880 -850 35890 -790
rect 35950 -850 35960 -790
rect 35880 -870 35960 -850
rect 35880 -930 35890 -870
rect 35950 -930 35960 -870
rect 35880 -940 35960 -930
rect 36120 -710 36200 -700
rect 36120 -770 36130 -710
rect 36190 -770 36200 -710
rect 36120 -790 36200 -770
rect 36120 -850 36130 -790
rect 36190 -850 36200 -790
rect 36120 -870 36200 -850
rect 36120 -930 36130 -870
rect 36190 -930 36200 -870
rect 36120 -940 36200 -930
rect 36360 -710 36440 -700
rect 36360 -770 36370 -710
rect 36430 -770 36440 -710
rect 36360 -790 36440 -770
rect 36360 -850 36370 -790
rect 36430 -850 36440 -790
rect 36360 -870 36440 -850
rect 36360 -930 36370 -870
rect 36430 -930 36440 -870
rect 36360 -940 36440 -930
rect 36600 -710 36680 -700
rect 36600 -770 36610 -710
rect 36670 -770 36680 -710
rect 36600 -790 36680 -770
rect 36600 -850 36610 -790
rect 36670 -850 36680 -790
rect 36600 -870 36680 -850
rect 36600 -930 36610 -870
rect 36670 -930 36680 -870
rect 36600 -940 36680 -930
rect 36840 -710 36920 -700
rect 36840 -770 36850 -710
rect 36910 -770 36920 -710
rect 36840 -790 36920 -770
rect 36840 -850 36850 -790
rect 36910 -850 36920 -790
rect 36840 -870 36920 -850
rect 36840 -930 36850 -870
rect 36910 -930 36920 -870
rect 36840 -940 36920 -930
rect 37080 -710 37160 -700
rect 37080 -770 37090 -710
rect 37150 -770 37160 -710
rect 37080 -790 37160 -770
rect 37080 -850 37090 -790
rect 37150 -850 37160 -790
rect 37080 -870 37160 -850
rect 37080 -930 37090 -870
rect 37150 -930 37160 -870
rect 37080 -940 37160 -930
rect 37320 -710 37400 -700
rect 37320 -770 37330 -710
rect 37390 -770 37400 -710
rect 37320 -790 37400 -770
rect 37320 -850 37330 -790
rect 37390 -850 37400 -790
rect 37320 -870 37400 -850
rect 37320 -930 37330 -870
rect 37390 -930 37400 -870
rect 37320 -940 37400 -930
rect 37560 -710 37640 -700
rect 37560 -770 37570 -710
rect 37630 -770 37640 -710
rect 37560 -790 37640 -770
rect 37560 -850 37570 -790
rect 37630 -850 37640 -790
rect 37560 -870 37640 -850
rect 37560 -930 37570 -870
rect 37630 -930 37640 -870
rect 37560 -940 37640 -930
rect 37800 -710 37880 -700
rect 37800 -770 37810 -710
rect 37870 -770 37880 -710
rect 37800 -790 37880 -770
rect 37800 -850 37810 -790
rect 37870 -850 37880 -790
rect 37800 -870 37880 -850
rect 37800 -930 37810 -870
rect 37870 -930 37880 -870
rect 37800 -940 37880 -930
rect 38040 -710 38120 -700
rect 38040 -770 38050 -710
rect 38110 -770 38120 -710
rect 38040 -790 38120 -770
rect 38040 -850 38050 -790
rect 38110 -850 38120 -790
rect 38040 -870 38120 -850
rect 38040 -930 38050 -870
rect 38110 -930 38120 -870
rect 38040 -940 38120 -930
rect 38280 -710 38360 -700
rect 38280 -770 38290 -710
rect 38350 -770 38360 -710
rect 38280 -790 38360 -770
rect 38280 -850 38290 -790
rect 38350 -850 38360 -790
rect 38280 -870 38360 -850
rect 38280 -930 38290 -870
rect 38350 -930 38360 -870
rect 38280 -940 38360 -930
rect 35380 -1040 35390 -980
rect 35450 -1040 35460 -980
rect 35380 -1050 35460 -1040
rect 35740 -980 35820 -970
rect 35740 -1040 35750 -980
rect 35810 -1040 35820 -980
rect 35740 -1050 35820 -1040
rect 35890 -990 35950 -940
rect 35890 -1030 35900 -990
rect 35940 -1030 35950 -990
rect 35250 -1150 35260 -1110
rect 35300 -1150 35310 -1110
rect 35250 -1210 35310 -1150
rect 35250 -1250 35260 -1210
rect 35300 -1250 35310 -1210
rect 35250 -1270 35310 -1250
rect 35070 -1330 35130 -1310
rect 35070 -1370 35080 -1330
rect 35120 -1370 35130 -1330
rect 35070 -1430 35130 -1370
rect 34160 -1440 34240 -1430
rect 34160 -1500 34170 -1440
rect 34230 -1500 34240 -1440
rect 34160 -1520 34240 -1500
rect 34160 -1580 34170 -1520
rect 34230 -1580 34240 -1520
rect 34160 -1600 34240 -1580
rect 34160 -1660 34170 -1600
rect 34230 -1660 34240 -1600
rect 34160 -1670 34240 -1660
rect 34400 -1440 34480 -1430
rect 34400 -1500 34410 -1440
rect 34470 -1500 34480 -1440
rect 34400 -1520 34480 -1500
rect 34400 -1580 34410 -1520
rect 34470 -1580 34480 -1520
rect 34400 -1600 34480 -1580
rect 34400 -1660 34410 -1600
rect 34470 -1660 34480 -1600
rect 34400 -1670 34480 -1660
rect 34640 -1440 34720 -1430
rect 34640 -1500 34650 -1440
rect 34710 -1500 34720 -1440
rect 34640 -1520 34720 -1500
rect 34640 -1580 34650 -1520
rect 34710 -1580 34720 -1520
rect 34640 -1600 34720 -1580
rect 34640 -1660 34650 -1600
rect 34710 -1660 34720 -1600
rect 34640 -1670 34720 -1660
rect 34880 -1440 34960 -1430
rect 34880 -1500 34890 -1440
rect 34950 -1500 34960 -1440
rect 34880 -1520 34960 -1500
rect 34880 -1580 34890 -1520
rect 34950 -1580 34960 -1520
rect 34880 -1600 34960 -1580
rect 34880 -1660 34890 -1600
rect 34950 -1660 34960 -1600
rect 34880 -1670 34960 -1660
rect 35060 -1440 35140 -1430
rect 35060 -1500 35070 -1440
rect 35130 -1500 35140 -1440
rect 35060 -1520 35140 -1500
rect 35060 -1580 35070 -1520
rect 35130 -1580 35140 -1520
rect 35060 -1600 35140 -1580
rect 35060 -1660 35070 -1600
rect 35130 -1660 35140 -1600
rect 35060 -1670 35140 -1660
rect 34160 -1710 34240 -1700
rect 34160 -1770 34170 -1710
rect 34230 -1770 34240 -1710
rect 34160 -1780 34240 -1770
rect 34640 -1710 34720 -1700
rect 34640 -1770 34650 -1710
rect 34710 -1770 34720 -1710
rect 34640 -1780 34720 -1770
rect 33920 -1880 33930 -1820
rect 33990 -1880 34000 -1820
rect 33920 -1890 34000 -1880
rect 33852 -1930 33910 -1920
rect 33852 -1982 33856 -1930
rect 33908 -1982 33910 -1930
rect 33852 -1990 33910 -1982
rect 33940 -2030 33980 -1890
rect 34010 -1930 34068 -1920
rect 34010 -1982 34014 -1930
rect 34066 -1982 34068 -1930
rect 34010 -1990 34068 -1982
rect 34180 -2030 34220 -1780
rect 34400 -1820 34480 -1810
rect 34400 -1880 34410 -1820
rect 34470 -1880 34480 -1820
rect 34400 -1890 34480 -1880
rect 34334 -1930 34392 -1920
rect 34334 -1982 34338 -1930
rect 34390 -1982 34392 -1930
rect 34334 -1990 34392 -1982
rect 34420 -2030 34460 -1890
rect 34488 -1930 34546 -1920
rect 34488 -1982 34492 -1930
rect 34544 -1982 34546 -1930
rect 34488 -1990 34546 -1982
rect 34660 -2030 34700 -1780
rect 34880 -1820 34960 -1810
rect 34880 -1880 34890 -1820
rect 34950 -1880 34960 -1820
rect 34880 -1890 34960 -1880
rect 34812 -1930 34870 -1920
rect 34812 -1982 34816 -1930
rect 34868 -1982 34870 -1930
rect 34812 -1990 34870 -1982
rect 34900 -2030 34940 -1890
rect 35120 -1970 35200 -1960
rect 35120 -2030 35130 -1970
rect 35190 -2030 35200 -1970
rect 33690 -2090 33700 -2050
rect 33740 -2090 33750 -2050
rect 33690 -2110 33750 -2090
rect 33810 -2050 33870 -2030
rect 33810 -2090 33820 -2050
rect 33860 -2090 33870 -2050
rect 33810 -2110 33870 -2090
rect 33930 -2050 33990 -2030
rect 33930 -2090 33940 -2050
rect 33980 -2090 33990 -2050
rect 33930 -2110 33990 -2090
rect 34050 -2050 34110 -2030
rect 34050 -2090 34060 -2050
rect 34100 -2090 34110 -2050
rect 34050 -2110 34110 -2090
rect 34170 -2050 34230 -2030
rect 34170 -2090 34180 -2050
rect 34220 -2090 34230 -2050
rect 34170 -2110 34230 -2090
rect 34290 -2050 34350 -2030
rect 34290 -2090 34300 -2050
rect 34340 -2090 34350 -2050
rect 34290 -2110 34350 -2090
rect 34410 -2050 34470 -2030
rect 34410 -2090 34420 -2050
rect 34460 -2090 34470 -2050
rect 34410 -2110 34470 -2090
rect 34530 -2050 34590 -2030
rect 34530 -2090 34540 -2050
rect 34580 -2090 34590 -2050
rect 34530 -2110 34590 -2090
rect 34650 -2050 34710 -2030
rect 34650 -2090 34660 -2050
rect 34700 -2090 34710 -2050
rect 34650 -2110 34710 -2090
rect 34770 -2050 34830 -2030
rect 34770 -2090 34780 -2050
rect 34820 -2090 34830 -2050
rect 34770 -2110 34830 -2090
rect 34890 -2050 34950 -2030
rect 34890 -2090 34900 -2050
rect 34940 -2090 34950 -2050
rect 34890 -2110 34950 -2090
rect 35120 -2050 35200 -2030
rect 35120 -2110 35130 -2050
rect 35190 -2110 35200 -2050
rect 32650 -2150 32730 -2140
rect 32650 -2210 32660 -2150
rect 32720 -2210 32730 -2150
rect 32650 -2220 32730 -2210
rect 33751 -2158 33809 -2150
rect 33751 -2210 33753 -2158
rect 33805 -2210 33809 -2158
rect 33751 -2220 33809 -2210
rect 32670 -3990 32710 -2220
rect 33840 -2250 33870 -2110
rect 34050 -2250 34080 -2110
rect 34111 -2158 34169 -2150
rect 34111 -2210 34113 -2158
rect 34165 -2210 34169 -2158
rect 34111 -2220 34169 -2210
rect 34231 -2158 34289 -2150
rect 34231 -2210 34233 -2158
rect 34285 -2210 34289 -2158
rect 34231 -2220 34289 -2210
rect 34320 -2250 34350 -2110
rect 34530 -2250 34560 -2110
rect 34591 -2158 34649 -2150
rect 34591 -2210 34593 -2158
rect 34645 -2210 34649 -2158
rect 34591 -2220 34649 -2210
rect 34711 -2158 34769 -2150
rect 34711 -2210 34713 -2158
rect 34765 -2210 34769 -2158
rect 34711 -2220 34769 -2210
rect 34800 -2250 34830 -2110
rect 35120 -2130 35200 -2110
rect 35120 -2190 35130 -2130
rect 35190 -2190 35200 -2130
rect 35120 -2200 35200 -2190
rect 33060 -2260 33140 -2250
rect 33060 -2320 33070 -2260
rect 33130 -2320 33140 -2260
rect 33060 -2330 33140 -2320
rect 33810 -2260 33890 -2250
rect 33810 -2320 33820 -2260
rect 33880 -2320 33890 -2260
rect 33810 -2330 33890 -2320
rect 34030 -2260 34110 -2250
rect 34030 -2320 34040 -2260
rect 34100 -2320 34110 -2260
rect 34030 -2330 34110 -2320
rect 34290 -2260 34370 -2250
rect 34290 -2320 34300 -2260
rect 34360 -2320 34370 -2260
rect 34290 -2330 34370 -2320
rect 34510 -2260 34590 -2250
rect 34510 -2320 34520 -2260
rect 34580 -2320 34590 -2260
rect 34510 -2330 34590 -2320
rect 34770 -2260 34850 -2250
rect 34770 -2320 34780 -2260
rect 34840 -2320 34850 -2260
rect 34770 -2330 34850 -2320
rect 33070 -2660 33130 -2330
rect 33240 -2370 33320 -2360
rect 33240 -2430 33250 -2370
rect 33310 -2430 33320 -2370
rect 33240 -2450 33320 -2430
rect 33240 -2510 33250 -2450
rect 33310 -2510 33320 -2450
rect 33240 -2530 33320 -2510
rect 33240 -2590 33250 -2530
rect 33310 -2590 33320 -2530
rect 33240 -2600 33320 -2590
rect 33480 -2370 33560 -2360
rect 33480 -2430 33490 -2370
rect 33550 -2430 33560 -2370
rect 33480 -2450 33560 -2430
rect 33480 -2510 33490 -2450
rect 33550 -2510 33560 -2450
rect 33480 -2530 33560 -2510
rect 33480 -2590 33490 -2530
rect 33550 -2590 33560 -2530
rect 33480 -2600 33560 -2590
rect 33720 -2370 33800 -2360
rect 33720 -2430 33730 -2370
rect 33790 -2430 33800 -2370
rect 33720 -2450 33800 -2430
rect 33720 -2510 33730 -2450
rect 33790 -2510 33800 -2450
rect 33720 -2530 33800 -2510
rect 33720 -2590 33730 -2530
rect 33790 -2590 33800 -2530
rect 33720 -2600 33800 -2590
rect 33960 -2370 34040 -2360
rect 33960 -2430 33970 -2370
rect 34030 -2430 34040 -2370
rect 33960 -2450 34040 -2430
rect 33960 -2510 33970 -2450
rect 34030 -2510 34040 -2450
rect 33960 -2530 34040 -2510
rect 33960 -2590 33970 -2530
rect 34030 -2590 34040 -2530
rect 33960 -2600 34040 -2590
rect 34600 -2370 34680 -2360
rect 34600 -2430 34610 -2370
rect 34670 -2430 34680 -2370
rect 34600 -2450 34680 -2430
rect 34600 -2510 34610 -2450
rect 34670 -2510 34680 -2450
rect 34600 -2530 34680 -2510
rect 34600 -2590 34610 -2530
rect 34670 -2590 34680 -2530
rect 34600 -2600 34680 -2590
rect 34840 -2370 34920 -2360
rect 34840 -2430 34850 -2370
rect 34910 -2430 34920 -2370
rect 34840 -2450 34920 -2430
rect 34840 -2510 34850 -2450
rect 34910 -2510 34920 -2450
rect 34840 -2530 34920 -2510
rect 34840 -2590 34850 -2530
rect 34910 -2590 34920 -2530
rect 34840 -2600 34920 -2590
rect 35080 -2370 35160 -2360
rect 35080 -2430 35090 -2370
rect 35150 -2430 35160 -2370
rect 35080 -2450 35160 -2430
rect 35080 -2510 35090 -2450
rect 35150 -2510 35160 -2450
rect 35080 -2530 35160 -2510
rect 35080 -2590 35090 -2530
rect 35150 -2590 35160 -2530
rect 35080 -2600 35160 -2590
rect 35390 -2570 35450 -1050
rect 35390 -2610 35400 -2570
rect 35440 -2610 35450 -2570
rect 35390 -2630 35450 -2610
rect 35480 -1970 35720 -1960
rect 35480 -2030 35490 -1970
rect 35550 -2030 35570 -1970
rect 35630 -2030 35650 -1970
rect 35710 -2030 35720 -1970
rect 35480 -2050 35720 -2030
rect 35480 -2110 35490 -2050
rect 35550 -2110 35570 -2050
rect 35630 -2110 35650 -2050
rect 35710 -2110 35720 -2050
rect 35480 -2130 35720 -2110
rect 35480 -2190 35490 -2130
rect 35550 -2190 35570 -2130
rect 35630 -2190 35650 -2130
rect 35710 -2190 35720 -2130
rect 33070 -2700 33080 -2660
rect 33120 -2700 33130 -2660
rect 33070 -2760 33130 -2700
rect 33070 -2800 33080 -2760
rect 33120 -2800 33130 -2760
rect 33070 -2860 33130 -2800
rect 33070 -2900 33080 -2860
rect 33120 -2900 33130 -2860
rect 33070 -2960 33130 -2900
rect 33070 -3000 33080 -2960
rect 33120 -3000 33130 -2960
rect 33070 -3060 33130 -3000
rect 33070 -3100 33080 -3060
rect 33120 -3100 33130 -3060
rect 33070 -3120 33130 -3100
rect 34220 -3170 34300 -3160
rect 34220 -3230 34230 -3170
rect 34290 -3230 34300 -3170
rect 34220 -3250 34300 -3230
rect 34220 -3310 34230 -3250
rect 34290 -3310 34300 -3250
rect 34220 -3330 34300 -3310
rect 34220 -3390 34230 -3330
rect 34290 -3390 34300 -3330
rect 34220 -3400 34300 -3390
rect 35480 -3170 35720 -2190
rect 35750 -2570 35810 -1050
rect 35890 -1110 35950 -1030
rect 36000 -980 36080 -970
rect 36000 -1040 36010 -980
rect 36070 -1040 36080 -980
rect 36000 -1050 36080 -1040
rect 35890 -1150 35900 -1110
rect 35940 -1150 35950 -1110
rect 35890 -1210 35950 -1150
rect 35890 -1250 35900 -1210
rect 35940 -1250 35950 -1210
rect 35890 -1270 35950 -1250
rect 36010 -1110 36070 -1050
rect 36010 -1150 36020 -1110
rect 36060 -1150 36070 -1110
rect 36010 -1210 36070 -1150
rect 36010 -1250 36020 -1210
rect 36060 -1250 36070 -1210
rect 36010 -1270 36070 -1250
rect 36130 -1110 36190 -940
rect 36130 -1150 36140 -1110
rect 36180 -1150 36190 -1110
rect 36130 -1210 36190 -1150
rect 36130 -1250 36140 -1210
rect 36180 -1250 36190 -1210
rect 36130 -1270 36190 -1250
rect 36250 -1110 36310 -1090
rect 36250 -1150 36260 -1110
rect 36300 -1150 36310 -1110
rect 36250 -1210 36310 -1150
rect 36250 -1250 36260 -1210
rect 36300 -1250 36310 -1210
rect 36070 -1330 36130 -1310
rect 36070 -1370 36080 -1330
rect 36120 -1370 36130 -1330
rect 36070 -1430 36130 -1370
rect 36250 -1430 36310 -1250
rect 36370 -1110 36430 -940
rect 36370 -1150 36380 -1110
rect 36420 -1150 36430 -1110
rect 36370 -1210 36430 -1150
rect 36370 -1250 36380 -1210
rect 36420 -1250 36430 -1210
rect 36370 -1270 36430 -1250
rect 36490 -1110 36550 -1090
rect 36490 -1150 36500 -1110
rect 36540 -1150 36550 -1110
rect 36490 -1210 36550 -1150
rect 36490 -1250 36500 -1210
rect 36540 -1250 36550 -1210
rect 36490 -1310 36550 -1250
rect 36610 -1110 36670 -940
rect 36720 -980 36800 -970
rect 36720 -1040 36730 -980
rect 36790 -1040 36800 -980
rect 36720 -1050 36800 -1040
rect 36610 -1150 36620 -1110
rect 36660 -1150 36670 -1110
rect 36610 -1210 36670 -1150
rect 36610 -1250 36620 -1210
rect 36660 -1250 36670 -1210
rect 36610 -1270 36670 -1250
rect 36730 -1110 36790 -1050
rect 36730 -1150 36740 -1110
rect 36780 -1150 36790 -1110
rect 36730 -1210 36790 -1150
rect 36730 -1250 36740 -1210
rect 36780 -1250 36790 -1210
rect 36730 -1270 36790 -1250
rect 36850 -1110 36910 -940
rect 36850 -1150 36860 -1110
rect 36900 -1150 36910 -1110
rect 36850 -1210 36910 -1150
rect 36850 -1250 36860 -1210
rect 36900 -1250 36910 -1210
rect 36850 -1270 36910 -1250
rect 36970 -1110 37030 -1090
rect 36970 -1150 36980 -1110
rect 37020 -1150 37030 -1110
rect 36970 -1210 37030 -1150
rect 36970 -1250 36980 -1210
rect 37020 -1250 37030 -1210
rect 36480 -1320 36560 -1310
rect 36480 -1380 36490 -1320
rect 36550 -1380 36560 -1320
rect 36480 -1390 36560 -1380
rect 36730 -1330 36790 -1310
rect 36730 -1370 36740 -1330
rect 36780 -1370 36790 -1330
rect 36730 -1430 36790 -1370
rect 36970 -1430 37030 -1250
rect 37090 -1110 37150 -940
rect 37090 -1150 37100 -1110
rect 37140 -1150 37150 -1110
rect 37090 -1210 37150 -1150
rect 37090 -1250 37100 -1210
rect 37140 -1250 37150 -1210
rect 37090 -1270 37150 -1250
rect 37210 -1110 37270 -1090
rect 37210 -1150 37220 -1110
rect 37260 -1150 37270 -1110
rect 37210 -1210 37270 -1150
rect 37210 -1250 37220 -1210
rect 37260 -1250 37270 -1210
rect 37210 -1310 37270 -1250
rect 37330 -1110 37390 -940
rect 37440 -980 37520 -970
rect 37440 -1040 37450 -980
rect 37510 -1040 37520 -980
rect 37440 -1050 37520 -1040
rect 37330 -1150 37340 -1110
rect 37380 -1150 37390 -1110
rect 37330 -1210 37390 -1150
rect 37330 -1250 37340 -1210
rect 37380 -1250 37390 -1210
rect 37330 -1270 37390 -1250
rect 37450 -1110 37510 -1050
rect 37450 -1150 37460 -1110
rect 37500 -1150 37510 -1110
rect 37450 -1210 37510 -1150
rect 37450 -1250 37460 -1210
rect 37500 -1250 37510 -1210
rect 37450 -1270 37510 -1250
rect 37570 -1110 37630 -940
rect 37570 -1150 37580 -1110
rect 37620 -1150 37630 -1110
rect 37570 -1210 37630 -1150
rect 37570 -1250 37580 -1210
rect 37620 -1250 37630 -1210
rect 37570 -1270 37630 -1250
rect 37690 -1110 37750 -1090
rect 37690 -1150 37700 -1110
rect 37740 -1150 37750 -1110
rect 37690 -1210 37750 -1150
rect 37690 -1250 37700 -1210
rect 37740 -1250 37750 -1210
rect 37200 -1320 37280 -1310
rect 37200 -1380 37210 -1320
rect 37270 -1380 37280 -1320
rect 36060 -1440 36140 -1430
rect 36060 -1500 36070 -1440
rect 36130 -1500 36140 -1440
rect 36060 -1510 36140 -1500
rect 36240 -1440 36320 -1430
rect 36240 -1500 36250 -1440
rect 36310 -1500 36320 -1440
rect 36240 -1510 36320 -1500
rect 36720 -1440 36800 -1430
rect 36720 -1500 36730 -1440
rect 36790 -1500 36800 -1440
rect 36720 -1510 36800 -1500
rect 36960 -1440 37040 -1430
rect 36960 -1500 36970 -1440
rect 37030 -1500 37040 -1440
rect 36960 -1510 37040 -1500
rect 36480 -1710 36560 -1700
rect 36480 -1770 36490 -1710
rect 36550 -1770 36560 -1710
rect 36480 -1780 36560 -1770
rect 36960 -1710 37040 -1700
rect 36960 -1770 36970 -1710
rect 37030 -1770 37040 -1710
rect 36960 -1780 37040 -1770
rect 36240 -1820 36320 -1810
rect 36240 -1880 36250 -1820
rect 36310 -1880 36320 -1820
rect 36240 -1890 36320 -1880
rect 36000 -1970 36080 -1960
rect 36000 -2030 36010 -1970
rect 36070 -2030 36080 -1970
rect 36260 -2030 36300 -1890
rect 36330 -1930 36388 -1920
rect 36330 -1982 36332 -1930
rect 36384 -1982 36388 -1930
rect 36330 -1990 36388 -1982
rect 36500 -2030 36540 -1780
rect 36720 -1820 36800 -1810
rect 36720 -1880 36730 -1820
rect 36790 -1880 36800 -1820
rect 36720 -1890 36800 -1880
rect 36654 -1930 36712 -1920
rect 36654 -1982 36656 -1930
rect 36708 -1982 36712 -1930
rect 36654 -1990 36712 -1982
rect 36740 -2030 36780 -1890
rect 36808 -1930 36866 -1920
rect 36808 -1982 36810 -1930
rect 36862 -1982 36866 -1930
rect 36808 -1990 36866 -1982
rect 36980 -2030 37020 -1780
rect 37200 -1820 37280 -1380
rect 37450 -1330 37510 -1310
rect 37450 -1370 37460 -1330
rect 37500 -1370 37510 -1330
rect 37450 -1430 37510 -1370
rect 37690 -1430 37750 -1250
rect 37810 -1110 37870 -940
rect 37810 -1150 37820 -1110
rect 37860 -1150 37870 -1110
rect 37810 -1210 37870 -1150
rect 37810 -1250 37820 -1210
rect 37860 -1250 37870 -1210
rect 37810 -1270 37870 -1250
rect 37930 -1110 37990 -1090
rect 37930 -1150 37940 -1110
rect 37980 -1150 37990 -1110
rect 37930 -1210 37990 -1150
rect 37930 -1250 37940 -1210
rect 37980 -1250 37990 -1210
rect 37930 -1310 37990 -1250
rect 38050 -1110 38110 -940
rect 38160 -980 38240 -970
rect 38160 -1040 38170 -980
rect 38230 -1040 38240 -980
rect 38160 -1050 38240 -1040
rect 38290 -990 38350 -940
rect 38290 -1030 38300 -990
rect 38340 -1030 38350 -990
rect 38050 -1150 38060 -1110
rect 38100 -1150 38110 -1110
rect 38050 -1210 38110 -1150
rect 38050 -1250 38060 -1210
rect 38100 -1250 38110 -1210
rect 38050 -1270 38110 -1250
rect 38170 -1110 38230 -1050
rect 38170 -1150 38180 -1110
rect 38220 -1150 38230 -1110
rect 38170 -1210 38230 -1150
rect 38170 -1250 38180 -1210
rect 38220 -1250 38230 -1210
rect 38170 -1270 38230 -1250
rect 38290 -1110 38350 -1030
rect 38290 -1150 38300 -1110
rect 38340 -1150 38350 -1110
rect 38290 -1210 38350 -1150
rect 38290 -1250 38300 -1210
rect 38340 -1250 38350 -1210
rect 38290 -1270 38350 -1250
rect 37920 -1320 38000 -1310
rect 37920 -1380 37930 -1320
rect 37990 -1380 38000 -1320
rect 37920 -1390 38000 -1380
rect 38110 -1340 38170 -1320
rect 38110 -1380 38120 -1340
rect 38160 -1380 38170 -1340
rect 38110 -1430 38170 -1380
rect 37440 -1440 37520 -1430
rect 37440 -1500 37450 -1440
rect 37510 -1500 37520 -1440
rect 37440 -1710 37520 -1500
rect 37680 -1440 37760 -1430
rect 37680 -1500 37690 -1440
rect 37750 -1500 37760 -1440
rect 37680 -1510 37760 -1500
rect 38100 -1440 38260 -1430
rect 38100 -1500 38110 -1440
rect 38170 -1500 38190 -1440
rect 38250 -1500 38260 -1440
rect 38100 -1510 38260 -1500
rect 37440 -1770 37450 -1710
rect 37510 -1770 37520 -1710
rect 37440 -1780 37520 -1770
rect 37200 -1880 37210 -1820
rect 37270 -1880 37280 -1820
rect 37200 -1890 37280 -1880
rect 37132 -1930 37190 -1920
rect 37132 -1982 37134 -1930
rect 37186 -1982 37190 -1930
rect 37132 -1990 37190 -1982
rect 37220 -2030 37260 -1890
rect 37290 -1930 37348 -1920
rect 37290 -1982 37292 -1930
rect 37344 -1982 37348 -1930
rect 37290 -1990 37348 -1982
rect 36000 -2050 36080 -2030
rect 36000 -2110 36010 -2050
rect 36070 -2110 36080 -2050
rect 36250 -2050 36310 -2030
rect 36250 -2090 36260 -2050
rect 36300 -2090 36310 -2050
rect 36250 -2110 36310 -2090
rect 36370 -2050 36430 -2030
rect 36370 -2090 36380 -2050
rect 36420 -2090 36430 -2050
rect 36370 -2110 36430 -2090
rect 36490 -2050 36550 -2030
rect 36490 -2090 36500 -2050
rect 36540 -2090 36550 -2050
rect 36490 -2110 36550 -2090
rect 36610 -2050 36670 -2030
rect 36610 -2090 36620 -2050
rect 36660 -2090 36670 -2050
rect 36610 -2110 36670 -2090
rect 36730 -2050 36790 -2030
rect 36730 -2090 36740 -2050
rect 36780 -2090 36790 -2050
rect 36730 -2110 36790 -2090
rect 36850 -2050 36910 -2030
rect 36850 -2090 36860 -2050
rect 36900 -2090 36910 -2050
rect 36850 -2110 36910 -2090
rect 36970 -2050 37030 -2030
rect 36970 -2090 36980 -2050
rect 37020 -2090 37030 -2050
rect 36970 -2110 37030 -2090
rect 37090 -2050 37150 -2030
rect 37090 -2090 37100 -2050
rect 37140 -2090 37150 -2050
rect 37090 -2110 37150 -2090
rect 37210 -2050 37270 -2030
rect 37210 -2090 37220 -2050
rect 37260 -2090 37270 -2050
rect 37210 -2110 37270 -2090
rect 37330 -2050 37390 -2030
rect 37330 -2090 37340 -2050
rect 37380 -2090 37390 -2050
rect 37330 -2110 37390 -2090
rect 37450 -2050 37510 -1780
rect 37450 -2090 37460 -2050
rect 37500 -2090 37510 -2050
rect 37450 -2110 37510 -2090
rect 36000 -2130 36080 -2110
rect 36000 -2190 36010 -2130
rect 36070 -2190 36080 -2130
rect 36000 -2200 36080 -2190
rect 36370 -2250 36400 -2110
rect 36431 -2158 36489 -2150
rect 36431 -2210 36435 -2158
rect 36487 -2210 36489 -2158
rect 36431 -2220 36489 -2210
rect 36551 -2158 36609 -2150
rect 36551 -2210 36555 -2158
rect 36607 -2210 36609 -2158
rect 36551 -2220 36609 -2210
rect 36640 -2250 36670 -2110
rect 36850 -2250 36880 -2110
rect 36911 -2158 36969 -2150
rect 36911 -2210 36915 -2158
rect 36967 -2210 36969 -2158
rect 36911 -2220 36969 -2210
rect 37031 -2158 37089 -2150
rect 37031 -2210 37035 -2158
rect 37087 -2210 37089 -2158
rect 37031 -2220 37089 -2210
rect 37120 -2250 37150 -2110
rect 37330 -2250 37360 -2110
rect 37391 -2158 37449 -2150
rect 37391 -2210 37395 -2158
rect 37447 -2210 37449 -2158
rect 37391 -2220 37449 -2210
rect 36350 -2260 36430 -2250
rect 36350 -2320 36360 -2260
rect 36420 -2320 36430 -2260
rect 36350 -2330 36430 -2320
rect 36610 -2260 36690 -2250
rect 36610 -2320 36620 -2260
rect 36680 -2320 36690 -2260
rect 36610 -2330 36690 -2320
rect 36830 -2260 36910 -2250
rect 36830 -2320 36840 -2260
rect 36900 -2320 36910 -2260
rect 36830 -2330 36910 -2320
rect 37090 -2260 37170 -2250
rect 37090 -2320 37100 -2260
rect 37160 -2320 37170 -2260
rect 37090 -2330 37170 -2320
rect 37310 -2260 37390 -2250
rect 37310 -2320 37320 -2260
rect 37380 -2320 37390 -2260
rect 37310 -2330 37390 -2320
rect 38060 -2260 38140 -2250
rect 38060 -2320 38070 -2260
rect 38130 -2320 38140 -2260
rect 38060 -2330 38140 -2320
rect 35750 -2610 35760 -2570
rect 35800 -2610 35810 -2570
rect 36040 -2370 36120 -2360
rect 36040 -2430 36050 -2370
rect 36110 -2430 36120 -2370
rect 36040 -2450 36120 -2430
rect 36040 -2510 36050 -2450
rect 36110 -2510 36120 -2450
rect 36040 -2530 36120 -2510
rect 36040 -2590 36050 -2530
rect 36110 -2590 36120 -2530
rect 36040 -2600 36120 -2590
rect 36280 -2370 36360 -2360
rect 36280 -2430 36290 -2370
rect 36350 -2430 36360 -2370
rect 36280 -2450 36360 -2430
rect 36280 -2510 36290 -2450
rect 36350 -2510 36360 -2450
rect 36280 -2530 36360 -2510
rect 36280 -2590 36290 -2530
rect 36350 -2590 36360 -2530
rect 36280 -2600 36360 -2590
rect 36520 -2370 36600 -2360
rect 36520 -2430 36530 -2370
rect 36590 -2430 36600 -2370
rect 36520 -2450 36600 -2430
rect 36520 -2510 36530 -2450
rect 36590 -2510 36600 -2450
rect 36520 -2530 36600 -2510
rect 36520 -2590 36530 -2530
rect 36590 -2590 36600 -2530
rect 36520 -2600 36600 -2590
rect 37160 -2370 37240 -2360
rect 37160 -2430 37170 -2370
rect 37230 -2430 37240 -2370
rect 37160 -2450 37240 -2430
rect 37160 -2510 37170 -2450
rect 37230 -2510 37240 -2450
rect 37160 -2530 37240 -2510
rect 37160 -2590 37170 -2530
rect 37230 -2590 37240 -2530
rect 37160 -2600 37240 -2590
rect 37400 -2370 37480 -2360
rect 37400 -2430 37410 -2370
rect 37470 -2430 37480 -2370
rect 37400 -2450 37480 -2430
rect 37400 -2510 37410 -2450
rect 37470 -2510 37480 -2450
rect 37400 -2530 37480 -2510
rect 37400 -2590 37410 -2530
rect 37470 -2590 37480 -2530
rect 37400 -2600 37480 -2590
rect 37640 -2370 37720 -2360
rect 37640 -2430 37650 -2370
rect 37710 -2430 37720 -2370
rect 37640 -2450 37720 -2430
rect 37640 -2510 37650 -2450
rect 37710 -2510 37720 -2450
rect 37640 -2530 37720 -2510
rect 37640 -2590 37650 -2530
rect 37710 -2590 37720 -2530
rect 37640 -2600 37720 -2590
rect 37880 -2370 37960 -2360
rect 37880 -2430 37890 -2370
rect 37950 -2430 37960 -2370
rect 37880 -2450 37960 -2430
rect 37880 -2510 37890 -2450
rect 37950 -2510 37960 -2450
rect 37880 -2530 37960 -2510
rect 37880 -2590 37890 -2530
rect 37950 -2590 37960 -2530
rect 38080 -2560 38120 -2330
rect 37880 -2600 37960 -2590
rect 38060 -2580 38140 -2560
rect 35750 -2630 35810 -2610
rect 38060 -2620 38080 -2580
rect 38120 -2620 38140 -2580
rect 38060 -2640 38140 -2620
rect 35480 -3230 35490 -3170
rect 35550 -3230 35570 -3170
rect 35630 -3230 35650 -3170
rect 35710 -3230 35720 -3170
rect 35480 -3250 35720 -3230
rect 35480 -3310 35490 -3250
rect 35550 -3310 35570 -3250
rect 35630 -3310 35650 -3250
rect 35710 -3310 35720 -3250
rect 35480 -3330 35720 -3310
rect 35480 -3390 35490 -3330
rect 35550 -3390 35570 -3330
rect 35630 -3390 35650 -3330
rect 35710 -3390 35720 -3330
rect 35480 -3400 35720 -3390
rect 36900 -3170 36980 -3160
rect 36900 -3230 36910 -3170
rect 36970 -3230 36980 -3170
rect 36900 -3250 36980 -3230
rect 36900 -3310 36910 -3250
rect 36970 -3310 36980 -3250
rect 36900 -3330 36980 -3310
rect 36900 -3390 36910 -3330
rect 36970 -3390 36980 -3330
rect 36900 -3400 36980 -3390
rect 33640 -3440 33720 -3430
rect 33640 -3500 33650 -3440
rect 33710 -3500 33720 -3440
rect 33640 -3510 33720 -3500
rect 33800 -3440 33880 -3430
rect 33800 -3500 33810 -3440
rect 33870 -3500 33880 -3440
rect 33800 -3510 33880 -3500
rect 33960 -3440 34040 -3430
rect 33960 -3500 33970 -3440
rect 34030 -3500 34040 -3440
rect 33960 -3510 34040 -3500
rect 34120 -3440 34200 -3430
rect 34120 -3500 34130 -3440
rect 34190 -3500 34200 -3440
rect 34120 -3510 34200 -3500
rect 34280 -3440 34360 -3430
rect 34280 -3500 34290 -3440
rect 34350 -3500 34360 -3440
rect 34280 -3510 34360 -3500
rect 34440 -3440 34520 -3430
rect 34440 -3500 34450 -3440
rect 34510 -3500 34520 -3440
rect 34440 -3510 34520 -3500
rect 34600 -3440 34680 -3430
rect 34600 -3500 34610 -3440
rect 34670 -3500 34680 -3440
rect 34600 -3510 34680 -3500
rect 34760 -3440 34840 -3430
rect 34760 -3500 34770 -3440
rect 34830 -3500 34840 -3440
rect 34760 -3510 34840 -3500
rect 34920 -3440 35000 -3430
rect 34920 -3500 34930 -3440
rect 34990 -3500 35000 -3440
rect 34920 -3510 35000 -3500
rect 35080 -3440 35160 -3430
rect 35080 -3500 35090 -3440
rect 35150 -3500 35160 -3440
rect 35080 -3510 35160 -3500
rect 35240 -3440 35320 -3430
rect 35240 -3500 35250 -3440
rect 35310 -3500 35320 -3440
rect 35240 -3510 35320 -3500
rect 35400 -3440 35480 -3430
rect 35400 -3500 35410 -3440
rect 35470 -3500 35480 -3440
rect 35400 -3510 35480 -3500
rect 35560 -3440 35640 -3430
rect 35560 -3500 35570 -3440
rect 35630 -3500 35640 -3440
rect 35560 -3510 35640 -3500
rect 35720 -3440 35800 -3430
rect 35720 -3500 35730 -3440
rect 35790 -3500 35800 -3440
rect 35720 -3510 35800 -3500
rect 35880 -3440 35960 -3430
rect 35880 -3500 35890 -3440
rect 35950 -3500 35960 -3440
rect 35880 -3510 35960 -3500
rect 36040 -3440 36120 -3430
rect 36040 -3500 36050 -3440
rect 36110 -3500 36120 -3440
rect 36040 -3510 36120 -3500
rect 36200 -3440 36280 -3430
rect 36200 -3500 36210 -3440
rect 36270 -3500 36280 -3440
rect 36200 -3510 36280 -3500
rect 36360 -3440 36440 -3430
rect 36360 -3500 36370 -3440
rect 36430 -3500 36440 -3440
rect 36360 -3510 36440 -3500
rect 36520 -3440 36600 -3430
rect 36520 -3500 36530 -3440
rect 36590 -3500 36600 -3440
rect 36520 -3510 36600 -3500
rect 36680 -3440 36760 -3430
rect 36680 -3500 36690 -3440
rect 36750 -3500 36760 -3440
rect 36680 -3510 36760 -3500
rect 36840 -3440 36920 -3430
rect 36840 -3500 36850 -3440
rect 36910 -3500 36920 -3440
rect 36840 -3510 36920 -3500
rect 37000 -3440 37080 -3430
rect 37000 -3500 37010 -3440
rect 37070 -3500 37080 -3440
rect 37000 -3510 37080 -3500
rect 37160 -3440 37240 -3430
rect 37160 -3500 37170 -3440
rect 37230 -3500 37240 -3440
rect 37160 -3510 37240 -3500
rect 37320 -3440 37400 -3430
rect 37320 -3500 37330 -3440
rect 37390 -3500 37400 -3440
rect 37320 -3510 37400 -3500
rect 37480 -3440 37560 -3430
rect 37480 -3500 37490 -3440
rect 37550 -3500 37560 -3440
rect 37480 -3510 37560 -3500
rect 37640 -3440 37720 -3430
rect 37640 -3500 37650 -3440
rect 37710 -3500 37720 -3440
rect 37640 -3510 37720 -3500
rect 33330 -3570 33410 -3560
rect 33330 -3630 33340 -3570
rect 33400 -3630 33410 -3570
rect 33330 -3650 33410 -3630
rect 33330 -3710 33340 -3650
rect 33400 -3710 33410 -3650
rect 37720 -3610 37800 -3600
rect 37720 -3670 37730 -3610
rect 37790 -3670 37800 -3610
rect 37720 -3680 37800 -3670
rect 33330 -3720 33410 -3710
rect 37770 -3780 37850 -3770
rect 37770 -3840 37780 -3780
rect 37840 -3840 37850 -3780
rect 32990 -3890 33070 -3880
rect 32990 -3950 33000 -3890
rect 33060 -3950 33070 -3890
rect 32650 -4000 32730 -3990
rect 32650 -4060 32660 -4000
rect 32720 -4060 32730 -4000
rect 32650 -4070 32730 -4060
rect 32560 -4200 32640 -4190
rect 32560 -4260 32570 -4200
rect 32630 -4260 32640 -4200
rect 32560 -4270 32640 -4260
rect 32330 -6210 32340 -6150
rect 32400 -6210 32410 -6150
rect 32330 -6430 32410 -6210
rect 32340 -6442 32410 -6430
rect 32340 -6522 32410 -6512
rect 32990 -6640 33070 -3950
rect 34850 -4070 34860 -4000
rect 34930 -4070 34940 -4000
rect 36248 -4070 36258 -4000
rect 36328 -4070 36338 -4000
rect 37660 -4010 37740 -4000
rect 37660 -4070 37670 -4010
rect 37730 -4070 37740 -4010
rect 34850 -4120 34930 -4070
rect 34850 -4180 34860 -4120
rect 34920 -4180 34930 -4120
rect 34850 -4190 34930 -4180
rect 33110 -4200 33190 -4190
rect 33110 -4260 33120 -4200
rect 33180 -4260 33190 -4200
rect 33110 -4270 33190 -4260
rect 33460 -4200 33540 -4190
rect 33460 -4260 33470 -4200
rect 33530 -4260 33540 -4200
rect 33460 -4270 33540 -4260
rect 33130 -5790 33170 -4270
rect 33120 -5800 33190 -5790
rect 33120 -5880 33190 -5870
rect 33480 -6200 33520 -4270
rect 33890 -5230 37310 -4530
rect 33460 -6210 33540 -6200
rect 33460 -6270 33470 -6210
rect 33530 -6270 33540 -6210
rect 33460 -6280 33540 -6270
rect 33000 -6650 33070 -6640
rect 33000 -6730 33070 -6720
rect 33890 -7250 34590 -5230
rect 35250 -6210 35950 -5890
rect 35250 -6270 35570 -6210
rect 35630 -6270 35950 -6210
rect 35250 -6590 35950 -6270
rect 36610 -6210 37310 -5230
rect 36610 -6270 37240 -6210
rect 37300 -6270 37310 -6210
rect 36610 -7250 37310 -6270
rect 37660 -6210 37740 -4070
rect 37660 -6270 37670 -6210
rect 37730 -6270 37740 -6210
rect 37660 -6280 37740 -6270
rect 31950 -7790 32040 -7780
rect 31950 -7860 31960 -7790
rect 32030 -7860 32040 -7790
rect 31950 -7870 32040 -7860
rect 32340 -7788 32410 -7778
rect 32340 -7870 32410 -7858
rect 33000 -7788 33070 -7778
rect 31510 -8250 31590 -8240
rect 31510 -8310 31520 -8250
rect 31580 -8310 31590 -8250
rect 31510 -8590 31590 -8310
rect 33000 -8310 33070 -7858
rect 33360 -7938 33430 -7928
rect 33890 -7950 37310 -7250
rect 33360 -8310 33430 -8008
rect 33000 -8320 33080 -8310
rect 33000 -8380 33010 -8320
rect 33070 -8380 33080 -8320
rect 33000 -8400 33080 -8380
rect 33000 -8460 33010 -8400
rect 33070 -8460 33080 -8400
rect 33000 -8480 33080 -8460
rect 33000 -8540 33010 -8480
rect 33070 -8540 33080 -8480
rect 33000 -8550 33080 -8540
rect 33360 -8320 33440 -8310
rect 33360 -8380 33370 -8320
rect 33430 -8380 33440 -8320
rect 33360 -8400 33440 -8380
rect 33360 -8460 33370 -8400
rect 33430 -8460 33440 -8400
rect 33360 -8480 33440 -8460
rect 33360 -8540 33370 -8480
rect 33430 -8540 33440 -8480
rect 33360 -8550 33440 -8540
rect 35560 -8320 35640 -8310
rect 35560 -8380 35570 -8320
rect 35630 -8380 35640 -8320
rect 35560 -8400 35640 -8380
rect 35560 -8460 35570 -8400
rect 35630 -8460 35640 -8400
rect 35560 -8480 35640 -8460
rect 35560 -8540 35570 -8480
rect 35630 -8540 35640 -8480
rect 35560 -8550 35640 -8540
rect 31510 -8650 31520 -8590
rect 31580 -8650 31590 -8590
rect 31510 -8660 31590 -8650
rect 37770 -8660 37850 -3840
rect 38180 -3780 38260 -1510
rect 38180 -3840 38190 -3780
rect 38250 -3840 38260 -3780
rect 38180 -3850 38260 -3840
rect 38450 -2150 38530 1230
rect 38680 840 38760 850
rect 38680 780 38690 840
rect 38750 780 38760 840
rect 38450 -2210 38460 -2150
rect 38520 -2210 38530 -2150
rect 38450 -3890 38530 -2210
rect 38450 -3950 38460 -3890
rect 38520 -3950 38530 -3890
rect 38450 -3960 38530 -3950
rect 38560 -600 38640 -590
rect 38560 -660 38570 -600
rect 38630 -660 38640 -600
rect 38560 -1920 38640 -660
rect 38560 -1980 38570 -1920
rect 38630 -1980 38640 -1920
rect 38130 -4120 38210 -4110
rect 38130 -4180 38140 -4120
rect 38200 -4180 38210 -4120
rect 38130 -5790 38210 -4180
rect 38130 -5800 38200 -5790
rect 38130 -5880 38200 -5870
rect 38560 -6176 38640 -1980
rect 38680 -980 38760 780
rect 38680 -1040 38690 -980
rect 38750 -1040 38760 -980
rect 38560 -6180 38630 -6176
rect 38560 -6260 38630 -6250
rect 38680 -6230 38760 -1040
rect 38790 -490 38870 -480
rect 38790 -550 38800 -490
rect 38860 -550 38870 -490
rect 38790 -3610 38870 -550
rect 38790 -3670 38800 -3610
rect 38860 -3670 38870 -3610
rect 38790 -3680 38870 -3670
rect 38680 -6320 38750 -6300
rect 38680 -7578 38750 -7568
rect 38320 -7788 38390 -7778
rect 37890 -7938 37960 -7928
rect 37890 -8010 37960 -8008
rect 37880 -8320 37960 -8010
rect 37880 -8380 37890 -8320
rect 37950 -8380 37960 -8320
rect 37880 -8400 37960 -8380
rect 37880 -8460 37890 -8400
rect 37950 -8460 37960 -8400
rect 37880 -8480 37960 -8460
rect 37880 -8540 37890 -8480
rect 37950 -8540 37960 -8480
rect 37880 -8550 37960 -8540
rect 38310 -8320 38390 -7858
rect 38310 -8380 38320 -8320
rect 38380 -8380 38390 -8320
rect 38310 -8400 38390 -8380
rect 38310 -8460 38320 -8400
rect 38380 -8460 38390 -8400
rect 38310 -8480 38390 -8460
rect 38310 -8540 38320 -8480
rect 38380 -8540 38390 -8480
rect 38310 -8550 38390 -8540
rect 38680 -8590 38760 -7648
rect 38680 -8650 38690 -8590
rect 38750 -8650 38760 -8590
rect 38680 -8660 38760 -8650
<< via1 >>
rect 34070 1230 34130 1290
rect 34290 1230 34350 1290
rect 34510 1230 34570 1290
rect 34730 1230 34790 1290
rect 34950 1230 35010 1290
rect 35170 1230 35230 1290
rect 35970 1230 36030 1290
rect 36190 1230 36250 1290
rect 36410 1230 36470 1290
rect 36630 1230 36690 1290
rect 36850 1230 36910 1290
rect 37070 1230 37130 1290
rect 38460 1230 38520 1290
rect 33960 1170 34020 1180
rect 33960 1130 33970 1170
rect 33970 1130 34010 1170
rect 34010 1130 34020 1170
rect 33960 1120 34020 1130
rect 34180 1120 34240 1180
rect 34400 1120 34460 1180
rect 34620 1120 34680 1180
rect 34840 1120 34900 1180
rect 35060 1120 35120 1180
rect 35280 1170 35340 1180
rect 35280 1130 35290 1170
rect 35290 1130 35330 1170
rect 35330 1130 35340 1170
rect 35280 1120 35340 1130
rect 35860 1170 35920 1180
rect 35860 1130 35870 1170
rect 35870 1130 35910 1170
rect 35910 1130 35920 1170
rect 35860 1120 35920 1130
rect 36080 1120 36140 1180
rect 36300 1120 36360 1180
rect 36520 1120 36580 1180
rect 36740 1120 36800 1180
rect 36960 1120 37020 1180
rect 37180 1170 37240 1180
rect 37180 1130 37190 1170
rect 37190 1130 37230 1170
rect 37230 1130 37240 1170
rect 37180 1120 37240 1130
rect 34130 832 34182 842
rect 34130 798 34138 832
rect 34138 798 34172 832
rect 34172 798 34182 832
rect 34130 790 34182 798
rect 34240 832 34292 842
rect 34240 798 34248 832
rect 34248 798 34282 832
rect 34282 798 34292 832
rect 34240 790 34292 798
rect 34350 832 34402 842
rect 34350 798 34358 832
rect 34358 798 34392 832
rect 34392 798 34402 832
rect 34350 790 34402 798
rect 34460 832 34512 842
rect 34460 798 34468 832
rect 34468 798 34502 832
rect 34502 798 34512 832
rect 34460 790 34512 798
rect 34570 832 34622 842
rect 34570 798 34578 832
rect 34578 798 34612 832
rect 34612 798 34622 832
rect 34570 790 34622 798
rect 34680 832 34732 842
rect 34680 798 34688 832
rect 34688 798 34722 832
rect 34722 798 34732 832
rect 34680 790 34732 798
rect 34790 832 34842 842
rect 34790 798 34798 832
rect 34798 798 34832 832
rect 34832 798 34842 832
rect 34790 790 34842 798
rect 34900 832 34952 842
rect 34900 798 34908 832
rect 34908 798 34942 832
rect 34942 798 34952 832
rect 34900 790 34952 798
rect 35010 832 35062 842
rect 35010 798 35018 832
rect 35018 798 35052 832
rect 35052 798 35062 832
rect 35010 790 35062 798
rect 35120 832 35172 842
rect 35120 798 35128 832
rect 35128 798 35162 832
rect 35162 798 35172 832
rect 35120 790 35172 798
rect 36030 832 36082 842
rect 36030 798 36038 832
rect 36038 798 36072 832
rect 36072 798 36082 832
rect 36030 790 36082 798
rect 36140 832 36192 842
rect 36140 798 36148 832
rect 36148 798 36182 832
rect 36182 798 36192 832
rect 36140 790 36192 798
rect 36250 832 36302 842
rect 36250 798 36258 832
rect 36258 798 36292 832
rect 36292 798 36302 832
rect 36250 790 36302 798
rect 36360 832 36412 842
rect 36360 798 36368 832
rect 36368 798 36402 832
rect 36402 798 36412 832
rect 36360 790 36412 798
rect 36470 832 36522 842
rect 36470 798 36478 832
rect 36478 798 36512 832
rect 36512 798 36522 832
rect 36470 790 36522 798
rect 36580 832 36632 842
rect 36580 798 36588 832
rect 36588 798 36622 832
rect 36622 798 36632 832
rect 36580 790 36632 798
rect 36690 832 36742 842
rect 36690 798 36698 832
rect 36698 798 36732 832
rect 36732 798 36742 832
rect 36690 790 36742 798
rect 36800 832 36852 842
rect 36800 798 36808 832
rect 36808 798 36842 832
rect 36842 798 36852 832
rect 36800 790 36852 798
rect 36910 832 36962 842
rect 36910 798 36918 832
rect 36918 798 36952 832
rect 36952 798 36962 832
rect 36910 790 36962 798
rect 37020 832 37072 842
rect 37020 798 37028 832
rect 37028 798 37062 832
rect 37062 798 37072 832
rect 37020 790 37072 798
rect 32880 680 32940 740
rect 32880 600 32940 660
rect 32880 520 32940 580
rect 33320 680 33380 740
rect 33320 600 33380 660
rect 33320 520 33380 580
rect 33950 680 34010 740
rect 33950 600 34010 660
rect 33950 570 34010 580
rect 33950 530 33960 570
rect 33960 530 34000 570
rect 34000 530 34010 570
rect 33950 520 34010 530
rect 34310 680 34370 740
rect 34310 600 34370 660
rect 34310 570 34370 580
rect 34310 530 34320 570
rect 34320 530 34360 570
rect 34360 530 34370 570
rect 34310 520 34370 530
rect 34670 680 34730 740
rect 34670 600 34730 660
rect 34670 570 34730 580
rect 34670 530 34680 570
rect 34680 530 34720 570
rect 34720 530 34730 570
rect 34670 520 34730 530
rect 35030 680 35090 740
rect 35030 600 35090 660
rect 35030 570 35090 580
rect 35030 530 35040 570
rect 35040 530 35080 570
rect 35080 530 35090 570
rect 35030 520 35090 530
rect 35390 680 35450 740
rect 35390 600 35450 660
rect 35390 570 35450 580
rect 35390 530 35400 570
rect 35400 530 35440 570
rect 35440 530 35450 570
rect 35390 520 35450 530
rect 35750 680 35810 740
rect 35750 600 35810 660
rect 35750 570 35810 580
rect 35750 530 35760 570
rect 35760 530 35800 570
rect 35800 530 35810 570
rect 35750 520 35810 530
rect 36110 680 36170 740
rect 36110 600 36170 660
rect 36110 570 36170 580
rect 36110 530 36120 570
rect 36120 530 36160 570
rect 36160 530 36170 570
rect 36110 520 36170 530
rect 36470 680 36530 740
rect 36470 600 36530 660
rect 36470 570 36530 580
rect 36470 530 36480 570
rect 36480 530 36520 570
rect 36520 530 36530 570
rect 36470 520 36530 530
rect 36830 680 36890 740
rect 36830 600 36890 660
rect 36830 570 36890 580
rect 36830 530 36840 570
rect 36840 530 36880 570
rect 36880 530 36890 570
rect 36830 520 36890 530
rect 37190 680 37250 740
rect 37190 600 37250 660
rect 37190 570 37250 580
rect 37190 530 37200 570
rect 37200 530 37240 570
rect 37240 530 37250 570
rect 37190 520 37250 530
rect 33100 370 33160 380
rect 33100 330 33110 370
rect 33110 330 33150 370
rect 33150 330 33160 370
rect 33100 320 33160 330
rect 33570 320 33630 380
rect 32980 30 33040 40
rect 32980 -10 32990 30
rect 32990 -10 33030 30
rect 33030 -10 33040 30
rect 32980 -20 33040 -10
rect 32660 -330 32720 -270
rect 32570 -440 32630 -380
rect 32340 -1040 32400 -980
rect 32070 -1500 32130 -1440
rect 32150 -1500 32210 -1440
rect 32230 -1500 32290 -1440
rect 32070 -1580 32130 -1520
rect 32150 -1580 32210 -1520
rect 32230 -1580 32290 -1520
rect 32070 -1660 32130 -1600
rect 32150 -1660 32210 -1600
rect 32230 -1660 32290 -1600
rect 31840 -3840 31900 -3780
rect 31720 -4810 31780 -4750
rect 31720 -6210 31780 -6150
rect 31590 -6910 31650 -6850
rect 32070 -4810 32130 -4750
rect 32150 -4810 32210 -4750
rect 32230 -4810 32290 -4750
rect 31960 -5510 32020 -5450
rect 31840 -7610 31900 -7550
rect 32570 -1980 32630 -1920
rect 32850 -770 32910 -710
rect 32850 -850 32910 -790
rect 32850 -930 32910 -870
rect 33220 30 33280 40
rect 33220 -10 33230 30
rect 33230 -10 33270 30
rect 33270 -10 33280 30
rect 33220 -20 33280 -10
rect 33570 -440 33630 -380
rect 33100 -550 33160 -490
rect 34220 -170 34280 -160
rect 34220 -210 34230 -170
rect 34230 -210 34270 -170
rect 34270 -210 34280 -170
rect 34220 -220 34280 -210
rect 34400 -170 34460 -160
rect 34400 -210 34410 -170
rect 34410 -210 34450 -170
rect 34450 -210 34460 -170
rect 34400 -220 34460 -210
rect 34580 -170 34640 -160
rect 34580 -210 34590 -170
rect 34590 -210 34630 -170
rect 34630 -210 34640 -170
rect 34580 -220 34640 -210
rect 34760 -170 34820 -160
rect 34760 -210 34770 -170
rect 34770 -210 34810 -170
rect 34810 -210 34820 -170
rect 34760 -220 34820 -210
rect 34940 -170 35000 -160
rect 34940 -210 34950 -170
rect 34950 -210 34990 -170
rect 34990 -210 35000 -170
rect 34940 -220 35000 -210
rect 35120 -170 35180 -160
rect 35120 -210 35130 -170
rect 35130 -210 35170 -170
rect 35170 -210 35180 -170
rect 35120 -220 35180 -210
rect 35300 -170 35360 -160
rect 35300 -210 35310 -170
rect 35310 -210 35350 -170
rect 35350 -210 35360 -170
rect 35300 -220 35360 -210
rect 35390 -220 35450 -160
rect 35480 -170 35540 -160
rect 35480 -210 35490 -170
rect 35490 -210 35530 -170
rect 35530 -210 35540 -170
rect 35480 -220 35540 -210
rect 35210 -330 35270 -270
rect 34850 -440 34910 -380
rect 34490 -550 34550 -490
rect 34130 -660 34190 -600
rect 33090 -770 33150 -710
rect 33090 -850 33150 -790
rect 33090 -930 33150 -870
rect 33330 -770 33390 -710
rect 33330 -850 33390 -790
rect 33330 -930 33390 -870
rect 33570 -770 33630 -710
rect 33570 -850 33630 -790
rect 33570 -930 33630 -870
rect 33810 -770 33870 -710
rect 33810 -850 33870 -790
rect 33810 -930 33870 -870
rect 34050 -770 34110 -710
rect 34050 -850 34110 -790
rect 34050 -930 34110 -870
rect 34290 -770 34350 -710
rect 34290 -850 34350 -790
rect 34290 -930 34350 -870
rect 34530 -770 34590 -710
rect 34530 -850 34590 -790
rect 34530 -930 34590 -870
rect 34770 -770 34830 -710
rect 34770 -850 34830 -790
rect 34770 -930 34830 -870
rect 35010 -770 35070 -710
rect 35010 -850 35070 -790
rect 35010 -930 35070 -870
rect 35250 -770 35310 -710
rect 35250 -850 35310 -790
rect 35250 -930 35310 -870
rect 32970 -1040 33030 -980
rect 33210 -1330 33270 -1320
rect 33210 -1370 33220 -1330
rect 33220 -1370 33260 -1330
rect 33260 -1370 33270 -1330
rect 33210 -1380 33270 -1370
rect 33690 -1040 33750 -980
rect 33930 -1330 33990 -1320
rect 33930 -1370 33940 -1330
rect 33940 -1370 33980 -1330
rect 33980 -1370 33990 -1330
rect 33930 -1380 33990 -1370
rect 33030 -1500 33090 -1440
rect 33030 -1580 33090 -1520
rect 33030 -1660 33090 -1600
rect 33450 -1500 33510 -1440
rect 33450 -1580 33510 -1520
rect 33450 -1660 33510 -1600
rect 33690 -1500 33750 -1440
rect 33690 -1580 33750 -1520
rect 33690 -1660 33750 -1600
rect 33690 -1770 33750 -1710
rect 34410 -1040 34470 -980
rect 34650 -1330 34710 -1320
rect 34650 -1370 34660 -1330
rect 34660 -1370 34700 -1330
rect 34700 -1370 34710 -1330
rect 34650 -1380 34710 -1370
rect 35130 -1040 35190 -980
rect 35660 -170 35720 -160
rect 35660 -210 35670 -170
rect 35670 -210 35710 -170
rect 35710 -210 35720 -170
rect 35660 -220 35720 -210
rect 35840 -170 35900 -160
rect 35840 -210 35850 -170
rect 35850 -210 35890 -170
rect 35890 -210 35900 -170
rect 35840 -220 35900 -210
rect 36020 -170 36080 -160
rect 36020 -210 36030 -170
rect 36030 -210 36070 -170
rect 36070 -210 36080 -170
rect 36020 -220 36080 -210
rect 36200 -170 36260 -160
rect 36200 -210 36210 -170
rect 36210 -210 36250 -170
rect 36250 -210 36260 -170
rect 36200 -220 36260 -210
rect 35930 -330 35990 -270
rect 36380 -170 36440 -160
rect 36380 -210 36390 -170
rect 36390 -210 36430 -170
rect 36430 -210 36440 -170
rect 36380 -220 36440 -210
rect 36560 -170 36620 -160
rect 36560 -210 36570 -170
rect 36570 -210 36610 -170
rect 36610 -210 36620 -170
rect 36560 -220 36620 -210
rect 36290 -440 36350 -380
rect 36740 -170 36800 -160
rect 36740 -210 36750 -170
rect 36750 -210 36790 -170
rect 36790 -210 36800 -170
rect 36740 -220 36800 -210
rect 36920 -170 36980 -160
rect 36920 -210 36930 -170
rect 36930 -210 36970 -170
rect 36970 -210 36980 -170
rect 36920 -220 36980 -210
rect 36650 -550 36710 -490
rect 35570 -660 35630 -600
rect 37010 -660 37070 -600
rect 35890 -770 35950 -710
rect 35890 -850 35950 -790
rect 35890 -930 35950 -870
rect 36130 -770 36190 -710
rect 36130 -850 36190 -790
rect 36130 -930 36190 -870
rect 36370 -770 36430 -710
rect 36370 -850 36430 -790
rect 36370 -930 36430 -870
rect 36610 -770 36670 -710
rect 36610 -850 36670 -790
rect 36610 -930 36670 -870
rect 36850 -770 36910 -710
rect 36850 -850 36910 -790
rect 36850 -930 36910 -870
rect 37090 -770 37150 -710
rect 37090 -850 37150 -790
rect 37090 -930 37150 -870
rect 37330 -770 37390 -710
rect 37330 -850 37390 -790
rect 37330 -930 37390 -870
rect 37570 -770 37630 -710
rect 37570 -850 37630 -790
rect 37570 -930 37630 -870
rect 37810 -770 37870 -710
rect 37810 -850 37870 -790
rect 37810 -930 37870 -870
rect 38050 -770 38110 -710
rect 38050 -850 38110 -790
rect 38050 -930 38110 -870
rect 38290 -770 38350 -710
rect 38290 -850 38350 -790
rect 38290 -930 38350 -870
rect 35390 -1040 35450 -980
rect 35750 -1040 35810 -980
rect 34170 -1500 34230 -1440
rect 34170 -1580 34230 -1520
rect 34170 -1660 34230 -1600
rect 34410 -1500 34470 -1440
rect 34410 -1580 34470 -1520
rect 34410 -1660 34470 -1600
rect 34650 -1500 34710 -1440
rect 34650 -1580 34710 -1520
rect 34650 -1660 34710 -1600
rect 34890 -1500 34950 -1440
rect 34890 -1580 34950 -1520
rect 34890 -1660 34950 -1600
rect 35070 -1500 35130 -1440
rect 35070 -1580 35130 -1520
rect 35070 -1660 35130 -1600
rect 34170 -1770 34230 -1710
rect 34650 -1770 34710 -1710
rect 33930 -1880 33990 -1820
rect 33856 -1938 33908 -1930
rect 33856 -1972 33864 -1938
rect 33864 -1972 33898 -1938
rect 33898 -1972 33908 -1938
rect 33856 -1982 33908 -1972
rect 34014 -1938 34066 -1930
rect 34014 -1972 34022 -1938
rect 34022 -1972 34056 -1938
rect 34056 -1972 34066 -1938
rect 34014 -1982 34066 -1972
rect 34410 -1880 34470 -1820
rect 34338 -1938 34390 -1930
rect 34338 -1972 34346 -1938
rect 34346 -1972 34380 -1938
rect 34380 -1972 34390 -1938
rect 34338 -1982 34390 -1972
rect 34492 -1938 34544 -1930
rect 34492 -1972 34500 -1938
rect 34500 -1972 34534 -1938
rect 34534 -1972 34544 -1938
rect 34492 -1982 34544 -1972
rect 34890 -1880 34950 -1820
rect 34816 -1938 34868 -1930
rect 34816 -1972 34824 -1938
rect 34824 -1972 34858 -1938
rect 34858 -1972 34868 -1938
rect 34816 -1982 34868 -1972
rect 35130 -1980 35190 -1970
rect 35130 -2020 35140 -1980
rect 35140 -2020 35180 -1980
rect 35180 -2020 35190 -1980
rect 35130 -2030 35190 -2020
rect 35130 -2060 35190 -2050
rect 35130 -2100 35140 -2060
rect 35140 -2100 35180 -2060
rect 35180 -2100 35190 -2060
rect 35130 -2110 35190 -2100
rect 32660 -2210 32720 -2150
rect 33753 -2168 33805 -2158
rect 33753 -2202 33763 -2168
rect 33763 -2202 33797 -2168
rect 33797 -2202 33805 -2168
rect 33753 -2210 33805 -2202
rect 34113 -2168 34165 -2158
rect 34113 -2202 34123 -2168
rect 34123 -2202 34157 -2168
rect 34157 -2202 34165 -2168
rect 34113 -2210 34165 -2202
rect 34233 -2168 34285 -2158
rect 34233 -2202 34243 -2168
rect 34243 -2202 34277 -2168
rect 34277 -2202 34285 -2168
rect 34233 -2210 34285 -2202
rect 34593 -2168 34645 -2158
rect 34593 -2202 34603 -2168
rect 34603 -2202 34637 -2168
rect 34637 -2202 34645 -2168
rect 34593 -2210 34645 -2202
rect 34713 -2168 34765 -2158
rect 34713 -2202 34723 -2168
rect 34723 -2202 34757 -2168
rect 34757 -2202 34765 -2168
rect 34713 -2210 34765 -2202
rect 35130 -2140 35190 -2130
rect 35130 -2180 35140 -2140
rect 35140 -2180 35180 -2140
rect 35180 -2180 35190 -2140
rect 35130 -2190 35190 -2180
rect 33070 -2320 33130 -2260
rect 33820 -2320 33880 -2260
rect 34040 -2320 34100 -2260
rect 34300 -2320 34360 -2260
rect 34520 -2320 34580 -2260
rect 34780 -2320 34840 -2260
rect 33250 -2430 33310 -2370
rect 33250 -2510 33310 -2450
rect 33250 -2540 33310 -2530
rect 33250 -2580 33260 -2540
rect 33260 -2580 33300 -2540
rect 33300 -2580 33310 -2540
rect 33250 -2590 33310 -2580
rect 33490 -2430 33550 -2370
rect 33490 -2510 33550 -2450
rect 33490 -2540 33550 -2530
rect 33490 -2580 33500 -2540
rect 33500 -2580 33540 -2540
rect 33540 -2580 33550 -2540
rect 33490 -2590 33550 -2580
rect 33730 -2430 33790 -2370
rect 33730 -2510 33790 -2450
rect 33730 -2540 33790 -2530
rect 33730 -2580 33740 -2540
rect 33740 -2580 33780 -2540
rect 33780 -2580 33790 -2540
rect 33730 -2590 33790 -2580
rect 33970 -2430 34030 -2370
rect 33970 -2510 34030 -2450
rect 33970 -2540 34030 -2530
rect 33970 -2580 33980 -2540
rect 33980 -2580 34020 -2540
rect 34020 -2580 34030 -2540
rect 33970 -2590 34030 -2580
rect 34610 -2430 34670 -2370
rect 34610 -2510 34670 -2450
rect 34610 -2540 34670 -2530
rect 34610 -2580 34620 -2540
rect 34620 -2580 34660 -2540
rect 34660 -2580 34670 -2540
rect 34610 -2590 34670 -2580
rect 34850 -2430 34910 -2370
rect 34850 -2510 34910 -2450
rect 34850 -2540 34910 -2530
rect 34850 -2580 34860 -2540
rect 34860 -2580 34900 -2540
rect 34900 -2580 34910 -2540
rect 34850 -2590 34910 -2580
rect 35090 -2430 35150 -2370
rect 35090 -2510 35150 -2450
rect 35090 -2540 35150 -2530
rect 35090 -2580 35100 -2540
rect 35100 -2580 35140 -2540
rect 35140 -2580 35150 -2540
rect 35090 -2590 35150 -2580
rect 35490 -2030 35550 -1970
rect 35570 -2030 35630 -1970
rect 35650 -2030 35710 -1970
rect 35490 -2110 35550 -2050
rect 35570 -2110 35630 -2050
rect 35650 -2110 35710 -2050
rect 35490 -2190 35550 -2130
rect 35570 -2190 35630 -2130
rect 35650 -2190 35710 -2130
rect 34230 -3180 34290 -3170
rect 34230 -3220 34240 -3180
rect 34240 -3220 34280 -3180
rect 34280 -3220 34290 -3180
rect 34230 -3230 34290 -3220
rect 34230 -3310 34290 -3250
rect 34230 -3390 34290 -3330
rect 36010 -1040 36070 -980
rect 36730 -1040 36790 -980
rect 36490 -1330 36550 -1320
rect 36490 -1370 36500 -1330
rect 36500 -1370 36540 -1330
rect 36540 -1370 36550 -1330
rect 36490 -1380 36550 -1370
rect 37450 -1040 37510 -980
rect 37210 -1330 37270 -1320
rect 37210 -1370 37220 -1330
rect 37220 -1370 37260 -1330
rect 37260 -1370 37270 -1330
rect 37210 -1380 37270 -1370
rect 36070 -1500 36130 -1440
rect 36250 -1500 36310 -1440
rect 36730 -1500 36790 -1440
rect 36970 -1500 37030 -1440
rect 36490 -1770 36550 -1710
rect 36970 -1770 37030 -1710
rect 36250 -1880 36310 -1820
rect 36010 -1980 36070 -1970
rect 36010 -2020 36020 -1980
rect 36020 -2020 36060 -1980
rect 36060 -2020 36070 -1980
rect 36010 -2030 36070 -2020
rect 36332 -1938 36384 -1930
rect 36332 -1972 36342 -1938
rect 36342 -1972 36376 -1938
rect 36376 -1972 36384 -1938
rect 36332 -1982 36384 -1972
rect 36730 -1880 36790 -1820
rect 36656 -1938 36708 -1930
rect 36656 -1972 36666 -1938
rect 36666 -1972 36700 -1938
rect 36700 -1972 36708 -1938
rect 36656 -1982 36708 -1972
rect 36810 -1938 36862 -1930
rect 36810 -1972 36820 -1938
rect 36820 -1972 36854 -1938
rect 36854 -1972 36862 -1938
rect 36810 -1982 36862 -1972
rect 38170 -1040 38230 -980
rect 37930 -1330 37990 -1320
rect 37930 -1370 37940 -1330
rect 37940 -1370 37980 -1330
rect 37980 -1370 37990 -1330
rect 37930 -1380 37990 -1370
rect 37450 -1500 37510 -1440
rect 37690 -1500 37750 -1440
rect 38110 -1500 38170 -1440
rect 38190 -1500 38250 -1440
rect 37450 -1770 37510 -1710
rect 37210 -1880 37270 -1820
rect 37134 -1938 37186 -1930
rect 37134 -1972 37144 -1938
rect 37144 -1972 37178 -1938
rect 37178 -1972 37186 -1938
rect 37134 -1982 37186 -1972
rect 37292 -1938 37344 -1930
rect 37292 -1972 37302 -1938
rect 37302 -1972 37336 -1938
rect 37336 -1972 37344 -1938
rect 37292 -1982 37344 -1972
rect 36010 -2060 36070 -2050
rect 36010 -2100 36020 -2060
rect 36020 -2100 36060 -2060
rect 36060 -2100 36070 -2060
rect 36010 -2110 36070 -2100
rect 36010 -2140 36070 -2130
rect 36010 -2180 36020 -2140
rect 36020 -2180 36060 -2140
rect 36060 -2180 36070 -2140
rect 36010 -2190 36070 -2180
rect 36435 -2168 36487 -2158
rect 36435 -2202 36443 -2168
rect 36443 -2202 36477 -2168
rect 36477 -2202 36487 -2168
rect 36435 -2210 36487 -2202
rect 36555 -2168 36607 -2158
rect 36555 -2202 36563 -2168
rect 36563 -2202 36597 -2168
rect 36597 -2202 36607 -2168
rect 36555 -2210 36607 -2202
rect 36915 -2168 36967 -2158
rect 36915 -2202 36923 -2168
rect 36923 -2202 36957 -2168
rect 36957 -2202 36967 -2168
rect 36915 -2210 36967 -2202
rect 37035 -2168 37087 -2158
rect 37035 -2202 37043 -2168
rect 37043 -2202 37077 -2168
rect 37077 -2202 37087 -2168
rect 37035 -2210 37087 -2202
rect 37395 -2168 37447 -2158
rect 37395 -2202 37403 -2168
rect 37403 -2202 37437 -2168
rect 37437 -2202 37447 -2168
rect 37395 -2210 37447 -2202
rect 36360 -2320 36420 -2260
rect 36620 -2320 36680 -2260
rect 36840 -2320 36900 -2260
rect 37100 -2320 37160 -2260
rect 37320 -2320 37380 -2260
rect 38070 -2320 38130 -2260
rect 36050 -2430 36110 -2370
rect 36050 -2510 36110 -2450
rect 36050 -2540 36110 -2530
rect 36050 -2580 36060 -2540
rect 36060 -2580 36100 -2540
rect 36100 -2580 36110 -2540
rect 36050 -2590 36110 -2580
rect 36290 -2430 36350 -2370
rect 36290 -2510 36350 -2450
rect 36290 -2540 36350 -2530
rect 36290 -2580 36300 -2540
rect 36300 -2580 36340 -2540
rect 36340 -2580 36350 -2540
rect 36290 -2590 36350 -2580
rect 36530 -2430 36590 -2370
rect 36530 -2510 36590 -2450
rect 36530 -2540 36590 -2530
rect 36530 -2580 36540 -2540
rect 36540 -2580 36580 -2540
rect 36580 -2580 36590 -2540
rect 36530 -2590 36590 -2580
rect 37170 -2430 37230 -2370
rect 37170 -2510 37230 -2450
rect 37170 -2540 37230 -2530
rect 37170 -2580 37180 -2540
rect 37180 -2580 37220 -2540
rect 37220 -2580 37230 -2540
rect 37170 -2590 37230 -2580
rect 37410 -2430 37470 -2370
rect 37410 -2510 37470 -2450
rect 37410 -2540 37470 -2530
rect 37410 -2580 37420 -2540
rect 37420 -2580 37460 -2540
rect 37460 -2580 37470 -2540
rect 37410 -2590 37470 -2580
rect 37650 -2430 37710 -2370
rect 37650 -2510 37710 -2450
rect 37650 -2540 37710 -2530
rect 37650 -2580 37660 -2540
rect 37660 -2580 37700 -2540
rect 37700 -2580 37710 -2540
rect 37650 -2590 37710 -2580
rect 37890 -2430 37950 -2370
rect 37890 -2510 37950 -2450
rect 37890 -2540 37950 -2530
rect 37890 -2580 37900 -2540
rect 37900 -2580 37940 -2540
rect 37940 -2580 37950 -2540
rect 37890 -2590 37950 -2580
rect 35490 -3230 35550 -3170
rect 35570 -3230 35630 -3170
rect 35650 -3230 35710 -3170
rect 35490 -3310 35550 -3250
rect 35570 -3310 35630 -3250
rect 35650 -3310 35710 -3250
rect 35490 -3390 35550 -3330
rect 35570 -3390 35630 -3330
rect 35650 -3390 35710 -3330
rect 36910 -3180 36970 -3170
rect 36910 -3220 36920 -3180
rect 36920 -3220 36960 -3180
rect 36960 -3220 36970 -3180
rect 36910 -3230 36970 -3220
rect 36910 -3310 36970 -3250
rect 36910 -3390 36970 -3330
rect 33650 -3450 33710 -3440
rect 33650 -3490 33660 -3450
rect 33660 -3490 33700 -3450
rect 33700 -3490 33710 -3450
rect 33650 -3500 33710 -3490
rect 33810 -3450 33870 -3440
rect 33810 -3490 33820 -3450
rect 33820 -3490 33860 -3450
rect 33860 -3490 33870 -3450
rect 33810 -3500 33870 -3490
rect 33970 -3450 34030 -3440
rect 33970 -3490 33980 -3450
rect 33980 -3490 34020 -3450
rect 34020 -3490 34030 -3450
rect 33970 -3500 34030 -3490
rect 34130 -3450 34190 -3440
rect 34130 -3490 34140 -3450
rect 34140 -3490 34180 -3450
rect 34180 -3490 34190 -3450
rect 34130 -3500 34190 -3490
rect 34290 -3450 34350 -3440
rect 34290 -3490 34300 -3450
rect 34300 -3490 34340 -3450
rect 34340 -3490 34350 -3450
rect 34290 -3500 34350 -3490
rect 34450 -3450 34510 -3440
rect 34450 -3490 34460 -3450
rect 34460 -3490 34500 -3450
rect 34500 -3490 34510 -3450
rect 34450 -3500 34510 -3490
rect 34610 -3450 34670 -3440
rect 34610 -3490 34620 -3450
rect 34620 -3490 34660 -3450
rect 34660 -3490 34670 -3450
rect 34610 -3500 34670 -3490
rect 34770 -3450 34830 -3440
rect 34770 -3490 34780 -3450
rect 34780 -3490 34820 -3450
rect 34820 -3490 34830 -3450
rect 34770 -3500 34830 -3490
rect 34930 -3450 34990 -3440
rect 34930 -3490 34940 -3450
rect 34940 -3490 34980 -3450
rect 34980 -3490 34990 -3450
rect 34930 -3500 34990 -3490
rect 35090 -3450 35150 -3440
rect 35090 -3490 35100 -3450
rect 35100 -3490 35140 -3450
rect 35140 -3490 35150 -3450
rect 35090 -3500 35150 -3490
rect 35250 -3450 35310 -3440
rect 35250 -3490 35260 -3450
rect 35260 -3490 35300 -3450
rect 35300 -3490 35310 -3450
rect 35250 -3500 35310 -3490
rect 35410 -3450 35470 -3440
rect 35410 -3490 35420 -3450
rect 35420 -3490 35460 -3450
rect 35460 -3490 35470 -3450
rect 35410 -3500 35470 -3490
rect 35570 -3450 35630 -3440
rect 35570 -3490 35580 -3450
rect 35580 -3490 35620 -3450
rect 35620 -3490 35630 -3450
rect 35570 -3500 35630 -3490
rect 35730 -3450 35790 -3440
rect 35730 -3490 35740 -3450
rect 35740 -3490 35780 -3450
rect 35780 -3490 35790 -3450
rect 35730 -3500 35790 -3490
rect 35890 -3450 35950 -3440
rect 35890 -3490 35900 -3450
rect 35900 -3490 35940 -3450
rect 35940 -3490 35950 -3450
rect 35890 -3500 35950 -3490
rect 36050 -3450 36110 -3440
rect 36050 -3490 36060 -3450
rect 36060 -3490 36100 -3450
rect 36100 -3490 36110 -3450
rect 36050 -3500 36110 -3490
rect 36210 -3450 36270 -3440
rect 36210 -3490 36220 -3450
rect 36220 -3490 36260 -3450
rect 36260 -3490 36270 -3450
rect 36210 -3500 36270 -3490
rect 36370 -3450 36430 -3440
rect 36370 -3490 36380 -3450
rect 36380 -3490 36420 -3450
rect 36420 -3490 36430 -3450
rect 36370 -3500 36430 -3490
rect 36530 -3450 36590 -3440
rect 36530 -3490 36540 -3450
rect 36540 -3490 36580 -3450
rect 36580 -3490 36590 -3450
rect 36530 -3500 36590 -3490
rect 36690 -3450 36750 -3440
rect 36690 -3490 36700 -3450
rect 36700 -3490 36740 -3450
rect 36740 -3490 36750 -3450
rect 36690 -3500 36750 -3490
rect 36850 -3450 36910 -3440
rect 36850 -3490 36860 -3450
rect 36860 -3490 36900 -3450
rect 36900 -3490 36910 -3450
rect 36850 -3500 36910 -3490
rect 37010 -3450 37070 -3440
rect 37010 -3490 37020 -3450
rect 37020 -3490 37060 -3450
rect 37060 -3490 37070 -3450
rect 37010 -3500 37070 -3490
rect 37170 -3450 37230 -3440
rect 37170 -3490 37180 -3450
rect 37180 -3490 37220 -3450
rect 37220 -3490 37230 -3450
rect 37170 -3500 37230 -3490
rect 37330 -3450 37390 -3440
rect 37330 -3490 37340 -3450
rect 37340 -3490 37380 -3450
rect 37380 -3490 37390 -3450
rect 37330 -3500 37390 -3490
rect 37490 -3450 37550 -3440
rect 37490 -3490 37500 -3450
rect 37500 -3490 37540 -3450
rect 37540 -3490 37550 -3450
rect 37490 -3500 37550 -3490
rect 37650 -3450 37710 -3440
rect 37650 -3490 37660 -3450
rect 37660 -3490 37700 -3450
rect 37700 -3490 37710 -3450
rect 37650 -3500 37710 -3490
rect 33340 -3580 33400 -3570
rect 33340 -3620 33350 -3580
rect 33350 -3620 33390 -3580
rect 33390 -3620 33400 -3580
rect 33340 -3630 33400 -3620
rect 33340 -3660 33400 -3650
rect 33340 -3700 33350 -3660
rect 33350 -3700 33390 -3660
rect 33390 -3700 33400 -3660
rect 33340 -3710 33400 -3700
rect 37730 -3620 37790 -3610
rect 37730 -3660 37740 -3620
rect 37740 -3660 37780 -3620
rect 37780 -3660 37790 -3620
rect 37730 -3670 37790 -3660
rect 37780 -3840 37840 -3780
rect 33000 -3950 33060 -3890
rect 32660 -4060 32720 -4000
rect 32570 -4260 32630 -4200
rect 32340 -6210 32400 -6150
rect 32340 -6452 32410 -6442
rect 32340 -6502 32350 -6452
rect 32350 -6502 32400 -6452
rect 32400 -6502 32410 -6452
rect 32340 -6512 32410 -6502
rect 34860 -4010 34930 -4000
rect 34860 -4060 34870 -4010
rect 34870 -4060 34920 -4010
rect 34920 -4060 34930 -4010
rect 34860 -4070 34930 -4060
rect 36258 -4010 36328 -4000
rect 36258 -4060 36268 -4010
rect 36268 -4060 36318 -4010
rect 36318 -4060 36328 -4010
rect 36258 -4070 36328 -4060
rect 37670 -4070 37730 -4010
rect 34860 -4180 34920 -4120
rect 33120 -4260 33180 -4200
rect 33470 -4260 33530 -4200
rect 33120 -5810 33190 -5800
rect 33120 -5860 33130 -5810
rect 33130 -5860 33180 -5810
rect 33180 -5860 33190 -5810
rect 33120 -5870 33190 -5860
rect 33470 -6270 33530 -6210
rect 33000 -6660 33070 -6650
rect 33000 -6710 33010 -6660
rect 33010 -6710 33060 -6660
rect 33060 -6710 33070 -6660
rect 33000 -6720 33070 -6710
rect 35570 -6270 35630 -6210
rect 37240 -6270 37300 -6210
rect 37670 -6270 37730 -6210
rect 31960 -7860 32030 -7790
rect 32340 -7798 32410 -7788
rect 32340 -7848 32350 -7798
rect 32350 -7848 32400 -7798
rect 32400 -7848 32410 -7798
rect 32340 -7858 32410 -7848
rect 33000 -7798 33070 -7788
rect 33000 -7848 33010 -7798
rect 33010 -7848 33060 -7798
rect 33060 -7848 33070 -7798
rect 33000 -7858 33070 -7848
rect 31520 -8310 31580 -8250
rect 33360 -7948 33430 -7938
rect 33360 -7998 33370 -7948
rect 33370 -7998 33420 -7948
rect 33420 -7998 33430 -7948
rect 33360 -8008 33430 -7998
rect 33010 -8380 33070 -8320
rect 33010 -8460 33070 -8400
rect 33010 -8540 33070 -8480
rect 33370 -8380 33430 -8320
rect 33370 -8460 33430 -8400
rect 33370 -8540 33430 -8480
rect 35570 -8330 35630 -8320
rect 35570 -8370 35580 -8330
rect 35580 -8370 35620 -8330
rect 35620 -8370 35630 -8330
rect 35570 -8380 35630 -8370
rect 35570 -8410 35630 -8400
rect 35570 -8450 35580 -8410
rect 35580 -8450 35620 -8410
rect 35620 -8450 35630 -8410
rect 35570 -8460 35630 -8450
rect 35570 -8490 35630 -8480
rect 35570 -8530 35580 -8490
rect 35580 -8530 35620 -8490
rect 35620 -8530 35630 -8490
rect 35570 -8540 35630 -8530
rect 31520 -8650 31580 -8590
rect 38190 -3840 38250 -3780
rect 38690 780 38750 840
rect 38460 -2210 38520 -2150
rect 38460 -3950 38520 -3890
rect 38570 -660 38630 -600
rect 38570 -1980 38630 -1920
rect 38140 -4180 38200 -4120
rect 38130 -5810 38200 -5800
rect 38130 -5860 38140 -5810
rect 38140 -5860 38190 -5810
rect 38190 -5860 38200 -5810
rect 38130 -5870 38200 -5860
rect 38690 -1040 38750 -980
rect 38560 -6190 38630 -6180
rect 38560 -6240 38570 -6190
rect 38570 -6240 38620 -6190
rect 38620 -6240 38630 -6190
rect 38560 -6250 38630 -6240
rect 38800 -550 38860 -490
rect 38800 -3670 38860 -3610
rect 38680 -6240 38750 -6230
rect 38680 -6290 38690 -6240
rect 38690 -6290 38740 -6240
rect 38740 -6290 38750 -6240
rect 38680 -6300 38750 -6290
rect 38680 -7588 38750 -7578
rect 38680 -7638 38690 -7588
rect 38690 -7638 38740 -7588
rect 38740 -7638 38750 -7588
rect 38680 -7648 38750 -7638
rect 38320 -7798 38390 -7788
rect 38320 -7848 38330 -7798
rect 38330 -7848 38380 -7798
rect 38380 -7848 38390 -7798
rect 38320 -7858 38390 -7848
rect 37890 -7948 37960 -7938
rect 37890 -7998 37900 -7948
rect 37900 -7998 37950 -7948
rect 37950 -7998 37960 -7948
rect 37890 -8008 37960 -7998
rect 37890 -8380 37950 -8320
rect 37890 -8460 37950 -8400
rect 37890 -8540 37950 -8480
rect 38320 -8380 38380 -8320
rect 38320 -8460 38380 -8400
rect 38320 -8540 38380 -8480
rect 38690 -8650 38750 -8590
<< metal2 >>
rect 34060 1290 35240 1300
rect 34060 1230 34070 1290
rect 34130 1230 34290 1290
rect 34350 1230 34510 1290
rect 34570 1230 34730 1290
rect 34790 1230 34950 1290
rect 35010 1230 35170 1290
rect 35230 1230 35240 1290
rect 34060 1220 35240 1230
rect 35960 1290 38530 1300
rect 35960 1230 35970 1290
rect 36030 1230 36190 1290
rect 36250 1230 36410 1290
rect 36470 1230 36630 1290
rect 36690 1230 36850 1290
rect 36910 1230 37070 1290
rect 37130 1230 38460 1290
rect 38520 1230 38530 1290
rect 35960 1220 38530 1230
rect 32870 1180 37250 1190
rect 32870 1120 33960 1180
rect 34020 1120 34180 1180
rect 34240 1120 34400 1180
rect 34460 1120 34620 1180
rect 34680 1120 34840 1180
rect 34900 1120 35060 1180
rect 35120 1120 35280 1180
rect 35340 1120 35860 1180
rect 35920 1120 36080 1180
rect 36140 1120 36300 1180
rect 36360 1120 36520 1180
rect 36580 1120 36740 1180
rect 36800 1120 36960 1180
rect 37020 1120 37180 1180
rect 37240 1120 37250 1180
rect 32870 1110 37250 1120
rect 34126 842 38760 850
rect 34126 790 34130 842
rect 34182 790 34240 842
rect 34292 790 34350 842
rect 34402 790 34460 842
rect 34512 790 34570 842
rect 34622 790 34680 842
rect 34732 790 34790 842
rect 34842 790 34900 842
rect 34952 790 35010 842
rect 35062 790 35120 842
rect 35172 790 36030 842
rect 36082 790 36140 842
rect 36192 790 36250 842
rect 36302 790 36360 842
rect 36412 790 36470 842
rect 36522 790 36580 842
rect 36632 790 36690 842
rect 36742 790 36800 842
rect 36852 790 36910 842
rect 36962 790 37020 842
rect 37072 840 38760 842
rect 37072 790 38690 840
rect 34126 780 38690 790
rect 38750 780 38760 840
rect 32870 740 37260 750
rect 32870 680 32880 740
rect 32940 680 33320 740
rect 33380 680 33950 740
rect 34010 680 34310 740
rect 34370 680 34670 740
rect 34730 680 35030 740
rect 35090 680 35390 740
rect 35450 680 35750 740
rect 35810 680 36110 740
rect 36170 680 36470 740
rect 36530 680 36830 740
rect 36890 680 37190 740
rect 37250 680 37260 740
rect 32870 660 37260 680
rect 32870 600 32880 660
rect 32940 600 33320 660
rect 33380 600 33950 660
rect 34010 600 34310 660
rect 34370 600 34670 660
rect 34730 600 35030 660
rect 35090 600 35390 660
rect 35450 600 35750 660
rect 35810 600 36110 660
rect 36170 600 36470 660
rect 36530 600 36830 660
rect 36890 600 37190 660
rect 37250 600 37260 660
rect 32870 580 37260 600
rect 32870 520 32880 580
rect 32940 520 33320 580
rect 33380 520 33950 580
rect 34010 520 34310 580
rect 34370 520 34670 580
rect 34730 520 35030 580
rect 35090 520 35390 580
rect 35450 520 35750 580
rect 35810 520 36110 580
rect 36170 520 36470 580
rect 36530 520 36830 580
rect 36890 520 37190 580
rect 37250 520 37260 580
rect 32870 510 37260 520
rect 33090 380 33170 390
rect 33090 320 33100 380
rect 33160 370 33170 380
rect 33560 380 33640 390
rect 33560 370 33570 380
rect 33160 330 33570 370
rect 33160 320 33170 330
rect 33090 310 33170 320
rect 33560 320 33570 330
rect 33630 320 33640 380
rect 33560 310 33640 320
rect 32970 40 33290 50
rect 32970 -20 32980 40
rect 33040 -20 33220 40
rect 33280 -20 33290 40
rect 32970 -30 33290 -20
rect 34220 -160 36980 -150
rect 34280 -220 34400 -160
rect 34460 -220 34580 -160
rect 34640 -220 34760 -160
rect 34820 -220 34940 -160
rect 35000 -220 35120 -160
rect 35180 -220 35300 -160
rect 35360 -220 35390 -160
rect 35450 -220 35480 -160
rect 35540 -220 35660 -160
rect 35720 -220 35840 -160
rect 35900 -220 36020 -160
rect 36080 -220 36200 -160
rect 36260 -220 36380 -160
rect 36440 -220 36560 -160
rect 36620 -220 36740 -160
rect 36800 -220 36920 -160
rect 34220 -230 36980 -220
rect 32650 -270 36000 -260
rect 32650 -330 32660 -270
rect 32720 -330 35210 -270
rect 35270 -330 35930 -270
rect 35990 -330 36000 -270
rect 32650 -340 36000 -330
rect 32560 -380 36360 -370
rect 32560 -440 32570 -380
rect 32630 -440 33570 -380
rect 33630 -440 34850 -380
rect 34910 -440 36290 -380
rect 36350 -440 36360 -380
rect 32560 -450 36360 -440
rect 33090 -490 38870 -480
rect 33090 -550 33100 -490
rect 33160 -550 34490 -490
rect 34550 -550 36650 -490
rect 36710 -550 38800 -490
rect 38860 -550 38870 -490
rect 33090 -560 38870 -550
rect 34120 -600 38640 -590
rect 34120 -660 34130 -600
rect 34190 -660 35570 -600
rect 35630 -660 37010 -600
rect 37070 -660 38570 -600
rect 38630 -660 38640 -600
rect 34120 -670 38640 -660
rect 32840 -710 38360 -700
rect 32840 -770 32850 -710
rect 32910 -770 33090 -710
rect 33150 -770 33330 -710
rect 33390 -770 33570 -710
rect 33630 -770 33810 -710
rect 33870 -770 34050 -710
rect 34110 -770 34290 -710
rect 34350 -770 34530 -710
rect 34590 -770 34770 -710
rect 34830 -770 35010 -710
rect 35070 -770 35250 -710
rect 35310 -770 35890 -710
rect 35950 -770 36130 -710
rect 36190 -770 36370 -710
rect 36430 -770 36610 -710
rect 36670 -770 36850 -710
rect 36910 -770 37090 -710
rect 37150 -770 37330 -710
rect 37390 -770 37570 -710
rect 37630 -770 37810 -710
rect 37870 -770 38050 -710
rect 38110 -770 38290 -710
rect 38350 -770 38360 -710
rect 32840 -790 38360 -770
rect 32840 -850 32850 -790
rect 32910 -850 33090 -790
rect 33150 -850 33330 -790
rect 33390 -850 33570 -790
rect 33630 -850 33810 -790
rect 33870 -850 34050 -790
rect 34110 -850 34290 -790
rect 34350 -850 34530 -790
rect 34590 -850 34770 -790
rect 34830 -850 35010 -790
rect 35070 -850 35250 -790
rect 35310 -850 35890 -790
rect 35950 -850 36130 -790
rect 36190 -850 36370 -790
rect 36430 -850 36610 -790
rect 36670 -850 36850 -790
rect 36910 -850 37090 -790
rect 37150 -850 37330 -790
rect 37390 -850 37570 -790
rect 37630 -850 37810 -790
rect 37870 -850 38050 -790
rect 38110 -850 38290 -790
rect 38350 -850 38360 -790
rect 32840 -870 38360 -850
rect 32840 -930 32850 -870
rect 32910 -930 33090 -870
rect 33150 -930 33330 -870
rect 33390 -930 33570 -870
rect 33630 -930 33810 -870
rect 33870 -930 34050 -870
rect 34110 -930 34290 -870
rect 34350 -930 34530 -870
rect 34590 -930 34770 -870
rect 34830 -930 35010 -870
rect 35070 -930 35250 -870
rect 35310 -930 35890 -870
rect 35950 -930 36130 -870
rect 36190 -930 36370 -870
rect 36430 -930 36610 -870
rect 36670 -930 36850 -870
rect 36910 -930 37090 -870
rect 37150 -930 37330 -870
rect 37390 -930 37570 -870
rect 37630 -930 37810 -870
rect 37870 -930 38050 -870
rect 38110 -930 38290 -870
rect 38350 -930 38360 -870
rect 32840 -940 38360 -930
rect 32330 -980 35460 -970
rect 32330 -1040 32340 -980
rect 32400 -1040 32970 -980
rect 33030 -1040 33690 -980
rect 33750 -1040 34410 -980
rect 34470 -1040 35130 -980
rect 35190 -1040 35390 -980
rect 35450 -1040 35460 -980
rect 32330 -1050 35460 -1040
rect 35740 -980 38760 -970
rect 35740 -1040 35750 -980
rect 35810 -1040 36010 -980
rect 36070 -1040 36730 -980
rect 36790 -1040 37450 -980
rect 37510 -1040 38170 -980
rect 38230 -1040 38690 -980
rect 38750 -1040 38760 -980
rect 35740 -1050 38760 -1040
rect 33690 -1090 33750 -1050
rect 37450 -1080 37510 -1050
rect 33200 -1320 33280 -1310
rect 33200 -1380 33210 -1320
rect 33270 -1330 33280 -1320
rect 33920 -1320 34000 -1310
rect 33920 -1330 33930 -1320
rect 33270 -1370 33930 -1330
rect 33270 -1380 33280 -1370
rect 33200 -1390 33280 -1380
rect 33920 -1380 33930 -1370
rect 33990 -1330 34000 -1320
rect 34640 -1320 34720 -1310
rect 34640 -1330 34650 -1320
rect 33990 -1370 34650 -1330
rect 33990 -1380 34000 -1370
rect 33920 -1390 34000 -1380
rect 34640 -1380 34650 -1370
rect 34710 -1380 34720 -1320
rect 34640 -1390 34720 -1380
rect 36480 -1320 36560 -1310
rect 36480 -1380 36490 -1320
rect 36550 -1330 36560 -1320
rect 37200 -1320 37280 -1310
rect 37200 -1330 37210 -1320
rect 36550 -1370 37210 -1330
rect 36550 -1380 36560 -1370
rect 36480 -1390 36560 -1380
rect 37200 -1380 37210 -1370
rect 37270 -1330 37280 -1320
rect 37920 -1320 38000 -1310
rect 37920 -1330 37930 -1320
rect 37270 -1370 37930 -1330
rect 37270 -1380 37280 -1370
rect 37200 -1390 37280 -1380
rect 37920 -1380 37930 -1370
rect 37990 -1380 38000 -1320
rect 37920 -1390 38000 -1380
rect 32060 -1440 35140 -1430
rect 32060 -1500 32070 -1440
rect 32130 -1500 32150 -1440
rect 32210 -1500 32230 -1440
rect 32290 -1500 33030 -1440
rect 33090 -1500 33450 -1440
rect 33510 -1500 33690 -1440
rect 33750 -1500 34170 -1440
rect 34230 -1500 34410 -1440
rect 34470 -1500 34650 -1440
rect 34710 -1500 34890 -1440
rect 34950 -1500 35070 -1440
rect 35130 -1500 35140 -1440
rect 32060 -1520 35140 -1500
rect 36060 -1440 38260 -1430
rect 36060 -1500 36070 -1440
rect 36130 -1500 36250 -1440
rect 36310 -1500 36730 -1440
rect 36790 -1500 36970 -1440
rect 37030 -1500 37450 -1440
rect 37510 -1500 37690 -1440
rect 37750 -1500 38110 -1440
rect 38170 -1500 38190 -1440
rect 38250 -1500 38260 -1440
rect 36060 -1510 38260 -1500
rect 32060 -1580 32070 -1520
rect 32130 -1580 32150 -1520
rect 32210 -1580 32230 -1520
rect 32290 -1580 33030 -1520
rect 33090 -1580 33450 -1520
rect 33510 -1580 33690 -1520
rect 33750 -1580 34170 -1520
rect 34230 -1580 34410 -1520
rect 34470 -1580 34650 -1520
rect 34710 -1580 34890 -1520
rect 34950 -1580 35070 -1520
rect 35130 -1580 35140 -1520
rect 32060 -1600 35140 -1580
rect 32060 -1660 32070 -1600
rect 32130 -1660 32150 -1600
rect 32210 -1660 32230 -1600
rect 32290 -1660 33030 -1600
rect 33090 -1660 33450 -1600
rect 33510 -1660 33690 -1600
rect 33750 -1660 34170 -1600
rect 34230 -1660 34410 -1600
rect 34470 -1660 34650 -1600
rect 34710 -1660 34890 -1600
rect 34950 -1660 35070 -1600
rect 35130 -1660 35140 -1600
rect 32060 -1670 35140 -1660
rect 33680 -1710 34720 -1700
rect 33680 -1770 33690 -1710
rect 33750 -1770 34170 -1710
rect 34230 -1770 34650 -1710
rect 34710 -1770 34720 -1710
rect 33680 -1780 34720 -1770
rect 36480 -1710 37520 -1700
rect 36480 -1770 36490 -1710
rect 36550 -1770 36970 -1710
rect 37030 -1770 37450 -1710
rect 37510 -1770 37520 -1710
rect 36480 -1780 37520 -1770
rect 33920 -1820 34960 -1810
rect 33920 -1880 33930 -1820
rect 33990 -1880 34410 -1820
rect 34470 -1880 34890 -1820
rect 34950 -1880 34960 -1820
rect 33920 -1890 34960 -1880
rect 36240 -1820 37280 -1810
rect 36240 -1880 36250 -1820
rect 36310 -1880 36730 -1820
rect 36790 -1880 37210 -1820
rect 37270 -1880 37280 -1820
rect 36240 -1890 37280 -1880
rect 32560 -1920 32640 -1910
rect 38560 -1920 38640 -1910
rect 32560 -1980 32570 -1920
rect 32630 -1930 34870 -1920
rect 32630 -1980 33856 -1930
rect 32560 -1982 33856 -1980
rect 33908 -1982 34014 -1930
rect 34066 -1982 34338 -1930
rect 34390 -1982 34492 -1930
rect 34544 -1982 34816 -1930
rect 34868 -1982 34870 -1930
rect 36330 -1930 38570 -1920
rect 32560 -1990 34870 -1982
rect 35120 -1970 36080 -1960
rect 35120 -2030 35130 -1970
rect 35190 -2030 35490 -1970
rect 35550 -2030 35570 -1970
rect 35630 -2030 35650 -1970
rect 35710 -2030 36010 -1970
rect 36070 -2030 36080 -1970
rect 36330 -1982 36332 -1930
rect 36384 -1982 36656 -1930
rect 36708 -1982 36810 -1930
rect 36862 -1982 37134 -1930
rect 37186 -1982 37292 -1930
rect 37344 -1980 38570 -1930
rect 38630 -1980 38640 -1920
rect 37344 -1982 38640 -1980
rect 36330 -1990 38640 -1982
rect 35120 -2050 36080 -2030
rect 35120 -2110 35130 -2050
rect 35190 -2110 35490 -2050
rect 35550 -2110 35570 -2050
rect 35630 -2110 35650 -2050
rect 35710 -2110 36010 -2050
rect 36070 -2110 36080 -2050
rect 35120 -2130 36080 -2110
rect 32650 -2150 32730 -2140
rect 32650 -2210 32660 -2150
rect 32720 -2158 34769 -2150
rect 32720 -2210 33753 -2158
rect 33805 -2210 34113 -2158
rect 34165 -2210 34233 -2158
rect 34285 -2210 34593 -2158
rect 34645 -2210 34713 -2158
rect 34765 -2210 34769 -2158
rect 35120 -2190 35130 -2130
rect 35190 -2190 35490 -2130
rect 35550 -2190 35570 -2130
rect 35630 -2190 35650 -2130
rect 35710 -2190 36010 -2130
rect 36070 -2190 36080 -2130
rect 38450 -2150 38530 -2140
rect 35120 -2200 36080 -2190
rect 36431 -2158 38460 -2150
rect 32650 -2220 34769 -2210
rect 36431 -2210 36435 -2158
rect 36487 -2210 36555 -2158
rect 36607 -2210 36915 -2158
rect 36967 -2210 37035 -2158
rect 37087 -2210 37395 -2158
rect 37447 -2210 38460 -2158
rect 38520 -2210 38530 -2150
rect 36431 -2220 38530 -2210
rect 33060 -2260 34850 -2250
rect 33060 -2320 33070 -2260
rect 33130 -2320 33820 -2260
rect 33880 -2320 34040 -2260
rect 34100 -2320 34300 -2260
rect 34360 -2320 34520 -2260
rect 34580 -2320 34780 -2260
rect 34840 -2320 34850 -2260
rect 33060 -2330 34850 -2320
rect 36350 -2260 38140 -2250
rect 36350 -2320 36360 -2260
rect 36420 -2320 36620 -2260
rect 36680 -2320 36840 -2260
rect 36900 -2320 37100 -2260
rect 37160 -2320 37320 -2260
rect 37380 -2320 38070 -2260
rect 38130 -2320 38140 -2260
rect 36350 -2330 38140 -2320
rect 33240 -2370 37960 -2360
rect 33240 -2430 33250 -2370
rect 33310 -2430 33490 -2370
rect 33550 -2430 33730 -2370
rect 33790 -2430 33970 -2370
rect 34030 -2430 34610 -2370
rect 34670 -2430 34850 -2370
rect 34910 -2430 35090 -2370
rect 35150 -2430 36050 -2370
rect 36110 -2430 36290 -2370
rect 36350 -2430 36530 -2370
rect 36590 -2430 37170 -2370
rect 37230 -2430 37410 -2370
rect 37470 -2430 37650 -2370
rect 37710 -2430 37890 -2370
rect 37950 -2430 37960 -2370
rect 33240 -2450 37960 -2430
rect 33240 -2510 33250 -2450
rect 33310 -2510 33490 -2450
rect 33550 -2510 33730 -2450
rect 33790 -2510 33970 -2450
rect 34030 -2510 34610 -2450
rect 34670 -2510 34850 -2450
rect 34910 -2510 35090 -2450
rect 35150 -2510 36050 -2450
rect 36110 -2510 36290 -2450
rect 36350 -2510 36530 -2450
rect 36590 -2510 37170 -2450
rect 37230 -2510 37410 -2450
rect 37470 -2510 37650 -2450
rect 37710 -2510 37890 -2450
rect 37950 -2510 37960 -2450
rect 33240 -2530 37960 -2510
rect 33240 -2590 33250 -2530
rect 33310 -2590 33490 -2530
rect 33550 -2590 33730 -2530
rect 33790 -2590 33970 -2530
rect 34030 -2590 34610 -2530
rect 34670 -2590 34850 -2530
rect 34910 -2590 35090 -2530
rect 35150 -2590 36050 -2530
rect 36110 -2590 36290 -2530
rect 36350 -2590 36530 -2530
rect 36590 -2590 37170 -2530
rect 37230 -2590 37410 -2530
rect 37470 -2590 37650 -2530
rect 37710 -2590 37890 -2530
rect 37950 -2590 37960 -2530
rect 33240 -2600 37960 -2590
rect 34220 -3170 36980 -3160
rect 34220 -3230 34230 -3170
rect 34290 -3230 35490 -3170
rect 35550 -3230 35570 -3170
rect 35630 -3230 35650 -3170
rect 35710 -3230 36910 -3170
rect 36970 -3230 36980 -3170
rect 34220 -3250 36980 -3230
rect 34220 -3310 34230 -3250
rect 34290 -3310 35490 -3250
rect 35550 -3310 35570 -3250
rect 35630 -3310 35650 -3250
rect 35710 -3310 36910 -3250
rect 36970 -3310 36980 -3250
rect 34220 -3330 36980 -3310
rect 34220 -3390 34230 -3330
rect 34290 -3390 35490 -3330
rect 35550 -3390 35570 -3330
rect 35630 -3390 35650 -3330
rect 35710 -3390 36910 -3330
rect 36970 -3390 36980 -3330
rect 34220 -3400 36980 -3390
rect 33640 -3440 33720 -3430
rect 33640 -3500 33650 -3440
rect 33710 -3450 33720 -3440
rect 33800 -3440 33880 -3430
rect 33800 -3450 33810 -3440
rect 33710 -3490 33810 -3450
rect 33710 -3500 33720 -3490
rect 33640 -3510 33720 -3500
rect 33800 -3500 33810 -3490
rect 33870 -3450 33880 -3440
rect 33960 -3440 34040 -3430
rect 33960 -3450 33970 -3440
rect 33870 -3490 33970 -3450
rect 33870 -3500 33880 -3490
rect 33800 -3510 33880 -3500
rect 33960 -3500 33970 -3490
rect 34030 -3450 34040 -3440
rect 34120 -3440 34200 -3430
rect 34120 -3450 34130 -3440
rect 34030 -3490 34130 -3450
rect 34030 -3500 34040 -3490
rect 33960 -3510 34040 -3500
rect 34120 -3500 34130 -3490
rect 34190 -3450 34200 -3440
rect 34280 -3440 34360 -3430
rect 34280 -3450 34290 -3440
rect 34190 -3490 34290 -3450
rect 34190 -3500 34200 -3490
rect 34120 -3510 34200 -3500
rect 34280 -3500 34290 -3490
rect 34350 -3450 34360 -3440
rect 34440 -3440 34520 -3430
rect 34440 -3450 34450 -3440
rect 34350 -3490 34450 -3450
rect 34350 -3500 34360 -3490
rect 34280 -3510 34360 -3500
rect 34440 -3500 34450 -3490
rect 34510 -3450 34520 -3440
rect 34600 -3440 34680 -3430
rect 34600 -3450 34610 -3440
rect 34510 -3490 34610 -3450
rect 34510 -3500 34520 -3490
rect 34440 -3510 34520 -3500
rect 34600 -3500 34610 -3490
rect 34670 -3450 34680 -3440
rect 34760 -3440 34840 -3430
rect 34760 -3450 34770 -3440
rect 34670 -3490 34770 -3450
rect 34670 -3500 34680 -3490
rect 34600 -3510 34680 -3500
rect 34760 -3500 34770 -3490
rect 34830 -3450 34840 -3440
rect 34920 -3440 35000 -3430
rect 34920 -3450 34930 -3440
rect 34830 -3490 34930 -3450
rect 34830 -3500 34840 -3490
rect 34760 -3510 34840 -3500
rect 34920 -3500 34930 -3490
rect 34990 -3450 35000 -3440
rect 35080 -3440 35160 -3430
rect 35080 -3450 35090 -3440
rect 34990 -3490 35090 -3450
rect 34990 -3500 35000 -3490
rect 34920 -3510 35000 -3500
rect 35080 -3500 35090 -3490
rect 35150 -3450 35160 -3440
rect 35240 -3440 35320 -3430
rect 35240 -3450 35250 -3440
rect 35150 -3490 35250 -3450
rect 35150 -3500 35160 -3490
rect 35080 -3510 35160 -3500
rect 35240 -3500 35250 -3490
rect 35310 -3450 35320 -3440
rect 35400 -3440 35480 -3430
rect 35400 -3450 35410 -3440
rect 35310 -3490 35410 -3450
rect 35310 -3500 35320 -3490
rect 35240 -3510 35320 -3500
rect 35400 -3500 35410 -3490
rect 35470 -3450 35480 -3440
rect 35560 -3440 35640 -3430
rect 35560 -3450 35570 -3440
rect 35470 -3490 35570 -3450
rect 35470 -3500 35480 -3490
rect 35400 -3510 35480 -3500
rect 35560 -3500 35570 -3490
rect 35630 -3500 35640 -3440
rect 35560 -3510 35640 -3500
rect 35720 -3440 35800 -3430
rect 35720 -3500 35730 -3440
rect 35790 -3450 35800 -3440
rect 35880 -3440 35960 -3430
rect 35880 -3450 35890 -3440
rect 35790 -3490 35890 -3450
rect 35790 -3500 35800 -3490
rect 35720 -3510 35800 -3500
rect 35880 -3500 35890 -3490
rect 35950 -3450 35960 -3440
rect 36040 -3440 36120 -3430
rect 36040 -3450 36050 -3440
rect 35950 -3490 36050 -3450
rect 35950 -3500 35960 -3490
rect 35880 -3510 35960 -3500
rect 36040 -3500 36050 -3490
rect 36110 -3450 36120 -3440
rect 36200 -3440 36280 -3430
rect 36200 -3450 36210 -3440
rect 36110 -3490 36210 -3450
rect 36110 -3500 36120 -3490
rect 36040 -3510 36120 -3500
rect 36200 -3500 36210 -3490
rect 36270 -3450 36280 -3440
rect 36360 -3440 36440 -3430
rect 36360 -3450 36370 -3440
rect 36270 -3490 36370 -3450
rect 36270 -3500 36280 -3490
rect 36200 -3510 36280 -3500
rect 36360 -3500 36370 -3490
rect 36430 -3450 36440 -3440
rect 36520 -3440 36600 -3430
rect 36520 -3450 36530 -3440
rect 36430 -3490 36530 -3450
rect 36430 -3500 36440 -3490
rect 36360 -3510 36440 -3500
rect 36520 -3500 36530 -3490
rect 36590 -3450 36600 -3440
rect 36680 -3440 36760 -3430
rect 36680 -3450 36690 -3440
rect 36590 -3490 36690 -3450
rect 36590 -3500 36600 -3490
rect 36520 -3510 36600 -3500
rect 36680 -3500 36690 -3490
rect 36750 -3450 36760 -3440
rect 36840 -3440 36920 -3430
rect 36840 -3450 36850 -3440
rect 36750 -3490 36850 -3450
rect 36750 -3500 36760 -3490
rect 36680 -3510 36760 -3500
rect 36840 -3500 36850 -3490
rect 36910 -3450 36920 -3440
rect 37000 -3440 37080 -3430
rect 37000 -3450 37010 -3440
rect 36910 -3490 37010 -3450
rect 36910 -3500 36920 -3490
rect 36840 -3510 36920 -3500
rect 37000 -3500 37010 -3490
rect 37070 -3450 37080 -3440
rect 37160 -3440 37240 -3430
rect 37160 -3450 37170 -3440
rect 37070 -3490 37170 -3450
rect 37070 -3500 37080 -3490
rect 37000 -3510 37080 -3500
rect 37160 -3500 37170 -3490
rect 37230 -3450 37240 -3440
rect 37320 -3440 37400 -3430
rect 37320 -3450 37330 -3440
rect 37230 -3490 37330 -3450
rect 37230 -3500 37240 -3490
rect 37160 -3510 37240 -3500
rect 37320 -3500 37330 -3490
rect 37390 -3450 37400 -3440
rect 37480 -3440 37560 -3430
rect 37480 -3450 37490 -3440
rect 37390 -3490 37490 -3450
rect 37390 -3500 37400 -3490
rect 37320 -3510 37400 -3500
rect 37480 -3500 37490 -3490
rect 37550 -3450 37560 -3440
rect 37640 -3440 37720 -3430
rect 37640 -3450 37650 -3440
rect 37550 -3490 37650 -3450
rect 37550 -3500 37560 -3490
rect 37480 -3510 37560 -3500
rect 37640 -3500 37650 -3490
rect 37710 -3500 37720 -3440
rect 37640 -3510 37720 -3500
rect 33330 -3570 33410 -3560
rect 33330 -3630 33340 -3570
rect 33400 -3630 33410 -3570
rect 33330 -3650 33410 -3630
rect 33330 -3710 33340 -3650
rect 33400 -3710 33410 -3650
rect 37720 -3610 38870 -3600
rect 37720 -3670 37730 -3610
rect 37790 -3670 38800 -3610
rect 38860 -3670 38870 -3610
rect 37720 -3680 38870 -3670
rect 33330 -3720 33410 -3710
rect 31830 -3780 38260 -3770
rect 31830 -3840 31840 -3780
rect 31900 -3840 37780 -3780
rect 37840 -3840 38190 -3780
rect 38250 -3840 38260 -3780
rect 31830 -3850 38260 -3840
rect 32990 -3890 38530 -3880
rect 32990 -3950 33000 -3890
rect 33060 -3950 38460 -3890
rect 38520 -3950 38530 -3890
rect 32990 -3960 38530 -3950
rect 32650 -4000 32730 -3990
rect 32650 -4060 32660 -4000
rect 32720 -4010 32730 -4000
rect 34850 -4010 34860 -4000
rect 32720 -4050 34860 -4010
rect 32720 -4060 32730 -4050
rect 32650 -4070 32730 -4060
rect 34850 -4070 34860 -4050
rect 34930 -4070 34940 -4000
rect 36248 -4070 36258 -4000
rect 36328 -4010 37740 -4000
rect 36328 -4070 37670 -4010
rect 37730 -4070 37740 -4010
rect 36330 -4080 37740 -4070
rect 34850 -4120 38210 -4110
rect 34850 -4180 34860 -4120
rect 34920 -4180 38140 -4120
rect 38200 -4180 38210 -4120
rect 34850 -4190 38210 -4180
rect 32560 -4200 32640 -4190
rect 32560 -4260 32570 -4200
rect 32630 -4210 32640 -4200
rect 33110 -4200 33190 -4190
rect 33110 -4210 33120 -4200
rect 32630 -4250 33120 -4210
rect 32630 -4260 32640 -4250
rect 32560 -4270 32640 -4260
rect 33110 -4260 33120 -4250
rect 33180 -4210 33190 -4200
rect 33460 -4200 33540 -4190
rect 33460 -4210 33470 -4200
rect 33180 -4250 33470 -4210
rect 33180 -4260 33190 -4250
rect 33110 -4270 33190 -4260
rect 33460 -4260 33470 -4250
rect 33530 -4260 33540 -4200
rect 33460 -4270 33540 -4260
rect 31700 -4750 32300 -4730
rect 31700 -4810 31720 -4750
rect 31780 -4810 32070 -4750
rect 32130 -4810 32150 -4750
rect 32210 -4810 32230 -4750
rect 32290 -4810 32300 -4750
rect 31700 -4830 32300 -4810
rect 31510 -5450 32030 -5440
rect 31510 -5510 31520 -5450
rect 31580 -5510 31960 -5450
rect 32020 -5510 32030 -5450
rect 31510 -5520 32030 -5510
rect 33120 -5800 33190 -5790
rect 33120 -5880 33190 -5870
rect 38130 -5800 38200 -5790
rect 38130 -5880 38200 -5870
rect 31700 -6150 32410 -6130
rect 31700 -6210 31720 -6150
rect 31780 -6210 32340 -6150
rect 32400 -6210 32410 -6150
rect 38560 -6180 38630 -6170
rect 31700 -6230 32410 -6210
rect 33460 -6210 35640 -6200
rect 33460 -6270 33470 -6210
rect 33530 -6270 35570 -6210
rect 35630 -6270 35640 -6210
rect 33460 -6280 35640 -6270
rect 37230 -6210 37740 -6200
rect 37230 -6270 37240 -6210
rect 37300 -6270 37670 -6210
rect 37730 -6270 37740 -6210
rect 38560 -6260 38630 -6250
rect 38680 -6230 38750 -6220
rect 37230 -6280 37740 -6270
rect 38680 -6320 38750 -6300
rect 32340 -6442 32410 -6430
rect 32340 -6522 32410 -6512
rect 33000 -6650 33070 -6640
rect 33000 -6730 33070 -6720
rect 31580 -6850 31660 -6840
rect 31580 -6910 31590 -6850
rect 31650 -6910 31660 -6850
rect 31580 -6920 31660 -6910
rect 31820 -7550 31920 -7530
rect 31820 -7610 31840 -7550
rect 31900 -7610 31920 -7550
rect 31820 -7630 31920 -7610
rect 38680 -7578 38750 -7568
rect 38680 -7658 38750 -7648
rect 38700 -7660 38740 -7658
rect 32340 -7780 32410 -7778
rect 31950 -7788 32410 -7780
rect 31950 -7790 32340 -7788
rect 31950 -7860 31960 -7790
rect 32030 -7858 32340 -7790
rect 32030 -7860 32410 -7858
rect 31950 -7870 32410 -7860
rect 33000 -7788 33070 -7778
rect 33000 -7868 33070 -7858
rect 38320 -7788 38390 -7778
rect 38320 -7868 38390 -7858
rect 33020 -7870 33060 -7868
rect 38330 -7870 38370 -7868
rect 33360 -7938 33430 -7928
rect 33360 -8018 33430 -8008
rect 37890 -7938 37960 -7928
rect 37890 -8018 37960 -8008
rect 33380 -8020 33420 -8018
rect 37900 -8020 37940 -8018
rect 31510 -8250 31590 -8240
rect 31510 -8310 31520 -8250
rect 31580 -8310 31590 -8250
rect 31510 -8320 31590 -8310
rect 33000 -8320 38390 -8310
rect 33000 -8380 33010 -8320
rect 33070 -8380 33370 -8320
rect 33430 -8380 35570 -8320
rect 35630 -8380 37890 -8320
rect 37950 -8380 38320 -8320
rect 38380 -8380 38390 -8320
rect 33000 -8400 38390 -8380
rect 33000 -8460 33010 -8400
rect 33070 -8460 33370 -8400
rect 33430 -8460 35570 -8400
rect 35630 -8460 37890 -8400
rect 37950 -8460 38320 -8400
rect 38380 -8460 38390 -8400
rect 33000 -8480 38390 -8460
rect 33000 -8540 33010 -8480
rect 33070 -8540 33370 -8480
rect 33430 -8540 35570 -8480
rect 35630 -8540 37890 -8480
rect 37950 -8540 38320 -8480
rect 38380 -8540 38390 -8480
rect 33000 -8550 38390 -8540
rect 31510 -8590 38760 -8580
rect 31510 -8650 31520 -8590
rect 31580 -8650 38690 -8590
rect 38750 -8650 38760 -8590
rect 31510 -8660 38760 -8650
<< via2 >>
rect 31720 -4810 31780 -4750
rect 31520 -5510 31580 -5450
rect 31720 -6210 31780 -6150
rect 31590 -6910 31650 -6850
rect 31840 -7610 31900 -7550
rect 31520 -8310 31580 -8250
<< metal3 >>
rect 24700 -4730 25160 -4540
rect 25400 -4730 25860 -4540
rect 26100 -4730 26560 -4540
rect 26800 -4730 27260 -4540
rect 27500 -4730 27960 -4540
rect 28200 -4730 28660 -4540
rect 28900 -4730 29360 -4540
rect 29600 -4730 30060 -4540
rect 30300 -4730 30760 -4540
rect 31000 -4730 31460 -4540
rect 24700 -4830 31460 -4730
rect 31700 -4740 31800 -4730
rect 31700 -4820 31710 -4740
rect 31790 -4820 31800 -4740
rect 31700 -4830 31800 -4820
rect 24700 -5000 25160 -4830
rect 25400 -5000 25860 -4830
rect 26100 -5000 26560 -4830
rect 26800 -5000 27260 -4830
rect 27500 -5000 27960 -4830
rect 28200 -5000 28660 -4830
rect 28900 -5000 29360 -4830
rect 29600 -5000 30060 -4830
rect 30300 -5000 30760 -4830
rect 31000 -5000 31460 -4830
rect 24880 -5240 24980 -5000
rect 24700 -5430 25160 -5240
rect 25400 -5430 25860 -5240
rect 26100 -5430 26560 -5240
rect 26800 -5430 27260 -5240
rect 27500 -5430 27960 -5240
rect 28200 -5430 28660 -5240
rect 28900 -5430 29360 -5240
rect 29600 -5430 30060 -5240
rect 30300 -5430 30760 -5240
rect 31000 -5430 31460 -5240
rect 24700 -5440 31460 -5430
rect 24700 -5450 31590 -5440
rect 24700 -5510 31520 -5450
rect 31580 -5510 31590 -5450
rect 24700 -5520 31590 -5510
rect 24700 -5530 31460 -5520
rect 24700 -5700 25160 -5530
rect 25400 -5700 25860 -5530
rect 26100 -5700 26560 -5530
rect 26800 -5700 27260 -5530
rect 27500 -5700 27960 -5530
rect 28200 -5700 28660 -5530
rect 28900 -5700 29360 -5530
rect 29600 -5700 30060 -5530
rect 30300 -5700 30760 -5530
rect 31000 -5700 31460 -5530
rect 24700 -6130 25160 -5940
rect 25400 -6130 25860 -5940
rect 26100 -6130 26560 -5940
rect 26800 -6130 27260 -5940
rect 27500 -6130 27960 -5940
rect 28200 -6130 28660 -5940
rect 28900 -6130 29360 -5940
rect 29600 -6130 30060 -5940
rect 30300 -6130 30760 -5940
rect 31000 -6130 31460 -5940
rect 24700 -6230 31460 -6130
rect 31700 -6140 31800 -6130
rect 31700 -6220 31710 -6140
rect 31790 -6220 31800 -6140
rect 31700 -6230 31800 -6220
rect 24700 -6400 25160 -6230
rect 25400 -6400 25860 -6230
rect 26100 -6400 26560 -6230
rect 26800 -6400 27260 -6230
rect 27500 -6400 27960 -6230
rect 28200 -6400 28660 -6230
rect 28900 -6400 29360 -6230
rect 29600 -6400 30060 -6230
rect 30300 -6400 30760 -6230
rect 31000 -6400 31460 -6230
rect 24880 -6640 24980 -6400
rect 24700 -6830 25160 -6640
rect 25400 -6830 25860 -6640
rect 26100 -6830 26560 -6640
rect 26800 -6830 27260 -6640
rect 27500 -6830 27960 -6640
rect 28200 -6830 28660 -6640
rect 28900 -6830 29360 -6640
rect 29600 -6830 30060 -6640
rect 30300 -6830 30760 -6640
rect 31000 -6830 31460 -6640
rect 24700 -6840 31460 -6830
rect 24700 -6850 31660 -6840
rect 24700 -6910 31590 -6850
rect 31650 -6910 31660 -6850
rect 24700 -6920 31660 -6910
rect 24700 -6930 31460 -6920
rect 24700 -7100 25160 -6930
rect 25400 -7100 25860 -6930
rect 26100 -7100 26560 -6930
rect 26800 -7100 27260 -6930
rect 27500 -7100 27960 -6930
rect 28200 -7100 28660 -6930
rect 28900 -7100 29360 -6930
rect 29600 -7100 30060 -6930
rect 30300 -7100 30760 -6930
rect 31000 -7100 31460 -6930
rect 24700 -7530 25160 -7340
rect 25400 -7530 25860 -7340
rect 26100 -7530 26560 -7340
rect 26800 -7530 27260 -7340
rect 27500 -7530 27960 -7340
rect 28200 -7530 28660 -7340
rect 28900 -7530 29360 -7340
rect 29600 -7530 30060 -7340
rect 30300 -7530 30760 -7340
rect 31000 -7530 31460 -7340
rect 24700 -7630 31460 -7530
rect 31820 -7540 31920 -7530
rect 31820 -7620 31830 -7540
rect 31910 -7620 31920 -7540
rect 31820 -7630 31920 -7620
rect 24700 -7800 25160 -7630
rect 25400 -7800 25860 -7630
rect 26100 -7800 26560 -7630
rect 26800 -7800 27260 -7630
rect 27500 -7800 27960 -7630
rect 28200 -7800 28660 -7630
rect 28900 -7800 29360 -7630
rect 29600 -7800 30060 -7630
rect 30300 -7800 30760 -7630
rect 31000 -7800 31460 -7630
rect 24880 -8040 24980 -7800
rect 24700 -8230 25160 -8040
rect 25400 -8230 25860 -8040
rect 26100 -8230 26560 -8040
rect 26800 -8230 27260 -8040
rect 27500 -8230 27960 -8040
rect 28200 -8230 28660 -8040
rect 28900 -8230 29360 -8040
rect 29600 -8230 30060 -8040
rect 30300 -8230 30760 -8040
rect 31000 -8230 31460 -8040
rect 24700 -8240 31460 -8230
rect 24700 -8250 31590 -8240
rect 24700 -8310 31520 -8250
rect 31580 -8310 31590 -8250
rect 24700 -8320 31590 -8310
rect 24700 -8330 31460 -8320
rect 24700 -8500 25160 -8330
rect 25400 -8500 25860 -8330
rect 26100 -8500 26560 -8330
rect 26800 -8500 27260 -8330
rect 27500 -8500 27960 -8330
rect 28200 -8500 28660 -8330
rect 28900 -8500 29360 -8330
rect 29600 -8500 30060 -8330
rect 30300 -8500 30760 -8330
rect 31000 -8500 31460 -8330
<< via3 >>
rect 31710 -4750 31790 -4740
rect 31710 -4810 31720 -4750
rect 31720 -4810 31780 -4750
rect 31780 -4810 31790 -4750
rect 31710 -4820 31790 -4810
rect 31710 -6150 31790 -6140
rect 31710 -6210 31720 -6150
rect 31720 -6210 31780 -6150
rect 31780 -6210 31790 -6150
rect 31710 -6220 31790 -6210
rect 31830 -7550 31910 -7540
rect 31830 -7610 31840 -7550
rect 31840 -7610 31900 -7550
rect 31900 -7610 31910 -7550
rect 31830 -7620 31910 -7610
<< mimcap >>
rect 24730 -4740 25130 -4570
rect 24730 -4820 24890 -4740
rect 24970 -4820 25130 -4740
rect 24730 -4970 25130 -4820
rect 25430 -4740 25830 -4570
rect 25430 -4820 25590 -4740
rect 25670 -4820 25830 -4740
rect 25430 -4970 25830 -4820
rect 26130 -4740 26530 -4570
rect 26130 -4820 26290 -4740
rect 26370 -4820 26530 -4740
rect 26130 -4970 26530 -4820
rect 26830 -4740 27230 -4570
rect 26830 -4820 26990 -4740
rect 27070 -4820 27230 -4740
rect 26830 -4970 27230 -4820
rect 27530 -4740 27930 -4570
rect 27530 -4820 27690 -4740
rect 27770 -4820 27930 -4740
rect 27530 -4970 27930 -4820
rect 28230 -4740 28630 -4570
rect 28230 -4820 28390 -4740
rect 28470 -4820 28630 -4740
rect 28230 -4970 28630 -4820
rect 28930 -4740 29330 -4570
rect 28930 -4820 29090 -4740
rect 29170 -4820 29330 -4740
rect 28930 -4970 29330 -4820
rect 29630 -4740 30030 -4570
rect 29630 -4820 29790 -4740
rect 29870 -4820 30030 -4740
rect 29630 -4970 30030 -4820
rect 30330 -4740 30730 -4570
rect 30330 -4820 30490 -4740
rect 30570 -4820 30730 -4740
rect 30330 -4970 30730 -4820
rect 31030 -4740 31430 -4570
rect 31030 -4820 31180 -4740
rect 31260 -4820 31430 -4740
rect 31030 -4970 31430 -4820
rect 24730 -5440 25130 -5270
rect 24730 -5520 24890 -5440
rect 24970 -5520 25130 -5440
rect 24730 -5670 25130 -5520
rect 25430 -5440 25830 -5270
rect 25430 -5520 25590 -5440
rect 25670 -5520 25830 -5440
rect 25430 -5670 25830 -5520
rect 26130 -5440 26530 -5270
rect 26130 -5520 26290 -5440
rect 26370 -5520 26530 -5440
rect 26130 -5670 26530 -5520
rect 26830 -5440 27230 -5270
rect 26830 -5520 26990 -5440
rect 27070 -5520 27230 -5440
rect 26830 -5670 27230 -5520
rect 27530 -5440 27930 -5270
rect 27530 -5520 27690 -5440
rect 27770 -5520 27930 -5440
rect 27530 -5670 27930 -5520
rect 28230 -5440 28630 -5270
rect 28230 -5520 28390 -5440
rect 28470 -5520 28630 -5440
rect 28230 -5670 28630 -5520
rect 28930 -5440 29330 -5270
rect 28930 -5520 29090 -5440
rect 29170 -5520 29330 -5440
rect 28930 -5670 29330 -5520
rect 29630 -5440 30030 -5270
rect 29630 -5520 29790 -5440
rect 29870 -5520 30030 -5440
rect 29630 -5670 30030 -5520
rect 30330 -5440 30730 -5270
rect 30330 -5520 30490 -5440
rect 30570 -5520 30730 -5440
rect 30330 -5670 30730 -5520
rect 31030 -5440 31430 -5270
rect 31030 -5520 31180 -5440
rect 31260 -5520 31430 -5440
rect 31030 -5670 31430 -5520
rect 24730 -6140 25130 -5970
rect 24730 -6220 24890 -6140
rect 24970 -6220 25130 -6140
rect 24730 -6370 25130 -6220
rect 25430 -6140 25830 -5970
rect 25430 -6220 25590 -6140
rect 25670 -6220 25830 -6140
rect 25430 -6370 25830 -6220
rect 26130 -6140 26530 -5970
rect 26130 -6220 26290 -6140
rect 26370 -6220 26530 -6140
rect 26130 -6370 26530 -6220
rect 26830 -6140 27230 -5970
rect 26830 -6220 26990 -6140
rect 27070 -6220 27230 -6140
rect 26830 -6370 27230 -6220
rect 27530 -6140 27930 -5970
rect 27530 -6220 27690 -6140
rect 27770 -6220 27930 -6140
rect 27530 -6370 27930 -6220
rect 28230 -6140 28630 -5970
rect 28230 -6220 28390 -6140
rect 28470 -6220 28630 -6140
rect 28230 -6370 28630 -6220
rect 28930 -6140 29330 -5970
rect 28930 -6220 29090 -6140
rect 29170 -6220 29330 -6140
rect 28930 -6370 29330 -6220
rect 29630 -6140 30030 -5970
rect 29630 -6220 29790 -6140
rect 29870 -6220 30030 -6140
rect 29630 -6370 30030 -6220
rect 30330 -6140 30730 -5970
rect 30330 -6220 30490 -6140
rect 30570 -6220 30730 -6140
rect 30330 -6370 30730 -6220
rect 31030 -6140 31430 -5970
rect 31030 -6220 31180 -6140
rect 31260 -6220 31430 -6140
rect 31030 -6370 31430 -6220
rect 24730 -6840 25130 -6670
rect 24730 -6920 24890 -6840
rect 24970 -6920 25130 -6840
rect 24730 -7070 25130 -6920
rect 25430 -6840 25830 -6670
rect 25430 -6920 25590 -6840
rect 25670 -6920 25830 -6840
rect 25430 -7070 25830 -6920
rect 26130 -6840 26530 -6670
rect 26130 -6920 26290 -6840
rect 26370 -6920 26530 -6840
rect 26130 -7070 26530 -6920
rect 26830 -6840 27230 -6670
rect 26830 -6920 26990 -6840
rect 27070 -6920 27230 -6840
rect 26830 -7070 27230 -6920
rect 27530 -6840 27930 -6670
rect 27530 -6920 27690 -6840
rect 27770 -6920 27930 -6840
rect 27530 -7070 27930 -6920
rect 28230 -6840 28630 -6670
rect 28230 -6920 28390 -6840
rect 28470 -6920 28630 -6840
rect 28230 -7070 28630 -6920
rect 28930 -6840 29330 -6670
rect 28930 -6920 29090 -6840
rect 29170 -6920 29330 -6840
rect 28930 -7070 29330 -6920
rect 29630 -6840 30030 -6670
rect 29630 -6920 29790 -6840
rect 29870 -6920 30030 -6840
rect 29630 -7070 30030 -6920
rect 30330 -6840 30730 -6670
rect 30330 -6920 30490 -6840
rect 30570 -6920 30730 -6840
rect 30330 -7070 30730 -6920
rect 31030 -6840 31430 -6670
rect 31030 -6920 31180 -6840
rect 31260 -6920 31430 -6840
rect 31030 -7070 31430 -6920
rect 24730 -7540 25130 -7370
rect 24730 -7620 24890 -7540
rect 24970 -7620 25130 -7540
rect 24730 -7770 25130 -7620
rect 25430 -7540 25830 -7370
rect 25430 -7620 25590 -7540
rect 25670 -7620 25830 -7540
rect 25430 -7770 25830 -7620
rect 26130 -7540 26530 -7370
rect 26130 -7620 26290 -7540
rect 26370 -7620 26530 -7540
rect 26130 -7770 26530 -7620
rect 26830 -7540 27230 -7370
rect 26830 -7620 26990 -7540
rect 27070 -7620 27230 -7540
rect 26830 -7770 27230 -7620
rect 27530 -7540 27930 -7370
rect 27530 -7620 27690 -7540
rect 27770 -7620 27930 -7540
rect 27530 -7770 27930 -7620
rect 28230 -7540 28630 -7370
rect 28230 -7620 28390 -7540
rect 28470 -7620 28630 -7540
rect 28230 -7770 28630 -7620
rect 28930 -7540 29330 -7370
rect 28930 -7620 29090 -7540
rect 29170 -7620 29330 -7540
rect 28930 -7770 29330 -7620
rect 29630 -7540 30030 -7370
rect 29630 -7620 29790 -7540
rect 29870 -7620 30030 -7540
rect 29630 -7770 30030 -7620
rect 30330 -7540 30730 -7370
rect 30330 -7620 30490 -7540
rect 30570 -7620 30730 -7540
rect 30330 -7770 30730 -7620
rect 31030 -7540 31430 -7370
rect 31030 -7620 31180 -7540
rect 31260 -7620 31430 -7540
rect 31030 -7770 31430 -7620
rect 24730 -8240 25130 -8070
rect 24730 -8320 24890 -8240
rect 24970 -8320 25130 -8240
rect 24730 -8470 25130 -8320
rect 25430 -8240 25830 -8070
rect 25430 -8320 25590 -8240
rect 25670 -8320 25830 -8240
rect 25430 -8470 25830 -8320
rect 26130 -8240 26530 -8070
rect 26130 -8320 26290 -8240
rect 26370 -8320 26530 -8240
rect 26130 -8470 26530 -8320
rect 26830 -8240 27230 -8070
rect 26830 -8320 26990 -8240
rect 27070 -8320 27230 -8240
rect 26830 -8470 27230 -8320
rect 27530 -8240 27930 -8070
rect 27530 -8320 27690 -8240
rect 27770 -8320 27930 -8240
rect 27530 -8470 27930 -8320
rect 28230 -8240 28630 -8070
rect 28230 -8320 28390 -8240
rect 28470 -8320 28630 -8240
rect 28230 -8470 28630 -8320
rect 28930 -8240 29330 -8070
rect 28930 -8320 29090 -8240
rect 29170 -8320 29330 -8240
rect 28930 -8470 29330 -8320
rect 29630 -8240 30030 -8070
rect 29630 -8320 29790 -8240
rect 29870 -8320 30030 -8240
rect 29630 -8470 30030 -8320
rect 30330 -8240 30730 -8070
rect 30330 -8320 30490 -8240
rect 30570 -8320 30730 -8240
rect 30330 -8470 30730 -8320
rect 31030 -8240 31430 -8070
rect 31030 -8320 31180 -8240
rect 31260 -8320 31430 -8240
rect 31030 -8470 31430 -8320
<< mimcapcontact >>
rect 24890 -4820 24970 -4740
rect 25590 -4820 25670 -4740
rect 26290 -4820 26370 -4740
rect 26990 -4820 27070 -4740
rect 27690 -4820 27770 -4740
rect 28390 -4820 28470 -4740
rect 29090 -4820 29170 -4740
rect 29790 -4820 29870 -4740
rect 30490 -4820 30570 -4740
rect 31180 -4820 31260 -4740
rect 24890 -5520 24970 -5440
rect 25590 -5520 25670 -5440
rect 26290 -5520 26370 -5440
rect 26990 -5520 27070 -5440
rect 27690 -5520 27770 -5440
rect 28390 -5520 28470 -5440
rect 29090 -5520 29170 -5440
rect 29790 -5520 29870 -5440
rect 30490 -5520 30570 -5440
rect 31180 -5520 31260 -5440
rect 24890 -6220 24970 -6140
rect 25590 -6220 25670 -6140
rect 26290 -6220 26370 -6140
rect 26990 -6220 27070 -6140
rect 27690 -6220 27770 -6140
rect 28390 -6220 28470 -6140
rect 29090 -6220 29170 -6140
rect 29790 -6220 29870 -6140
rect 30490 -6220 30570 -6140
rect 31180 -6220 31260 -6140
rect 24890 -6920 24970 -6840
rect 25590 -6920 25670 -6840
rect 26290 -6920 26370 -6840
rect 26990 -6920 27070 -6840
rect 27690 -6920 27770 -6840
rect 28390 -6920 28470 -6840
rect 29090 -6920 29170 -6840
rect 29790 -6920 29870 -6840
rect 30490 -6920 30570 -6840
rect 31180 -6920 31260 -6840
rect 24890 -7620 24970 -7540
rect 25590 -7620 25670 -7540
rect 26290 -7620 26370 -7540
rect 26990 -7620 27070 -7540
rect 27690 -7620 27770 -7540
rect 28390 -7620 28470 -7540
rect 29090 -7620 29170 -7540
rect 29790 -7620 29870 -7540
rect 30490 -7620 30570 -7540
rect 31180 -7620 31260 -7540
rect 24890 -8320 24970 -8240
rect 25590 -8320 25670 -8240
rect 26290 -8320 26370 -8240
rect 26990 -8320 27070 -8240
rect 27690 -8320 27770 -8240
rect 28390 -8320 28470 -8240
rect 29090 -8320 29170 -8240
rect 29790 -8320 29870 -8240
rect 30490 -8320 30570 -8240
rect 31180 -8320 31260 -8240
<< metal4 >>
rect 24880 -4740 31800 -4730
rect 24880 -4820 24890 -4740
rect 24970 -4820 25590 -4740
rect 25670 -4820 26290 -4740
rect 26370 -4820 26990 -4740
rect 27070 -4820 27690 -4740
rect 27770 -4820 28390 -4740
rect 28470 -4820 29090 -4740
rect 29170 -4820 29790 -4740
rect 29870 -4820 30490 -4740
rect 30570 -4820 31180 -4740
rect 31260 -4820 31710 -4740
rect 31790 -4820 31800 -4740
rect 24880 -4830 31800 -4820
rect 24880 -5430 24980 -4830
rect 24880 -5440 31270 -5430
rect 24880 -5520 24890 -5440
rect 24970 -5520 25590 -5440
rect 25670 -5520 26290 -5440
rect 26370 -5520 26990 -5440
rect 27070 -5520 27690 -5440
rect 27770 -5520 28390 -5440
rect 28470 -5520 29090 -5440
rect 29170 -5520 29790 -5440
rect 29870 -5520 30490 -5440
rect 30570 -5520 31180 -5440
rect 31260 -5520 31270 -5440
rect 24880 -5530 31270 -5520
rect 24880 -6140 31800 -6130
rect 24880 -6220 24890 -6140
rect 24970 -6220 25590 -6140
rect 25670 -6220 26290 -6140
rect 26370 -6220 26990 -6140
rect 27070 -6220 27690 -6140
rect 27770 -6220 28390 -6140
rect 28470 -6220 29090 -6140
rect 29170 -6220 29790 -6140
rect 29870 -6220 30490 -6140
rect 30570 -6220 31180 -6140
rect 31260 -6220 31710 -6140
rect 31790 -6220 31800 -6140
rect 24880 -6230 31800 -6220
rect 24880 -6830 24980 -6230
rect 24880 -6840 31270 -6830
rect 24880 -6920 24890 -6840
rect 24970 -6920 25590 -6840
rect 25670 -6920 26290 -6840
rect 26370 -6920 26990 -6840
rect 27070 -6920 27690 -6840
rect 27770 -6920 28390 -6840
rect 28470 -6920 29090 -6840
rect 29170 -6920 29790 -6840
rect 29870 -6920 30490 -6840
rect 30570 -6920 31180 -6840
rect 31260 -6920 31270 -6840
rect 24880 -6930 31270 -6920
rect 24880 -7540 31920 -7530
rect 24880 -7620 24890 -7540
rect 24970 -7620 25590 -7540
rect 25670 -7620 26290 -7540
rect 26370 -7620 26990 -7540
rect 27070 -7620 27690 -7540
rect 27770 -7620 28390 -7540
rect 28470 -7620 29090 -7540
rect 29170 -7620 29790 -7540
rect 29870 -7620 30490 -7540
rect 30570 -7620 31180 -7540
rect 31260 -7620 31830 -7540
rect 31910 -7620 31920 -7540
rect 24880 -7630 31920 -7620
rect 24880 -8230 24980 -7630
rect 24880 -8240 31270 -8230
rect 24880 -8320 24890 -8240
rect 24970 -8320 25590 -8240
rect 25670 -8320 26290 -8240
rect 26370 -8320 26990 -8240
rect 27070 -8320 27690 -8240
rect 27770 -8320 28390 -8240
rect 28470 -8320 29090 -8240
rect 29170 -8320 29790 -8240
rect 29870 -8320 30490 -8240
rect 30570 -8320 31180 -8240
rect 31260 -8320 31270 -8240
rect 24880 -8330 31270 -8320
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8 $PDKPATH/libs.ref/sky130_fd_pr/mag
timestamp 1723858470
transform 1 0 36290 0 1 -5550
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_18
timestamp 1723858470
transform 1 0 33570 0 1 -5550
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_19
timestamp 1723858470
transform 1 0 34930 0 1 -5550
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_20
timestamp 1723858470
transform 1 0 36290 0 1 -8270
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_21
timestamp 1723858470
transform 1 0 36290 0 1 -6910
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_22
timestamp 1723858470
transform 1 0 34930 0 1 -8270
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_23
timestamp 1723858470
transform 1 0 34930 0 1 -6910
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_24
timestamp 1723858470
transform 1 0 33570 0 1 -8270
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25
timestamp 1723858470
transform 1 0 33570 0 1 -6910
box 0 0 1340 1340
<< labels >>
flabel metal2 31790 -8660 31790 -8660 5 FreeSans 800 0 0 -400 cap_res2
flabel metal2 31710 -5440 31710 -5440 1 FreeSans 800 0 0 400 cap_res1
flabel metal2 34370 -2330 34370 -2330 3 FreeSans 800 0 400 0 V_p_1
flabel metal2 36910 -2330 36910 -2330 3 FreeSans 800 180 400 0 V_p_2
flabel metal2 32780 -1970 32780 -1970 5 FreeSans 800 0 0 -160 Vin-
flabel metal2 32790 -2180 32790 -2180 1 FreeSans 800 0 0 160 Vin+
flabel metal2 36860 -170 36860 -170 5 FreeSans 800 0 0 -80 V_TOP
flabel metal2 35140 -1470 35140 -1470 3 FreeSans 480 0 240 0 1st_Vout_1
flabel metal2 33240 -1390 33240 -1390 5 FreeSans 800 0 0 -80 V_mir1
flabel metal2 36060 -1470 36060 -1470 7 FreeSans 480 0 -240 0 1st_Vout_2
flabel metal2 38140 -590 38140 -590 1 FreeSans 640 0 0 320 V1
flabel metal1 38760 -1450 38760 -1450 3 FreeSans 640 0 320 0 V2
flabel metal1 34760 1300 34760 1300 1 FreeSans 1600 0 800 0 CURRENT_OUTPUT
port 2 n
flabel metal1 33640 -3470 33640 -3470 7 FreeSans 800 180 -400 0 START_UP_NFET1
flabel metal2 38360 -2160 38360 -2160 1 FreeSans 800 0 0 160 V_CUR_REF_REG
<< end >>
