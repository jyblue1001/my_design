magic
tech sky130A
timestamp 1753589008
<< nwell >>
rect 56025 4340 56365 4730
rect 56495 4340 56835 4560
rect 56965 4340 57305 4730
rect 57435 4340 57775 4730
rect 54865 3670 55745 4060
rect 55945 3670 56825 4060
rect 56975 3670 57855 4060
rect 58055 3670 58940 4060
rect 57400 3665 57530 3670
rect 54895 2645 55715 3285
rect 56215 3185 57585 3275
rect 55970 2875 56790 2965
rect 57010 2875 57830 2965
rect 58090 2645 58910 3285
rect 54895 2150 55715 2390
rect 58090 2150 58910 2390
<< nmos >>
rect 56590 2535 56605 2585
rect 56645 2535 56660 2585
rect 56700 2535 56715 2585
rect 56755 2535 56770 2585
rect 56810 2535 56825 2585
rect 56865 2535 56880 2585
rect 56920 2535 56935 2585
rect 56975 2535 56990 2585
rect 57030 2535 57045 2585
rect 57085 2535 57100 2585
rect 57140 2535 57155 2585
rect 57195 2535 57210 2585
rect 56070 2030 56085 2180
rect 56125 2030 56140 2180
rect 56180 2030 56195 2180
rect 56235 2030 56250 2180
rect 56290 2030 56305 2180
rect 56345 2030 56360 2180
rect 56400 2030 56415 2180
rect 56455 2030 56470 2180
rect 56510 2030 56525 2180
rect 56565 2030 56580 2180
rect 56620 2030 56635 2180
rect 56675 2030 56690 2180
rect 57110 2030 57125 2180
rect 57165 2030 57180 2180
rect 57220 2030 57235 2180
rect 57275 2030 57290 2180
rect 57330 2030 57345 2180
rect 57385 2030 57400 2180
rect 57440 2030 57455 2180
rect 57495 2030 57510 2180
rect 57550 2030 57565 2180
rect 57605 2030 57620 2180
rect 57660 2030 57675 2180
rect 57715 2030 57730 2180
rect 54995 1610 55010 1910
rect 55050 1610 55065 1910
rect 55105 1610 55120 1910
rect 55160 1610 55175 1910
rect 55215 1610 55230 1910
rect 55270 1610 55285 1910
rect 55325 1610 55340 1910
rect 55380 1610 55395 1910
rect 55435 1610 55450 1910
rect 55490 1610 55505 1910
rect 55545 1610 55560 1910
rect 55600 1610 55615 1910
rect 56070 1560 56085 1710
rect 56125 1560 56140 1710
rect 56180 1560 56195 1710
rect 56235 1560 56250 1710
rect 56290 1560 56305 1710
rect 56345 1560 56360 1710
rect 56400 1560 56415 1710
rect 56455 1560 56470 1710
rect 56510 1560 56525 1710
rect 56565 1560 56580 1710
rect 56620 1560 56635 1710
rect 56675 1560 56690 1710
rect 56810 1560 56825 1710
rect 56865 1560 56880 1710
rect 56920 1560 56935 1710
rect 56975 1560 56990 1710
rect 57110 1560 57125 1710
rect 57165 1560 57180 1710
rect 57220 1560 57235 1710
rect 57275 1560 57290 1710
rect 57330 1560 57345 1710
rect 57385 1560 57400 1710
rect 57440 1560 57455 1710
rect 57495 1560 57510 1710
rect 57550 1560 57565 1710
rect 57605 1560 57620 1710
rect 57660 1560 57675 1710
rect 57715 1560 57730 1710
rect 58190 1610 58205 1910
rect 58245 1610 58260 1910
rect 58300 1610 58315 1910
rect 58355 1610 58370 1910
rect 58410 1610 58425 1910
rect 58465 1610 58480 1910
rect 58520 1610 58535 1910
rect 58575 1610 58590 1910
rect 58630 1610 58645 1910
rect 58685 1610 58700 1910
rect 58740 1610 58755 1910
rect 58795 1610 58810 1910
rect 55025 520 55085 1220
rect 55125 520 55185 1220
rect 55225 520 55285 1220
rect 55325 520 55385 1220
rect 55425 520 55485 1220
rect 55525 520 55585 1220
rect 56260 910 56275 1160
rect 56315 910 56330 1160
rect 56370 910 56385 1160
rect 56425 910 56440 1160
rect 56480 910 56495 1160
rect 56535 910 56550 1160
rect 56590 910 56605 1160
rect 56645 910 56660 1160
rect 56700 910 56715 1160
rect 56755 910 56770 1160
rect 56810 910 56825 1160
rect 56865 910 56880 1160
rect 56920 910 56935 1160
rect 56975 910 56990 1160
rect 57030 910 57045 1160
rect 57085 910 57100 1160
rect 57140 910 57155 1160
rect 57195 910 57210 1160
rect 57250 910 57265 1160
rect 57305 910 57320 1160
rect 57360 910 57375 1160
rect 57415 910 57430 1160
rect 57470 910 57485 1160
rect 56470 545 56485 695
rect 56525 545 56540 695
rect 56580 545 56595 695
rect 56635 545 56650 695
rect 56690 545 56705 695
rect 56745 545 56760 695
rect 56910 545 57210 695
rect 58220 520 58280 1220
rect 58320 520 58380 1220
rect 58420 520 58480 1220
rect 58520 520 58580 1220
rect 58620 520 58680 1220
rect 58720 520 58780 1220
<< pmos >>
rect 56125 4360 56145 4710
rect 56185 4360 56205 4710
rect 56245 4360 56265 4710
rect 56595 4360 56615 4540
rect 56655 4360 56675 4540
rect 56715 4360 56735 4540
rect 57065 4360 57085 4710
rect 57125 4360 57145 4710
rect 57185 4360 57205 4710
rect 57535 4360 57555 4710
rect 57595 4360 57615 4710
rect 57655 4360 57675 4710
rect 54965 3690 54985 4040
rect 55025 3690 55045 4040
rect 55085 3690 55105 4040
rect 55145 3690 55165 4040
rect 55205 3690 55225 4040
rect 55265 3690 55285 4040
rect 55325 3690 55345 4040
rect 55385 3690 55405 4040
rect 55445 3690 55465 4040
rect 55505 3690 55525 4040
rect 55565 3690 55585 4040
rect 55625 3690 55645 4040
rect 56045 3690 56065 4040
rect 56105 3690 56125 4040
rect 56165 3690 56185 4040
rect 56225 3690 56245 4040
rect 56285 3690 56305 4040
rect 56345 3690 56365 4040
rect 56405 3690 56425 4040
rect 56465 3690 56485 4040
rect 56525 3690 56545 4040
rect 56585 3690 56605 4040
rect 56645 3690 56665 4040
rect 56705 3690 56725 4040
rect 57075 3690 57095 4040
rect 57135 3690 57155 4040
rect 57195 3690 57215 4040
rect 57255 3690 57275 4040
rect 57315 3690 57335 4040
rect 57375 3690 57395 4040
rect 57435 3690 57455 4040
rect 57495 3690 57515 4040
rect 57555 3690 57575 4040
rect 57615 3690 57635 4040
rect 57675 3690 57695 4040
rect 57735 3690 57755 4040
rect 58160 3690 58180 4040
rect 58220 3690 58240 4040
rect 58280 3690 58300 4040
rect 58340 3690 58360 4040
rect 58400 3690 58420 4040
rect 58460 3690 58480 4040
rect 58520 3690 58540 4040
rect 58580 3690 58600 4040
rect 58640 3690 58660 4040
rect 58700 3690 58720 4040
rect 58760 3690 58780 4040
rect 58820 3690 58840 4040
rect 54995 2665 55010 3265
rect 55050 2665 55065 3265
rect 55105 2665 55120 3265
rect 55160 2665 55175 3265
rect 55215 2665 55230 3265
rect 55270 2665 55285 3265
rect 55325 2665 55340 3265
rect 55380 2665 55395 3265
rect 55435 2665 55450 3265
rect 55490 2665 55505 3265
rect 55545 2665 55560 3265
rect 55600 2665 55615 3265
rect 56315 3205 56330 3255
rect 56370 3205 56385 3255
rect 56425 3205 56440 3255
rect 56480 3205 56495 3255
rect 56535 3205 56550 3255
rect 56590 3205 56605 3255
rect 56645 3205 56660 3255
rect 56700 3205 56715 3255
rect 56755 3205 56770 3255
rect 56810 3205 56825 3255
rect 56865 3205 56880 3255
rect 56920 3205 56935 3255
rect 56975 3205 56990 3255
rect 57030 3205 57045 3255
rect 57085 3205 57100 3255
rect 57140 3205 57155 3255
rect 57195 3205 57210 3255
rect 57250 3205 57265 3255
rect 57305 3205 57320 3255
rect 57360 3205 57375 3255
rect 57415 3205 57430 3255
rect 57470 3205 57485 3255
rect 56070 2895 56085 2945
rect 56125 2895 56140 2945
rect 56180 2895 56195 2945
rect 56235 2895 56250 2945
rect 56290 2895 56305 2945
rect 56345 2895 56360 2945
rect 56400 2895 56415 2945
rect 56455 2895 56470 2945
rect 56510 2895 56525 2945
rect 56565 2895 56580 2945
rect 56620 2895 56635 2945
rect 56675 2895 56690 2945
rect 57110 2895 57125 2945
rect 57165 2895 57180 2945
rect 57220 2895 57235 2945
rect 57275 2895 57290 2945
rect 57330 2895 57345 2945
rect 57385 2895 57400 2945
rect 57440 2895 57455 2945
rect 57495 2895 57510 2945
rect 57550 2895 57565 2945
rect 57605 2895 57620 2945
rect 57660 2895 57675 2945
rect 57715 2895 57730 2945
rect 58190 2665 58205 3265
rect 58245 2665 58260 3265
rect 58300 2665 58315 3265
rect 58355 2665 58370 3265
rect 58410 2665 58425 3265
rect 58465 2665 58480 3265
rect 58520 2665 58535 3265
rect 58575 2665 58590 3265
rect 58630 2665 58645 3265
rect 58685 2665 58700 3265
rect 58740 2665 58755 3265
rect 58795 2665 58810 3265
rect 54995 2170 55010 2370
rect 55050 2170 55065 2370
rect 55105 2170 55120 2370
rect 55160 2170 55175 2370
rect 55215 2170 55230 2370
rect 55270 2170 55285 2370
rect 55325 2170 55340 2370
rect 55380 2170 55395 2370
rect 55435 2170 55450 2370
rect 55490 2170 55505 2370
rect 55545 2170 55560 2370
rect 55600 2170 55615 2370
rect 58190 2170 58205 2370
rect 58245 2170 58260 2370
rect 58300 2170 58315 2370
rect 58355 2170 58370 2370
rect 58410 2170 58425 2370
rect 58465 2170 58480 2370
rect 58520 2170 58535 2370
rect 58575 2170 58590 2370
rect 58630 2170 58645 2370
rect 58685 2170 58700 2370
rect 58740 2170 58755 2370
rect 58795 2170 58810 2370
<< ndiff >>
rect 56550 2570 56590 2585
rect 56550 2550 56560 2570
rect 56580 2550 56590 2570
rect 56550 2535 56590 2550
rect 56605 2570 56645 2585
rect 56605 2550 56615 2570
rect 56635 2550 56645 2570
rect 56605 2535 56645 2550
rect 56660 2570 56700 2585
rect 56660 2550 56670 2570
rect 56690 2550 56700 2570
rect 56660 2535 56700 2550
rect 56715 2570 56755 2585
rect 56715 2550 56725 2570
rect 56745 2550 56755 2570
rect 56715 2535 56755 2550
rect 56770 2570 56810 2585
rect 56770 2550 56780 2570
rect 56800 2550 56810 2570
rect 56770 2535 56810 2550
rect 56825 2570 56865 2585
rect 56825 2550 56835 2570
rect 56855 2550 56865 2570
rect 56825 2535 56865 2550
rect 56880 2570 56920 2585
rect 56880 2550 56890 2570
rect 56910 2550 56920 2570
rect 56880 2535 56920 2550
rect 56935 2570 56975 2585
rect 56935 2550 56945 2570
rect 56965 2550 56975 2570
rect 56935 2535 56975 2550
rect 56990 2570 57030 2585
rect 56990 2550 57000 2570
rect 57020 2550 57030 2570
rect 56990 2535 57030 2550
rect 57045 2570 57085 2585
rect 57045 2550 57055 2570
rect 57075 2550 57085 2570
rect 57045 2535 57085 2550
rect 57100 2570 57140 2585
rect 57100 2550 57110 2570
rect 57130 2550 57140 2570
rect 57100 2535 57140 2550
rect 57155 2570 57195 2585
rect 57155 2550 57165 2570
rect 57185 2550 57195 2570
rect 57155 2535 57195 2550
rect 57210 2570 57250 2585
rect 57210 2550 57220 2570
rect 57240 2550 57250 2570
rect 57210 2535 57250 2550
rect 56030 2165 56070 2180
rect 56030 2045 56040 2165
rect 56060 2045 56070 2165
rect 56030 2030 56070 2045
rect 56085 2165 56125 2180
rect 56085 2045 56095 2165
rect 56115 2045 56125 2165
rect 56085 2030 56125 2045
rect 56140 2165 56180 2180
rect 56140 2045 56150 2165
rect 56170 2045 56180 2165
rect 56140 2030 56180 2045
rect 56195 2165 56235 2180
rect 56195 2045 56205 2165
rect 56225 2045 56235 2165
rect 56195 2030 56235 2045
rect 56250 2165 56290 2180
rect 56250 2045 56260 2165
rect 56280 2045 56290 2165
rect 56250 2030 56290 2045
rect 56305 2165 56345 2180
rect 56305 2045 56315 2165
rect 56335 2045 56345 2165
rect 56305 2030 56345 2045
rect 56360 2165 56400 2180
rect 56360 2045 56370 2165
rect 56390 2045 56400 2165
rect 56360 2030 56400 2045
rect 56415 2165 56455 2180
rect 56415 2045 56425 2165
rect 56445 2045 56455 2165
rect 56415 2030 56455 2045
rect 56470 2165 56510 2180
rect 56470 2045 56480 2165
rect 56500 2045 56510 2165
rect 56470 2030 56510 2045
rect 56525 2165 56565 2180
rect 56525 2045 56535 2165
rect 56555 2045 56565 2165
rect 56525 2030 56565 2045
rect 56580 2165 56620 2180
rect 56580 2045 56590 2165
rect 56610 2045 56620 2165
rect 56580 2030 56620 2045
rect 56635 2165 56675 2180
rect 56635 2045 56645 2165
rect 56665 2045 56675 2165
rect 56635 2030 56675 2045
rect 56690 2165 56730 2180
rect 56690 2045 56700 2165
rect 56720 2045 56730 2165
rect 56690 2030 56730 2045
rect 57070 2165 57110 2180
rect 57070 2045 57080 2165
rect 57100 2045 57110 2165
rect 57070 2030 57110 2045
rect 57125 2165 57165 2180
rect 57125 2045 57135 2165
rect 57155 2045 57165 2165
rect 57125 2030 57165 2045
rect 57180 2165 57220 2180
rect 57180 2045 57190 2165
rect 57210 2045 57220 2165
rect 57180 2030 57220 2045
rect 57235 2165 57275 2180
rect 57235 2045 57245 2165
rect 57265 2045 57275 2165
rect 57235 2030 57275 2045
rect 57290 2165 57330 2180
rect 57290 2045 57300 2165
rect 57320 2045 57330 2165
rect 57290 2030 57330 2045
rect 57345 2165 57385 2180
rect 57345 2045 57355 2165
rect 57375 2045 57385 2165
rect 57345 2030 57385 2045
rect 57400 2165 57440 2180
rect 57400 2045 57410 2165
rect 57430 2045 57440 2165
rect 57400 2030 57440 2045
rect 57455 2165 57495 2180
rect 57455 2045 57465 2165
rect 57485 2045 57495 2165
rect 57455 2030 57495 2045
rect 57510 2165 57550 2180
rect 57510 2045 57520 2165
rect 57540 2045 57550 2165
rect 57510 2030 57550 2045
rect 57565 2165 57605 2180
rect 57565 2045 57575 2165
rect 57595 2045 57605 2165
rect 57565 2030 57605 2045
rect 57620 2165 57660 2180
rect 57620 2045 57630 2165
rect 57650 2045 57660 2165
rect 57620 2030 57660 2045
rect 57675 2165 57715 2180
rect 57675 2045 57685 2165
rect 57705 2045 57715 2165
rect 57675 2030 57715 2045
rect 57730 2165 57770 2180
rect 57730 2045 57740 2165
rect 57760 2045 57770 2165
rect 57730 2030 57770 2045
rect 54955 1895 54995 1910
rect 54955 1625 54965 1895
rect 54985 1625 54995 1895
rect 54955 1610 54995 1625
rect 55010 1895 55050 1910
rect 55010 1625 55020 1895
rect 55040 1625 55050 1895
rect 55010 1610 55050 1625
rect 55065 1895 55105 1910
rect 55065 1625 55075 1895
rect 55095 1625 55105 1895
rect 55065 1610 55105 1625
rect 55120 1895 55160 1910
rect 55120 1625 55130 1895
rect 55150 1625 55160 1895
rect 55120 1610 55160 1625
rect 55175 1895 55215 1910
rect 55175 1625 55185 1895
rect 55205 1625 55215 1895
rect 55175 1610 55215 1625
rect 55230 1895 55270 1910
rect 55230 1625 55240 1895
rect 55260 1625 55270 1895
rect 55230 1610 55270 1625
rect 55285 1895 55325 1910
rect 55285 1625 55295 1895
rect 55315 1625 55325 1895
rect 55285 1610 55325 1625
rect 55340 1895 55380 1910
rect 55340 1625 55350 1895
rect 55370 1625 55380 1895
rect 55340 1610 55380 1625
rect 55395 1895 55435 1910
rect 55395 1625 55405 1895
rect 55425 1625 55435 1895
rect 55395 1610 55435 1625
rect 55450 1895 55490 1910
rect 55450 1625 55460 1895
rect 55480 1625 55490 1895
rect 55450 1610 55490 1625
rect 55505 1895 55545 1910
rect 55505 1625 55515 1895
rect 55535 1625 55545 1895
rect 55505 1610 55545 1625
rect 55560 1895 55600 1910
rect 55560 1625 55570 1895
rect 55590 1625 55600 1895
rect 55560 1610 55600 1625
rect 55615 1895 55655 1910
rect 55615 1625 55625 1895
rect 55645 1625 55655 1895
rect 58150 1895 58190 1910
rect 55615 1610 55655 1625
rect 56030 1695 56070 1710
rect 56030 1575 56040 1695
rect 56060 1575 56070 1695
rect 56030 1560 56070 1575
rect 56085 1695 56125 1710
rect 56085 1575 56095 1695
rect 56115 1575 56125 1695
rect 56085 1560 56125 1575
rect 56140 1695 56180 1710
rect 56140 1575 56150 1695
rect 56170 1575 56180 1695
rect 56140 1560 56180 1575
rect 56195 1695 56235 1710
rect 56195 1575 56205 1695
rect 56225 1575 56235 1695
rect 56195 1560 56235 1575
rect 56250 1695 56290 1710
rect 56250 1575 56260 1695
rect 56280 1575 56290 1695
rect 56250 1560 56290 1575
rect 56305 1695 56345 1710
rect 56305 1575 56315 1695
rect 56335 1575 56345 1695
rect 56305 1560 56345 1575
rect 56360 1695 56400 1710
rect 56360 1575 56370 1695
rect 56390 1575 56400 1695
rect 56360 1560 56400 1575
rect 56415 1695 56455 1710
rect 56415 1575 56425 1695
rect 56445 1575 56455 1695
rect 56415 1560 56455 1575
rect 56470 1695 56510 1710
rect 56470 1575 56480 1695
rect 56500 1575 56510 1695
rect 56470 1560 56510 1575
rect 56525 1695 56565 1710
rect 56525 1575 56535 1695
rect 56555 1575 56565 1695
rect 56525 1560 56565 1575
rect 56580 1695 56620 1710
rect 56580 1575 56590 1695
rect 56610 1575 56620 1695
rect 56580 1560 56620 1575
rect 56635 1695 56675 1710
rect 56635 1575 56645 1695
rect 56665 1575 56675 1695
rect 56635 1560 56675 1575
rect 56690 1695 56730 1710
rect 56770 1695 56810 1710
rect 56690 1575 56700 1695
rect 56720 1575 56730 1695
rect 56770 1575 56780 1695
rect 56800 1575 56810 1695
rect 56690 1560 56730 1575
rect 56770 1560 56810 1575
rect 56825 1695 56865 1710
rect 56825 1575 56835 1695
rect 56855 1575 56865 1695
rect 56825 1560 56865 1575
rect 56880 1695 56920 1710
rect 56880 1575 56890 1695
rect 56910 1575 56920 1695
rect 56880 1560 56920 1575
rect 56935 1695 56975 1710
rect 56935 1575 56945 1695
rect 56965 1575 56975 1695
rect 56935 1560 56975 1575
rect 56990 1695 57030 1710
rect 57070 1695 57110 1710
rect 56990 1575 57000 1695
rect 57020 1575 57030 1695
rect 57070 1575 57080 1695
rect 57100 1575 57110 1695
rect 56990 1560 57030 1575
rect 57070 1560 57110 1575
rect 57125 1695 57165 1710
rect 57125 1575 57135 1695
rect 57155 1575 57165 1695
rect 57125 1560 57165 1575
rect 57180 1695 57220 1710
rect 57180 1575 57190 1695
rect 57210 1575 57220 1695
rect 57180 1560 57220 1575
rect 57235 1695 57275 1710
rect 57235 1575 57245 1695
rect 57265 1575 57275 1695
rect 57235 1560 57275 1575
rect 57290 1695 57330 1710
rect 57290 1575 57300 1695
rect 57320 1575 57330 1695
rect 57290 1560 57330 1575
rect 57345 1695 57385 1710
rect 57345 1575 57355 1695
rect 57375 1575 57385 1695
rect 57345 1560 57385 1575
rect 57400 1695 57440 1710
rect 57400 1575 57410 1695
rect 57430 1575 57440 1695
rect 57400 1560 57440 1575
rect 57455 1695 57495 1710
rect 57455 1575 57465 1695
rect 57485 1575 57495 1695
rect 57455 1560 57495 1575
rect 57510 1695 57550 1710
rect 57510 1575 57520 1695
rect 57540 1575 57550 1695
rect 57510 1560 57550 1575
rect 57565 1695 57605 1710
rect 57565 1575 57575 1695
rect 57595 1575 57605 1695
rect 57565 1560 57605 1575
rect 57620 1695 57660 1710
rect 57620 1575 57630 1695
rect 57650 1575 57660 1695
rect 57620 1560 57660 1575
rect 57675 1695 57715 1710
rect 57675 1575 57685 1695
rect 57705 1575 57715 1695
rect 57675 1560 57715 1575
rect 57730 1695 57770 1710
rect 57730 1575 57740 1695
rect 57760 1575 57770 1695
rect 58150 1625 58160 1895
rect 58180 1625 58190 1895
rect 58150 1610 58190 1625
rect 58205 1895 58245 1910
rect 58205 1625 58215 1895
rect 58235 1625 58245 1895
rect 58205 1610 58245 1625
rect 58260 1895 58300 1910
rect 58260 1625 58270 1895
rect 58290 1625 58300 1895
rect 58260 1610 58300 1625
rect 58315 1895 58355 1910
rect 58315 1625 58325 1895
rect 58345 1625 58355 1895
rect 58315 1610 58355 1625
rect 58370 1895 58410 1910
rect 58370 1625 58380 1895
rect 58400 1625 58410 1895
rect 58370 1610 58410 1625
rect 58425 1895 58465 1910
rect 58425 1625 58435 1895
rect 58455 1625 58465 1895
rect 58425 1610 58465 1625
rect 58480 1895 58520 1910
rect 58480 1625 58490 1895
rect 58510 1625 58520 1895
rect 58480 1610 58520 1625
rect 58535 1895 58575 1910
rect 58535 1625 58545 1895
rect 58565 1625 58575 1895
rect 58535 1610 58575 1625
rect 58590 1895 58630 1910
rect 58590 1625 58600 1895
rect 58620 1625 58630 1895
rect 58590 1610 58630 1625
rect 58645 1895 58685 1910
rect 58645 1625 58655 1895
rect 58675 1625 58685 1895
rect 58645 1610 58685 1625
rect 58700 1895 58740 1910
rect 58700 1625 58710 1895
rect 58730 1625 58740 1895
rect 58700 1610 58740 1625
rect 58755 1895 58795 1910
rect 58755 1625 58765 1895
rect 58785 1625 58795 1895
rect 58755 1610 58795 1625
rect 58810 1895 58850 1910
rect 58810 1625 58820 1895
rect 58840 1625 58850 1895
rect 58810 1610 58850 1625
rect 57730 1560 57770 1575
rect 54985 1205 55025 1220
rect 54985 535 54995 1205
rect 55015 535 55025 1205
rect 54985 520 55025 535
rect 55085 1205 55125 1220
rect 55085 535 55095 1205
rect 55115 535 55125 1205
rect 55085 520 55125 535
rect 55185 1205 55225 1220
rect 55185 535 55195 1205
rect 55215 535 55225 1205
rect 55185 520 55225 535
rect 55285 1205 55325 1220
rect 55285 535 55295 1205
rect 55315 535 55325 1205
rect 55285 520 55325 535
rect 55385 1205 55425 1220
rect 55385 535 55395 1205
rect 55415 535 55425 1205
rect 55385 520 55425 535
rect 55485 1205 55525 1220
rect 55485 535 55495 1205
rect 55515 535 55525 1205
rect 55485 520 55525 535
rect 55585 1205 55625 1220
rect 55585 535 55595 1205
rect 55615 535 55625 1205
rect 58180 1205 58220 1220
rect 56220 1145 56260 1160
rect 56220 925 56230 1145
rect 56250 925 56260 1145
rect 56220 910 56260 925
rect 56275 1145 56315 1160
rect 56275 925 56285 1145
rect 56305 925 56315 1145
rect 56275 910 56315 925
rect 56330 1145 56370 1160
rect 56330 925 56340 1145
rect 56360 925 56370 1145
rect 56330 910 56370 925
rect 56385 1145 56425 1160
rect 56385 925 56395 1145
rect 56415 925 56425 1145
rect 56385 910 56425 925
rect 56440 1145 56480 1160
rect 56440 925 56450 1145
rect 56470 925 56480 1145
rect 56440 910 56480 925
rect 56495 1145 56535 1160
rect 56495 925 56505 1145
rect 56525 925 56535 1145
rect 56495 910 56535 925
rect 56550 1145 56590 1160
rect 56550 925 56560 1145
rect 56580 925 56590 1145
rect 56550 910 56590 925
rect 56605 1145 56645 1160
rect 56605 925 56615 1145
rect 56635 925 56645 1145
rect 56605 910 56645 925
rect 56660 1145 56700 1160
rect 56660 925 56670 1145
rect 56690 925 56700 1145
rect 56660 910 56700 925
rect 56715 1145 56755 1160
rect 56715 925 56725 1145
rect 56745 925 56755 1145
rect 56715 910 56755 925
rect 56770 1145 56810 1160
rect 56770 925 56780 1145
rect 56800 925 56810 1145
rect 56770 910 56810 925
rect 56825 1145 56865 1160
rect 56825 925 56835 1145
rect 56855 925 56865 1145
rect 56825 910 56865 925
rect 56880 1145 56920 1160
rect 56880 925 56890 1145
rect 56910 925 56920 1145
rect 56880 910 56920 925
rect 56935 1145 56975 1160
rect 56935 925 56945 1145
rect 56965 925 56975 1145
rect 56935 910 56975 925
rect 56990 1145 57030 1160
rect 56990 925 57000 1145
rect 57020 925 57030 1145
rect 56990 910 57030 925
rect 57045 1145 57085 1160
rect 57045 925 57055 1145
rect 57075 925 57085 1145
rect 57045 910 57085 925
rect 57100 1145 57140 1160
rect 57100 925 57110 1145
rect 57130 925 57140 1145
rect 57100 910 57140 925
rect 57155 1145 57195 1160
rect 57155 925 57165 1145
rect 57185 925 57195 1145
rect 57155 910 57195 925
rect 57210 1145 57250 1160
rect 57210 925 57220 1145
rect 57240 925 57250 1145
rect 57210 910 57250 925
rect 57265 1145 57305 1160
rect 57265 925 57275 1145
rect 57295 925 57305 1145
rect 57265 910 57305 925
rect 57320 1145 57360 1160
rect 57320 925 57330 1145
rect 57350 925 57360 1145
rect 57320 910 57360 925
rect 57375 1145 57415 1160
rect 57375 925 57385 1145
rect 57405 925 57415 1145
rect 57375 910 57415 925
rect 57430 1145 57470 1160
rect 57430 925 57440 1145
rect 57460 925 57470 1145
rect 57430 910 57470 925
rect 57485 1145 57525 1160
rect 57485 925 57495 1145
rect 57515 925 57525 1145
rect 57485 910 57525 925
rect 56430 680 56470 695
rect 56430 560 56440 680
rect 56460 560 56470 680
rect 56430 545 56470 560
rect 56485 680 56525 695
rect 56485 560 56495 680
rect 56515 560 56525 680
rect 56485 545 56525 560
rect 56540 680 56580 695
rect 56540 560 56550 680
rect 56570 560 56580 680
rect 56540 545 56580 560
rect 56595 680 56635 695
rect 56595 560 56605 680
rect 56625 560 56635 680
rect 56595 545 56635 560
rect 56650 680 56690 695
rect 56650 560 56660 680
rect 56680 560 56690 680
rect 56650 545 56690 560
rect 56705 680 56745 695
rect 56705 560 56715 680
rect 56735 560 56745 680
rect 56705 545 56745 560
rect 56760 680 56800 695
rect 56760 560 56770 680
rect 56790 560 56800 680
rect 56760 545 56800 560
rect 56870 680 56910 695
rect 56870 560 56880 680
rect 56900 560 56910 680
rect 56870 545 56910 560
rect 57210 680 57250 695
rect 57210 560 57220 680
rect 57240 560 57250 680
rect 57210 545 57250 560
rect 55585 520 55625 535
rect 58180 535 58190 1205
rect 58210 535 58220 1205
rect 58180 520 58220 535
rect 58280 1205 58320 1220
rect 58280 535 58290 1205
rect 58310 535 58320 1205
rect 58280 520 58320 535
rect 58380 1205 58420 1220
rect 58380 535 58390 1205
rect 58410 535 58420 1205
rect 58380 520 58420 535
rect 58480 1205 58520 1220
rect 58480 535 58490 1205
rect 58510 535 58520 1205
rect 58480 520 58520 535
rect 58580 1205 58620 1220
rect 58580 535 58590 1205
rect 58610 535 58620 1205
rect 58580 520 58620 535
rect 58680 1205 58720 1220
rect 58680 535 58690 1205
rect 58710 535 58720 1205
rect 58680 520 58720 535
rect 58780 1205 58820 1220
rect 58780 535 58790 1205
rect 58810 535 58820 1205
rect 58780 520 58820 535
<< pdiff >>
rect 56085 4695 56125 4710
rect 56085 4375 56095 4695
rect 56115 4375 56125 4695
rect 56085 4360 56125 4375
rect 56145 4695 56185 4710
rect 56145 4375 56155 4695
rect 56175 4375 56185 4695
rect 56145 4360 56185 4375
rect 56205 4695 56245 4710
rect 56205 4375 56215 4695
rect 56235 4375 56245 4695
rect 56205 4360 56245 4375
rect 56265 4695 56305 4710
rect 56265 4375 56275 4695
rect 56295 4375 56305 4695
rect 57025 4695 57065 4710
rect 56265 4360 56305 4375
rect 56555 4525 56595 4540
rect 56555 4375 56565 4525
rect 56585 4375 56595 4525
rect 56555 4360 56595 4375
rect 56615 4525 56655 4540
rect 56615 4375 56625 4525
rect 56645 4375 56655 4525
rect 56615 4360 56655 4375
rect 56675 4525 56715 4540
rect 56675 4375 56685 4525
rect 56705 4375 56715 4525
rect 56675 4360 56715 4375
rect 56735 4525 56775 4540
rect 56735 4375 56745 4525
rect 56765 4375 56775 4525
rect 56735 4360 56775 4375
rect 57025 4375 57035 4695
rect 57055 4375 57065 4695
rect 57025 4360 57065 4375
rect 57085 4695 57125 4710
rect 57085 4375 57095 4695
rect 57115 4375 57125 4695
rect 57085 4360 57125 4375
rect 57145 4695 57185 4710
rect 57145 4375 57155 4695
rect 57175 4375 57185 4695
rect 57145 4360 57185 4375
rect 57205 4695 57245 4710
rect 57205 4375 57215 4695
rect 57235 4375 57245 4695
rect 57205 4360 57245 4375
rect 57495 4695 57535 4710
rect 57495 4375 57505 4695
rect 57525 4375 57535 4695
rect 57495 4360 57535 4375
rect 57555 4695 57595 4710
rect 57555 4375 57565 4695
rect 57585 4375 57595 4695
rect 57555 4360 57595 4375
rect 57615 4695 57655 4710
rect 57615 4375 57625 4695
rect 57645 4375 57655 4695
rect 57615 4360 57655 4375
rect 57675 4695 57715 4710
rect 57675 4375 57685 4695
rect 57705 4375 57715 4695
rect 57675 4360 57715 4375
rect 54925 4025 54965 4040
rect 54925 3705 54935 4025
rect 54955 3705 54965 4025
rect 54925 3690 54965 3705
rect 54985 4025 55025 4040
rect 54985 3705 54995 4025
rect 55015 3705 55025 4025
rect 54985 3690 55025 3705
rect 55045 4025 55085 4040
rect 55045 3705 55055 4025
rect 55075 3705 55085 4025
rect 55045 3690 55085 3705
rect 55105 4025 55145 4040
rect 55105 3705 55115 4025
rect 55135 3705 55145 4025
rect 55105 3690 55145 3705
rect 55165 4025 55205 4040
rect 55165 3705 55175 4025
rect 55195 3705 55205 4025
rect 55165 3690 55205 3705
rect 55225 4025 55265 4040
rect 55225 3705 55235 4025
rect 55255 3705 55265 4025
rect 55225 3690 55265 3705
rect 55285 4025 55325 4040
rect 55285 3705 55295 4025
rect 55315 3705 55325 4025
rect 55285 3690 55325 3705
rect 55345 4025 55385 4040
rect 55345 3705 55355 4025
rect 55375 3705 55385 4025
rect 55345 3690 55385 3705
rect 55405 4025 55445 4040
rect 55405 3705 55415 4025
rect 55435 3705 55445 4025
rect 55405 3690 55445 3705
rect 55465 4025 55505 4040
rect 55465 3705 55475 4025
rect 55495 3705 55505 4025
rect 55465 3690 55505 3705
rect 55525 4025 55565 4040
rect 55525 3705 55535 4025
rect 55555 3705 55565 4025
rect 55525 3690 55565 3705
rect 55585 4025 55625 4040
rect 55585 3705 55595 4025
rect 55615 3705 55625 4025
rect 55585 3690 55625 3705
rect 55645 4025 55685 4040
rect 55645 3705 55655 4025
rect 55675 3705 55685 4025
rect 55645 3690 55685 3705
rect 56005 4025 56045 4040
rect 56005 3705 56015 4025
rect 56035 3705 56045 4025
rect 56005 3690 56045 3705
rect 56065 4025 56105 4040
rect 56065 3705 56075 4025
rect 56095 3705 56105 4025
rect 56065 3690 56105 3705
rect 56125 4025 56165 4040
rect 56125 3705 56135 4025
rect 56155 3705 56165 4025
rect 56125 3690 56165 3705
rect 56185 4025 56225 4040
rect 56185 3705 56195 4025
rect 56215 3705 56225 4025
rect 56185 3690 56225 3705
rect 56245 4025 56285 4040
rect 56245 3705 56255 4025
rect 56275 3705 56285 4025
rect 56245 3690 56285 3705
rect 56305 4025 56345 4040
rect 56305 3705 56315 4025
rect 56335 3705 56345 4025
rect 56305 3690 56345 3705
rect 56365 4025 56405 4040
rect 56365 3705 56375 4025
rect 56395 3705 56405 4025
rect 56365 3690 56405 3705
rect 56425 4025 56465 4040
rect 56425 3705 56435 4025
rect 56455 3705 56465 4025
rect 56425 3690 56465 3705
rect 56485 4025 56525 4040
rect 56485 3705 56495 4025
rect 56515 3705 56525 4025
rect 56485 3690 56525 3705
rect 56545 4025 56585 4040
rect 56545 3705 56555 4025
rect 56575 3705 56585 4025
rect 56545 3690 56585 3705
rect 56605 4025 56645 4040
rect 56605 3705 56615 4025
rect 56635 3705 56645 4025
rect 56605 3690 56645 3705
rect 56665 4025 56705 4040
rect 56665 3705 56675 4025
rect 56695 3705 56705 4025
rect 56665 3690 56705 3705
rect 56725 4025 56765 4040
rect 56725 3705 56735 4025
rect 56755 3705 56765 4025
rect 56725 3690 56765 3705
rect 57035 4025 57075 4040
rect 57035 3705 57045 4025
rect 57065 3705 57075 4025
rect 57035 3690 57075 3705
rect 57095 4025 57135 4040
rect 57095 3705 57105 4025
rect 57125 3705 57135 4025
rect 57095 3690 57135 3705
rect 57155 4025 57195 4040
rect 57155 3705 57165 4025
rect 57185 3705 57195 4025
rect 57155 3690 57195 3705
rect 57215 4025 57255 4040
rect 57215 3705 57225 4025
rect 57245 3705 57255 4025
rect 57215 3690 57255 3705
rect 57275 4025 57315 4040
rect 57275 3705 57285 4025
rect 57305 3705 57315 4025
rect 57275 3690 57315 3705
rect 57335 4025 57375 4040
rect 57335 3705 57345 4025
rect 57365 3705 57375 4025
rect 57335 3690 57375 3705
rect 57395 4025 57435 4040
rect 57395 3705 57405 4025
rect 57425 3705 57435 4025
rect 57395 3690 57435 3705
rect 57455 4025 57495 4040
rect 57455 3705 57465 4025
rect 57485 3705 57495 4025
rect 57455 3690 57495 3705
rect 57515 4025 57555 4040
rect 57515 3705 57525 4025
rect 57545 3705 57555 4025
rect 57515 3690 57555 3705
rect 57575 4025 57615 4040
rect 57575 3705 57585 4025
rect 57605 3705 57615 4025
rect 57575 3690 57615 3705
rect 57635 4025 57675 4040
rect 57635 3705 57645 4025
rect 57665 3705 57675 4025
rect 57635 3690 57675 3705
rect 57695 4025 57735 4040
rect 57695 3705 57705 4025
rect 57725 3705 57735 4025
rect 57695 3690 57735 3705
rect 57755 4025 57795 4040
rect 57755 3705 57765 4025
rect 57785 3705 57795 4025
rect 57755 3690 57795 3705
rect 58120 4025 58160 4040
rect 58120 3705 58130 4025
rect 58150 3705 58160 4025
rect 58120 3690 58160 3705
rect 58180 4025 58220 4040
rect 58180 3705 58190 4025
rect 58210 3705 58220 4025
rect 58180 3690 58220 3705
rect 58240 4025 58280 4040
rect 58240 3705 58250 4025
rect 58270 3705 58280 4025
rect 58240 3690 58280 3705
rect 58300 4025 58340 4040
rect 58300 3705 58310 4025
rect 58330 3705 58340 4025
rect 58300 3690 58340 3705
rect 58360 4025 58400 4040
rect 58360 3705 58370 4025
rect 58390 3705 58400 4025
rect 58360 3690 58400 3705
rect 58420 4025 58460 4040
rect 58420 3705 58430 4025
rect 58450 3705 58460 4025
rect 58420 3690 58460 3705
rect 58480 4025 58520 4040
rect 58480 3705 58490 4025
rect 58510 3705 58520 4025
rect 58480 3690 58520 3705
rect 58540 4025 58580 4040
rect 58540 3705 58550 4025
rect 58570 3705 58580 4025
rect 58540 3690 58580 3705
rect 58600 4025 58640 4040
rect 58600 3705 58610 4025
rect 58630 3705 58640 4025
rect 58600 3690 58640 3705
rect 58660 4025 58700 4040
rect 58660 3705 58670 4025
rect 58690 3705 58700 4025
rect 58660 3690 58700 3705
rect 58720 4025 58760 4040
rect 58720 3705 58730 4025
rect 58750 3705 58760 4025
rect 58720 3690 58760 3705
rect 58780 4025 58820 4040
rect 58780 3705 58790 4025
rect 58810 3705 58820 4025
rect 58780 3690 58820 3705
rect 58840 4025 58880 4040
rect 58840 3705 58850 4025
rect 58870 3705 58880 4025
rect 58840 3690 58880 3705
rect 54955 3250 54995 3265
rect 54955 2680 54965 3250
rect 54985 2680 54995 3250
rect 54955 2665 54995 2680
rect 55010 3250 55050 3265
rect 55010 2680 55020 3250
rect 55040 2680 55050 3250
rect 55010 2665 55050 2680
rect 55065 3250 55105 3265
rect 55065 2680 55075 3250
rect 55095 2680 55105 3250
rect 55065 2665 55105 2680
rect 55120 3250 55160 3265
rect 55120 2680 55130 3250
rect 55150 2680 55160 3250
rect 55120 2665 55160 2680
rect 55175 3250 55215 3265
rect 55175 2680 55185 3250
rect 55205 2680 55215 3250
rect 55175 2665 55215 2680
rect 55230 3250 55270 3265
rect 55230 2680 55240 3250
rect 55260 2680 55270 3250
rect 55230 2665 55270 2680
rect 55285 3250 55325 3265
rect 55285 2680 55295 3250
rect 55315 2680 55325 3250
rect 55285 2665 55325 2680
rect 55340 3250 55380 3265
rect 55340 2680 55350 3250
rect 55370 2680 55380 3250
rect 55340 2665 55380 2680
rect 55395 3250 55435 3265
rect 55395 2680 55405 3250
rect 55425 2680 55435 3250
rect 55395 2665 55435 2680
rect 55450 3250 55490 3265
rect 55450 2680 55460 3250
rect 55480 2680 55490 3250
rect 55450 2665 55490 2680
rect 55505 3250 55545 3265
rect 55505 2680 55515 3250
rect 55535 2680 55545 3250
rect 55505 2665 55545 2680
rect 55560 3250 55600 3265
rect 55560 2680 55570 3250
rect 55590 2680 55600 3250
rect 55560 2665 55600 2680
rect 55615 3250 55655 3265
rect 55615 2680 55625 3250
rect 55645 2680 55655 3250
rect 56275 3240 56315 3255
rect 56275 3220 56285 3240
rect 56305 3220 56315 3240
rect 56275 3205 56315 3220
rect 56330 3240 56370 3255
rect 56330 3220 56340 3240
rect 56360 3220 56370 3240
rect 56330 3205 56370 3220
rect 56385 3240 56425 3255
rect 56385 3220 56395 3240
rect 56415 3220 56425 3240
rect 56385 3205 56425 3220
rect 56440 3240 56480 3255
rect 56440 3220 56450 3240
rect 56470 3220 56480 3240
rect 56440 3205 56480 3220
rect 56495 3240 56535 3255
rect 56495 3220 56505 3240
rect 56525 3220 56535 3240
rect 56495 3205 56535 3220
rect 56550 3240 56590 3255
rect 56550 3220 56560 3240
rect 56580 3220 56590 3240
rect 56550 3205 56590 3220
rect 56605 3240 56645 3255
rect 56605 3220 56615 3240
rect 56635 3220 56645 3240
rect 56605 3205 56645 3220
rect 56660 3240 56700 3255
rect 56660 3220 56670 3240
rect 56690 3220 56700 3240
rect 56660 3205 56700 3220
rect 56715 3240 56755 3255
rect 56715 3220 56725 3240
rect 56745 3220 56755 3240
rect 56715 3205 56755 3220
rect 56770 3240 56810 3255
rect 56770 3220 56780 3240
rect 56800 3220 56810 3240
rect 56770 3205 56810 3220
rect 56825 3240 56865 3255
rect 56825 3220 56835 3240
rect 56855 3220 56865 3240
rect 56825 3205 56865 3220
rect 56880 3240 56920 3255
rect 56880 3220 56890 3240
rect 56910 3220 56920 3240
rect 56880 3205 56920 3220
rect 56935 3240 56975 3255
rect 56935 3220 56945 3240
rect 56965 3220 56975 3240
rect 56935 3205 56975 3220
rect 56990 3240 57030 3255
rect 56990 3220 57000 3240
rect 57020 3220 57030 3240
rect 56990 3205 57030 3220
rect 57045 3240 57085 3255
rect 57045 3220 57055 3240
rect 57075 3220 57085 3240
rect 57045 3205 57085 3220
rect 57100 3240 57140 3255
rect 57100 3220 57110 3240
rect 57130 3220 57140 3240
rect 57100 3205 57140 3220
rect 57155 3240 57195 3255
rect 57155 3220 57165 3240
rect 57185 3220 57195 3240
rect 57155 3205 57195 3220
rect 57210 3240 57250 3255
rect 57210 3220 57220 3240
rect 57240 3220 57250 3240
rect 57210 3205 57250 3220
rect 57265 3240 57305 3255
rect 57265 3220 57275 3240
rect 57295 3220 57305 3240
rect 57265 3205 57305 3220
rect 57320 3240 57360 3255
rect 57320 3220 57330 3240
rect 57350 3220 57360 3240
rect 57320 3205 57360 3220
rect 57375 3240 57415 3255
rect 57375 3220 57385 3240
rect 57405 3220 57415 3240
rect 57375 3205 57415 3220
rect 57430 3240 57470 3255
rect 57430 3220 57440 3240
rect 57460 3220 57470 3240
rect 57430 3205 57470 3220
rect 57485 3240 57525 3255
rect 57485 3220 57495 3240
rect 57515 3220 57525 3240
rect 57485 3205 57525 3220
rect 58150 3250 58190 3265
rect 56030 2930 56070 2945
rect 56030 2910 56040 2930
rect 56060 2910 56070 2930
rect 56030 2895 56070 2910
rect 56085 2930 56125 2945
rect 56085 2910 56095 2930
rect 56115 2910 56125 2930
rect 56085 2895 56125 2910
rect 56140 2930 56180 2945
rect 56140 2910 56150 2930
rect 56170 2910 56180 2930
rect 56140 2895 56180 2910
rect 56195 2930 56235 2945
rect 56195 2910 56205 2930
rect 56225 2910 56235 2930
rect 56195 2895 56235 2910
rect 56250 2930 56290 2945
rect 56250 2910 56260 2930
rect 56280 2910 56290 2930
rect 56250 2895 56290 2910
rect 56305 2930 56345 2945
rect 56305 2910 56315 2930
rect 56335 2910 56345 2930
rect 56305 2895 56345 2910
rect 56360 2930 56400 2945
rect 56360 2910 56370 2930
rect 56390 2910 56400 2930
rect 56360 2895 56400 2910
rect 56415 2930 56455 2945
rect 56415 2910 56425 2930
rect 56445 2910 56455 2930
rect 56415 2895 56455 2910
rect 56470 2930 56510 2945
rect 56470 2910 56480 2930
rect 56500 2910 56510 2930
rect 56470 2895 56510 2910
rect 56525 2930 56565 2945
rect 56525 2910 56535 2930
rect 56555 2910 56565 2930
rect 56525 2895 56565 2910
rect 56580 2930 56620 2945
rect 56580 2910 56590 2930
rect 56610 2910 56620 2930
rect 56580 2895 56620 2910
rect 56635 2930 56675 2945
rect 56635 2910 56645 2930
rect 56665 2910 56675 2930
rect 56635 2895 56675 2910
rect 56690 2930 56730 2945
rect 56690 2910 56700 2930
rect 56720 2910 56730 2930
rect 56690 2895 56730 2910
rect 57070 2930 57110 2945
rect 57070 2910 57080 2930
rect 57100 2910 57110 2930
rect 57070 2895 57110 2910
rect 57125 2930 57165 2945
rect 57125 2910 57135 2930
rect 57155 2910 57165 2930
rect 57125 2895 57165 2910
rect 57180 2930 57220 2945
rect 57180 2910 57190 2930
rect 57210 2910 57220 2930
rect 57180 2895 57220 2910
rect 57235 2930 57275 2945
rect 57235 2910 57245 2930
rect 57265 2910 57275 2930
rect 57235 2895 57275 2910
rect 57290 2930 57330 2945
rect 57290 2910 57300 2930
rect 57320 2910 57330 2930
rect 57290 2895 57330 2910
rect 57345 2930 57385 2945
rect 57345 2910 57355 2930
rect 57375 2910 57385 2930
rect 57345 2895 57385 2910
rect 57400 2930 57440 2945
rect 57400 2910 57410 2930
rect 57430 2910 57440 2930
rect 57400 2895 57440 2910
rect 57455 2930 57495 2945
rect 57455 2910 57465 2930
rect 57485 2910 57495 2930
rect 57455 2895 57495 2910
rect 57510 2930 57550 2945
rect 57510 2910 57520 2930
rect 57540 2910 57550 2930
rect 57510 2895 57550 2910
rect 57565 2930 57605 2945
rect 57565 2910 57575 2930
rect 57595 2910 57605 2930
rect 57565 2895 57605 2910
rect 57620 2930 57660 2945
rect 57620 2910 57630 2930
rect 57650 2910 57660 2930
rect 57620 2895 57660 2910
rect 57675 2930 57715 2945
rect 57675 2910 57685 2930
rect 57705 2910 57715 2930
rect 57675 2895 57715 2910
rect 57730 2930 57770 2945
rect 57730 2910 57740 2930
rect 57760 2910 57770 2930
rect 57730 2895 57770 2910
rect 55615 2665 55655 2680
rect 58150 2680 58160 3250
rect 58180 2680 58190 3250
rect 58150 2665 58190 2680
rect 58205 3250 58245 3265
rect 58205 2680 58215 3250
rect 58235 2680 58245 3250
rect 58205 2665 58245 2680
rect 58260 3250 58300 3265
rect 58260 2680 58270 3250
rect 58290 2680 58300 3250
rect 58260 2665 58300 2680
rect 58315 3250 58355 3265
rect 58315 2680 58325 3250
rect 58345 2680 58355 3250
rect 58315 2665 58355 2680
rect 58370 3250 58410 3265
rect 58370 2680 58380 3250
rect 58400 2680 58410 3250
rect 58370 2665 58410 2680
rect 58425 3250 58465 3265
rect 58425 2680 58435 3250
rect 58455 2680 58465 3250
rect 58425 2665 58465 2680
rect 58480 3250 58520 3265
rect 58480 2680 58490 3250
rect 58510 2680 58520 3250
rect 58480 2665 58520 2680
rect 58535 3250 58575 3265
rect 58535 2680 58545 3250
rect 58565 2680 58575 3250
rect 58535 2665 58575 2680
rect 58590 3250 58630 3265
rect 58590 2680 58600 3250
rect 58620 2680 58630 3250
rect 58590 2665 58630 2680
rect 58645 3250 58685 3265
rect 58645 2680 58655 3250
rect 58675 2680 58685 3250
rect 58645 2665 58685 2680
rect 58700 3250 58740 3265
rect 58700 2680 58710 3250
rect 58730 2680 58740 3250
rect 58700 2665 58740 2680
rect 58755 3250 58795 3265
rect 58755 2680 58765 3250
rect 58785 2680 58795 3250
rect 58755 2665 58795 2680
rect 58810 3250 58850 3265
rect 58810 2680 58820 3250
rect 58840 2680 58850 3250
rect 58810 2665 58850 2680
rect 54955 2355 54995 2370
rect 54955 2185 54965 2355
rect 54985 2185 54995 2355
rect 54955 2170 54995 2185
rect 55010 2355 55050 2370
rect 55010 2185 55020 2355
rect 55040 2185 55050 2355
rect 55010 2170 55050 2185
rect 55065 2355 55105 2370
rect 55065 2185 55075 2355
rect 55095 2185 55105 2355
rect 55065 2170 55105 2185
rect 55120 2355 55160 2370
rect 55120 2185 55130 2355
rect 55150 2185 55160 2355
rect 55120 2170 55160 2185
rect 55175 2355 55215 2370
rect 55175 2185 55185 2355
rect 55205 2185 55215 2355
rect 55175 2170 55215 2185
rect 55230 2355 55270 2370
rect 55230 2185 55240 2355
rect 55260 2185 55270 2355
rect 55230 2170 55270 2185
rect 55285 2355 55325 2370
rect 55285 2185 55295 2355
rect 55315 2185 55325 2355
rect 55285 2170 55325 2185
rect 55340 2355 55380 2370
rect 55340 2185 55350 2355
rect 55370 2185 55380 2355
rect 55340 2170 55380 2185
rect 55395 2355 55435 2370
rect 55395 2185 55405 2355
rect 55425 2185 55435 2355
rect 55395 2170 55435 2185
rect 55450 2355 55490 2370
rect 55450 2185 55460 2355
rect 55480 2185 55490 2355
rect 55450 2170 55490 2185
rect 55505 2355 55545 2370
rect 55505 2185 55515 2355
rect 55535 2185 55545 2355
rect 55505 2170 55545 2185
rect 55560 2355 55600 2370
rect 55560 2185 55570 2355
rect 55590 2185 55600 2355
rect 55560 2170 55600 2185
rect 55615 2355 55655 2370
rect 55615 2185 55625 2355
rect 55645 2185 55655 2355
rect 58150 2355 58190 2370
rect 55615 2170 55655 2185
rect 58150 2185 58160 2355
rect 58180 2185 58190 2355
rect 58150 2170 58190 2185
rect 58205 2355 58245 2370
rect 58205 2185 58215 2355
rect 58235 2185 58245 2355
rect 58205 2170 58245 2185
rect 58260 2355 58300 2370
rect 58260 2185 58270 2355
rect 58290 2185 58300 2355
rect 58260 2170 58300 2185
rect 58315 2355 58355 2370
rect 58315 2185 58325 2355
rect 58345 2185 58355 2355
rect 58315 2170 58355 2185
rect 58370 2355 58410 2370
rect 58370 2185 58380 2355
rect 58400 2185 58410 2355
rect 58370 2170 58410 2185
rect 58425 2355 58465 2370
rect 58425 2185 58435 2355
rect 58455 2185 58465 2355
rect 58425 2170 58465 2185
rect 58480 2355 58520 2370
rect 58480 2185 58490 2355
rect 58510 2185 58520 2355
rect 58480 2170 58520 2185
rect 58535 2355 58575 2370
rect 58535 2185 58545 2355
rect 58565 2185 58575 2355
rect 58535 2170 58575 2185
rect 58590 2355 58630 2370
rect 58590 2185 58600 2355
rect 58620 2185 58630 2355
rect 58590 2170 58630 2185
rect 58645 2355 58685 2370
rect 58645 2185 58655 2355
rect 58675 2185 58685 2355
rect 58645 2170 58685 2185
rect 58700 2355 58740 2370
rect 58700 2185 58710 2355
rect 58730 2185 58740 2355
rect 58700 2170 58740 2185
rect 58755 2355 58795 2370
rect 58755 2185 58765 2355
rect 58785 2185 58795 2355
rect 58755 2170 58795 2185
rect 58810 2355 58850 2370
rect 58810 2185 58820 2355
rect 58840 2185 58850 2355
rect 58810 2170 58850 2185
<< ndiffc >>
rect 56560 2550 56580 2570
rect 56615 2550 56635 2570
rect 56670 2550 56690 2570
rect 56725 2550 56745 2570
rect 56780 2550 56800 2570
rect 56835 2550 56855 2570
rect 56890 2550 56910 2570
rect 56945 2550 56965 2570
rect 57000 2550 57020 2570
rect 57055 2550 57075 2570
rect 57110 2550 57130 2570
rect 57165 2550 57185 2570
rect 57220 2550 57240 2570
rect 56040 2045 56060 2165
rect 56095 2045 56115 2165
rect 56150 2045 56170 2165
rect 56205 2045 56225 2165
rect 56260 2045 56280 2165
rect 56315 2045 56335 2165
rect 56370 2045 56390 2165
rect 56425 2045 56445 2165
rect 56480 2045 56500 2165
rect 56535 2045 56555 2165
rect 56590 2045 56610 2165
rect 56645 2045 56665 2165
rect 56700 2045 56720 2165
rect 57080 2045 57100 2165
rect 57135 2045 57155 2165
rect 57190 2045 57210 2165
rect 57245 2045 57265 2165
rect 57300 2045 57320 2165
rect 57355 2045 57375 2165
rect 57410 2045 57430 2165
rect 57465 2045 57485 2165
rect 57520 2045 57540 2165
rect 57575 2045 57595 2165
rect 57630 2045 57650 2165
rect 57685 2045 57705 2165
rect 57740 2045 57760 2165
rect 54965 1625 54985 1895
rect 55020 1625 55040 1895
rect 55075 1625 55095 1895
rect 55130 1625 55150 1895
rect 55185 1625 55205 1895
rect 55240 1625 55260 1895
rect 55295 1625 55315 1895
rect 55350 1625 55370 1895
rect 55405 1625 55425 1895
rect 55460 1625 55480 1895
rect 55515 1625 55535 1895
rect 55570 1625 55590 1895
rect 55625 1625 55645 1895
rect 56040 1575 56060 1695
rect 56095 1575 56115 1695
rect 56150 1575 56170 1695
rect 56205 1575 56225 1695
rect 56260 1575 56280 1695
rect 56315 1575 56335 1695
rect 56370 1575 56390 1695
rect 56425 1575 56445 1695
rect 56480 1575 56500 1695
rect 56535 1575 56555 1695
rect 56590 1575 56610 1695
rect 56645 1575 56665 1695
rect 56700 1575 56720 1695
rect 56780 1575 56800 1695
rect 56835 1575 56855 1695
rect 56890 1575 56910 1695
rect 56945 1575 56965 1695
rect 57000 1575 57020 1695
rect 57080 1575 57100 1695
rect 57135 1575 57155 1695
rect 57190 1575 57210 1695
rect 57245 1575 57265 1695
rect 57300 1575 57320 1695
rect 57355 1575 57375 1695
rect 57410 1575 57430 1695
rect 57465 1575 57485 1695
rect 57520 1575 57540 1695
rect 57575 1575 57595 1695
rect 57630 1575 57650 1695
rect 57685 1575 57705 1695
rect 57740 1575 57760 1695
rect 58160 1625 58180 1895
rect 58215 1625 58235 1895
rect 58270 1625 58290 1895
rect 58325 1625 58345 1895
rect 58380 1625 58400 1895
rect 58435 1625 58455 1895
rect 58490 1625 58510 1895
rect 58545 1625 58565 1895
rect 58600 1625 58620 1895
rect 58655 1625 58675 1895
rect 58710 1625 58730 1895
rect 58765 1625 58785 1895
rect 58820 1625 58840 1895
rect 54995 535 55015 1205
rect 55095 535 55115 1205
rect 55195 535 55215 1205
rect 55295 535 55315 1205
rect 55395 535 55415 1205
rect 55495 535 55515 1205
rect 55595 535 55615 1205
rect 56230 925 56250 1145
rect 56285 925 56305 1145
rect 56340 925 56360 1145
rect 56395 925 56415 1145
rect 56450 925 56470 1145
rect 56505 925 56525 1145
rect 56560 925 56580 1145
rect 56615 925 56635 1145
rect 56670 925 56690 1145
rect 56725 925 56745 1145
rect 56780 925 56800 1145
rect 56835 925 56855 1145
rect 56890 925 56910 1145
rect 56945 925 56965 1145
rect 57000 925 57020 1145
rect 57055 925 57075 1145
rect 57110 925 57130 1145
rect 57165 925 57185 1145
rect 57220 925 57240 1145
rect 57275 925 57295 1145
rect 57330 925 57350 1145
rect 57385 925 57405 1145
rect 57440 925 57460 1145
rect 57495 925 57515 1145
rect 56440 560 56460 680
rect 56495 560 56515 680
rect 56550 560 56570 680
rect 56605 560 56625 680
rect 56660 560 56680 680
rect 56715 560 56735 680
rect 56770 560 56790 680
rect 56880 560 56900 680
rect 57220 560 57240 680
rect 58190 535 58210 1205
rect 58290 535 58310 1205
rect 58390 535 58410 1205
rect 58490 535 58510 1205
rect 58590 535 58610 1205
rect 58690 535 58710 1205
rect 58790 535 58810 1205
<< pdiffc >>
rect 56095 4375 56115 4695
rect 56155 4375 56175 4695
rect 56215 4375 56235 4695
rect 56275 4375 56295 4695
rect 56565 4375 56585 4525
rect 56625 4375 56645 4525
rect 56685 4375 56705 4525
rect 56745 4375 56765 4525
rect 57035 4375 57055 4695
rect 57095 4375 57115 4695
rect 57155 4375 57175 4695
rect 57215 4375 57235 4695
rect 57505 4375 57525 4695
rect 57565 4375 57585 4695
rect 57625 4375 57645 4695
rect 57685 4375 57705 4695
rect 54935 3705 54955 4025
rect 54995 3705 55015 4025
rect 55055 3705 55075 4025
rect 55115 3705 55135 4025
rect 55175 3705 55195 4025
rect 55235 3705 55255 4025
rect 55295 3705 55315 4025
rect 55355 3705 55375 4025
rect 55415 3705 55435 4025
rect 55475 3705 55495 4025
rect 55535 3705 55555 4025
rect 55595 3705 55615 4025
rect 55655 3705 55675 4025
rect 56015 3705 56035 4025
rect 56075 3705 56095 4025
rect 56135 3705 56155 4025
rect 56195 3705 56215 4025
rect 56255 3705 56275 4025
rect 56315 3705 56335 4025
rect 56375 3705 56395 4025
rect 56435 3705 56455 4025
rect 56495 3705 56515 4025
rect 56555 3705 56575 4025
rect 56615 3705 56635 4025
rect 56675 3705 56695 4025
rect 56735 3705 56755 4025
rect 57045 3705 57065 4025
rect 57105 3705 57125 4025
rect 57165 3705 57185 4025
rect 57225 3705 57245 4025
rect 57285 3705 57305 4025
rect 57345 3705 57365 4025
rect 57405 3705 57425 4025
rect 57465 3705 57485 4025
rect 57525 3705 57545 4025
rect 57585 3705 57605 4025
rect 57645 3705 57665 4025
rect 57705 3705 57725 4025
rect 57765 3705 57785 4025
rect 58130 3705 58150 4025
rect 58190 3705 58210 4025
rect 58250 3705 58270 4025
rect 58310 3705 58330 4025
rect 58370 3705 58390 4025
rect 58430 3705 58450 4025
rect 58490 3705 58510 4025
rect 58550 3705 58570 4025
rect 58610 3705 58630 4025
rect 58670 3705 58690 4025
rect 58730 3705 58750 4025
rect 58790 3705 58810 4025
rect 58850 3705 58870 4025
rect 54965 2680 54985 3250
rect 55020 2680 55040 3250
rect 55075 2680 55095 3250
rect 55130 2680 55150 3250
rect 55185 2680 55205 3250
rect 55240 2680 55260 3250
rect 55295 2680 55315 3250
rect 55350 2680 55370 3250
rect 55405 2680 55425 3250
rect 55460 2680 55480 3250
rect 55515 2680 55535 3250
rect 55570 2680 55590 3250
rect 55625 2680 55645 3250
rect 56285 3220 56305 3240
rect 56340 3220 56360 3240
rect 56395 3220 56415 3240
rect 56450 3220 56470 3240
rect 56505 3220 56525 3240
rect 56560 3220 56580 3240
rect 56615 3220 56635 3240
rect 56670 3220 56690 3240
rect 56725 3220 56745 3240
rect 56780 3220 56800 3240
rect 56835 3220 56855 3240
rect 56890 3220 56910 3240
rect 56945 3220 56965 3240
rect 57000 3220 57020 3240
rect 57055 3220 57075 3240
rect 57110 3220 57130 3240
rect 57165 3220 57185 3240
rect 57220 3220 57240 3240
rect 57275 3220 57295 3240
rect 57330 3220 57350 3240
rect 57385 3220 57405 3240
rect 57440 3220 57460 3240
rect 57495 3220 57515 3240
rect 56040 2910 56060 2930
rect 56095 2910 56115 2930
rect 56150 2910 56170 2930
rect 56205 2910 56225 2930
rect 56260 2910 56280 2930
rect 56315 2910 56335 2930
rect 56370 2910 56390 2930
rect 56425 2910 56445 2930
rect 56480 2910 56500 2930
rect 56535 2910 56555 2930
rect 56590 2910 56610 2930
rect 56645 2910 56665 2930
rect 56700 2910 56720 2930
rect 57080 2910 57100 2930
rect 57135 2910 57155 2930
rect 57190 2910 57210 2930
rect 57245 2910 57265 2930
rect 57300 2910 57320 2930
rect 57355 2910 57375 2930
rect 57410 2910 57430 2930
rect 57465 2910 57485 2930
rect 57520 2910 57540 2930
rect 57575 2910 57595 2930
rect 57630 2910 57650 2930
rect 57685 2910 57705 2930
rect 57740 2910 57760 2930
rect 58160 2680 58180 3250
rect 58215 2680 58235 3250
rect 58270 2680 58290 3250
rect 58325 2680 58345 3250
rect 58380 2680 58400 3250
rect 58435 2680 58455 3250
rect 58490 2680 58510 3250
rect 58545 2680 58565 3250
rect 58600 2680 58620 3250
rect 58655 2680 58675 3250
rect 58710 2680 58730 3250
rect 58765 2680 58785 3250
rect 58820 2680 58840 3250
rect 54965 2185 54985 2355
rect 55020 2185 55040 2355
rect 55075 2185 55095 2355
rect 55130 2185 55150 2355
rect 55185 2185 55205 2355
rect 55240 2185 55260 2355
rect 55295 2185 55315 2355
rect 55350 2185 55370 2355
rect 55405 2185 55425 2355
rect 55460 2185 55480 2355
rect 55515 2185 55535 2355
rect 55570 2185 55590 2355
rect 55625 2185 55645 2355
rect 58160 2185 58180 2355
rect 58215 2185 58235 2355
rect 58270 2185 58290 2355
rect 58325 2185 58345 2355
rect 58380 2185 58400 2355
rect 58435 2185 58455 2355
rect 58490 2185 58510 2355
rect 58545 2185 58565 2355
rect 58600 2185 58620 2355
rect 58655 2185 58675 2355
rect 58710 2185 58730 2355
rect 58765 2185 58785 2355
rect 58820 2185 58840 2355
<< psubdiff >>
rect 56510 2570 56550 2585
rect 56510 2550 56520 2570
rect 56540 2550 56550 2570
rect 56510 2535 56550 2550
rect 57250 2570 57290 2585
rect 57250 2550 57260 2570
rect 57280 2550 57290 2570
rect 57250 2535 57290 2550
rect 55990 2165 56030 2180
rect 55990 2045 56000 2165
rect 56020 2045 56030 2165
rect 55990 2030 56030 2045
rect 56730 2165 56770 2180
rect 56730 2045 56740 2165
rect 56760 2045 56770 2165
rect 56730 2030 56770 2045
rect 57030 2165 57070 2180
rect 57030 2045 57040 2165
rect 57060 2045 57070 2165
rect 57030 2030 57070 2045
rect 57770 2165 57810 2180
rect 57770 2045 57780 2165
rect 57800 2045 57810 2165
rect 57770 2030 57810 2045
rect 54915 1895 54955 1910
rect 54915 1625 54925 1895
rect 54945 1625 54955 1895
rect 54915 1610 54955 1625
rect 55655 1895 55695 1910
rect 55655 1625 55665 1895
rect 55685 1625 55695 1895
rect 58110 1895 58150 1910
rect 55655 1610 55695 1625
rect 55990 1695 56030 1710
rect 55990 1575 56000 1695
rect 56020 1575 56030 1695
rect 55990 1560 56030 1575
rect 56730 1695 56770 1710
rect 56730 1575 56740 1695
rect 56760 1575 56770 1695
rect 56730 1560 56770 1575
rect 57030 1695 57070 1710
rect 57030 1575 57040 1695
rect 57060 1575 57070 1695
rect 57030 1560 57070 1575
rect 57770 1695 57810 1710
rect 57770 1575 57780 1695
rect 57800 1575 57810 1695
rect 58110 1625 58120 1895
rect 58140 1625 58150 1895
rect 58110 1610 58150 1625
rect 58850 1895 58890 1910
rect 58850 1625 58860 1895
rect 58880 1625 58890 1895
rect 58850 1610 58890 1625
rect 57770 1560 57810 1575
rect 54945 1205 54985 1220
rect 54945 535 54955 1205
rect 54975 535 54985 1205
rect 54945 520 54985 535
rect 55625 1205 55665 1220
rect 55625 535 55635 1205
rect 55655 535 55665 1205
rect 58140 1205 58180 1220
rect 56180 1145 56220 1160
rect 56180 925 56190 1145
rect 56210 925 56220 1145
rect 56180 910 56220 925
rect 57525 1145 57565 1160
rect 57525 925 57535 1145
rect 57555 925 57565 1145
rect 57525 910 57565 925
rect 56390 680 56430 695
rect 56390 560 56400 680
rect 56420 560 56430 680
rect 56390 545 56430 560
rect 56800 680 56840 695
rect 56800 560 56810 680
rect 56830 560 56840 680
rect 56800 545 56840 560
rect 55625 520 55665 535
rect 58140 535 58150 1205
rect 58170 535 58180 1205
rect 58140 520 58180 535
rect 58820 1205 58860 1220
rect 58820 535 58830 1205
rect 58850 535 58860 1205
rect 58820 520 58860 535
<< nsubdiff >>
rect 56045 4695 56085 4710
rect 56045 4375 56055 4695
rect 56075 4375 56085 4695
rect 56045 4360 56085 4375
rect 56305 4695 56345 4710
rect 56305 4375 56315 4695
rect 56335 4375 56345 4695
rect 56985 4695 57025 4710
rect 56305 4360 56345 4375
rect 56515 4525 56555 4540
rect 56515 4375 56525 4525
rect 56545 4375 56555 4525
rect 56515 4360 56555 4375
rect 56775 4525 56815 4540
rect 56775 4375 56785 4525
rect 56805 4375 56815 4525
rect 56775 4360 56815 4375
rect 56985 4375 56995 4695
rect 57015 4375 57025 4695
rect 56985 4360 57025 4375
rect 57245 4695 57285 4710
rect 57245 4375 57255 4695
rect 57275 4375 57285 4695
rect 57245 4360 57285 4375
rect 57455 4695 57495 4710
rect 57455 4375 57465 4695
rect 57485 4375 57495 4695
rect 57455 4360 57495 4375
rect 57715 4695 57755 4710
rect 57715 4375 57725 4695
rect 57745 4375 57755 4695
rect 57715 4360 57755 4375
rect 54885 4025 54925 4040
rect 54885 3705 54895 4025
rect 54915 3705 54925 4025
rect 54885 3690 54925 3705
rect 55685 4025 55725 4040
rect 55685 3705 55695 4025
rect 55715 3705 55725 4025
rect 55685 3690 55725 3705
rect 55965 4025 56005 4040
rect 55965 3705 55975 4025
rect 55995 3705 56005 4025
rect 55965 3690 56005 3705
rect 56765 4025 56805 4040
rect 56765 3705 56775 4025
rect 56795 3705 56805 4025
rect 56765 3690 56805 3705
rect 56995 4025 57035 4040
rect 56995 3705 57005 4025
rect 57025 3705 57035 4025
rect 56995 3690 57035 3705
rect 57795 4025 57835 4040
rect 57795 3705 57805 4025
rect 57825 3705 57835 4025
rect 57795 3690 57835 3705
rect 58080 4025 58120 4040
rect 58080 3705 58090 4025
rect 58110 3705 58120 4025
rect 58080 3690 58120 3705
rect 58880 4025 58920 4040
rect 58880 3705 58890 4025
rect 58910 3705 58920 4025
rect 58880 3690 58920 3705
rect 54915 3250 54955 3265
rect 54915 2680 54925 3250
rect 54945 2680 54955 3250
rect 54915 2665 54955 2680
rect 55655 3250 55695 3265
rect 55655 2680 55665 3250
rect 55685 2680 55695 3250
rect 56235 3240 56275 3255
rect 56235 3220 56245 3240
rect 56265 3220 56275 3240
rect 56235 3205 56275 3220
rect 57525 3240 57565 3255
rect 57525 3220 57535 3240
rect 57555 3220 57565 3240
rect 57525 3205 57565 3220
rect 58110 3250 58150 3265
rect 55990 2930 56030 2945
rect 55990 2910 56000 2930
rect 56020 2910 56030 2930
rect 55990 2895 56030 2910
rect 56730 2930 56770 2945
rect 56730 2910 56740 2930
rect 56760 2910 56770 2930
rect 56730 2895 56770 2910
rect 57030 2930 57070 2945
rect 57030 2910 57040 2930
rect 57060 2910 57070 2930
rect 57030 2895 57070 2910
rect 57770 2930 57810 2945
rect 57770 2910 57780 2930
rect 57800 2910 57810 2930
rect 57770 2895 57810 2910
rect 55655 2665 55695 2680
rect 58110 2680 58120 3250
rect 58140 2680 58150 3250
rect 58110 2665 58150 2680
rect 58850 3250 58890 3265
rect 58850 2680 58860 3250
rect 58880 2680 58890 3250
rect 58850 2665 58890 2680
rect 54915 2355 54955 2370
rect 54915 2185 54925 2355
rect 54945 2185 54955 2355
rect 54915 2170 54955 2185
rect 55655 2355 55695 2370
rect 55655 2185 55665 2355
rect 55685 2185 55695 2355
rect 58110 2355 58150 2370
rect 55655 2170 55695 2185
rect 58110 2185 58120 2355
rect 58140 2185 58150 2355
rect 58110 2170 58150 2185
rect 58850 2355 58890 2370
rect 58850 2185 58860 2355
rect 58880 2185 58890 2355
rect 58850 2170 58890 2185
<< psubdiffcont >>
rect 56520 2550 56540 2570
rect 57260 2550 57280 2570
rect 56000 2045 56020 2165
rect 56740 2045 56760 2165
rect 57040 2045 57060 2165
rect 57780 2045 57800 2165
rect 54925 1625 54945 1895
rect 55665 1625 55685 1895
rect 56000 1575 56020 1695
rect 56740 1575 56760 1695
rect 57040 1575 57060 1695
rect 57780 1575 57800 1695
rect 58120 1625 58140 1895
rect 58860 1625 58880 1895
rect 54955 535 54975 1205
rect 55635 535 55655 1205
rect 56190 925 56210 1145
rect 57535 925 57555 1145
rect 56400 560 56420 680
rect 56810 560 56830 680
rect 58150 535 58170 1205
rect 58830 535 58850 1205
<< nsubdiffcont >>
rect 56055 4375 56075 4695
rect 56315 4375 56335 4695
rect 56525 4375 56545 4525
rect 56785 4375 56805 4525
rect 56995 4375 57015 4695
rect 57255 4375 57275 4695
rect 57465 4375 57485 4695
rect 57725 4375 57745 4695
rect 54895 3705 54915 4025
rect 55695 3705 55715 4025
rect 55975 3705 55995 4025
rect 56775 3705 56795 4025
rect 57005 3705 57025 4025
rect 57805 3705 57825 4025
rect 58090 3705 58110 4025
rect 58890 3705 58910 4025
rect 54925 2680 54945 3250
rect 55665 2680 55685 3250
rect 56245 3220 56265 3240
rect 57535 3220 57555 3240
rect 56000 2910 56020 2930
rect 56740 2910 56760 2930
rect 57040 2910 57060 2930
rect 57780 2910 57800 2930
rect 58120 2680 58140 3250
rect 58860 2680 58880 3250
rect 54925 2185 54945 2355
rect 55665 2185 55685 2355
rect 58120 2185 58140 2355
rect 58860 2185 58880 2355
<< poly >>
rect 56085 4755 56125 4765
rect 56085 4735 56095 4755
rect 56115 4740 56125 4755
rect 56265 4755 56305 4765
rect 56265 4740 56275 4755
rect 56115 4735 56145 4740
rect 56085 4725 56145 4735
rect 56245 4735 56275 4740
rect 56295 4735 56305 4755
rect 56245 4725 56305 4735
rect 57025 4755 57065 4765
rect 57025 4735 57035 4755
rect 57055 4740 57065 4755
rect 57205 4755 57245 4765
rect 57205 4740 57215 4755
rect 57055 4735 57085 4740
rect 57025 4725 57085 4735
rect 57185 4735 57215 4740
rect 57235 4735 57245 4755
rect 57185 4725 57245 4735
rect 57495 4755 57535 4765
rect 57495 4735 57505 4755
rect 57525 4740 57535 4755
rect 57675 4755 57715 4765
rect 57675 4740 57685 4755
rect 57525 4735 57555 4740
rect 57495 4725 57555 4735
rect 57655 4735 57685 4740
rect 57705 4735 57715 4755
rect 57655 4725 57715 4735
rect 56125 4710 56145 4725
rect 56185 4710 56205 4725
rect 56245 4710 56265 4725
rect 57065 4710 57085 4725
rect 57125 4710 57145 4725
rect 57185 4710 57205 4725
rect 57535 4710 57555 4725
rect 57595 4710 57615 4725
rect 57655 4710 57675 4725
rect 56555 4585 56595 4595
rect 56555 4565 56565 4585
rect 56585 4570 56595 4585
rect 56735 4585 56775 4595
rect 56735 4570 56745 4585
rect 56585 4565 56615 4570
rect 56555 4555 56615 4565
rect 56715 4565 56745 4570
rect 56765 4565 56775 4585
rect 56715 4555 56775 4565
rect 56595 4540 56615 4555
rect 56655 4540 56675 4555
rect 56715 4540 56735 4555
rect 56125 4345 56145 4360
rect 56185 4315 56205 4360
rect 56245 4345 56265 4360
rect 56595 4345 56615 4360
rect 56655 4315 56675 4360
rect 56715 4345 56735 4360
rect 57065 4345 57085 4360
rect 56150 4305 56205 4315
rect 56150 4285 56160 4305
rect 56180 4285 56205 4305
rect 56150 4275 56205 4285
rect 56630 4305 56675 4315
rect 56630 4285 56635 4305
rect 56655 4300 56675 4305
rect 57125 4315 57145 4360
rect 57185 4345 57205 4360
rect 57535 4345 57555 4360
rect 57125 4305 57170 4315
rect 57595 4305 57615 4360
rect 57655 4345 57675 4360
rect 57125 4300 57145 4305
rect 56655 4285 56660 4300
rect 56630 4275 56660 4285
rect 57140 4285 57145 4300
rect 57165 4285 57170 4305
rect 57140 4275 57170 4285
rect 57576 4295 57615 4305
rect 57576 4275 57581 4295
rect 57601 4290 57615 4295
rect 57601 4275 57606 4290
rect 57576 4265 57606 4275
rect 54965 4040 54985 4055
rect 55025 4040 55045 4055
rect 55085 4040 55105 4055
rect 55145 4040 55165 4055
rect 55205 4040 55225 4055
rect 55265 4040 55285 4055
rect 55325 4040 55345 4055
rect 55385 4040 55405 4055
rect 55445 4040 55465 4055
rect 55505 4040 55525 4055
rect 55565 4040 55585 4055
rect 55625 4040 55645 4055
rect 56045 4040 56065 4055
rect 56105 4040 56125 4055
rect 56165 4040 56185 4055
rect 56225 4040 56245 4055
rect 56285 4040 56305 4055
rect 56345 4040 56365 4055
rect 56405 4040 56425 4055
rect 56465 4040 56485 4055
rect 56525 4040 56545 4055
rect 56585 4040 56605 4055
rect 56645 4040 56665 4055
rect 56705 4040 56725 4055
rect 57075 4040 57095 4055
rect 57135 4040 57155 4055
rect 57195 4040 57215 4055
rect 57255 4040 57275 4055
rect 57315 4040 57335 4055
rect 57375 4040 57395 4055
rect 57435 4040 57455 4055
rect 57495 4040 57515 4055
rect 57555 4040 57575 4055
rect 57615 4040 57635 4055
rect 57675 4040 57695 4055
rect 57735 4040 57755 4055
rect 58160 4040 58180 4055
rect 58220 4040 58240 4055
rect 58280 4040 58300 4055
rect 58340 4040 58360 4055
rect 58400 4040 58420 4055
rect 58460 4040 58480 4055
rect 58520 4040 58540 4055
rect 58580 4040 58600 4055
rect 58640 4040 58660 4055
rect 58700 4040 58720 4055
rect 58760 4040 58780 4055
rect 58820 4040 58840 4055
rect 54965 3675 54985 3690
rect 54930 3665 54985 3675
rect 55025 3680 55045 3690
rect 55085 3680 55105 3690
rect 55145 3680 55165 3690
rect 55205 3680 55225 3690
rect 55265 3680 55285 3690
rect 55325 3680 55345 3690
rect 55385 3680 55405 3690
rect 55445 3680 55465 3690
rect 55505 3680 55525 3690
rect 55565 3680 55585 3690
rect 55025 3665 55585 3680
rect 55625 3675 55645 3690
rect 56045 3675 56065 3690
rect 55625 3665 55680 3675
rect 54930 3645 54935 3665
rect 54955 3660 54985 3665
rect 54955 3645 54960 3660
rect 54930 3635 54960 3645
rect 55290 3645 55295 3665
rect 55315 3645 55320 3665
rect 55625 3660 55655 3665
rect 55290 3635 55320 3645
rect 55650 3645 55655 3660
rect 55675 3645 55680 3665
rect 55650 3635 55680 3645
rect 56010 3665 56065 3675
rect 56105 3680 56125 3690
rect 56165 3680 56185 3690
rect 56225 3680 56245 3690
rect 56285 3680 56305 3690
rect 56345 3680 56365 3690
rect 56405 3680 56425 3690
rect 56465 3680 56485 3690
rect 56525 3680 56545 3690
rect 56585 3680 56605 3690
rect 56645 3680 56665 3690
rect 56105 3665 56665 3680
rect 56705 3675 56725 3690
rect 57075 3675 57095 3690
rect 56705 3665 56760 3675
rect 56010 3645 56015 3665
rect 56035 3660 56065 3665
rect 56035 3645 56040 3660
rect 56010 3635 56040 3645
rect 56370 3645 56375 3665
rect 56395 3645 56400 3665
rect 56705 3660 56735 3665
rect 56370 3635 56400 3645
rect 56730 3645 56735 3660
rect 56755 3645 56760 3665
rect 56730 3635 56760 3645
rect 57040 3665 57095 3675
rect 57135 3680 57155 3690
rect 57195 3680 57215 3690
rect 57255 3680 57275 3690
rect 57315 3680 57335 3690
rect 57375 3680 57395 3690
rect 57435 3680 57455 3690
rect 57495 3680 57515 3690
rect 57555 3680 57575 3690
rect 57615 3680 57635 3690
rect 57675 3680 57695 3690
rect 57135 3665 57695 3680
rect 57735 3675 57755 3690
rect 58160 3675 58180 3690
rect 57735 3665 57790 3675
rect 57040 3645 57045 3665
rect 57065 3660 57095 3665
rect 57065 3645 57070 3660
rect 57040 3635 57070 3645
rect 57400 3645 57405 3665
rect 57425 3645 57430 3665
rect 57735 3660 57765 3665
rect 57400 3635 57430 3645
rect 57760 3645 57765 3660
rect 57785 3645 57790 3665
rect 57760 3635 57790 3645
rect 58125 3665 58180 3675
rect 58220 3680 58240 3690
rect 58280 3680 58300 3690
rect 58340 3680 58360 3690
rect 58400 3680 58420 3690
rect 58460 3680 58480 3690
rect 58520 3680 58540 3690
rect 58580 3680 58600 3690
rect 58640 3680 58660 3690
rect 58700 3680 58720 3690
rect 58760 3680 58780 3690
rect 58220 3665 58780 3680
rect 58820 3675 58840 3690
rect 58820 3665 58875 3675
rect 58125 3645 58130 3665
rect 58150 3660 58180 3665
rect 58150 3645 58155 3660
rect 58125 3635 58155 3645
rect 58485 3645 58490 3665
rect 58510 3645 58515 3665
rect 58820 3660 58850 3665
rect 58485 3635 58515 3645
rect 58845 3645 58850 3660
rect 58870 3645 58875 3665
rect 58845 3635 58875 3645
rect 55295 3565 55315 3635
rect 56375 3610 56395 3635
rect 57405 3610 57425 3635
rect 56365 3600 56405 3610
rect 56365 3580 56375 3600
rect 56395 3580 56405 3600
rect 56365 3570 56405 3580
rect 57395 3600 57435 3610
rect 57395 3580 57405 3600
rect 57425 3580 57435 3600
rect 57395 3570 57435 3580
rect 58490 3565 58510 3635
rect 55285 3555 55325 3565
rect 55285 3535 55295 3555
rect 55315 3535 55325 3555
rect 55285 3525 55325 3535
rect 58480 3555 58520 3565
rect 58480 3535 58490 3555
rect 58510 3535 58520 3555
rect 58480 3525 58520 3535
rect 54960 3310 54990 3320
rect 54960 3290 54965 3310
rect 54985 3295 54990 3310
rect 55620 3310 55650 3320
rect 55620 3295 55625 3310
rect 54985 3290 55010 3295
rect 54960 3280 55010 3290
rect 55600 3290 55625 3295
rect 55645 3290 55650 3310
rect 55600 3280 55650 3290
rect 58155 3310 58185 3320
rect 58155 3290 58160 3310
rect 58180 3295 58185 3310
rect 58815 3310 58845 3320
rect 58815 3295 58820 3310
rect 58180 3290 58205 3295
rect 58155 3280 58205 3290
rect 58795 3290 58820 3295
rect 58840 3290 58845 3310
rect 58795 3280 58845 3290
rect 54995 3265 55010 3280
rect 55050 3265 55065 3280
rect 55105 3265 55120 3280
rect 55160 3265 55175 3280
rect 55215 3265 55230 3280
rect 55270 3265 55285 3280
rect 55325 3265 55340 3280
rect 55380 3265 55395 3280
rect 55435 3265 55450 3280
rect 55490 3265 55505 3280
rect 55545 3265 55560 3280
rect 55600 3265 55615 3280
rect 56315 3255 56330 3270
rect 56370 3255 56385 3270
rect 56425 3255 56440 3270
rect 56480 3255 56495 3270
rect 56535 3255 56550 3270
rect 56590 3255 56605 3270
rect 56645 3255 56660 3270
rect 56700 3255 56715 3270
rect 56755 3255 56770 3270
rect 56810 3255 56825 3270
rect 56865 3255 56880 3270
rect 56920 3255 56935 3270
rect 56975 3255 56990 3270
rect 57030 3255 57045 3270
rect 57085 3255 57100 3270
rect 57140 3255 57155 3270
rect 57195 3255 57210 3270
rect 57250 3255 57265 3270
rect 57305 3255 57320 3270
rect 57360 3255 57375 3270
rect 57415 3255 57430 3270
rect 57470 3255 57485 3270
rect 58190 3265 58205 3280
rect 58245 3265 58260 3280
rect 58300 3265 58315 3280
rect 58355 3265 58370 3280
rect 58410 3265 58425 3280
rect 58465 3265 58480 3280
rect 58520 3265 58535 3280
rect 58575 3265 58590 3280
rect 58630 3265 58645 3280
rect 58685 3265 58700 3280
rect 58740 3265 58755 3280
rect 58795 3265 58810 3280
rect 56315 3190 56330 3205
rect 56280 3180 56330 3190
rect 56370 3195 56385 3205
rect 56425 3195 56440 3205
rect 56480 3195 56495 3205
rect 56535 3195 56550 3205
rect 56590 3195 56605 3205
rect 56645 3195 56660 3205
rect 56700 3195 56715 3205
rect 56755 3195 56770 3205
rect 56810 3195 56825 3205
rect 56865 3195 56880 3205
rect 56920 3195 56935 3205
rect 56975 3195 56990 3205
rect 57030 3195 57045 3205
rect 57085 3195 57100 3205
rect 57140 3195 57155 3205
rect 57195 3195 57210 3205
rect 57250 3195 57265 3205
rect 57305 3195 57320 3205
rect 57360 3195 57375 3205
rect 57415 3195 57430 3205
rect 56370 3180 57430 3195
rect 57470 3190 57485 3205
rect 57470 3180 57520 3190
rect 56280 3160 56285 3180
rect 56305 3175 56330 3180
rect 56305 3160 56310 3175
rect 56280 3150 56310 3160
rect 56390 3160 56395 3180
rect 56415 3160 56420 3180
rect 56390 3150 56420 3160
rect 56830 3160 56835 3180
rect 56855 3160 56860 3180
rect 57470 3175 57495 3180
rect 56830 3150 56860 3160
rect 57490 3160 57495 3175
rect 57515 3160 57520 3180
rect 57490 3150 57520 3160
rect 56040 3015 56070 3025
rect 56040 2995 56045 3015
rect 56065 3000 56070 3015
rect 56690 3015 56720 3025
rect 56690 3000 56695 3015
rect 56065 2995 56695 3000
rect 56715 2995 56720 3015
rect 56040 2985 56720 2995
rect 57080 3015 57110 3025
rect 57080 2995 57085 3015
rect 57105 3000 57110 3015
rect 57730 3015 57760 3025
rect 57730 3000 57735 3015
rect 57105 2995 57735 3000
rect 57755 2995 57760 3015
rect 57080 2985 57760 2995
rect 56070 2945 56085 2960
rect 56125 2945 56140 2960
rect 56180 2945 56195 2985
rect 56235 2945 56250 2985
rect 56290 2945 56305 2960
rect 56345 2945 56360 2960
rect 56400 2945 56415 2985
rect 56455 2945 56470 2985
rect 56510 2945 56525 2960
rect 56565 2945 56580 2960
rect 56620 2945 56635 2985
rect 56675 2945 56690 2960
rect 57110 2945 57125 2960
rect 57165 2945 57180 2985
rect 57220 2945 57235 2960
rect 57275 2945 57290 2960
rect 57330 2945 57345 2985
rect 57385 2945 57400 2985
rect 57440 2945 57455 2960
rect 57495 2945 57510 2960
rect 57550 2945 57565 2985
rect 57605 2945 57620 2985
rect 57660 2945 57675 2960
rect 57715 2945 57730 2960
rect 56070 2880 56085 2895
rect 56035 2870 56085 2880
rect 56035 2850 56040 2870
rect 56060 2865 56085 2870
rect 56060 2850 56065 2865
rect 56035 2840 56065 2850
rect 56125 2855 56140 2895
rect 56180 2880 56195 2895
rect 56235 2880 56250 2895
rect 56290 2855 56305 2895
rect 56345 2855 56360 2895
rect 56400 2880 56415 2895
rect 56455 2880 56470 2895
rect 56510 2855 56525 2895
rect 56565 2855 56580 2895
rect 56620 2880 56635 2895
rect 56675 2880 56690 2895
rect 57110 2880 57125 2895
rect 57165 2880 57180 2895
rect 56675 2870 56725 2880
rect 56675 2865 56700 2870
rect 56125 2840 56580 2855
rect 56695 2850 56700 2865
rect 56720 2850 56725 2870
rect 56695 2840 56725 2850
rect 57075 2870 57125 2880
rect 57075 2850 57080 2870
rect 57100 2865 57125 2870
rect 57100 2850 57105 2865
rect 57075 2840 57105 2850
rect 57220 2855 57235 2895
rect 57275 2855 57290 2895
rect 57330 2880 57345 2895
rect 57385 2880 57400 2895
rect 57440 2855 57455 2895
rect 57495 2855 57510 2895
rect 57550 2880 57565 2895
rect 57605 2880 57620 2895
rect 57660 2855 57675 2895
rect 57715 2880 57730 2895
rect 57715 2870 57765 2880
rect 57715 2865 57740 2870
rect 57220 2840 57675 2855
rect 57735 2850 57740 2865
rect 57760 2850 57765 2870
rect 57735 2840 57765 2850
rect 56125 2795 56140 2840
rect 56095 2785 56140 2795
rect 56095 2765 56100 2785
rect 56120 2775 56140 2785
rect 56565 2795 56580 2840
rect 57220 2795 57235 2840
rect 56565 2785 56610 2795
rect 56565 2775 56585 2785
rect 56120 2765 56125 2775
rect 56095 2755 56125 2765
rect 56580 2765 56585 2775
rect 56605 2765 56610 2785
rect 56580 2755 56610 2765
rect 57190 2785 57235 2795
rect 57190 2765 57195 2785
rect 57215 2775 57235 2785
rect 57215 2765 57220 2775
rect 57190 2755 57220 2765
rect 54995 2650 55010 2665
rect 55050 2655 55065 2665
rect 55105 2655 55120 2665
rect 55160 2655 55175 2665
rect 55215 2655 55230 2665
rect 55270 2655 55285 2665
rect 55325 2655 55340 2665
rect 55380 2655 55395 2665
rect 55435 2655 55450 2665
rect 55490 2655 55505 2665
rect 55545 2655 55560 2665
rect 55050 2640 55560 2655
rect 55600 2650 55615 2665
rect 58190 2650 58205 2665
rect 58245 2655 58260 2665
rect 58300 2655 58315 2665
rect 58355 2655 58370 2665
rect 58410 2655 58425 2665
rect 58465 2655 58480 2665
rect 58520 2655 58535 2665
rect 58575 2655 58590 2665
rect 58630 2655 58645 2665
rect 58685 2655 58700 2665
rect 58740 2655 58755 2665
rect 58245 2640 58755 2655
rect 58795 2650 58810 2665
rect 55180 2620 55185 2640
rect 55205 2620 55210 2640
rect 55180 2610 55210 2620
rect 56715 2630 56755 2640
rect 56715 2610 56725 2630
rect 56745 2610 56755 2630
rect 56935 2630 56975 2640
rect 56935 2610 56945 2630
rect 56965 2610 56975 2630
rect 58595 2620 58600 2640
rect 58620 2620 58625 2640
rect 58595 2610 58625 2620
rect 55185 2585 55205 2610
rect 56590 2585 56605 2600
rect 56645 2595 57155 2610
rect 56645 2585 56660 2595
rect 56700 2585 56715 2595
rect 56755 2585 56770 2595
rect 56810 2585 56825 2595
rect 56865 2585 56880 2595
rect 56920 2585 56935 2595
rect 56975 2585 56990 2595
rect 57030 2585 57045 2595
rect 57085 2585 57100 2595
rect 57140 2585 57155 2595
rect 57195 2585 57210 2600
rect 58600 2585 58620 2610
rect 55175 2580 55215 2585
rect 55175 2560 55185 2580
rect 55205 2560 55215 2580
rect 55175 2555 55215 2560
rect 58590 2580 58630 2585
rect 58590 2560 58600 2580
rect 58620 2560 58630 2580
rect 58590 2555 58630 2560
rect 56590 2520 56605 2535
rect 56645 2520 56660 2535
rect 56700 2520 56715 2535
rect 56755 2520 56770 2535
rect 56810 2520 56825 2535
rect 56865 2520 56880 2535
rect 56920 2520 56935 2535
rect 56975 2520 56990 2535
rect 57030 2520 57045 2535
rect 57085 2520 57100 2535
rect 57140 2520 57155 2535
rect 57195 2520 57210 2535
rect 56550 2510 56605 2520
rect 56550 2490 56560 2510
rect 56580 2505 56605 2510
rect 57195 2510 57250 2520
rect 57195 2505 57220 2510
rect 56580 2490 56590 2505
rect 56550 2480 56590 2490
rect 57210 2490 57220 2505
rect 57240 2490 57250 2510
rect 57210 2480 57250 2490
rect 54960 2415 54990 2425
rect 54960 2395 54965 2415
rect 54985 2400 54990 2415
rect 55620 2415 55650 2425
rect 55620 2400 55625 2415
rect 54985 2395 55010 2400
rect 54960 2385 55010 2395
rect 55600 2395 55625 2400
rect 55645 2395 55650 2415
rect 55600 2385 55650 2395
rect 58155 2415 58185 2425
rect 58155 2395 58160 2415
rect 58180 2400 58185 2415
rect 58815 2415 58845 2425
rect 58815 2400 58820 2415
rect 58180 2395 58205 2400
rect 58155 2385 58205 2395
rect 58795 2395 58820 2400
rect 58840 2395 58845 2415
rect 58795 2385 58845 2395
rect 54995 2370 55010 2385
rect 55050 2370 55065 2385
rect 55105 2370 55120 2385
rect 55160 2370 55175 2385
rect 55215 2370 55230 2385
rect 55270 2370 55285 2385
rect 55325 2370 55340 2385
rect 55380 2370 55395 2385
rect 55435 2370 55450 2385
rect 55490 2370 55505 2385
rect 55545 2370 55560 2385
rect 55600 2370 55615 2385
rect 58190 2370 58205 2385
rect 58245 2370 58260 2385
rect 58300 2370 58315 2385
rect 58355 2370 58370 2385
rect 58410 2370 58425 2385
rect 58465 2370 58480 2385
rect 58520 2370 58535 2385
rect 58575 2370 58590 2385
rect 58630 2370 58645 2385
rect 58685 2370 58700 2385
rect 58740 2370 58755 2385
rect 58795 2370 58810 2385
rect 56095 2265 56125 2275
rect 56095 2245 56100 2265
rect 56120 2250 56125 2265
rect 56635 2265 56665 2275
rect 56635 2250 56640 2265
rect 56120 2245 56140 2250
rect 56095 2235 56140 2245
rect 56125 2205 56140 2235
rect 56620 2245 56640 2250
rect 56660 2245 56665 2265
rect 56620 2235 56665 2245
rect 57135 2265 57165 2275
rect 57135 2245 57140 2265
rect 57160 2250 57165 2265
rect 57160 2245 57180 2250
rect 57135 2235 57180 2245
rect 56620 2205 56635 2235
rect 56070 2180 56085 2195
rect 56125 2190 56635 2205
rect 57165 2205 57180 2235
rect 56125 2180 56140 2190
rect 56180 2180 56195 2190
rect 56235 2180 56250 2190
rect 56290 2180 56305 2190
rect 56345 2180 56360 2190
rect 56400 2180 56415 2190
rect 56455 2180 56470 2190
rect 56510 2180 56525 2190
rect 56565 2180 56580 2190
rect 56620 2180 56635 2190
rect 56675 2180 56690 2195
rect 57110 2180 57125 2195
rect 57165 2190 57675 2205
rect 57165 2180 57180 2190
rect 57220 2180 57235 2190
rect 57275 2180 57290 2190
rect 57330 2180 57345 2190
rect 57385 2180 57400 2190
rect 57440 2180 57455 2190
rect 57495 2180 57510 2190
rect 57550 2180 57565 2190
rect 57605 2180 57620 2190
rect 57660 2180 57675 2190
rect 57715 2180 57730 2195
rect 54995 2155 55010 2170
rect 55050 2160 55065 2170
rect 55105 2160 55120 2170
rect 55160 2160 55175 2170
rect 55215 2160 55230 2170
rect 55270 2160 55285 2170
rect 55325 2160 55340 2170
rect 55380 2160 55395 2170
rect 55435 2160 55450 2170
rect 55490 2160 55505 2170
rect 55545 2160 55560 2170
rect 55050 2145 55560 2160
rect 55600 2155 55615 2170
rect 55455 2125 55460 2145
rect 55480 2125 55485 2145
rect 55455 2115 55485 2125
rect 55460 2060 55480 2115
rect 55450 2050 55490 2060
rect 55450 2030 55460 2050
rect 55480 2030 55490 2050
rect 58190 2155 58205 2170
rect 58245 2160 58260 2170
rect 58300 2160 58315 2170
rect 58355 2160 58370 2170
rect 58410 2160 58425 2170
rect 58465 2160 58480 2170
rect 58520 2160 58535 2170
rect 58575 2160 58590 2170
rect 58630 2160 58645 2170
rect 58685 2160 58700 2170
rect 58740 2160 58755 2170
rect 58245 2145 58755 2160
rect 58795 2155 58810 2170
rect 58320 2125 58325 2145
rect 58345 2125 58350 2145
rect 58320 2115 58350 2125
rect 58325 2060 58345 2115
rect 58315 2050 58355 2060
rect 58315 2030 58325 2050
rect 58345 2030 58355 2050
rect 55450 2020 55490 2030
rect 55460 1965 55480 2020
rect 56070 2015 56085 2030
rect 56125 2015 56140 2030
rect 56180 2015 56195 2030
rect 56235 2015 56250 2030
rect 56290 2015 56305 2030
rect 56345 2015 56360 2030
rect 56400 2015 56415 2030
rect 56455 2015 56470 2030
rect 56510 2015 56525 2030
rect 56565 2015 56580 2030
rect 56620 2015 56635 2030
rect 56675 2015 56690 2030
rect 57110 2015 57125 2030
rect 57165 2015 57180 2030
rect 57220 2015 57235 2030
rect 57275 2015 57290 2030
rect 57330 2015 57345 2030
rect 57385 2015 57400 2030
rect 57440 2015 57455 2030
rect 57495 2015 57510 2030
rect 57550 2015 57565 2030
rect 57605 2015 57620 2030
rect 57660 2015 57675 2030
rect 57715 2015 57730 2030
rect 58315 2020 58355 2030
rect 56035 2005 56085 2015
rect 56035 1985 56040 2005
rect 56060 2000 56085 2005
rect 56675 2005 56725 2015
rect 56675 2000 56700 2005
rect 56060 1985 56065 2000
rect 56035 1975 56065 1985
rect 56695 1985 56700 2000
rect 56720 1985 56725 2005
rect 56695 1975 56725 1985
rect 57075 2005 57125 2015
rect 57075 1985 57080 2005
rect 57100 2000 57125 2005
rect 57715 2005 57765 2015
rect 57715 2000 57740 2005
rect 57100 1985 57105 2000
rect 57075 1975 57105 1985
rect 57735 1985 57740 2000
rect 57760 1985 57765 2005
rect 57735 1975 57765 1985
rect 58325 1965 58345 2020
rect 55455 1955 55485 1965
rect 55455 1935 55460 1955
rect 55480 1935 55485 1955
rect 58320 1955 58350 1965
rect 58320 1935 58325 1955
rect 58345 1935 58350 1955
rect 54995 1910 55010 1925
rect 55050 1920 55560 1935
rect 55050 1910 55065 1920
rect 55105 1910 55120 1920
rect 55160 1910 55175 1920
rect 55215 1910 55230 1920
rect 55270 1910 55285 1920
rect 55325 1910 55340 1920
rect 55380 1910 55395 1920
rect 55435 1910 55450 1920
rect 55490 1910 55505 1920
rect 55545 1910 55560 1920
rect 55600 1910 55615 1925
rect 58190 1910 58205 1925
rect 58245 1920 58755 1935
rect 58245 1910 58260 1920
rect 58300 1910 58315 1920
rect 58355 1910 58370 1920
rect 58410 1910 58425 1920
rect 58465 1910 58480 1920
rect 58520 1910 58535 1920
rect 58575 1910 58590 1920
rect 58630 1910 58645 1920
rect 58685 1910 58700 1920
rect 58740 1910 58755 1920
rect 58795 1910 58810 1925
rect 56040 1780 56070 1790
rect 56040 1760 56045 1780
rect 56065 1765 56070 1780
rect 56690 1780 56720 1790
rect 56690 1765 56695 1780
rect 56065 1760 56140 1765
rect 56040 1750 56140 1760
rect 56125 1735 56140 1750
rect 56620 1760 56695 1765
rect 56715 1760 56720 1780
rect 56620 1750 56720 1760
rect 56850 1780 56880 1790
rect 56850 1760 56855 1780
rect 56875 1760 56880 1780
rect 56850 1750 56880 1760
rect 56903 1780 56933 1790
rect 56903 1760 56908 1780
rect 56928 1760 56933 1780
rect 57080 1780 57110 1790
rect 57080 1760 57085 1780
rect 57105 1765 57110 1780
rect 57730 1780 57760 1790
rect 57730 1765 57735 1780
rect 57105 1760 57180 1765
rect 56903 1750 56935 1760
rect 57080 1750 57180 1760
rect 56620 1735 56635 1750
rect 56070 1710 56085 1725
rect 56125 1720 56635 1735
rect 56125 1710 56140 1720
rect 56180 1710 56195 1720
rect 56235 1710 56250 1720
rect 56290 1710 56305 1720
rect 56345 1710 56360 1720
rect 56400 1710 56415 1720
rect 56455 1710 56470 1720
rect 56510 1710 56525 1720
rect 56565 1710 56580 1720
rect 56620 1710 56635 1720
rect 56675 1710 56690 1725
rect 56810 1710 56825 1725
rect 56865 1710 56880 1750
rect 56920 1710 56935 1750
rect 57165 1735 57180 1750
rect 57660 1760 57735 1765
rect 57755 1760 57760 1780
rect 57660 1750 57760 1760
rect 57660 1735 57675 1750
rect 56975 1710 56990 1725
rect 57110 1710 57125 1725
rect 57165 1720 57675 1735
rect 57165 1710 57180 1720
rect 57220 1710 57235 1720
rect 57275 1710 57290 1720
rect 57330 1710 57345 1720
rect 57385 1710 57400 1720
rect 57440 1710 57455 1720
rect 57495 1710 57510 1720
rect 57550 1710 57565 1720
rect 57605 1710 57620 1720
rect 57660 1710 57675 1720
rect 57715 1710 57730 1725
rect 54995 1595 55010 1610
rect 55050 1595 55065 1610
rect 55105 1595 55120 1610
rect 55160 1595 55175 1610
rect 55215 1595 55230 1610
rect 55270 1595 55285 1610
rect 55325 1595 55340 1610
rect 55380 1595 55395 1610
rect 55435 1595 55450 1610
rect 55490 1595 55505 1610
rect 55545 1595 55560 1610
rect 55600 1595 55615 1610
rect 54960 1585 55010 1595
rect 54960 1565 54965 1585
rect 54985 1580 55010 1585
rect 55600 1585 55650 1595
rect 55600 1580 55625 1585
rect 54985 1565 54990 1580
rect 54960 1555 54990 1565
rect 55620 1565 55625 1580
rect 55645 1565 55650 1585
rect 55620 1555 55650 1565
rect 58190 1595 58205 1610
rect 58245 1595 58260 1610
rect 58300 1595 58315 1610
rect 58355 1595 58370 1610
rect 58410 1595 58425 1610
rect 58465 1595 58480 1610
rect 58520 1595 58535 1610
rect 58575 1595 58590 1610
rect 58630 1595 58645 1610
rect 58685 1595 58700 1610
rect 58740 1595 58755 1610
rect 58795 1595 58810 1610
rect 58155 1585 58205 1595
rect 58155 1565 58160 1585
rect 58180 1580 58205 1585
rect 58795 1585 58845 1595
rect 58795 1580 58820 1585
rect 58180 1565 58185 1580
rect 56070 1545 56085 1560
rect 56125 1545 56140 1560
rect 56180 1545 56195 1560
rect 56235 1545 56250 1560
rect 56290 1545 56305 1560
rect 56345 1545 56360 1560
rect 56400 1545 56415 1560
rect 56455 1545 56470 1560
rect 56510 1545 56525 1560
rect 56565 1545 56580 1560
rect 56620 1545 56635 1560
rect 56675 1545 56690 1560
rect 56810 1545 56825 1560
rect 56865 1545 56880 1560
rect 56920 1545 56935 1560
rect 56975 1545 56990 1560
rect 57110 1545 57125 1560
rect 57165 1545 57180 1560
rect 57220 1545 57235 1560
rect 57275 1545 57290 1560
rect 57330 1545 57345 1560
rect 57385 1545 57400 1560
rect 57440 1545 57455 1560
rect 57495 1545 57510 1560
rect 57550 1545 57565 1560
rect 57605 1545 57620 1560
rect 57660 1545 57675 1560
rect 57715 1545 57730 1560
rect 58155 1555 58185 1565
rect 58815 1565 58820 1580
rect 58840 1565 58845 1585
rect 58815 1555 58845 1565
rect 56035 1535 56085 1545
rect 56035 1515 56040 1535
rect 56060 1530 56085 1535
rect 56675 1535 56825 1545
rect 56675 1530 56740 1535
rect 56060 1515 56065 1530
rect 56035 1505 56065 1515
rect 56735 1515 56740 1530
rect 56760 1530 56825 1535
rect 56975 1535 57125 1545
rect 56975 1530 57040 1535
rect 56760 1515 56765 1530
rect 56735 1505 56765 1515
rect 57035 1515 57040 1530
rect 57060 1530 57125 1535
rect 57715 1535 57765 1545
rect 57715 1530 57740 1535
rect 57060 1515 57065 1530
rect 57035 1505 57065 1515
rect 57735 1515 57740 1530
rect 57760 1515 57765 1535
rect 57735 1505 57765 1515
rect 55385 1265 55425 1275
rect 55385 1245 55395 1265
rect 55415 1245 55425 1265
rect 57405 1260 57445 1270
rect 55025 1220 55085 1235
rect 55125 1230 55485 1245
rect 57405 1240 57415 1260
rect 57435 1240 57445 1260
rect 58435 1265 58465 1275
rect 58435 1245 58440 1265
rect 58460 1245 58465 1265
rect 55125 1220 55185 1230
rect 55225 1220 55285 1230
rect 55325 1220 55385 1230
rect 55425 1220 55485 1230
rect 55525 1220 55585 1235
rect 57405 1230 57445 1240
rect 56830 1205 56860 1215
rect 56830 1185 56835 1205
rect 56855 1185 56860 1205
rect 56260 1160 56275 1175
rect 56315 1170 57375 1185
rect 56315 1160 56330 1170
rect 56370 1160 56385 1170
rect 56425 1160 56440 1170
rect 56480 1160 56495 1170
rect 56535 1160 56550 1170
rect 56590 1160 56605 1170
rect 56645 1160 56660 1170
rect 56700 1160 56715 1170
rect 56755 1160 56770 1170
rect 56810 1160 56825 1170
rect 56865 1160 56880 1170
rect 56920 1160 56935 1170
rect 56975 1160 56990 1170
rect 57030 1160 57045 1170
rect 57085 1160 57100 1170
rect 57140 1160 57155 1170
rect 57195 1160 57210 1170
rect 57250 1160 57265 1170
rect 57305 1160 57320 1170
rect 57360 1160 57375 1170
rect 57415 1160 57430 1230
rect 58220 1220 58280 1235
rect 58320 1230 58680 1245
rect 58320 1220 58380 1230
rect 58420 1220 58480 1230
rect 58520 1220 58580 1230
rect 58620 1220 58680 1230
rect 58720 1220 58780 1235
rect 57470 1160 57485 1175
rect 56260 895 56275 910
rect 56315 895 56330 910
rect 56370 895 56385 910
rect 56425 895 56440 910
rect 56480 895 56495 910
rect 56535 895 56550 910
rect 56590 895 56605 910
rect 56645 895 56660 910
rect 56700 895 56715 910
rect 56755 895 56770 910
rect 56810 895 56825 910
rect 56865 895 56880 910
rect 56920 895 56935 910
rect 56975 895 56990 910
rect 57030 895 57045 910
rect 57085 895 57100 910
rect 57140 895 57155 910
rect 57195 895 57210 910
rect 57250 895 57265 910
rect 57305 895 57320 910
rect 57360 895 57375 910
rect 57415 895 57430 910
rect 57470 895 57485 910
rect 56220 885 56275 895
rect 56220 865 56230 885
rect 56250 880 56275 885
rect 57470 885 57525 895
rect 57470 880 57495 885
rect 56250 865 56260 880
rect 56220 855 56260 865
rect 57485 865 57495 880
rect 57515 865 57525 885
rect 57485 855 57525 865
rect 56595 740 56635 750
rect 56595 720 56605 740
rect 56625 720 56635 740
rect 57040 740 57080 750
rect 57040 720 57050 740
rect 57070 720 57080 740
rect 56470 695 56485 710
rect 56525 705 56705 720
rect 57040 710 57080 720
rect 56525 695 56540 705
rect 56580 695 56595 705
rect 56635 695 56650 705
rect 56690 695 56705 705
rect 56745 695 56760 710
rect 56910 695 57210 710
rect 56470 530 56485 545
rect 56525 530 56540 545
rect 56580 530 56595 545
rect 56635 530 56650 545
rect 56690 530 56705 545
rect 56745 530 56760 545
rect 56910 530 57210 545
rect 56435 520 56485 530
rect 55025 505 55085 520
rect 55125 505 55185 520
rect 55225 505 55285 520
rect 55325 505 55385 520
rect 55425 505 55485 520
rect 55525 505 55585 520
rect 54990 495 55085 505
rect 54990 475 54995 495
rect 55015 490 55085 495
rect 55525 495 55620 505
rect 55525 490 55595 495
rect 55015 475 55020 490
rect 54990 465 55020 475
rect 55590 475 55595 490
rect 55615 475 55620 495
rect 56435 500 56440 520
rect 56460 515 56485 520
rect 56745 520 56795 530
rect 56745 515 56770 520
rect 56460 500 56465 515
rect 56435 490 56465 500
rect 56765 500 56770 515
rect 56790 500 56795 520
rect 58220 505 58280 520
rect 58320 505 58380 520
rect 58420 505 58480 520
rect 58520 505 58580 520
rect 58620 505 58680 520
rect 58720 505 58780 520
rect 56765 490 56795 500
rect 58185 495 58280 505
rect 55590 465 55620 475
rect 58185 475 58190 495
rect 58210 490 58280 495
rect 58720 495 58815 505
rect 58720 490 58790 495
rect 58210 475 58215 490
rect 58185 465 58215 475
rect 58785 475 58790 490
rect 58810 475 58815 495
rect 58785 465 58815 475
<< polycont >>
rect 56095 4735 56115 4755
rect 56275 4735 56295 4755
rect 57035 4735 57055 4755
rect 57215 4735 57235 4755
rect 57505 4735 57525 4755
rect 57685 4735 57705 4755
rect 56565 4565 56585 4585
rect 56745 4565 56765 4585
rect 56160 4285 56180 4305
rect 56635 4285 56655 4305
rect 57145 4285 57165 4305
rect 57581 4275 57601 4295
rect 54935 3645 54955 3665
rect 55295 3645 55315 3665
rect 55655 3645 55675 3665
rect 56015 3645 56035 3665
rect 56375 3645 56395 3665
rect 56735 3645 56755 3665
rect 57045 3645 57065 3665
rect 57405 3645 57425 3665
rect 57765 3645 57785 3665
rect 58130 3645 58150 3665
rect 58490 3645 58510 3665
rect 58850 3645 58870 3665
rect 56375 3580 56395 3600
rect 57405 3580 57425 3600
rect 55295 3535 55315 3555
rect 58490 3535 58510 3555
rect 54965 3290 54985 3310
rect 55625 3290 55645 3310
rect 58160 3290 58180 3310
rect 58820 3290 58840 3310
rect 56285 3160 56305 3180
rect 56395 3160 56415 3180
rect 56835 3160 56855 3180
rect 57495 3160 57515 3180
rect 56045 2995 56065 3015
rect 56695 2995 56715 3015
rect 57085 2995 57105 3015
rect 57735 2995 57755 3015
rect 56040 2850 56060 2870
rect 56700 2850 56720 2870
rect 57080 2850 57100 2870
rect 57740 2850 57760 2870
rect 56100 2765 56120 2785
rect 56585 2765 56605 2785
rect 57195 2765 57215 2785
rect 55185 2620 55205 2640
rect 56725 2610 56745 2630
rect 56945 2610 56965 2630
rect 58600 2620 58620 2640
rect 55185 2560 55205 2580
rect 58600 2560 58620 2580
rect 56560 2490 56580 2510
rect 57220 2490 57240 2510
rect 54965 2395 54985 2415
rect 55625 2395 55645 2415
rect 58160 2395 58180 2415
rect 58820 2395 58840 2415
rect 56100 2245 56120 2265
rect 56640 2245 56660 2265
rect 57140 2245 57160 2265
rect 55460 2125 55480 2145
rect 55460 2030 55480 2050
rect 58325 2125 58345 2145
rect 58325 2030 58345 2050
rect 56040 1985 56060 2005
rect 56700 1985 56720 2005
rect 57080 1985 57100 2005
rect 57740 1985 57760 2005
rect 55460 1935 55480 1955
rect 58325 1935 58345 1955
rect 56045 1760 56065 1780
rect 56695 1760 56715 1780
rect 56855 1760 56875 1780
rect 56908 1760 56928 1780
rect 57085 1760 57105 1780
rect 57735 1760 57755 1780
rect 54965 1565 54985 1585
rect 55625 1565 55645 1585
rect 58160 1565 58180 1585
rect 58820 1565 58840 1585
rect 56040 1515 56060 1535
rect 56740 1515 56760 1535
rect 57040 1515 57060 1535
rect 57740 1515 57760 1535
rect 55395 1245 55415 1265
rect 57415 1240 57435 1260
rect 58440 1245 58460 1265
rect 56835 1185 56855 1205
rect 56230 865 56250 885
rect 57495 865 57515 885
rect 56605 720 56625 740
rect 57050 720 57070 740
rect 54995 475 55015 495
rect 55595 475 55615 495
rect 56440 500 56460 520
rect 56770 500 56790 520
rect 58190 475 58210 495
rect 58790 475 58810 495
<< xpolycontact >>
rect 54554 3065 54695 3285
rect 54554 2720 54695 2940
rect 59105 3065 59246 3285
rect 59105 2720 59246 2940
rect 54450 1979 54485 2199
rect 54450 1600 54485 1820
rect 54510 1979 54545 2199
rect 54510 1600 54545 1820
rect 54570 1979 54605 2199
rect 54570 1600 54605 1820
rect 54630 1979 54665 2199
rect 59135 1929 59170 2149
rect 54630 1600 54665 1820
rect 59135 1550 59170 1770
rect 59195 1929 59230 2149
rect 59195 1550 59230 1770
rect 59255 1929 59290 2149
rect 59255 1550 59290 1770
rect 59315 1929 59350 2149
rect 59315 1550 59350 1770
rect 54710 935 54745 1155
rect 54710 468 54745 688
rect 54770 935 54805 1155
rect 54770 468 54805 688
rect 58975 940 59010 1160
rect 58975 473 59010 693
rect 59035 940 59070 1160
rect 59035 473 59070 693
<< ppolyres >>
rect 54554 2940 54695 3065
rect 59105 2940 59246 3065
<< xpolyres >>
rect 54450 1820 54485 1979
rect 54510 1820 54545 1979
rect 54570 1820 54605 1979
rect 54630 1820 54665 1979
rect 59135 1770 59170 1929
rect 59195 1770 59230 1929
rect 59255 1770 59290 1929
rect 59315 1770 59350 1929
rect 54710 688 54745 935
rect 54770 688 54805 935
rect 58975 693 59010 940
rect 59035 693 59070 940
<< locali >>
rect 56085 4755 56125 4765
rect 56085 4735 56095 4755
rect 56115 4735 56125 4755
rect 56085 4725 56125 4735
rect 56265 4755 56305 4765
rect 56265 4735 56275 4755
rect 56295 4735 56305 4755
rect 56265 4725 56305 4735
rect 57025 4755 57065 4765
rect 57025 4735 57035 4755
rect 57055 4735 57065 4755
rect 57025 4725 57065 4735
rect 57205 4755 57245 4765
rect 57205 4735 57215 4755
rect 57235 4735 57245 4755
rect 57205 4725 57245 4735
rect 57495 4755 57535 4765
rect 57495 4735 57505 4755
rect 57525 4735 57535 4755
rect 57495 4725 57535 4735
rect 57675 4755 57715 4765
rect 57675 4735 57685 4755
rect 57705 4735 57715 4755
rect 57675 4725 57715 4735
rect 56050 4695 56120 4705
rect 56050 4375 56055 4695
rect 56075 4375 56095 4695
rect 56115 4375 56120 4695
rect 56050 4365 56120 4375
rect 56150 4695 56180 4705
rect 56150 4375 56155 4695
rect 56175 4375 56180 4695
rect 56150 4365 56180 4375
rect 56210 4695 56240 4705
rect 56210 4375 56215 4695
rect 56235 4375 56240 4695
rect 56210 4365 56240 4375
rect 56270 4695 56340 4705
rect 56270 4375 56275 4695
rect 56295 4375 56315 4695
rect 56335 4375 56340 4695
rect 56990 4695 57060 4705
rect 56555 4585 56595 4595
rect 56555 4565 56565 4585
rect 56585 4565 56595 4585
rect 56555 4555 56595 4565
rect 56735 4585 56775 4595
rect 56735 4565 56745 4585
rect 56765 4565 56775 4585
rect 56735 4555 56775 4565
rect 56270 4365 56340 4375
rect 56520 4525 56590 4535
rect 56520 4375 56525 4525
rect 56545 4375 56565 4525
rect 56585 4375 56590 4525
rect 56520 4365 56590 4375
rect 56620 4525 56650 4535
rect 56620 4375 56625 4525
rect 56645 4375 56650 4525
rect 56620 4365 56650 4375
rect 56680 4525 56710 4535
rect 56680 4375 56685 4525
rect 56705 4375 56710 4525
rect 56680 4365 56710 4375
rect 56740 4525 56810 4535
rect 56740 4375 56745 4525
rect 56765 4375 56785 4525
rect 56805 4375 56810 4525
rect 56740 4365 56810 4375
rect 56990 4375 56995 4695
rect 57015 4375 57035 4695
rect 57055 4375 57060 4695
rect 56990 4365 57060 4375
rect 57090 4695 57120 4705
rect 57090 4375 57095 4695
rect 57115 4375 57120 4695
rect 57090 4365 57120 4375
rect 57150 4695 57180 4705
rect 57150 4375 57155 4695
rect 57175 4375 57180 4695
rect 57150 4365 57180 4375
rect 57210 4695 57280 4705
rect 57210 4375 57215 4695
rect 57235 4375 57255 4695
rect 57275 4375 57280 4695
rect 57210 4365 57280 4375
rect 57460 4695 57530 4705
rect 57460 4375 57465 4695
rect 57485 4375 57505 4695
rect 57525 4375 57530 4695
rect 57460 4365 57530 4375
rect 57560 4695 57590 4705
rect 57560 4375 57565 4695
rect 57585 4375 57590 4695
rect 57560 4365 57590 4375
rect 57620 4695 57650 4705
rect 57620 4375 57625 4695
rect 57645 4375 57650 4695
rect 57620 4365 57650 4375
rect 57680 4695 57750 4705
rect 57680 4375 57685 4695
rect 57705 4375 57725 4695
rect 57745 4375 57750 4695
rect 57680 4365 57750 4375
rect 56150 4305 56190 4315
rect 56150 4285 56160 4305
rect 56180 4285 56190 4305
rect 56150 4275 56190 4285
rect 56630 4305 56660 4315
rect 56630 4285 56635 4305
rect 56655 4285 56660 4305
rect 56630 4275 56660 4285
rect 57140 4305 57170 4315
rect 57140 4285 57145 4305
rect 57165 4285 57170 4305
rect 57140 4275 57170 4285
rect 57576 4295 57606 4305
rect 57576 4275 57581 4295
rect 57601 4275 57606 4295
rect 57576 4265 57606 4275
rect 54890 4025 54960 4035
rect 54890 3705 54895 4025
rect 54915 3705 54935 4025
rect 54955 3705 54960 4025
rect 54890 3695 54960 3705
rect 54990 4025 55020 4035
rect 54990 3705 54995 4025
rect 55015 3705 55020 4025
rect 54990 3695 55020 3705
rect 55050 4025 55080 4035
rect 55050 3705 55055 4025
rect 55075 3705 55080 4025
rect 55050 3695 55080 3705
rect 55110 4025 55140 4035
rect 55110 3705 55115 4025
rect 55135 3705 55140 4025
rect 55110 3695 55140 3705
rect 55170 4025 55200 4035
rect 55170 3705 55175 4025
rect 55195 3705 55200 4025
rect 55170 3695 55200 3705
rect 55230 4025 55260 4035
rect 55230 3705 55235 4025
rect 55255 3705 55260 4025
rect 55230 3695 55260 3705
rect 55290 4025 55320 4035
rect 55290 3705 55295 4025
rect 55315 3705 55320 4025
rect 55290 3695 55320 3705
rect 55350 4025 55380 4035
rect 55350 3705 55355 4025
rect 55375 3705 55380 4025
rect 55350 3695 55380 3705
rect 55410 4025 55440 4035
rect 55410 3705 55415 4025
rect 55435 3705 55440 4025
rect 55410 3695 55440 3705
rect 55470 4025 55500 4035
rect 55470 3705 55475 4025
rect 55495 3705 55500 4025
rect 55470 3695 55500 3705
rect 55530 4025 55560 4035
rect 55530 3705 55535 4025
rect 55555 3705 55560 4025
rect 55530 3695 55560 3705
rect 55590 4025 55620 4035
rect 55590 3705 55595 4025
rect 55615 3705 55620 4025
rect 55590 3695 55620 3705
rect 55650 4025 55720 4035
rect 55650 3705 55655 4025
rect 55675 3705 55695 4025
rect 55715 3705 55720 4025
rect 55650 3695 55720 3705
rect 55970 4025 56040 4035
rect 55970 3705 55975 4025
rect 55995 3705 56015 4025
rect 56035 3705 56040 4025
rect 55970 3695 56040 3705
rect 56070 4025 56100 4035
rect 56070 3705 56075 4025
rect 56095 3705 56100 4025
rect 56070 3695 56100 3705
rect 56130 4025 56160 4035
rect 56130 3705 56135 4025
rect 56155 3705 56160 4025
rect 56130 3695 56160 3705
rect 56190 4025 56220 4035
rect 56190 3705 56195 4025
rect 56215 3705 56220 4025
rect 56190 3695 56220 3705
rect 56250 4025 56280 4035
rect 56250 3705 56255 4025
rect 56275 3705 56280 4025
rect 56250 3695 56280 3705
rect 56310 4025 56340 4035
rect 56310 3705 56315 4025
rect 56335 3705 56340 4025
rect 56310 3695 56340 3705
rect 56370 4025 56400 4035
rect 56370 3705 56375 4025
rect 56395 3705 56400 4025
rect 56370 3695 56400 3705
rect 56430 4025 56460 4035
rect 56430 3705 56435 4025
rect 56455 3705 56460 4025
rect 56430 3695 56460 3705
rect 56490 4025 56520 4035
rect 56490 3705 56495 4025
rect 56515 3705 56520 4025
rect 56490 3695 56520 3705
rect 56550 4025 56580 4035
rect 56550 3705 56555 4025
rect 56575 3705 56580 4025
rect 56550 3695 56580 3705
rect 56610 4025 56640 4035
rect 56610 3705 56615 4025
rect 56635 3705 56640 4025
rect 56610 3695 56640 3705
rect 56670 4025 56700 4035
rect 56670 3705 56675 4025
rect 56695 3705 56700 4025
rect 56670 3695 56700 3705
rect 56730 4025 56800 4035
rect 56730 3705 56735 4025
rect 56755 3705 56775 4025
rect 56795 3705 56800 4025
rect 56730 3695 56800 3705
rect 57000 4025 57070 4035
rect 57000 3705 57005 4025
rect 57025 3705 57045 4025
rect 57065 3705 57070 4025
rect 57000 3695 57070 3705
rect 57100 4025 57130 4035
rect 57100 3705 57105 4025
rect 57125 3705 57130 4025
rect 57100 3695 57130 3705
rect 57160 4025 57190 4035
rect 57160 3705 57165 4025
rect 57185 3705 57190 4025
rect 57160 3695 57190 3705
rect 57220 4025 57250 4035
rect 57220 3705 57225 4025
rect 57245 3705 57250 4025
rect 57220 3695 57250 3705
rect 57280 4025 57310 4035
rect 57280 3705 57285 4025
rect 57305 3705 57310 4025
rect 57280 3695 57310 3705
rect 57340 4025 57370 4035
rect 57340 3705 57345 4025
rect 57365 3705 57370 4025
rect 57340 3695 57370 3705
rect 57400 4025 57430 4035
rect 57400 3705 57405 4025
rect 57425 3705 57430 4025
rect 57400 3695 57430 3705
rect 57460 4025 57490 4035
rect 57460 3705 57465 4025
rect 57485 3705 57490 4025
rect 57460 3695 57490 3705
rect 57520 4025 57550 4035
rect 57520 3705 57525 4025
rect 57545 3705 57550 4025
rect 57520 3695 57550 3705
rect 57580 4025 57610 4035
rect 57580 3705 57585 4025
rect 57605 3705 57610 4025
rect 57580 3695 57610 3705
rect 57640 4025 57670 4035
rect 57640 3705 57645 4025
rect 57665 3705 57670 4025
rect 57640 3695 57670 3705
rect 57700 4025 57730 4035
rect 57700 3705 57705 4025
rect 57725 3705 57730 4025
rect 57700 3695 57730 3705
rect 57760 4025 57830 4035
rect 57760 3705 57765 4025
rect 57785 3705 57805 4025
rect 57825 3705 57830 4025
rect 57760 3695 57830 3705
rect 58085 4025 58155 4035
rect 58085 3705 58090 4025
rect 58110 3705 58130 4025
rect 58150 3705 58155 4025
rect 58085 3695 58155 3705
rect 58185 4025 58215 4035
rect 58185 3705 58190 4025
rect 58210 3705 58215 4025
rect 58185 3695 58215 3705
rect 58245 4025 58275 4035
rect 58245 3705 58250 4025
rect 58270 3705 58275 4025
rect 58245 3695 58275 3705
rect 58305 4025 58335 4035
rect 58305 3705 58310 4025
rect 58330 3705 58335 4025
rect 58305 3695 58335 3705
rect 58365 4025 58395 4035
rect 58365 3705 58370 4025
rect 58390 3705 58395 4025
rect 58365 3695 58395 3705
rect 58425 4025 58455 4035
rect 58425 3705 58430 4025
rect 58450 3705 58455 4025
rect 58425 3695 58455 3705
rect 58485 4025 58515 4035
rect 58485 3705 58490 4025
rect 58510 3705 58515 4025
rect 58485 3695 58515 3705
rect 58545 4025 58575 4035
rect 58545 3705 58550 4025
rect 58570 3705 58575 4025
rect 58545 3695 58575 3705
rect 58605 4025 58635 4035
rect 58605 3705 58610 4025
rect 58630 3705 58635 4025
rect 58605 3695 58635 3705
rect 58665 4025 58695 4035
rect 58665 3705 58670 4025
rect 58690 3705 58695 4025
rect 58665 3695 58695 3705
rect 58725 4025 58755 4035
rect 58725 3705 58730 4025
rect 58750 3705 58755 4025
rect 58725 3695 58755 3705
rect 58785 4025 58815 4035
rect 58785 3705 58790 4025
rect 58810 3705 58815 4025
rect 58785 3695 58815 3705
rect 58845 4025 58915 4035
rect 58845 3705 58850 4025
rect 58870 3705 58890 4025
rect 58910 3705 58915 4025
rect 58845 3695 58915 3705
rect 54930 3665 54960 3675
rect 54930 3645 54935 3665
rect 54955 3645 54960 3665
rect 54930 3635 54960 3645
rect 55290 3665 55320 3675
rect 55290 3645 55295 3665
rect 55315 3645 55320 3665
rect 55290 3635 55320 3645
rect 55650 3665 55680 3675
rect 55650 3645 55655 3665
rect 55675 3645 55680 3665
rect 55650 3635 55680 3645
rect 56010 3665 56040 3675
rect 56010 3645 56015 3665
rect 56035 3645 56040 3665
rect 56010 3635 56040 3645
rect 56370 3665 56400 3675
rect 56370 3645 56375 3665
rect 56395 3645 56400 3665
rect 56370 3635 56400 3645
rect 56730 3665 56760 3675
rect 56730 3645 56735 3665
rect 56755 3645 56760 3665
rect 56730 3635 56760 3645
rect 57040 3665 57070 3675
rect 57040 3645 57045 3665
rect 57065 3645 57070 3665
rect 57040 3635 57070 3645
rect 57400 3665 57430 3675
rect 57400 3645 57405 3665
rect 57425 3645 57430 3665
rect 57400 3635 57430 3645
rect 57760 3665 57790 3675
rect 57760 3645 57765 3665
rect 57785 3645 57790 3665
rect 57760 3635 57790 3645
rect 58125 3665 58155 3675
rect 58125 3645 58130 3665
rect 58150 3645 58155 3665
rect 58125 3635 58155 3645
rect 58485 3665 58515 3675
rect 58485 3645 58490 3665
rect 58510 3645 58515 3665
rect 58485 3635 58515 3645
rect 58845 3665 58875 3675
rect 58845 3645 58850 3665
rect 58870 3645 58875 3665
rect 58845 3635 58875 3645
rect 56365 3600 56405 3610
rect 56365 3580 56375 3600
rect 56395 3580 56405 3600
rect 56365 3570 56405 3580
rect 57395 3600 57435 3610
rect 57395 3580 57405 3600
rect 57425 3580 57435 3600
rect 57395 3570 57435 3580
rect 55285 3555 55325 3565
rect 55285 3535 55295 3555
rect 55315 3535 55325 3555
rect 55285 3525 55325 3535
rect 58480 3555 58520 3565
rect 58480 3535 58490 3555
rect 58510 3535 58520 3555
rect 58480 3525 58520 3535
rect 54554 3315 54695 3325
rect 54554 3295 54560 3315
rect 54580 3295 54615 3315
rect 54635 3295 54670 3315
rect 54690 3295 54695 3315
rect 54554 3285 54695 3295
rect 54960 3310 54990 3320
rect 54960 3290 54965 3310
rect 54985 3290 54990 3310
rect 54960 3280 54990 3290
rect 55620 3310 55650 3320
rect 55620 3290 55625 3310
rect 55645 3290 55650 3310
rect 55620 3280 55650 3290
rect 58155 3310 58185 3320
rect 58155 3290 58160 3310
rect 58180 3290 58185 3310
rect 58155 3280 58185 3290
rect 58815 3310 58845 3320
rect 58815 3290 58820 3310
rect 58840 3290 58845 3310
rect 58815 3280 58845 3290
rect 59105 3315 59246 3325
rect 59105 3295 59110 3315
rect 59130 3295 59165 3315
rect 59185 3295 59220 3315
rect 59240 3295 59246 3315
rect 59105 3285 59246 3295
rect 54920 3250 54990 3260
rect 54554 2710 54695 2720
rect 54554 2690 54560 2710
rect 54580 2690 54615 2710
rect 54635 2690 54670 2710
rect 54690 2690 54695 2710
rect 54554 2680 54695 2690
rect 54920 2680 54925 3250
rect 54945 2680 54965 3250
rect 54985 2680 54990 3250
rect 54920 2670 54990 2680
rect 55015 3250 55045 3260
rect 55015 2680 55020 3250
rect 55040 2680 55045 3250
rect 55015 2670 55045 2680
rect 55070 3250 55100 3260
rect 55070 2680 55075 3250
rect 55095 2680 55100 3250
rect 55070 2670 55100 2680
rect 55125 3250 55155 3260
rect 55125 2680 55130 3250
rect 55150 2680 55155 3250
rect 55125 2670 55155 2680
rect 55180 3250 55210 3260
rect 55180 2680 55185 3250
rect 55205 2680 55210 3250
rect 55180 2670 55210 2680
rect 55235 3250 55265 3260
rect 55235 2680 55240 3250
rect 55260 2680 55265 3250
rect 55235 2670 55265 2680
rect 55290 3250 55320 3260
rect 55290 2680 55295 3250
rect 55315 2680 55320 3250
rect 55290 2670 55320 2680
rect 55345 3250 55375 3260
rect 55345 2680 55350 3250
rect 55370 2680 55375 3250
rect 55345 2670 55375 2680
rect 55400 3250 55430 3260
rect 55400 2680 55405 3250
rect 55425 2680 55430 3250
rect 55400 2670 55430 2680
rect 55455 3250 55485 3260
rect 55455 2680 55460 3250
rect 55480 2680 55485 3250
rect 55455 2670 55485 2680
rect 55510 3250 55540 3260
rect 55510 2680 55515 3250
rect 55535 2680 55540 3250
rect 55510 2670 55540 2680
rect 55565 3250 55595 3260
rect 55565 2680 55570 3250
rect 55590 2680 55595 3250
rect 55565 2670 55595 2680
rect 55620 3250 55690 3260
rect 58115 3250 58185 3260
rect 55620 2680 55625 3250
rect 55645 2680 55665 3250
rect 55685 2680 55690 3250
rect 56240 3240 56310 3250
rect 56240 3220 56245 3240
rect 56265 3220 56285 3240
rect 56305 3220 56310 3240
rect 56240 3210 56310 3220
rect 56335 3240 56365 3250
rect 56335 3220 56340 3240
rect 56360 3220 56365 3240
rect 56335 3210 56365 3220
rect 56390 3240 56420 3250
rect 56390 3220 56395 3240
rect 56415 3220 56420 3240
rect 56390 3210 56420 3220
rect 56445 3240 56475 3250
rect 56445 3220 56450 3240
rect 56470 3220 56475 3240
rect 56445 3210 56475 3220
rect 56500 3240 56530 3250
rect 56500 3220 56505 3240
rect 56525 3220 56530 3240
rect 56500 3210 56530 3220
rect 56555 3240 56585 3250
rect 56555 3220 56560 3240
rect 56580 3220 56585 3240
rect 56555 3210 56585 3220
rect 56610 3240 56640 3250
rect 56610 3220 56615 3240
rect 56635 3220 56640 3240
rect 56610 3210 56640 3220
rect 56665 3240 56695 3250
rect 56665 3220 56670 3240
rect 56690 3220 56695 3240
rect 56665 3210 56695 3220
rect 56720 3240 56750 3250
rect 56720 3220 56725 3240
rect 56745 3220 56750 3240
rect 56720 3210 56750 3220
rect 56775 3240 56805 3250
rect 56775 3220 56780 3240
rect 56800 3220 56805 3240
rect 56775 3210 56805 3220
rect 56830 3240 56860 3250
rect 56830 3220 56835 3240
rect 56855 3220 56860 3240
rect 56830 3210 56860 3220
rect 56885 3240 56915 3250
rect 56885 3220 56890 3240
rect 56910 3220 56915 3240
rect 56885 3210 56915 3220
rect 56940 3240 56970 3250
rect 56940 3220 56945 3240
rect 56965 3220 56970 3240
rect 56940 3210 56970 3220
rect 56995 3240 57025 3250
rect 56995 3220 57000 3240
rect 57020 3220 57025 3240
rect 56995 3210 57025 3220
rect 57050 3240 57080 3250
rect 57050 3220 57055 3240
rect 57075 3220 57080 3240
rect 57050 3210 57080 3220
rect 57105 3240 57135 3250
rect 57105 3220 57110 3240
rect 57130 3220 57135 3240
rect 57105 3210 57135 3220
rect 57160 3240 57190 3250
rect 57160 3220 57165 3240
rect 57185 3220 57190 3240
rect 57160 3210 57190 3220
rect 57215 3240 57245 3250
rect 57215 3220 57220 3240
rect 57240 3220 57245 3240
rect 57215 3210 57245 3220
rect 57270 3240 57300 3250
rect 57270 3220 57275 3240
rect 57295 3220 57300 3240
rect 57270 3210 57300 3220
rect 57325 3240 57355 3250
rect 57325 3220 57330 3240
rect 57350 3220 57355 3240
rect 57325 3210 57355 3220
rect 57380 3240 57410 3250
rect 57380 3220 57385 3240
rect 57405 3220 57410 3240
rect 57380 3210 57410 3220
rect 57435 3240 57465 3250
rect 57435 3220 57440 3240
rect 57460 3220 57465 3240
rect 57435 3210 57465 3220
rect 57490 3240 57560 3250
rect 57490 3220 57495 3240
rect 57515 3220 57535 3240
rect 57555 3220 57560 3240
rect 57490 3210 57560 3220
rect 56280 3180 56310 3190
rect 56280 3160 56285 3180
rect 56305 3160 56310 3180
rect 56280 3150 56310 3160
rect 56390 3180 56420 3190
rect 56390 3160 56395 3180
rect 56415 3160 56420 3180
rect 56390 3150 56420 3160
rect 56830 3180 56860 3190
rect 56830 3160 56835 3180
rect 56855 3160 56860 3180
rect 56830 3150 56860 3160
rect 57490 3180 57520 3190
rect 57490 3160 57495 3180
rect 57515 3160 57520 3180
rect 57490 3150 57520 3160
rect 56040 3015 56070 3025
rect 56040 2995 56045 3015
rect 56065 2995 56070 3015
rect 56040 2985 56070 2995
rect 56690 3015 56720 3025
rect 56690 2995 56695 3015
rect 56715 2995 56720 3015
rect 56690 2985 56720 2995
rect 57080 3015 57110 3025
rect 57080 2995 57085 3015
rect 57105 2995 57110 3015
rect 57080 2985 57110 2995
rect 57730 3015 57760 3025
rect 57730 2995 57735 3015
rect 57755 2995 57760 3015
rect 57730 2985 57760 2995
rect 55995 2930 56065 2940
rect 55995 2910 56000 2930
rect 56020 2910 56040 2930
rect 56060 2910 56065 2930
rect 55995 2900 56065 2910
rect 56090 2930 56120 2940
rect 56090 2910 56095 2930
rect 56115 2910 56120 2930
rect 56090 2900 56120 2910
rect 56145 2930 56175 2940
rect 56145 2910 56150 2930
rect 56170 2910 56175 2930
rect 56145 2900 56175 2910
rect 56200 2930 56230 2940
rect 56200 2910 56205 2930
rect 56225 2910 56230 2930
rect 56200 2900 56230 2910
rect 56255 2930 56285 2940
rect 56255 2910 56260 2930
rect 56280 2910 56285 2930
rect 56255 2900 56285 2910
rect 56310 2930 56340 2940
rect 56310 2910 56315 2930
rect 56335 2910 56340 2930
rect 56310 2900 56340 2910
rect 56365 2930 56395 2940
rect 56365 2910 56370 2930
rect 56390 2910 56395 2930
rect 56365 2900 56395 2910
rect 56420 2930 56450 2940
rect 56420 2910 56425 2930
rect 56445 2910 56450 2930
rect 56420 2900 56450 2910
rect 56475 2930 56505 2940
rect 56475 2910 56480 2930
rect 56500 2910 56505 2930
rect 56475 2900 56505 2910
rect 56530 2930 56560 2940
rect 56530 2910 56535 2930
rect 56555 2910 56560 2930
rect 56530 2900 56560 2910
rect 56585 2930 56615 2940
rect 56585 2910 56590 2930
rect 56610 2910 56615 2930
rect 56585 2900 56615 2910
rect 56640 2930 56670 2940
rect 56640 2910 56645 2930
rect 56665 2910 56670 2930
rect 56640 2900 56670 2910
rect 56695 2930 56765 2940
rect 56695 2910 56700 2930
rect 56720 2910 56740 2930
rect 56760 2910 56765 2930
rect 56695 2900 56765 2910
rect 57035 2930 57105 2940
rect 57035 2910 57040 2930
rect 57060 2910 57080 2930
rect 57100 2910 57105 2930
rect 57035 2900 57105 2910
rect 57130 2930 57160 2940
rect 57130 2910 57135 2930
rect 57155 2910 57160 2930
rect 57130 2900 57160 2910
rect 57185 2930 57215 2940
rect 57185 2910 57190 2930
rect 57210 2910 57215 2930
rect 57185 2900 57215 2910
rect 57240 2930 57270 2940
rect 57240 2910 57245 2930
rect 57265 2910 57270 2930
rect 57240 2900 57270 2910
rect 57295 2930 57325 2940
rect 57295 2910 57300 2930
rect 57320 2910 57325 2930
rect 57295 2900 57325 2910
rect 57350 2930 57380 2940
rect 57350 2910 57355 2930
rect 57375 2910 57380 2930
rect 57350 2900 57380 2910
rect 57405 2930 57435 2940
rect 57405 2910 57410 2930
rect 57430 2910 57435 2930
rect 57405 2900 57435 2910
rect 57460 2930 57490 2940
rect 57460 2910 57465 2930
rect 57485 2910 57490 2930
rect 57460 2900 57490 2910
rect 57515 2930 57545 2940
rect 57515 2910 57520 2930
rect 57540 2910 57545 2930
rect 57515 2900 57545 2910
rect 57570 2930 57600 2940
rect 57570 2910 57575 2930
rect 57595 2910 57600 2930
rect 57570 2900 57600 2910
rect 57625 2930 57655 2940
rect 57625 2910 57630 2930
rect 57650 2910 57655 2930
rect 57625 2900 57655 2910
rect 57680 2930 57710 2940
rect 57680 2910 57685 2930
rect 57705 2910 57710 2930
rect 57680 2900 57710 2910
rect 57735 2930 57805 2940
rect 57735 2910 57740 2930
rect 57760 2910 57780 2930
rect 57800 2910 57805 2930
rect 57735 2900 57805 2910
rect 56035 2870 56065 2880
rect 56035 2850 56040 2870
rect 56060 2850 56065 2870
rect 56035 2840 56065 2850
rect 56695 2870 56725 2880
rect 56695 2850 56700 2870
rect 56720 2850 56725 2870
rect 56695 2840 56725 2850
rect 57075 2870 57105 2880
rect 57075 2850 57080 2870
rect 57100 2850 57105 2870
rect 57075 2840 57105 2850
rect 57735 2870 57765 2880
rect 57735 2850 57740 2870
rect 57760 2850 57765 2870
rect 57735 2840 57765 2850
rect 56095 2785 56125 2795
rect 56095 2765 56100 2785
rect 56120 2765 56125 2785
rect 56095 2755 56125 2765
rect 56580 2785 56610 2795
rect 56580 2765 56585 2785
rect 56605 2765 56610 2785
rect 56580 2755 56610 2765
rect 57190 2785 57220 2795
rect 57190 2765 57195 2785
rect 57215 2765 57220 2785
rect 57190 2755 57220 2765
rect 55620 2670 55690 2680
rect 58115 2680 58120 3250
rect 58140 2680 58160 3250
rect 58180 2680 58185 3250
rect 58115 2670 58185 2680
rect 58210 3250 58240 3260
rect 58210 2680 58215 3250
rect 58235 2680 58240 3250
rect 58210 2670 58240 2680
rect 58265 3250 58295 3260
rect 58265 2680 58270 3250
rect 58290 2680 58295 3250
rect 58265 2670 58295 2680
rect 58320 3250 58350 3260
rect 58320 2680 58325 3250
rect 58345 2680 58350 3250
rect 58320 2670 58350 2680
rect 58375 3250 58405 3260
rect 58375 2680 58380 3250
rect 58400 2680 58405 3250
rect 58375 2670 58405 2680
rect 58430 3250 58460 3260
rect 58430 2680 58435 3250
rect 58455 2680 58460 3250
rect 58430 2670 58460 2680
rect 58485 3250 58515 3260
rect 58485 2680 58490 3250
rect 58510 2680 58515 3250
rect 58485 2670 58515 2680
rect 58540 3250 58570 3260
rect 58540 2680 58545 3250
rect 58565 2680 58570 3250
rect 58540 2670 58570 2680
rect 58595 3250 58625 3260
rect 58595 2680 58600 3250
rect 58620 2680 58625 3250
rect 58595 2670 58625 2680
rect 58650 3250 58680 3260
rect 58650 2680 58655 3250
rect 58675 2680 58680 3250
rect 58650 2670 58680 2680
rect 58705 3250 58735 3260
rect 58705 2680 58710 3250
rect 58730 2680 58735 3250
rect 58705 2670 58735 2680
rect 58760 3250 58790 3260
rect 58760 2680 58765 3250
rect 58785 2680 58790 3250
rect 58760 2670 58790 2680
rect 58815 3250 58885 3260
rect 58815 2680 58820 3250
rect 58840 2680 58860 3250
rect 58880 2680 58885 3250
rect 59105 2710 59246 2720
rect 59105 2690 59110 2710
rect 59130 2690 59165 2710
rect 59185 2690 59220 2710
rect 59240 2690 59246 2710
rect 59105 2680 59246 2690
rect 58815 2670 58885 2680
rect 55180 2640 55210 2650
rect 58595 2640 58625 2650
rect 55180 2620 55185 2640
rect 55205 2620 55210 2640
rect 55180 2610 55210 2620
rect 56715 2630 56755 2640
rect 56715 2610 56725 2630
rect 56745 2610 56755 2630
rect 56715 2600 56755 2610
rect 56935 2630 56975 2640
rect 56935 2610 56945 2630
rect 56965 2610 56975 2630
rect 58595 2620 58600 2640
rect 58620 2620 58625 2640
rect 58595 2610 58625 2620
rect 56935 2600 56975 2610
rect 55175 2580 55215 2585
rect 58590 2580 58630 2585
rect 55175 2560 55185 2580
rect 55205 2560 55215 2580
rect 55175 2555 55215 2560
rect 56515 2570 56585 2580
rect 56515 2550 56520 2570
rect 56540 2550 56560 2570
rect 56580 2550 56585 2570
rect 56515 2540 56585 2550
rect 56610 2570 56640 2580
rect 56610 2550 56615 2570
rect 56635 2550 56640 2570
rect 56610 2540 56640 2550
rect 56665 2570 56695 2580
rect 56665 2550 56670 2570
rect 56690 2550 56695 2570
rect 56665 2540 56695 2550
rect 56720 2570 56750 2580
rect 56720 2550 56725 2570
rect 56745 2550 56750 2570
rect 56720 2540 56750 2550
rect 56775 2570 56805 2580
rect 56775 2550 56780 2570
rect 56800 2550 56805 2570
rect 56775 2540 56805 2550
rect 56830 2570 56860 2580
rect 56830 2550 56835 2570
rect 56855 2550 56860 2570
rect 56830 2540 56860 2550
rect 56885 2570 56915 2580
rect 56885 2550 56890 2570
rect 56910 2550 56915 2570
rect 56885 2540 56915 2550
rect 56940 2570 56970 2580
rect 56940 2550 56945 2570
rect 56965 2550 56970 2570
rect 56940 2540 56970 2550
rect 56995 2570 57025 2580
rect 56995 2550 57000 2570
rect 57020 2550 57025 2570
rect 56995 2540 57025 2550
rect 57050 2570 57080 2580
rect 57050 2550 57055 2570
rect 57075 2550 57080 2570
rect 57050 2540 57080 2550
rect 57105 2570 57135 2580
rect 57105 2550 57110 2570
rect 57130 2550 57135 2570
rect 57105 2540 57135 2550
rect 57160 2570 57190 2580
rect 57160 2550 57165 2570
rect 57185 2550 57190 2570
rect 57160 2540 57190 2550
rect 57215 2570 57285 2580
rect 57215 2550 57220 2570
rect 57240 2550 57260 2570
rect 57280 2550 57285 2570
rect 58590 2560 58600 2580
rect 58620 2560 58630 2580
rect 58590 2555 58630 2560
rect 57215 2540 57285 2550
rect 56550 2510 56590 2520
rect 56550 2490 56560 2510
rect 56580 2490 56590 2510
rect 56550 2480 56590 2490
rect 57210 2510 57250 2520
rect 57210 2490 57220 2510
rect 57240 2490 57250 2510
rect 57210 2480 57250 2490
rect 54960 2415 54990 2425
rect 54960 2395 54965 2415
rect 54985 2395 54990 2415
rect 54960 2385 54990 2395
rect 55620 2415 55650 2425
rect 55620 2395 55625 2415
rect 55645 2395 55650 2415
rect 55620 2385 55650 2395
rect 58155 2415 58185 2425
rect 58155 2395 58160 2415
rect 58180 2395 58185 2415
rect 58155 2385 58185 2395
rect 58815 2415 58845 2425
rect 58815 2395 58820 2415
rect 58840 2395 58845 2415
rect 58815 2385 58845 2395
rect 54920 2355 54990 2365
rect 54450 2216 54665 2236
rect 54450 2199 54485 2216
rect 54630 2199 54665 2216
rect 54545 2149 54570 2199
rect 54920 2185 54925 2355
rect 54945 2185 54965 2355
rect 54985 2185 54990 2355
rect 54920 2175 54990 2185
rect 55015 2355 55045 2365
rect 55015 2185 55020 2355
rect 55040 2185 55045 2355
rect 55015 2175 55045 2185
rect 55070 2355 55100 2365
rect 55070 2185 55075 2355
rect 55095 2185 55100 2355
rect 55070 2175 55100 2185
rect 55125 2355 55155 2365
rect 55125 2185 55130 2355
rect 55150 2185 55155 2355
rect 55125 2175 55155 2185
rect 55180 2355 55210 2365
rect 55180 2185 55185 2355
rect 55205 2185 55210 2355
rect 55180 2175 55210 2185
rect 55235 2355 55265 2365
rect 55235 2185 55240 2355
rect 55260 2185 55265 2355
rect 55235 2175 55265 2185
rect 55290 2355 55320 2365
rect 55290 2185 55295 2355
rect 55315 2185 55320 2355
rect 55290 2175 55320 2185
rect 55345 2355 55375 2365
rect 55345 2185 55350 2355
rect 55370 2185 55375 2355
rect 55345 2175 55375 2185
rect 55400 2355 55430 2365
rect 55400 2185 55405 2355
rect 55425 2185 55430 2355
rect 55400 2175 55430 2185
rect 55455 2355 55485 2365
rect 55455 2185 55460 2355
rect 55480 2185 55485 2355
rect 55455 2175 55485 2185
rect 55510 2355 55540 2365
rect 55510 2185 55515 2355
rect 55535 2185 55540 2355
rect 55510 2175 55540 2185
rect 55565 2355 55595 2365
rect 55565 2185 55570 2355
rect 55590 2185 55595 2355
rect 55565 2175 55595 2185
rect 55620 2355 55690 2365
rect 55620 2185 55625 2355
rect 55645 2185 55665 2355
rect 55685 2185 55690 2355
rect 58115 2355 58185 2365
rect 56095 2265 56125 2275
rect 56095 2245 56100 2265
rect 56120 2245 56125 2265
rect 56095 2235 56125 2245
rect 56635 2265 56665 2275
rect 56635 2245 56640 2265
rect 56660 2245 56665 2265
rect 56635 2235 56665 2245
rect 57135 2265 57165 2275
rect 57135 2245 57140 2265
rect 57160 2245 57165 2265
rect 57135 2235 57165 2245
rect 55620 2175 55690 2185
rect 58115 2185 58120 2355
rect 58140 2185 58160 2355
rect 58180 2185 58185 2355
rect 58115 2175 58185 2185
rect 58210 2355 58240 2365
rect 58210 2185 58215 2355
rect 58235 2185 58240 2355
rect 58210 2175 58240 2185
rect 58265 2355 58295 2365
rect 58265 2185 58270 2355
rect 58290 2185 58295 2355
rect 58265 2175 58295 2185
rect 58320 2355 58350 2365
rect 58320 2185 58325 2355
rect 58345 2185 58350 2355
rect 58320 2175 58350 2185
rect 58375 2355 58405 2365
rect 58375 2185 58380 2355
rect 58400 2185 58405 2355
rect 58375 2175 58405 2185
rect 58430 2355 58460 2365
rect 58430 2185 58435 2355
rect 58455 2185 58460 2355
rect 58430 2175 58460 2185
rect 58485 2355 58515 2365
rect 58485 2185 58490 2355
rect 58510 2185 58515 2355
rect 58485 2175 58515 2185
rect 58540 2355 58570 2365
rect 58540 2185 58545 2355
rect 58565 2185 58570 2355
rect 58540 2175 58570 2185
rect 58595 2355 58625 2365
rect 58595 2185 58600 2355
rect 58620 2185 58625 2355
rect 58595 2175 58625 2185
rect 58650 2355 58680 2365
rect 58650 2185 58655 2355
rect 58675 2185 58680 2355
rect 58650 2175 58680 2185
rect 58705 2355 58735 2365
rect 58705 2185 58710 2355
rect 58730 2185 58735 2355
rect 58705 2175 58735 2185
rect 58760 2355 58790 2365
rect 58760 2185 58765 2355
rect 58785 2185 58790 2355
rect 58760 2175 58790 2185
rect 58815 2355 58885 2365
rect 58815 2185 58820 2355
rect 58840 2185 58860 2355
rect 58880 2185 58885 2355
rect 58815 2175 58885 2185
rect 55995 2165 56065 2175
rect 55065 2145 55105 2155
rect 55065 2125 55075 2145
rect 55095 2125 55105 2145
rect 55065 2115 55105 2125
rect 55175 2145 55215 2155
rect 55175 2125 55185 2145
rect 55205 2125 55215 2145
rect 55175 2115 55215 2125
rect 55285 2145 55325 2155
rect 55285 2125 55295 2145
rect 55315 2125 55325 2145
rect 55285 2115 55325 2125
rect 55395 2145 55435 2155
rect 55395 2125 55405 2145
rect 55425 2125 55435 2145
rect 55395 2115 55435 2125
rect 55455 2145 55485 2155
rect 55455 2125 55460 2145
rect 55480 2125 55485 2145
rect 55455 2115 55485 2125
rect 55505 2145 55545 2155
rect 55505 2125 55515 2145
rect 55535 2125 55545 2145
rect 55505 2115 55545 2125
rect 55450 2050 55490 2060
rect 55450 2030 55460 2050
rect 55480 2030 55490 2050
rect 55995 2045 56000 2165
rect 56020 2045 56040 2165
rect 56060 2045 56065 2165
rect 55995 2035 56065 2045
rect 56090 2165 56120 2175
rect 56090 2045 56095 2165
rect 56115 2045 56120 2165
rect 56090 2035 56120 2045
rect 56145 2165 56175 2175
rect 56145 2045 56150 2165
rect 56170 2045 56175 2165
rect 56145 2035 56175 2045
rect 56200 2165 56230 2175
rect 56200 2045 56205 2165
rect 56225 2045 56230 2165
rect 56200 2035 56230 2045
rect 56255 2165 56285 2175
rect 56255 2045 56260 2165
rect 56280 2045 56285 2165
rect 56255 2035 56285 2045
rect 56310 2165 56340 2175
rect 56310 2045 56315 2165
rect 56335 2045 56340 2165
rect 56310 2035 56340 2045
rect 56365 2165 56395 2175
rect 56365 2045 56370 2165
rect 56390 2045 56395 2165
rect 56365 2035 56395 2045
rect 56420 2165 56450 2175
rect 56420 2045 56425 2165
rect 56445 2045 56450 2165
rect 56420 2035 56450 2045
rect 56475 2165 56505 2175
rect 56475 2045 56480 2165
rect 56500 2045 56505 2165
rect 56475 2035 56505 2045
rect 56530 2165 56560 2175
rect 56530 2045 56535 2165
rect 56555 2045 56560 2165
rect 56530 2035 56560 2045
rect 56585 2165 56615 2175
rect 56585 2045 56590 2165
rect 56610 2045 56615 2165
rect 56585 2035 56615 2045
rect 56640 2165 56670 2175
rect 56640 2045 56645 2165
rect 56665 2045 56670 2165
rect 56640 2035 56670 2045
rect 56695 2165 56765 2175
rect 56695 2045 56700 2165
rect 56720 2045 56740 2165
rect 56760 2045 56765 2165
rect 56695 2035 56765 2045
rect 57035 2165 57105 2175
rect 57035 2045 57040 2165
rect 57060 2045 57080 2165
rect 57100 2045 57105 2165
rect 57035 2035 57105 2045
rect 57130 2165 57160 2175
rect 57130 2045 57135 2165
rect 57155 2045 57160 2165
rect 57130 2035 57160 2045
rect 57185 2165 57215 2175
rect 57185 2045 57190 2165
rect 57210 2045 57215 2165
rect 57185 2035 57215 2045
rect 57240 2165 57270 2175
rect 57240 2045 57245 2165
rect 57265 2045 57270 2165
rect 57240 2035 57270 2045
rect 57295 2165 57325 2175
rect 57295 2045 57300 2165
rect 57320 2045 57325 2165
rect 57295 2035 57325 2045
rect 57350 2165 57380 2175
rect 57350 2045 57355 2165
rect 57375 2045 57380 2165
rect 57350 2035 57380 2045
rect 57405 2165 57435 2175
rect 57405 2045 57410 2165
rect 57430 2045 57435 2165
rect 57405 2035 57435 2045
rect 57460 2165 57490 2175
rect 57460 2045 57465 2165
rect 57485 2045 57490 2165
rect 57460 2035 57490 2045
rect 57515 2165 57545 2175
rect 57515 2045 57520 2165
rect 57540 2045 57545 2165
rect 57515 2035 57545 2045
rect 57570 2165 57600 2175
rect 57570 2045 57575 2165
rect 57595 2045 57600 2165
rect 57570 2035 57600 2045
rect 57625 2165 57655 2175
rect 57625 2045 57630 2165
rect 57650 2045 57655 2165
rect 57625 2035 57655 2045
rect 57680 2165 57710 2175
rect 57680 2045 57685 2165
rect 57705 2045 57710 2165
rect 57680 2035 57710 2045
rect 57735 2165 57805 2175
rect 57735 2045 57740 2165
rect 57760 2045 57780 2165
rect 57800 2045 57805 2165
rect 59135 2166 59350 2186
rect 58260 2145 58300 2155
rect 58260 2125 58270 2145
rect 58290 2125 58300 2145
rect 58260 2115 58300 2125
rect 58320 2145 58350 2155
rect 58320 2125 58325 2145
rect 58345 2125 58350 2145
rect 58320 2115 58350 2125
rect 58370 2145 58410 2155
rect 58370 2125 58380 2145
rect 58400 2125 58410 2145
rect 58370 2115 58410 2125
rect 58480 2145 58520 2155
rect 58480 2125 58490 2145
rect 58510 2125 58520 2145
rect 58480 2115 58520 2125
rect 58590 2145 58630 2155
rect 58590 2125 58600 2145
rect 58620 2125 58630 2145
rect 58590 2115 58630 2125
rect 58700 2145 58740 2155
rect 58700 2125 58710 2145
rect 58730 2125 58740 2145
rect 58700 2115 58740 2125
rect 59135 2149 59170 2166
rect 59315 2149 59350 2166
rect 57735 2035 57805 2045
rect 58315 2050 58355 2060
rect 55450 2020 55490 2030
rect 56035 2005 56065 2035
rect 56035 1985 56040 2005
rect 56060 1985 56065 2005
rect 56035 1975 56065 1985
rect 56695 2005 56725 2015
rect 56695 1985 56700 2005
rect 56720 1985 56725 2005
rect 56695 1975 56725 1985
rect 57075 2005 57105 2015
rect 57075 1985 57080 2005
rect 57100 1985 57105 2005
rect 57075 1975 57105 1985
rect 57735 2005 57765 2035
rect 58315 2030 58325 2050
rect 58345 2030 58355 2050
rect 58315 2020 58355 2030
rect 57735 1985 57740 2005
rect 57760 1985 57765 2005
rect 57735 1975 57765 1985
rect 55455 1955 55485 1965
rect 55455 1935 55460 1955
rect 55480 1935 55485 1955
rect 55455 1925 55485 1935
rect 58320 1955 58350 1965
rect 58320 1935 58325 1955
rect 58345 1935 58350 1955
rect 58320 1925 58350 1935
rect 59230 2099 59255 2149
rect 54920 1895 54990 1905
rect 54450 1590 54485 1600
rect 54450 1565 54455 1590
rect 54480 1565 54485 1590
rect 54450 1555 54485 1565
rect 54510 1590 54545 1600
rect 54510 1565 54515 1590
rect 54540 1565 54545 1590
rect 54510 1555 54545 1565
rect 54570 1590 54605 1600
rect 54570 1565 54575 1590
rect 54600 1565 54605 1590
rect 54570 1555 54605 1565
rect 54920 1625 54925 1895
rect 54945 1625 54965 1895
rect 54985 1625 54990 1895
rect 54920 1615 54990 1625
rect 55015 1895 55045 1905
rect 55015 1625 55020 1895
rect 55040 1625 55045 1895
rect 55015 1615 55045 1625
rect 55070 1895 55100 1905
rect 55070 1625 55075 1895
rect 55095 1625 55100 1895
rect 55070 1615 55100 1625
rect 55125 1895 55155 1905
rect 55125 1625 55130 1895
rect 55150 1625 55155 1895
rect 55125 1615 55155 1625
rect 55180 1895 55210 1905
rect 55180 1625 55185 1895
rect 55205 1625 55210 1895
rect 55180 1615 55210 1625
rect 55235 1895 55265 1905
rect 55235 1625 55240 1895
rect 55260 1625 55265 1895
rect 55235 1615 55265 1625
rect 55290 1895 55320 1905
rect 55290 1625 55295 1895
rect 55315 1625 55320 1895
rect 55290 1615 55320 1625
rect 55345 1895 55375 1905
rect 55345 1625 55350 1895
rect 55370 1625 55375 1895
rect 55345 1615 55375 1625
rect 55400 1895 55430 1905
rect 55400 1625 55405 1895
rect 55425 1625 55430 1895
rect 55400 1615 55430 1625
rect 55455 1895 55485 1905
rect 55455 1625 55460 1895
rect 55480 1625 55485 1895
rect 55455 1615 55485 1625
rect 55510 1895 55540 1905
rect 55510 1625 55515 1895
rect 55535 1625 55540 1895
rect 55510 1615 55540 1625
rect 55565 1895 55595 1905
rect 55565 1625 55570 1895
rect 55590 1625 55595 1895
rect 55565 1615 55595 1625
rect 55620 1895 55690 1905
rect 55620 1625 55625 1895
rect 55645 1625 55665 1895
rect 55685 1625 55690 1895
rect 58115 1895 58185 1905
rect 56040 1780 56070 1790
rect 56040 1760 56045 1780
rect 56065 1760 56070 1780
rect 56040 1750 56070 1760
rect 56690 1780 56720 1790
rect 56690 1760 56695 1780
rect 56715 1760 56720 1780
rect 56690 1750 56720 1760
rect 56850 1780 56880 1790
rect 56850 1760 56855 1780
rect 56875 1760 56880 1780
rect 56850 1750 56880 1760
rect 56903 1780 56933 1790
rect 56903 1760 56908 1780
rect 56928 1760 56933 1780
rect 56903 1750 56933 1760
rect 57080 1780 57110 1790
rect 57080 1760 57085 1780
rect 57105 1760 57110 1780
rect 57080 1750 57110 1760
rect 57730 1780 57760 1790
rect 57730 1760 57735 1780
rect 57755 1760 57760 1780
rect 57730 1750 57760 1760
rect 55620 1615 55690 1625
rect 55995 1695 56065 1705
rect 54630 1590 54665 1600
rect 54630 1565 54635 1590
rect 54660 1565 54665 1590
rect 54630 1555 54665 1565
rect 54960 1585 54990 1595
rect 54960 1565 54965 1585
rect 54985 1565 54990 1585
rect 54960 1555 54990 1565
rect 55620 1585 55650 1595
rect 55620 1565 55625 1585
rect 55645 1565 55650 1585
rect 55995 1575 56000 1695
rect 56020 1575 56040 1695
rect 56060 1575 56065 1695
rect 55995 1565 56065 1575
rect 56090 1695 56120 1705
rect 56090 1575 56095 1695
rect 56115 1575 56120 1695
rect 56090 1565 56120 1575
rect 56145 1695 56175 1705
rect 56145 1575 56150 1695
rect 56170 1575 56175 1695
rect 56145 1565 56175 1575
rect 56200 1695 56230 1705
rect 56200 1575 56205 1695
rect 56225 1575 56230 1695
rect 56200 1565 56230 1575
rect 56255 1695 56285 1705
rect 56255 1575 56260 1695
rect 56280 1575 56285 1695
rect 56255 1565 56285 1575
rect 56310 1695 56340 1705
rect 56310 1575 56315 1695
rect 56335 1575 56340 1695
rect 56310 1565 56340 1575
rect 56365 1695 56395 1705
rect 56365 1575 56370 1695
rect 56390 1575 56395 1695
rect 56365 1565 56395 1575
rect 56420 1695 56450 1705
rect 56420 1575 56425 1695
rect 56445 1575 56450 1695
rect 56420 1565 56450 1575
rect 56475 1695 56505 1705
rect 56475 1575 56480 1695
rect 56500 1575 56505 1695
rect 56475 1565 56505 1575
rect 56530 1695 56560 1705
rect 56530 1575 56535 1695
rect 56555 1575 56560 1695
rect 56530 1565 56560 1575
rect 56585 1695 56615 1705
rect 56585 1575 56590 1695
rect 56610 1575 56615 1695
rect 56585 1565 56615 1575
rect 56640 1695 56670 1705
rect 56640 1575 56645 1695
rect 56665 1575 56670 1695
rect 56640 1565 56670 1575
rect 56695 1695 56805 1705
rect 56695 1575 56700 1695
rect 56720 1575 56740 1695
rect 56760 1575 56780 1695
rect 56800 1575 56805 1695
rect 56695 1565 56805 1575
rect 56830 1695 56860 1705
rect 56830 1575 56835 1695
rect 56855 1575 56860 1695
rect 56830 1565 56860 1575
rect 56885 1695 56915 1705
rect 56885 1575 56890 1695
rect 56910 1575 56915 1695
rect 56885 1565 56915 1575
rect 56940 1695 56970 1705
rect 56940 1575 56945 1695
rect 56965 1575 56970 1695
rect 56940 1565 56970 1575
rect 56995 1695 57105 1705
rect 56995 1575 57000 1695
rect 57020 1575 57040 1695
rect 57060 1575 57080 1695
rect 57100 1575 57105 1695
rect 56995 1565 57105 1575
rect 57130 1695 57160 1705
rect 57130 1575 57135 1695
rect 57155 1575 57160 1695
rect 57130 1565 57160 1575
rect 57185 1695 57215 1705
rect 57185 1575 57190 1695
rect 57210 1575 57215 1695
rect 57185 1565 57215 1575
rect 57240 1695 57270 1705
rect 57240 1575 57245 1695
rect 57265 1575 57270 1695
rect 57240 1565 57270 1575
rect 57295 1695 57325 1705
rect 57295 1575 57300 1695
rect 57320 1575 57325 1695
rect 57295 1565 57325 1575
rect 57350 1695 57380 1705
rect 57350 1575 57355 1695
rect 57375 1575 57380 1695
rect 57350 1565 57380 1575
rect 57405 1695 57435 1705
rect 57405 1575 57410 1695
rect 57430 1575 57435 1695
rect 57405 1565 57435 1575
rect 57460 1695 57490 1705
rect 57460 1575 57465 1695
rect 57485 1575 57490 1695
rect 57460 1565 57490 1575
rect 57515 1695 57545 1705
rect 57515 1575 57520 1695
rect 57540 1575 57545 1695
rect 57515 1565 57545 1575
rect 57570 1695 57600 1705
rect 57570 1575 57575 1695
rect 57595 1575 57600 1695
rect 57570 1565 57600 1575
rect 57625 1695 57655 1705
rect 57625 1575 57630 1695
rect 57650 1575 57655 1695
rect 57625 1565 57655 1575
rect 57680 1695 57710 1705
rect 57680 1575 57685 1695
rect 57705 1575 57710 1695
rect 57680 1565 57710 1575
rect 57735 1695 57805 1705
rect 57735 1575 57740 1695
rect 57760 1575 57780 1695
rect 57800 1575 57805 1695
rect 58115 1625 58120 1895
rect 58140 1625 58160 1895
rect 58180 1625 58185 1895
rect 58115 1615 58185 1625
rect 58210 1895 58240 1905
rect 58210 1625 58215 1895
rect 58235 1625 58240 1895
rect 58210 1615 58240 1625
rect 58265 1895 58295 1905
rect 58265 1625 58270 1895
rect 58290 1625 58295 1895
rect 58265 1615 58295 1625
rect 58320 1895 58350 1905
rect 58320 1625 58325 1895
rect 58345 1625 58350 1895
rect 58320 1615 58350 1625
rect 58375 1895 58405 1905
rect 58375 1625 58380 1895
rect 58400 1625 58405 1895
rect 58375 1615 58405 1625
rect 58430 1895 58460 1905
rect 58430 1625 58435 1895
rect 58455 1625 58460 1895
rect 58430 1615 58460 1625
rect 58485 1895 58515 1905
rect 58485 1625 58490 1895
rect 58510 1625 58515 1895
rect 58485 1615 58515 1625
rect 58540 1895 58570 1905
rect 58540 1625 58545 1895
rect 58565 1625 58570 1895
rect 58540 1615 58570 1625
rect 58595 1895 58625 1905
rect 58595 1625 58600 1895
rect 58620 1625 58625 1895
rect 58595 1615 58625 1625
rect 58650 1895 58680 1905
rect 58650 1625 58655 1895
rect 58675 1625 58680 1895
rect 58650 1615 58680 1625
rect 58705 1895 58735 1905
rect 58705 1625 58710 1895
rect 58730 1625 58735 1895
rect 58705 1615 58735 1625
rect 58760 1895 58790 1905
rect 58760 1625 58765 1895
rect 58785 1625 58790 1895
rect 58760 1615 58790 1625
rect 58815 1895 58885 1905
rect 58815 1625 58820 1895
rect 58840 1625 58860 1895
rect 58880 1625 58885 1895
rect 58815 1615 58885 1625
rect 57735 1565 57805 1575
rect 58155 1585 58185 1595
rect 58155 1565 58160 1585
rect 58180 1565 58185 1585
rect 55620 1555 55650 1565
rect 56040 1545 56065 1565
rect 56035 1535 56065 1545
rect 56035 1515 56040 1535
rect 56060 1515 56065 1535
rect 56035 1505 56065 1515
rect 56735 1535 56765 1545
rect 56735 1515 56740 1535
rect 56760 1515 56765 1535
rect 56735 1505 56765 1515
rect 57035 1535 57065 1545
rect 57035 1515 57040 1535
rect 57060 1515 57065 1535
rect 57035 1505 57065 1515
rect 57735 1535 57765 1565
rect 58155 1555 58185 1565
rect 58815 1585 58845 1595
rect 58815 1565 58820 1585
rect 58840 1565 58845 1585
rect 58815 1555 58845 1565
rect 57735 1515 57740 1535
rect 57760 1515 57765 1535
rect 57735 1505 57765 1515
rect 59135 1540 59170 1550
rect 59135 1515 59140 1540
rect 59165 1515 59170 1540
rect 59135 1505 59170 1515
rect 59195 1540 59230 1550
rect 59195 1515 59200 1540
rect 59225 1515 59230 1540
rect 59195 1505 59230 1515
rect 59255 1540 59290 1550
rect 59255 1515 59260 1540
rect 59285 1515 59290 1540
rect 59255 1505 59290 1515
rect 59315 1540 59350 1550
rect 59315 1515 59320 1540
rect 59345 1515 59350 1540
rect 59315 1505 59350 1515
rect 55385 1265 55425 1275
rect 55385 1245 55395 1265
rect 55415 1245 55425 1265
rect 55385 1235 55425 1245
rect 57405 1260 57445 1270
rect 57405 1240 57415 1260
rect 57435 1240 57445 1260
rect 57405 1230 57445 1240
rect 58435 1265 58465 1275
rect 58435 1245 58440 1265
rect 58460 1245 58465 1265
rect 58435 1235 58465 1245
rect 54950 1205 55020 1215
rect 54710 1190 54745 1200
rect 54710 1165 54715 1190
rect 54740 1165 54745 1190
rect 54710 1155 54745 1165
rect 54770 1190 54805 1200
rect 54770 1165 54775 1190
rect 54800 1165 54805 1190
rect 54770 1155 54805 1165
rect 54745 468 54770 518
rect 54950 535 54955 1205
rect 54975 535 54995 1205
rect 55015 535 55020 1205
rect 54950 525 55020 535
rect 55090 1205 55120 1215
rect 55090 535 55095 1205
rect 55115 535 55120 1205
rect 55090 525 55120 535
rect 55190 1205 55220 1215
rect 55190 535 55195 1205
rect 55215 535 55220 1205
rect 55190 525 55220 535
rect 55290 1205 55320 1215
rect 55290 535 55295 1205
rect 55315 535 55320 1205
rect 55290 525 55320 535
rect 55390 1205 55420 1215
rect 55390 535 55395 1205
rect 55415 535 55420 1205
rect 55390 525 55420 535
rect 55490 1205 55520 1215
rect 55490 535 55495 1205
rect 55515 535 55520 1205
rect 55490 525 55520 535
rect 55590 1205 55660 1215
rect 55590 535 55595 1205
rect 55615 535 55635 1205
rect 55655 535 55660 1205
rect 56830 1205 56860 1215
rect 56830 1185 56835 1205
rect 56855 1185 56860 1205
rect 56830 1175 56860 1185
rect 58145 1205 58215 1215
rect 56185 1145 56255 1155
rect 56185 925 56190 1145
rect 56210 925 56230 1145
rect 56250 925 56255 1145
rect 56185 915 56255 925
rect 56280 1145 56310 1155
rect 56280 925 56285 1145
rect 56305 925 56310 1145
rect 56280 915 56310 925
rect 56335 1145 56365 1155
rect 56335 925 56340 1145
rect 56360 925 56365 1145
rect 56335 915 56365 925
rect 56390 1145 56420 1155
rect 56390 925 56395 1145
rect 56415 925 56420 1145
rect 56390 915 56420 925
rect 56445 1145 56475 1155
rect 56445 925 56450 1145
rect 56470 925 56475 1145
rect 56445 915 56475 925
rect 56500 1145 56530 1155
rect 56500 925 56505 1145
rect 56525 925 56530 1145
rect 56500 915 56530 925
rect 56555 1145 56585 1155
rect 56555 925 56560 1145
rect 56580 925 56585 1145
rect 56555 915 56585 925
rect 56610 1145 56640 1155
rect 56610 925 56615 1145
rect 56635 925 56640 1145
rect 56610 915 56640 925
rect 56665 1145 56695 1155
rect 56665 925 56670 1145
rect 56690 925 56695 1145
rect 56665 915 56695 925
rect 56720 1145 56750 1155
rect 56720 925 56725 1145
rect 56745 925 56750 1145
rect 56720 915 56750 925
rect 56775 1145 56805 1155
rect 56775 925 56780 1145
rect 56800 925 56805 1145
rect 56775 915 56805 925
rect 56830 1145 56860 1155
rect 56830 925 56835 1145
rect 56855 925 56860 1145
rect 56830 915 56860 925
rect 56885 1145 56915 1155
rect 56885 925 56890 1145
rect 56910 925 56915 1145
rect 56885 915 56915 925
rect 56940 1145 56970 1155
rect 56940 925 56945 1145
rect 56965 925 56970 1145
rect 56940 915 56970 925
rect 56995 1145 57025 1155
rect 56995 925 57000 1145
rect 57020 925 57025 1145
rect 56995 915 57025 925
rect 57050 1145 57080 1155
rect 57050 925 57055 1145
rect 57075 925 57080 1145
rect 57050 915 57080 925
rect 57105 1145 57135 1155
rect 57105 925 57110 1145
rect 57130 925 57135 1145
rect 57105 915 57135 925
rect 57160 1145 57190 1155
rect 57160 925 57165 1145
rect 57185 925 57190 1145
rect 57160 915 57190 925
rect 57215 1145 57245 1155
rect 57215 925 57220 1145
rect 57240 925 57245 1145
rect 57215 915 57245 925
rect 57270 1145 57300 1155
rect 57270 925 57275 1145
rect 57295 925 57300 1145
rect 57270 915 57300 925
rect 57325 1145 57355 1155
rect 57325 925 57330 1145
rect 57350 925 57355 1145
rect 57325 915 57355 925
rect 57380 1145 57410 1155
rect 57380 925 57385 1145
rect 57405 925 57410 1145
rect 57380 915 57410 925
rect 57435 1145 57465 1155
rect 57435 925 57440 1145
rect 57460 925 57465 1145
rect 57435 915 57465 925
rect 57490 1145 57560 1155
rect 57490 925 57495 1145
rect 57515 925 57535 1145
rect 57555 925 57560 1145
rect 57490 915 57560 925
rect 56220 885 56260 895
rect 56220 865 56230 885
rect 56250 865 56260 885
rect 56220 855 56260 865
rect 57485 885 57525 895
rect 57485 865 57495 885
rect 57515 865 57525 885
rect 57485 855 57525 865
rect 56595 740 56635 750
rect 56595 720 56605 740
rect 56625 720 56635 740
rect 56595 710 56635 720
rect 57040 740 57080 750
rect 57040 720 57050 740
rect 57070 720 57080 740
rect 57040 710 57080 720
rect 56395 680 56465 690
rect 56395 560 56400 680
rect 56420 560 56440 680
rect 56460 560 56465 680
rect 56395 550 56465 560
rect 56490 680 56520 690
rect 56490 560 56495 680
rect 56515 560 56520 680
rect 56490 550 56520 560
rect 56545 680 56575 690
rect 56545 560 56550 680
rect 56570 560 56575 680
rect 56545 550 56575 560
rect 56600 680 56630 690
rect 56600 560 56605 680
rect 56625 560 56630 680
rect 56600 550 56630 560
rect 56655 680 56685 690
rect 56655 560 56660 680
rect 56680 560 56685 680
rect 56655 550 56685 560
rect 56710 680 56740 690
rect 56710 560 56715 680
rect 56735 560 56740 680
rect 56710 550 56740 560
rect 56765 680 56835 690
rect 56765 560 56770 680
rect 56790 560 56810 680
rect 56830 560 56835 680
rect 56765 550 56835 560
rect 56875 680 56905 690
rect 56875 560 56880 680
rect 56900 560 56905 680
rect 56875 550 56905 560
rect 57215 680 57245 690
rect 57215 560 57220 680
rect 57240 560 57245 680
rect 57215 550 57245 560
rect 55590 525 55660 535
rect 58145 535 58150 1205
rect 58170 535 58190 1205
rect 58210 535 58215 1205
rect 56435 520 56465 530
rect 54990 495 55020 505
rect 54990 475 54995 495
rect 55015 475 55020 495
rect 54990 465 55020 475
rect 55590 495 55620 505
rect 55590 475 55595 495
rect 55615 475 55620 495
rect 56435 500 56440 520
rect 56460 500 56465 520
rect 56435 490 56465 500
rect 56765 520 56795 530
rect 58145 525 58215 535
rect 58285 1205 58315 1215
rect 58285 535 58290 1205
rect 58310 535 58315 1205
rect 58285 525 58315 535
rect 58385 1205 58415 1215
rect 58385 535 58390 1205
rect 58410 535 58415 1205
rect 58385 525 58415 535
rect 58485 1205 58515 1215
rect 58485 535 58490 1205
rect 58510 535 58515 1205
rect 58485 525 58515 535
rect 58585 1205 58615 1215
rect 58585 535 58590 1205
rect 58610 535 58615 1205
rect 58585 525 58615 535
rect 58685 1205 58715 1215
rect 58685 535 58690 1205
rect 58710 535 58715 1205
rect 58685 525 58715 535
rect 58785 1205 58855 1215
rect 58785 535 58790 1205
rect 58810 535 58830 1205
rect 58850 535 58855 1205
rect 58975 1195 59010 1205
rect 58975 1170 58980 1195
rect 59005 1170 59010 1195
rect 58975 1160 59010 1170
rect 59035 1195 59070 1205
rect 59035 1170 59040 1195
rect 59065 1170 59070 1195
rect 59035 1160 59070 1170
rect 58785 525 58855 535
rect 56765 500 56770 520
rect 56790 500 56795 520
rect 56765 490 56795 500
rect 58185 495 58215 505
rect 55590 465 55620 475
rect 58185 475 58190 495
rect 58210 475 58215 495
rect 58185 465 58215 475
rect 58785 495 58815 505
rect 58785 475 58790 495
rect 58810 475 58815 495
rect 58785 465 58815 475
rect 59010 473 59035 523
<< viali >>
rect 56095 4735 56115 4755
rect 56275 4735 56295 4755
rect 57035 4735 57055 4755
rect 57215 4735 57235 4755
rect 57505 4735 57525 4755
rect 57685 4735 57705 4755
rect 56095 4375 56115 4695
rect 56155 4375 56175 4695
rect 56215 4375 56235 4695
rect 56275 4375 56295 4695
rect 56565 4565 56585 4585
rect 56745 4565 56765 4585
rect 56565 4375 56585 4525
rect 56625 4375 56645 4525
rect 56685 4375 56705 4525
rect 56745 4375 56765 4525
rect 57035 4375 57055 4695
rect 57095 4375 57115 4695
rect 57155 4375 57175 4695
rect 57215 4375 57235 4695
rect 57505 4375 57525 4695
rect 57565 4375 57585 4695
rect 57625 4375 57645 4695
rect 57685 4375 57705 4695
rect 56160 4285 56180 4305
rect 56635 4285 56655 4305
rect 57145 4285 57165 4305
rect 57581 4275 57601 4295
rect 54935 3705 54955 4025
rect 54995 3705 55015 4025
rect 55055 3705 55075 4025
rect 55115 3705 55135 4025
rect 55175 3705 55195 4025
rect 55235 3705 55255 4025
rect 55295 3705 55315 4025
rect 55355 3705 55375 4025
rect 55415 3705 55435 4025
rect 55475 3705 55495 4025
rect 55535 3705 55555 4025
rect 55595 3705 55615 4025
rect 55655 3705 55675 4025
rect 56015 3705 56035 4025
rect 56075 3705 56095 4025
rect 56135 3705 56155 4025
rect 56195 3705 56215 4025
rect 56255 3705 56275 4025
rect 56315 3705 56335 4025
rect 56375 3705 56395 4025
rect 56435 3705 56455 4025
rect 56495 3705 56515 4025
rect 56555 3705 56575 4025
rect 56615 3705 56635 4025
rect 56675 3705 56695 4025
rect 56735 3705 56755 4025
rect 57045 3705 57065 4025
rect 57105 3705 57125 4025
rect 57165 3705 57185 4025
rect 57225 3705 57245 4025
rect 57285 3705 57305 4025
rect 57345 3705 57365 4025
rect 57405 3705 57425 4025
rect 57465 3705 57485 4025
rect 57525 3705 57545 4025
rect 57585 3705 57605 4025
rect 57645 3705 57665 4025
rect 57705 3705 57725 4025
rect 57765 3705 57785 4025
rect 58130 3705 58150 4025
rect 58190 3705 58210 4025
rect 58250 3705 58270 4025
rect 58310 3705 58330 4025
rect 58370 3705 58390 4025
rect 58430 3705 58450 4025
rect 58490 3705 58510 4025
rect 58550 3705 58570 4025
rect 58610 3705 58630 4025
rect 58670 3705 58690 4025
rect 58730 3705 58750 4025
rect 58790 3705 58810 4025
rect 58850 3705 58870 4025
rect 54935 3645 54955 3665
rect 55655 3645 55675 3665
rect 56015 3645 56035 3665
rect 56735 3645 56755 3665
rect 57045 3645 57065 3665
rect 57765 3645 57785 3665
rect 58130 3645 58150 3665
rect 58850 3645 58870 3665
rect 56375 3580 56395 3600
rect 57405 3580 57425 3600
rect 55295 3535 55315 3555
rect 58490 3535 58510 3555
rect 54560 3295 54580 3315
rect 54615 3295 54635 3315
rect 54670 3295 54690 3315
rect 54965 3290 54985 3310
rect 55625 3290 55645 3310
rect 58160 3290 58180 3310
rect 58820 3290 58840 3310
rect 59110 3295 59130 3315
rect 59165 3295 59185 3315
rect 59220 3295 59240 3315
rect 54560 2690 54580 2710
rect 54615 2690 54635 2710
rect 54670 2690 54690 2710
rect 54965 2680 54985 3250
rect 55020 2680 55040 3250
rect 55075 2680 55095 3250
rect 55130 2680 55150 3250
rect 55185 2680 55205 3250
rect 55240 2680 55260 3250
rect 55295 2680 55315 3250
rect 55350 2680 55370 3250
rect 55405 2680 55425 3250
rect 55460 2680 55480 3250
rect 55515 2680 55535 3250
rect 55570 2680 55590 3250
rect 55625 2680 55645 3250
rect 56285 3220 56305 3240
rect 56340 3220 56360 3240
rect 56395 3220 56415 3240
rect 56450 3220 56470 3240
rect 56505 3220 56525 3240
rect 56560 3220 56580 3240
rect 56615 3220 56635 3240
rect 56670 3220 56690 3240
rect 56725 3220 56745 3240
rect 56780 3220 56800 3240
rect 56835 3220 56855 3240
rect 56890 3220 56910 3240
rect 56945 3220 56965 3240
rect 57000 3220 57020 3240
rect 57055 3220 57075 3240
rect 57110 3220 57130 3240
rect 57165 3220 57185 3240
rect 57220 3220 57240 3240
rect 57275 3220 57295 3240
rect 57330 3220 57350 3240
rect 57385 3220 57405 3240
rect 57440 3220 57460 3240
rect 57495 3220 57515 3240
rect 56285 3160 56305 3180
rect 56395 3160 56415 3180
rect 56835 3160 56855 3180
rect 57495 3160 57515 3180
rect 56045 2995 56065 3015
rect 56695 2995 56715 3015
rect 57085 2995 57105 3015
rect 57735 2995 57755 3015
rect 56040 2910 56060 2930
rect 56095 2910 56115 2930
rect 56150 2910 56170 2930
rect 56205 2910 56225 2930
rect 56260 2910 56280 2930
rect 56315 2910 56335 2930
rect 56370 2910 56390 2930
rect 56425 2910 56445 2930
rect 56480 2910 56500 2930
rect 56535 2910 56555 2930
rect 56590 2910 56610 2930
rect 56645 2910 56665 2930
rect 56700 2910 56720 2930
rect 57080 2910 57100 2930
rect 57135 2910 57155 2930
rect 57190 2910 57210 2930
rect 57245 2910 57265 2930
rect 57300 2910 57320 2930
rect 57355 2910 57375 2930
rect 57410 2910 57430 2930
rect 57465 2910 57485 2930
rect 57520 2910 57540 2930
rect 57575 2910 57595 2930
rect 57630 2910 57650 2930
rect 57685 2910 57705 2930
rect 57740 2910 57760 2930
rect 56040 2850 56060 2870
rect 56700 2850 56720 2870
rect 57080 2850 57100 2870
rect 57740 2850 57760 2870
rect 56100 2765 56120 2785
rect 56585 2765 56605 2785
rect 57195 2765 57215 2785
rect 58160 2680 58180 3250
rect 58215 2680 58235 3250
rect 58270 2680 58290 3250
rect 58325 2680 58345 3250
rect 58380 2680 58400 3250
rect 58435 2680 58455 3250
rect 58490 2680 58510 3250
rect 58545 2680 58565 3250
rect 58600 2680 58620 3250
rect 58655 2680 58675 3250
rect 58710 2680 58730 3250
rect 58765 2680 58785 3250
rect 58820 2680 58840 3250
rect 59110 2690 59130 2710
rect 59165 2690 59185 2710
rect 59220 2690 59240 2710
rect 56725 2610 56745 2630
rect 56945 2610 56965 2630
rect 55185 2560 55205 2580
rect 56560 2550 56580 2570
rect 56615 2550 56635 2570
rect 56670 2550 56690 2570
rect 56725 2550 56745 2570
rect 56780 2550 56800 2570
rect 56835 2550 56855 2570
rect 56890 2550 56910 2570
rect 56945 2550 56965 2570
rect 57000 2550 57020 2570
rect 57055 2550 57075 2570
rect 57110 2550 57130 2570
rect 57165 2550 57185 2570
rect 57220 2550 57240 2570
rect 58600 2560 58620 2580
rect 56560 2490 56580 2510
rect 57220 2490 57240 2510
rect 54965 2395 54985 2415
rect 55625 2395 55645 2415
rect 58160 2395 58180 2415
rect 58820 2395 58840 2415
rect 54965 2185 54985 2355
rect 55020 2185 55040 2355
rect 55075 2185 55095 2355
rect 55130 2185 55150 2355
rect 55185 2185 55205 2355
rect 55240 2185 55260 2355
rect 55295 2185 55315 2355
rect 55350 2185 55370 2355
rect 55405 2185 55425 2355
rect 55460 2185 55480 2355
rect 55515 2185 55535 2355
rect 55570 2185 55590 2355
rect 55625 2185 55645 2355
rect 56100 2245 56120 2265
rect 56640 2245 56660 2265
rect 57140 2245 57160 2265
rect 58160 2185 58180 2355
rect 58215 2185 58235 2355
rect 58270 2185 58290 2355
rect 58325 2185 58345 2355
rect 58380 2185 58400 2355
rect 58435 2185 58455 2355
rect 58490 2185 58510 2355
rect 58545 2185 58565 2355
rect 58600 2185 58620 2355
rect 58655 2185 58675 2355
rect 58710 2185 58730 2355
rect 58765 2185 58785 2355
rect 58820 2185 58840 2355
rect 55075 2125 55095 2145
rect 55185 2125 55205 2145
rect 55295 2125 55315 2145
rect 55405 2125 55425 2145
rect 55515 2125 55535 2145
rect 55460 2030 55480 2050
rect 56040 2045 56060 2165
rect 56095 2045 56115 2165
rect 56150 2045 56170 2165
rect 56205 2045 56225 2165
rect 56260 2045 56280 2165
rect 56315 2045 56335 2165
rect 56370 2045 56390 2165
rect 56425 2045 56445 2165
rect 56480 2045 56500 2165
rect 56535 2045 56555 2165
rect 56590 2045 56610 2165
rect 56645 2045 56665 2165
rect 56700 2045 56720 2165
rect 57080 2045 57100 2165
rect 57135 2045 57155 2165
rect 57190 2045 57210 2165
rect 57245 2045 57265 2165
rect 57300 2045 57320 2165
rect 57355 2045 57375 2165
rect 57410 2045 57430 2165
rect 57465 2045 57485 2165
rect 57520 2045 57540 2165
rect 57575 2045 57595 2165
rect 57630 2045 57650 2165
rect 57685 2045 57705 2165
rect 57740 2045 57760 2165
rect 58270 2125 58290 2145
rect 58380 2125 58400 2145
rect 58490 2125 58510 2145
rect 58600 2125 58620 2145
rect 58710 2125 58730 2145
rect 56040 1985 56060 2005
rect 56700 1985 56720 2005
rect 57080 1985 57100 2005
rect 58325 2030 58345 2050
rect 57740 1985 57760 2005
rect 54455 1565 54480 1590
rect 54515 1565 54540 1590
rect 54575 1565 54600 1590
rect 54965 1625 54985 1895
rect 55020 1625 55040 1895
rect 55075 1625 55095 1895
rect 55130 1625 55150 1895
rect 55185 1625 55205 1895
rect 55240 1625 55260 1895
rect 55295 1625 55315 1895
rect 55350 1625 55370 1895
rect 55405 1625 55425 1895
rect 55460 1625 55480 1895
rect 55515 1625 55535 1895
rect 55570 1625 55590 1895
rect 55625 1625 55645 1895
rect 56045 1760 56065 1780
rect 56695 1760 56715 1780
rect 56855 1760 56875 1780
rect 56908 1760 56928 1780
rect 57085 1760 57105 1780
rect 57735 1760 57755 1780
rect 54635 1565 54660 1590
rect 54965 1565 54985 1585
rect 55625 1565 55645 1585
rect 56040 1575 56060 1695
rect 56095 1575 56115 1695
rect 56150 1575 56170 1695
rect 56205 1575 56225 1695
rect 56260 1575 56280 1695
rect 56315 1575 56335 1695
rect 56370 1575 56390 1695
rect 56425 1575 56445 1695
rect 56480 1575 56500 1695
rect 56535 1575 56555 1695
rect 56590 1575 56610 1695
rect 56645 1575 56665 1695
rect 56700 1575 56720 1695
rect 56780 1575 56800 1695
rect 56835 1575 56855 1695
rect 56890 1575 56910 1695
rect 56945 1575 56965 1695
rect 57000 1575 57020 1695
rect 57080 1575 57100 1695
rect 57135 1575 57155 1695
rect 57190 1575 57210 1695
rect 57245 1575 57265 1695
rect 57300 1575 57320 1695
rect 57355 1575 57375 1695
rect 57410 1575 57430 1695
rect 57465 1575 57485 1695
rect 57520 1575 57540 1695
rect 57575 1575 57595 1695
rect 57630 1575 57650 1695
rect 57685 1575 57705 1695
rect 57740 1575 57760 1695
rect 58160 1625 58180 1895
rect 58215 1625 58235 1895
rect 58270 1625 58290 1895
rect 58325 1625 58345 1895
rect 58380 1625 58400 1895
rect 58435 1625 58455 1895
rect 58490 1625 58510 1895
rect 58545 1625 58565 1895
rect 58600 1625 58620 1895
rect 58655 1625 58675 1895
rect 58710 1625 58730 1895
rect 58765 1625 58785 1895
rect 58820 1625 58840 1895
rect 58160 1565 58180 1585
rect 56040 1515 56060 1535
rect 56740 1515 56760 1535
rect 57040 1515 57060 1535
rect 58820 1565 58840 1585
rect 57740 1515 57760 1535
rect 59140 1515 59165 1540
rect 59200 1515 59225 1540
rect 59260 1515 59285 1540
rect 59320 1515 59345 1540
rect 55395 1245 55415 1265
rect 57415 1240 57435 1260
rect 58440 1245 58460 1265
rect 54715 1165 54740 1190
rect 54775 1165 54800 1190
rect 54995 535 55015 1205
rect 55095 535 55115 1205
rect 55195 535 55215 1205
rect 55295 535 55315 1205
rect 55395 535 55415 1205
rect 55495 535 55515 1205
rect 55595 535 55615 1205
rect 56835 1185 56855 1205
rect 56230 925 56250 1145
rect 56285 925 56305 1145
rect 56340 925 56360 1145
rect 56395 925 56415 1145
rect 56450 925 56470 1145
rect 56505 925 56525 1145
rect 56560 925 56580 1145
rect 56615 925 56635 1145
rect 56670 925 56690 1145
rect 56725 925 56745 1145
rect 56780 925 56800 1145
rect 56835 925 56855 1145
rect 56890 925 56910 1145
rect 56945 925 56965 1145
rect 57000 925 57020 1145
rect 57055 925 57075 1145
rect 57110 925 57130 1145
rect 57165 925 57185 1145
rect 57220 925 57240 1145
rect 57275 925 57295 1145
rect 57330 925 57350 1145
rect 57385 925 57405 1145
rect 57440 925 57460 1145
rect 57495 925 57515 1145
rect 56230 865 56250 885
rect 57495 865 57515 885
rect 56605 720 56625 740
rect 57050 720 57070 740
rect 56440 560 56460 680
rect 56495 560 56515 680
rect 56550 560 56570 680
rect 56605 560 56625 680
rect 56660 560 56680 680
rect 56715 560 56735 680
rect 56770 560 56790 680
rect 56880 560 56900 680
rect 57220 560 57240 680
rect 58190 535 58210 1205
rect 54995 475 55015 495
rect 55595 475 55615 495
rect 56440 500 56460 520
rect 58290 535 58310 1205
rect 58390 535 58410 1205
rect 58490 535 58510 1205
rect 58590 535 58610 1205
rect 58690 535 58710 1205
rect 58790 535 58810 1205
rect 58980 1170 59005 1195
rect 59040 1170 59065 1195
rect 56770 500 56790 520
rect 58190 475 58210 495
rect 58790 475 58810 495
<< metal1 >>
rect 56205 4815 56245 4820
rect 56205 4785 56210 4815
rect 56240 4785 56245 4815
rect 56085 4760 56125 4765
rect 56085 4730 56090 4760
rect 56120 4730 56125 4760
rect 56085 4725 56125 4730
rect 56205 4760 56245 4785
rect 56675 4815 56715 4820
rect 56675 4785 56680 4815
rect 56710 4785 56715 4815
rect 56675 4780 56715 4785
rect 56205 4730 56210 4760
rect 56240 4730 56245 4760
rect 56205 4725 56245 4730
rect 56265 4760 56305 4765
rect 56265 4730 56270 4760
rect 56300 4730 56305 4760
rect 56265 4725 56305 4730
rect 56090 4695 56120 4725
rect 56090 4375 56095 4695
rect 56115 4375 56120 4695
rect 56090 4365 56120 4375
rect 56150 4695 56180 4705
rect 56150 4375 56155 4695
rect 56175 4375 56180 4695
rect 56150 4315 56180 4375
rect 56210 4695 56240 4725
rect 56210 4375 56215 4695
rect 56235 4375 56240 4695
rect 56210 4360 56240 4375
rect 56270 4695 56300 4725
rect 56270 4375 56275 4695
rect 56295 4375 56300 4695
rect 56555 4590 56595 4595
rect 56555 4560 56560 4590
rect 56590 4560 56595 4590
rect 56555 4555 56595 4560
rect 56615 4590 56655 4595
rect 56615 4560 56620 4590
rect 56650 4560 56655 4590
rect 56615 4555 56655 4560
rect 56270 4365 56300 4375
rect 56560 4525 56590 4555
rect 56560 4375 56565 4525
rect 56585 4375 56590 4525
rect 56560 4365 56590 4375
rect 56620 4525 56650 4555
rect 56620 4375 56625 4525
rect 56645 4375 56650 4525
rect 56620 4365 56650 4375
rect 56680 4525 56710 4780
rect 56890 4765 56910 6101
rect 57085 4815 57125 4820
rect 57085 4785 57090 4815
rect 57120 4785 57125 4815
rect 57085 4780 57125 4785
rect 57555 4815 57595 4820
rect 57555 4785 57560 4815
rect 57590 4785 57595 4815
rect 56880 4760 56920 4765
rect 56880 4730 56885 4760
rect 56915 4730 56920 4760
rect 56880 4725 56920 4730
rect 57025 4760 57065 4765
rect 57025 4730 57030 4760
rect 57060 4730 57065 4760
rect 57025 4725 57065 4730
rect 56890 4595 56910 4725
rect 57030 4695 57060 4725
rect 56735 4590 56775 4595
rect 56735 4560 56740 4590
rect 56770 4560 56775 4590
rect 56735 4555 56775 4560
rect 56880 4590 56920 4595
rect 56880 4560 56885 4590
rect 56915 4560 56920 4590
rect 56880 4555 56920 4560
rect 56680 4375 56685 4525
rect 56705 4375 56710 4525
rect 56680 4360 56710 4375
rect 56740 4525 56770 4555
rect 56740 4375 56745 4525
rect 56765 4375 56770 4525
rect 56740 4365 56770 4375
rect 56205 4355 56245 4360
rect 56205 4325 56210 4355
rect 56240 4325 56245 4355
rect 56205 4320 56245 4325
rect 56675 4355 56715 4360
rect 56675 4325 56680 4355
rect 56710 4325 56715 4355
rect 56675 4320 56715 4325
rect 56150 4310 56190 4315
rect 56150 4280 56155 4310
rect 56185 4280 56190 4310
rect 56150 4275 56190 4280
rect 56630 4310 56660 4315
rect 56630 4275 56660 4280
rect 56825 4310 56865 4315
rect 56825 4280 56830 4310
rect 56860 4280 56865 4310
rect 56825 4275 56865 4280
rect 55285 4200 55325 4205
rect 55285 4170 55290 4200
rect 55320 4170 55325 4200
rect 55285 4165 55325 4170
rect 55760 4200 55800 4205
rect 55760 4170 55765 4200
rect 55795 4170 55800 4200
rect 55760 4165 55800 4170
rect 55295 4125 55315 4165
rect 54925 4120 54965 4125
rect 54925 4090 54930 4120
rect 54960 4090 54965 4120
rect 54925 4085 54965 4090
rect 55045 4120 55085 4125
rect 55045 4090 55050 4120
rect 55080 4090 55085 4120
rect 55045 4085 55085 4090
rect 55165 4120 55205 4125
rect 55165 4090 55170 4120
rect 55200 4090 55205 4120
rect 55165 4085 55205 4090
rect 55285 4120 55325 4125
rect 55285 4090 55290 4120
rect 55320 4090 55325 4120
rect 55285 4085 55325 4090
rect 55405 4120 55445 4125
rect 55405 4090 55410 4120
rect 55440 4090 55445 4120
rect 55405 4085 55445 4090
rect 55525 4120 55565 4125
rect 55525 4090 55530 4120
rect 55560 4090 55565 4120
rect 55525 4085 55565 4090
rect 55645 4120 55685 4125
rect 55645 4090 55650 4120
rect 55680 4090 55685 4120
rect 55645 4085 55685 4090
rect 54930 4025 54960 4085
rect 54985 4075 55025 4080
rect 54985 4045 54990 4075
rect 55020 4045 55025 4075
rect 54985 4040 55025 4045
rect 54930 3705 54935 4025
rect 54955 3705 54960 4025
rect 54930 3665 54960 3705
rect 54990 4025 55020 4040
rect 54990 3705 54995 4025
rect 55015 3705 55020 4025
rect 54990 3690 55020 3705
rect 55050 4025 55080 4085
rect 55105 4075 55145 4080
rect 55105 4045 55110 4075
rect 55140 4045 55145 4075
rect 55105 4040 55145 4045
rect 55050 3705 55055 4025
rect 55075 3705 55080 4025
rect 55050 3695 55080 3705
rect 55110 4025 55140 4040
rect 55110 3705 55115 4025
rect 55135 3705 55140 4025
rect 55110 3690 55140 3705
rect 55170 4025 55200 4085
rect 55225 4075 55265 4080
rect 55225 4045 55230 4075
rect 55260 4045 55265 4075
rect 55225 4040 55265 4045
rect 55170 3705 55175 4025
rect 55195 3705 55200 4025
rect 55170 3695 55200 3705
rect 55230 4025 55260 4040
rect 55230 3705 55235 4025
rect 55255 3705 55260 4025
rect 55230 3690 55260 3705
rect 55290 4025 55320 4085
rect 55345 4075 55385 4080
rect 55345 4045 55350 4075
rect 55380 4045 55385 4075
rect 55345 4040 55385 4045
rect 55290 3705 55295 4025
rect 55315 3705 55320 4025
rect 55290 3695 55320 3705
rect 55350 4025 55380 4040
rect 55350 3705 55355 4025
rect 55375 3705 55380 4025
rect 55350 3690 55380 3705
rect 55410 4025 55440 4085
rect 55465 4075 55505 4080
rect 55465 4045 55470 4075
rect 55500 4045 55505 4075
rect 55465 4040 55505 4045
rect 55410 3705 55415 4025
rect 55435 3705 55440 4025
rect 55410 3695 55440 3705
rect 55470 4025 55500 4040
rect 55470 3705 55475 4025
rect 55495 3705 55500 4025
rect 55470 3690 55500 3705
rect 55530 4025 55560 4085
rect 55585 4075 55625 4080
rect 55585 4045 55590 4075
rect 55620 4045 55625 4075
rect 55585 4040 55625 4045
rect 55530 3705 55535 4025
rect 55555 3705 55560 4025
rect 55530 3695 55560 3705
rect 55590 4025 55620 4040
rect 55590 3705 55595 4025
rect 55615 3705 55620 4025
rect 55590 3690 55620 3705
rect 55650 4025 55680 4085
rect 55650 3705 55655 4025
rect 55675 3705 55680 4025
rect 54930 3645 54935 3665
rect 54955 3645 54960 3665
rect 54985 3685 55025 3690
rect 54985 3655 54990 3685
rect 55020 3655 55025 3685
rect 54985 3650 55025 3655
rect 55105 3685 55145 3690
rect 55105 3655 55110 3685
rect 55140 3655 55145 3685
rect 55105 3650 55145 3655
rect 55225 3685 55265 3690
rect 55225 3655 55230 3685
rect 55260 3655 55265 3685
rect 55225 3650 55265 3655
rect 55345 3685 55385 3690
rect 55345 3655 55350 3685
rect 55380 3655 55385 3685
rect 55345 3650 55385 3655
rect 55465 3685 55505 3690
rect 55465 3655 55470 3685
rect 55500 3655 55505 3685
rect 55465 3650 55505 3655
rect 55585 3685 55625 3690
rect 55585 3655 55590 3685
rect 55620 3655 55625 3685
rect 55585 3650 55625 3655
rect 55650 3665 55680 3705
rect 54930 3635 54960 3645
rect 55650 3645 55655 3665
rect 55675 3645 55680 3665
rect 55650 3635 55680 3645
rect 55285 3560 55325 3565
rect 55285 3530 55290 3560
rect 55320 3530 55325 3560
rect 55285 3525 55325 3530
rect 54605 3400 54645 3405
rect 54605 3370 54610 3400
rect 54640 3370 54645 3400
rect 55770 3385 55790 4165
rect 55910 4120 55950 4125
rect 55910 4090 55915 4120
rect 55945 4090 55950 4120
rect 55910 4085 55950 4090
rect 56005 4120 56045 4125
rect 56005 4090 56010 4120
rect 56040 4090 56045 4120
rect 56005 4085 56045 4090
rect 56125 4120 56165 4125
rect 56125 4090 56130 4120
rect 56160 4090 56165 4120
rect 56125 4085 56165 4090
rect 56245 4120 56285 4125
rect 56245 4090 56250 4120
rect 56280 4090 56285 4120
rect 56245 4085 56285 4090
rect 56365 4120 56405 4125
rect 56365 4090 56370 4120
rect 56400 4090 56405 4120
rect 56365 4085 56405 4090
rect 56485 4120 56525 4125
rect 56485 4090 56490 4120
rect 56520 4090 56525 4120
rect 56485 4085 56525 4090
rect 56605 4120 56645 4125
rect 56605 4090 56610 4120
rect 56640 4090 56645 4120
rect 56605 4085 56645 4090
rect 56725 4120 56765 4125
rect 56725 4090 56730 4120
rect 56760 4090 56765 4120
rect 56725 4085 56765 4090
rect 55920 3690 55940 4085
rect 56010 4025 56040 4085
rect 56065 4075 56105 4080
rect 56065 4045 56070 4075
rect 56100 4045 56105 4075
rect 56065 4040 56105 4045
rect 56010 3705 56015 4025
rect 56035 3705 56040 4025
rect 55910 3685 55950 3690
rect 55910 3655 55915 3685
rect 55945 3655 55950 3685
rect 55910 3650 55950 3655
rect 56010 3665 56040 3705
rect 56070 4025 56100 4040
rect 56070 3705 56075 4025
rect 56095 3705 56100 4025
rect 56070 3690 56100 3705
rect 56130 4025 56160 4085
rect 56185 4075 56225 4080
rect 56185 4045 56190 4075
rect 56220 4045 56225 4075
rect 56185 4040 56225 4045
rect 56130 3705 56135 4025
rect 56155 3705 56160 4025
rect 56130 3695 56160 3705
rect 56190 4025 56220 4040
rect 56190 3705 56195 4025
rect 56215 3705 56220 4025
rect 56190 3690 56220 3705
rect 56250 4025 56280 4085
rect 56305 4075 56345 4080
rect 56305 4045 56310 4075
rect 56340 4045 56345 4075
rect 56305 4040 56345 4045
rect 56250 3705 56255 4025
rect 56275 3705 56280 4025
rect 56250 3695 56280 3705
rect 56310 4025 56340 4040
rect 56310 3705 56315 4025
rect 56335 3705 56340 4025
rect 56310 3690 56340 3705
rect 56370 4025 56400 4085
rect 56425 4075 56465 4080
rect 56425 4045 56430 4075
rect 56460 4045 56465 4075
rect 56425 4040 56465 4045
rect 56370 3705 56375 4025
rect 56395 3705 56400 4025
rect 56370 3695 56400 3705
rect 56430 4025 56460 4040
rect 56430 3705 56435 4025
rect 56455 3705 56460 4025
rect 56430 3690 56460 3705
rect 56490 4025 56520 4085
rect 56545 4075 56585 4080
rect 56545 4045 56550 4075
rect 56580 4045 56585 4075
rect 56545 4040 56585 4045
rect 56490 3705 56495 4025
rect 56515 3705 56520 4025
rect 56490 3695 56520 3705
rect 56550 4025 56580 4040
rect 56550 3705 56555 4025
rect 56575 3705 56580 4025
rect 56550 3690 56580 3705
rect 56610 4025 56640 4085
rect 56665 4075 56705 4080
rect 56665 4045 56670 4075
rect 56700 4045 56705 4075
rect 56665 4040 56705 4045
rect 56610 3705 56615 4025
rect 56635 3705 56640 4025
rect 56610 3695 56640 3705
rect 56670 4025 56700 4040
rect 56670 3705 56675 4025
rect 56695 3705 56700 4025
rect 56670 3690 56700 3705
rect 56730 4025 56760 4085
rect 56730 3705 56735 4025
rect 56755 3705 56760 4025
rect 56010 3645 56015 3665
rect 56035 3645 56040 3665
rect 56065 3685 56105 3690
rect 56065 3655 56070 3685
rect 56100 3655 56105 3685
rect 56065 3650 56105 3655
rect 56185 3685 56225 3690
rect 56185 3655 56190 3685
rect 56220 3655 56225 3685
rect 56185 3650 56225 3655
rect 56305 3685 56345 3690
rect 56305 3655 56310 3685
rect 56340 3655 56345 3685
rect 56305 3650 56345 3655
rect 56425 3685 56465 3690
rect 56425 3655 56430 3685
rect 56460 3655 56465 3685
rect 56425 3650 56465 3655
rect 56545 3685 56585 3690
rect 56545 3655 56550 3685
rect 56580 3655 56585 3685
rect 56545 3650 56585 3655
rect 56665 3685 56705 3690
rect 56665 3655 56670 3685
rect 56700 3655 56705 3685
rect 56665 3650 56705 3655
rect 56730 3665 56760 3705
rect 56010 3635 56040 3645
rect 54605 3365 54645 3370
rect 54955 3380 54995 3385
rect 54615 3325 54635 3365
rect 54955 3350 54960 3380
rect 54990 3350 54995 3380
rect 54955 3345 54995 3350
rect 55065 3380 55105 3385
rect 55065 3350 55070 3380
rect 55100 3350 55105 3380
rect 55065 3345 55105 3350
rect 55175 3380 55215 3385
rect 55175 3350 55180 3380
rect 55210 3350 55215 3380
rect 55175 3345 55215 3350
rect 55285 3380 55325 3385
rect 55285 3350 55290 3380
rect 55320 3350 55325 3380
rect 55285 3345 55325 3350
rect 55395 3380 55435 3385
rect 55395 3350 55400 3380
rect 55430 3350 55435 3380
rect 55395 3345 55435 3350
rect 55505 3380 55545 3385
rect 55505 3350 55510 3380
rect 55540 3350 55545 3380
rect 55505 3345 55545 3350
rect 55615 3380 55655 3385
rect 55615 3350 55620 3380
rect 55650 3350 55655 3380
rect 55615 3345 55655 3350
rect 55760 3380 55800 3385
rect 55760 3350 55765 3380
rect 55795 3350 55800 3380
rect 55760 3345 55800 3350
rect 54554 3315 54695 3325
rect 54554 3295 54560 3315
rect 54580 3295 54615 3315
rect 54635 3295 54670 3315
rect 54690 3295 54695 3315
rect 54554 3285 54695 3295
rect 54960 3310 54990 3345
rect 54960 3290 54965 3310
rect 54985 3290 54990 3310
rect 54960 3250 54990 3290
rect 55010 3300 55050 3305
rect 55010 3270 55015 3300
rect 55045 3270 55050 3300
rect 55010 3265 55050 3270
rect 54554 2710 54695 2720
rect 54554 2690 54560 2710
rect 54580 2690 54615 2710
rect 54635 2690 54670 2710
rect 54690 2690 54695 2710
rect 54554 2680 54695 2690
rect 54960 2680 54965 3250
rect 54985 2680 54990 3250
rect 54615 2595 54635 2680
rect 54960 2670 54990 2680
rect 55015 3250 55045 3265
rect 55015 2680 55020 3250
rect 55040 2680 55045 3250
rect 55015 2665 55045 2680
rect 55070 3250 55100 3345
rect 55120 3300 55160 3305
rect 55120 3270 55125 3300
rect 55155 3270 55160 3300
rect 55120 3265 55160 3270
rect 55070 2680 55075 3250
rect 55095 2680 55100 3250
rect 55070 2670 55100 2680
rect 55125 3250 55155 3265
rect 55125 2680 55130 3250
rect 55150 2680 55155 3250
rect 55125 2665 55155 2680
rect 55180 3250 55210 3345
rect 55230 3300 55270 3305
rect 55230 3270 55235 3300
rect 55265 3270 55270 3300
rect 55230 3265 55270 3270
rect 55180 2680 55185 3250
rect 55205 2680 55210 3250
rect 55180 2670 55210 2680
rect 55235 3250 55265 3265
rect 55235 2680 55240 3250
rect 55260 2680 55265 3250
rect 55235 2665 55265 2680
rect 55290 3250 55320 3345
rect 55340 3300 55380 3305
rect 55340 3270 55345 3300
rect 55375 3270 55380 3300
rect 55340 3265 55380 3270
rect 55290 2680 55295 3250
rect 55315 2680 55320 3250
rect 55290 2670 55320 2680
rect 55345 3250 55375 3265
rect 55345 2680 55350 3250
rect 55370 2680 55375 3250
rect 55345 2665 55375 2680
rect 55400 3250 55430 3345
rect 55450 3300 55490 3305
rect 55450 3270 55455 3300
rect 55485 3270 55490 3300
rect 55450 3265 55490 3270
rect 55400 2680 55405 3250
rect 55425 2680 55430 3250
rect 55400 2670 55430 2680
rect 55455 3250 55485 3265
rect 55455 2680 55460 3250
rect 55480 2680 55485 3250
rect 55455 2665 55485 2680
rect 55510 3250 55540 3345
rect 55620 3310 55650 3345
rect 55560 3300 55600 3305
rect 55560 3270 55565 3300
rect 55595 3270 55600 3300
rect 55560 3265 55600 3270
rect 55620 3290 55625 3310
rect 55645 3290 55650 3310
rect 55715 3325 55755 3330
rect 55715 3295 55720 3325
rect 55750 3295 55755 3325
rect 55715 3290 55755 3295
rect 55510 2680 55515 3250
rect 55535 2680 55540 3250
rect 55510 2670 55540 2680
rect 55565 3250 55595 3265
rect 55565 2680 55570 3250
rect 55590 2680 55595 3250
rect 55565 2665 55595 2680
rect 55620 3250 55650 3290
rect 55620 2680 55625 3250
rect 55645 2680 55650 3250
rect 55620 2670 55650 2680
rect 55010 2660 55050 2665
rect 55010 2630 55015 2660
rect 55045 2630 55050 2660
rect 55010 2625 55050 2630
rect 55120 2660 55160 2665
rect 55120 2630 55125 2660
rect 55155 2630 55160 2660
rect 55120 2625 55160 2630
rect 55230 2660 55270 2665
rect 55230 2630 55235 2660
rect 55265 2630 55270 2660
rect 55230 2625 55270 2630
rect 55340 2660 55380 2665
rect 55340 2630 55345 2660
rect 55375 2630 55380 2660
rect 55340 2625 55380 2630
rect 55450 2660 55490 2665
rect 55450 2630 55455 2660
rect 55485 2630 55490 2660
rect 55450 2625 55490 2630
rect 55560 2660 55600 2665
rect 55560 2630 55565 2660
rect 55595 2630 55600 2660
rect 55560 2625 55600 2630
rect 54605 2590 54645 2595
rect 54605 2560 54610 2590
rect 54640 2560 54645 2590
rect 54605 2555 54645 2560
rect 55175 2555 55180 2585
rect 55210 2555 55215 2585
rect 55460 2550 55480 2625
rect 55725 2595 55745 3290
rect 55770 2750 55790 3345
rect 56075 3330 56095 3650
rect 56730 3645 56735 3665
rect 56755 3645 56760 3665
rect 56730 3635 56760 3645
rect 56845 3610 56865 4275
rect 56890 4205 56910 4555
rect 57030 4375 57035 4695
rect 57055 4375 57060 4695
rect 57030 4365 57060 4375
rect 57090 4695 57120 4780
rect 57145 4760 57185 4765
rect 57145 4730 57150 4760
rect 57180 4730 57185 4760
rect 57145 4725 57185 4730
rect 57205 4760 57245 4765
rect 57205 4730 57210 4760
rect 57240 4730 57245 4760
rect 57205 4725 57245 4730
rect 57495 4760 57535 4765
rect 57495 4730 57500 4760
rect 57530 4730 57535 4760
rect 57495 4725 57535 4730
rect 57555 4760 57595 4785
rect 57555 4730 57560 4760
rect 57590 4730 57595 4760
rect 57555 4725 57595 4730
rect 57675 4760 57715 4765
rect 57675 4730 57680 4760
rect 57710 4730 57715 4760
rect 57675 4725 57715 4730
rect 57090 4375 57095 4695
rect 57115 4375 57120 4695
rect 57090 4360 57120 4375
rect 57150 4695 57180 4725
rect 57150 4375 57155 4695
rect 57175 4375 57180 4695
rect 57150 4365 57180 4375
rect 57210 4695 57240 4725
rect 57210 4375 57215 4695
rect 57235 4375 57240 4695
rect 57210 4365 57240 4375
rect 57500 4695 57530 4725
rect 57500 4375 57505 4695
rect 57525 4375 57530 4695
rect 57500 4365 57530 4375
rect 57560 4695 57590 4725
rect 57560 4375 57565 4695
rect 57585 4375 57590 4695
rect 57560 4360 57590 4375
rect 57620 4695 57650 4705
rect 57620 4375 57625 4695
rect 57645 4375 57650 4695
rect 57085 4355 57125 4360
rect 57085 4325 57090 4355
rect 57120 4325 57125 4355
rect 57085 4320 57125 4325
rect 57555 4355 57595 4360
rect 57555 4325 57560 4355
rect 57590 4325 57595 4355
rect 57555 4320 57595 4325
rect 57140 4305 57170 4315
rect 57140 4285 57145 4305
rect 57165 4285 57170 4305
rect 56935 4255 56975 4260
rect 56935 4225 56940 4255
rect 56970 4225 56975 4255
rect 57140 4250 57170 4285
rect 57576 4300 57606 4305
rect 57576 4265 57606 4270
rect 57620 4250 57650 4375
rect 57680 4695 57710 4725
rect 57680 4375 57685 4695
rect 57705 4375 57710 4695
rect 57680 4365 57710 4375
rect 56935 4220 56975 4225
rect 57135 4245 57175 4250
rect 56880 4200 56920 4205
rect 56880 4170 56885 4200
rect 56915 4170 56920 4200
rect 56880 4165 56920 4170
rect 56365 3605 56405 3610
rect 56365 3575 56370 3605
rect 56400 3575 56405 3605
rect 56365 3570 56405 3575
rect 56835 3605 56875 3610
rect 56835 3575 56840 3605
rect 56870 3575 56875 3605
rect 56835 3570 56875 3575
rect 56935 3565 56955 4220
rect 57135 4215 57140 4245
rect 57170 4215 57175 4245
rect 57135 4210 57175 4215
rect 57615 4245 57655 4250
rect 57615 4215 57620 4245
rect 57650 4215 57655 4245
rect 57615 4210 57655 4215
rect 58005 4200 58045 4205
rect 58005 4170 58010 4200
rect 58040 4170 58045 4200
rect 58005 4165 58045 4170
rect 58480 4200 58520 4205
rect 58480 4170 58485 4200
rect 58515 4170 58520 4200
rect 58480 4165 58520 4170
rect 57035 4120 57075 4125
rect 57035 4090 57040 4120
rect 57070 4090 57075 4120
rect 57035 4085 57075 4090
rect 57155 4120 57195 4125
rect 57155 4090 57160 4120
rect 57190 4090 57195 4120
rect 57155 4085 57195 4090
rect 57275 4120 57315 4125
rect 57275 4090 57280 4120
rect 57310 4090 57315 4120
rect 57275 4085 57315 4090
rect 57395 4120 57435 4125
rect 57395 4090 57400 4120
rect 57430 4090 57435 4120
rect 57395 4085 57435 4090
rect 57515 4120 57555 4125
rect 57515 4090 57520 4120
rect 57550 4090 57555 4120
rect 57515 4085 57555 4090
rect 57635 4120 57675 4125
rect 57635 4090 57640 4120
rect 57670 4090 57675 4120
rect 57635 4085 57675 4090
rect 57755 4120 57795 4125
rect 57755 4090 57760 4120
rect 57790 4090 57795 4120
rect 57755 4085 57795 4090
rect 57850 4120 57890 4125
rect 57850 4090 57855 4120
rect 57885 4090 57890 4120
rect 57850 4085 57890 4090
rect 57040 4025 57070 4085
rect 57095 4075 57135 4080
rect 57095 4045 57100 4075
rect 57130 4045 57135 4075
rect 57095 4040 57135 4045
rect 57040 3705 57045 4025
rect 57065 3705 57070 4025
rect 57040 3665 57070 3705
rect 57100 4025 57130 4040
rect 57100 3705 57105 4025
rect 57125 3705 57130 4025
rect 57100 3690 57130 3705
rect 57160 4025 57190 4085
rect 57215 4075 57255 4080
rect 57215 4045 57220 4075
rect 57250 4045 57255 4075
rect 57215 4040 57255 4045
rect 57160 3705 57165 4025
rect 57185 3705 57190 4025
rect 57160 3695 57190 3705
rect 57220 4025 57250 4040
rect 57220 3705 57225 4025
rect 57245 3705 57250 4025
rect 57220 3690 57250 3705
rect 57280 4025 57310 4085
rect 57335 4075 57375 4080
rect 57335 4045 57340 4075
rect 57370 4045 57375 4075
rect 57335 4040 57375 4045
rect 57280 3705 57285 4025
rect 57305 3705 57310 4025
rect 57280 3695 57310 3705
rect 57340 4025 57370 4040
rect 57340 3705 57345 4025
rect 57365 3705 57370 4025
rect 57340 3690 57370 3705
rect 57400 4025 57430 4085
rect 57455 4075 57495 4080
rect 57455 4045 57460 4075
rect 57490 4045 57495 4075
rect 57455 4040 57495 4045
rect 57400 3705 57405 4025
rect 57425 3705 57430 4025
rect 57400 3695 57430 3705
rect 57460 4025 57490 4040
rect 57460 3705 57465 4025
rect 57485 3705 57490 4025
rect 57460 3690 57490 3705
rect 57520 4025 57550 4085
rect 57575 4075 57615 4080
rect 57575 4045 57580 4075
rect 57610 4045 57615 4075
rect 57575 4040 57615 4045
rect 57520 3705 57525 4025
rect 57545 3705 57550 4025
rect 57520 3695 57550 3705
rect 57580 4025 57610 4040
rect 57580 3705 57585 4025
rect 57605 3705 57610 4025
rect 57580 3690 57610 3705
rect 57640 4025 57670 4085
rect 57695 4075 57735 4080
rect 57695 4045 57700 4075
rect 57730 4045 57735 4075
rect 57695 4040 57735 4045
rect 57640 3705 57645 4025
rect 57665 3705 57670 4025
rect 57640 3695 57670 3705
rect 57700 4025 57730 4040
rect 57700 3705 57705 4025
rect 57725 3705 57730 4025
rect 57700 3690 57730 3705
rect 57760 4025 57790 4085
rect 57760 3705 57765 4025
rect 57785 3705 57790 4025
rect 57040 3645 57045 3665
rect 57065 3645 57070 3665
rect 57095 3685 57135 3690
rect 57095 3655 57100 3685
rect 57130 3655 57135 3685
rect 57095 3650 57135 3655
rect 57215 3685 57255 3690
rect 57215 3655 57220 3685
rect 57250 3655 57255 3685
rect 57215 3650 57255 3655
rect 57335 3685 57375 3690
rect 57335 3655 57340 3685
rect 57370 3655 57375 3685
rect 57335 3650 57375 3655
rect 57455 3685 57495 3690
rect 57455 3655 57460 3685
rect 57490 3655 57495 3685
rect 57455 3650 57495 3655
rect 57575 3685 57615 3690
rect 57575 3655 57580 3685
rect 57610 3655 57615 3685
rect 57575 3650 57615 3655
rect 57695 3685 57735 3690
rect 57695 3655 57700 3685
rect 57730 3655 57735 3685
rect 57695 3650 57735 3655
rect 57760 3665 57790 3705
rect 57860 3690 57880 4085
rect 57040 3635 57070 3645
rect 57395 3605 57435 3610
rect 57395 3575 57400 3605
rect 57430 3575 57435 3605
rect 57395 3570 57435 3575
rect 56925 3560 56965 3565
rect 56925 3530 56930 3560
rect 56960 3530 56965 3560
rect 56925 3525 56965 3530
rect 56275 3380 56315 3385
rect 56275 3350 56280 3380
rect 56310 3350 56315 3380
rect 56275 3345 56315 3350
rect 56385 3380 56425 3385
rect 56385 3350 56390 3380
rect 56420 3350 56425 3380
rect 56385 3345 56425 3350
rect 56495 3380 56535 3385
rect 56495 3350 56500 3380
rect 56530 3350 56535 3380
rect 56495 3345 56535 3350
rect 56605 3380 56645 3385
rect 56605 3350 56610 3380
rect 56640 3350 56645 3380
rect 56605 3345 56645 3350
rect 56715 3380 56755 3385
rect 56715 3350 56720 3380
rect 56750 3350 56755 3380
rect 56715 3345 56755 3350
rect 56825 3380 56865 3385
rect 56825 3350 56830 3380
rect 56860 3350 56865 3380
rect 56825 3345 56865 3350
rect 56935 3380 56975 3385
rect 56935 3350 56940 3380
rect 56970 3350 56975 3380
rect 56935 3345 56975 3350
rect 57045 3380 57085 3385
rect 57045 3350 57050 3380
rect 57080 3350 57085 3380
rect 57045 3345 57085 3350
rect 57155 3380 57195 3385
rect 57155 3350 57160 3380
rect 57190 3350 57195 3380
rect 57155 3345 57195 3350
rect 57265 3380 57305 3385
rect 57265 3350 57270 3380
rect 57300 3350 57305 3380
rect 57265 3345 57305 3350
rect 57375 3380 57415 3385
rect 57375 3350 57380 3380
rect 57410 3350 57415 3380
rect 57375 3345 57415 3350
rect 57485 3380 57525 3385
rect 57485 3350 57490 3380
rect 57520 3350 57525 3380
rect 57485 3345 57525 3350
rect 56065 3325 56105 3330
rect 56065 3295 56070 3325
rect 56100 3295 56105 3325
rect 56065 3290 56105 3295
rect 56280 3240 56310 3345
rect 56330 3335 56370 3340
rect 56330 3305 56335 3335
rect 56365 3305 56370 3335
rect 56330 3300 56370 3305
rect 56280 3220 56285 3240
rect 56305 3220 56310 3240
rect 56280 3180 56310 3220
rect 56335 3240 56365 3300
rect 56335 3220 56340 3240
rect 56360 3220 56365 3240
rect 56335 3205 56365 3220
rect 56390 3240 56420 3345
rect 56440 3290 56480 3295
rect 56440 3260 56445 3290
rect 56475 3260 56480 3290
rect 56440 3255 56480 3260
rect 56390 3220 56395 3240
rect 56415 3220 56420 3240
rect 56390 3210 56420 3220
rect 56445 3240 56475 3255
rect 56445 3220 56450 3240
rect 56470 3220 56475 3240
rect 56280 3160 56285 3180
rect 56305 3160 56310 3180
rect 56330 3200 56370 3205
rect 56330 3170 56335 3200
rect 56365 3170 56370 3200
rect 56330 3165 56370 3170
rect 56390 3180 56420 3190
rect 56280 3150 56310 3160
rect 56390 3160 56395 3180
rect 56415 3160 56420 3180
rect 56390 3150 56420 3160
rect 56445 3135 56475 3220
rect 56500 3240 56530 3345
rect 56550 3335 56590 3340
rect 56550 3305 56555 3335
rect 56585 3305 56590 3335
rect 56550 3300 56590 3305
rect 56500 3220 56505 3240
rect 56525 3220 56530 3240
rect 56500 3210 56530 3220
rect 56555 3240 56585 3300
rect 56555 3220 56560 3240
rect 56580 3220 56585 3240
rect 56555 3205 56585 3220
rect 56610 3240 56640 3345
rect 56660 3290 56700 3295
rect 56660 3260 56665 3290
rect 56695 3260 56700 3290
rect 56660 3255 56700 3260
rect 56610 3220 56615 3240
rect 56635 3220 56640 3240
rect 56610 3210 56640 3220
rect 56665 3240 56695 3255
rect 56665 3220 56670 3240
rect 56690 3220 56695 3240
rect 56550 3200 56590 3205
rect 56550 3170 56555 3200
rect 56585 3170 56590 3200
rect 56550 3165 56590 3170
rect 56665 3135 56695 3220
rect 56720 3240 56750 3345
rect 56770 3335 56810 3340
rect 56770 3305 56775 3335
rect 56805 3305 56810 3335
rect 56770 3300 56810 3305
rect 56720 3220 56725 3240
rect 56745 3220 56750 3240
rect 56720 3210 56750 3220
rect 56775 3240 56805 3300
rect 56775 3220 56780 3240
rect 56800 3220 56805 3240
rect 56775 3205 56805 3220
rect 56830 3240 56860 3345
rect 56880 3290 56920 3295
rect 56880 3260 56885 3290
rect 56915 3260 56920 3290
rect 56880 3255 56920 3260
rect 56830 3220 56835 3240
rect 56855 3220 56860 3240
rect 56830 3210 56860 3220
rect 56885 3240 56915 3255
rect 56885 3220 56890 3240
rect 56910 3220 56915 3240
rect 56770 3200 56810 3205
rect 56770 3170 56775 3200
rect 56805 3170 56810 3200
rect 56770 3165 56810 3170
rect 56830 3180 56860 3190
rect 56830 3160 56835 3180
rect 56855 3160 56860 3180
rect 56830 3150 56860 3160
rect 56440 3130 56490 3135
rect 56440 3100 56445 3130
rect 56475 3100 56490 3130
rect 56440 3095 56490 3100
rect 56660 3130 56700 3135
rect 56660 3100 56665 3130
rect 56695 3100 56700 3130
rect 56660 3095 56700 3100
rect 56470 3030 56490 3095
rect 56140 3025 56180 3030
rect 55940 3020 55980 3025
rect 55940 2990 55945 3020
rect 55975 2990 55980 3020
rect 55940 2985 55980 2990
rect 56040 3020 56070 3025
rect 56140 2995 56145 3025
rect 56175 2995 56180 3025
rect 56140 2990 56180 2995
rect 56250 3025 56290 3030
rect 56250 2995 56255 3025
rect 56285 2995 56290 3025
rect 56250 2990 56290 2995
rect 56360 3025 56400 3030
rect 56360 2995 56365 3025
rect 56395 2995 56400 3025
rect 56360 2990 56400 2995
rect 56470 3025 56510 3030
rect 56470 2995 56475 3025
rect 56505 2995 56510 3025
rect 56470 2990 56510 2995
rect 56580 3025 56620 3030
rect 56580 2995 56585 3025
rect 56615 2995 56620 3025
rect 56580 2990 56620 2995
rect 56690 3020 56720 3025
rect 56040 2985 56070 2990
rect 55760 2745 55800 2750
rect 55760 2715 55765 2745
rect 55795 2715 55800 2745
rect 55760 2710 55800 2715
rect 55715 2590 55755 2595
rect 55715 2560 55720 2590
rect 55750 2560 55755 2590
rect 55715 2555 55755 2560
rect 54295 2545 54335 2550
rect 54295 2515 54300 2545
rect 54330 2515 54335 2545
rect 54295 2510 54335 2515
rect 55450 2545 55490 2550
rect 55450 2515 55455 2545
rect 55485 2515 55490 2545
rect 55450 2510 55490 2515
rect 54245 2450 54285 2455
rect 54245 2420 54250 2450
rect 54280 2420 54285 2450
rect 54245 2415 54285 2420
rect 54255 400 54275 2415
rect 54305 1920 54325 2510
rect 54955 2495 54995 2500
rect 54955 2465 54960 2495
rect 54990 2465 54995 2495
rect 54955 2460 54995 2465
rect 55615 2495 55655 2500
rect 55615 2465 55620 2495
rect 55650 2465 55655 2495
rect 55615 2460 55655 2465
rect 54960 2415 54990 2460
rect 55010 2450 55050 2455
rect 55010 2420 55015 2450
rect 55045 2420 55050 2450
rect 55010 2415 55050 2420
rect 55120 2450 55160 2455
rect 55120 2420 55125 2450
rect 55155 2420 55160 2450
rect 55120 2415 55160 2420
rect 55230 2450 55270 2455
rect 55230 2420 55235 2450
rect 55265 2420 55270 2450
rect 55230 2415 55270 2420
rect 55340 2450 55380 2455
rect 55340 2420 55345 2450
rect 55375 2420 55380 2450
rect 55340 2415 55380 2420
rect 55450 2450 55490 2455
rect 55450 2420 55455 2450
rect 55485 2420 55490 2450
rect 55450 2415 55490 2420
rect 55560 2450 55600 2455
rect 55560 2420 55565 2450
rect 55595 2420 55600 2450
rect 55560 2415 55600 2420
rect 55620 2415 55650 2460
rect 54960 2395 54965 2415
rect 54985 2395 54990 2415
rect 54960 2355 54990 2395
rect 54960 2185 54965 2355
rect 54985 2185 54990 2355
rect 54960 2175 54990 2185
rect 55015 2355 55045 2415
rect 55065 2405 55105 2410
rect 55065 2375 55070 2405
rect 55100 2375 55105 2405
rect 55065 2370 55105 2375
rect 55015 2185 55020 2355
rect 55040 2185 55045 2355
rect 55015 2175 55045 2185
rect 55070 2355 55100 2370
rect 55070 2185 55075 2355
rect 55095 2185 55100 2355
rect 55070 2155 55100 2185
rect 55125 2355 55155 2415
rect 55175 2405 55215 2410
rect 55175 2375 55180 2405
rect 55210 2375 55215 2405
rect 55175 2370 55215 2375
rect 55125 2185 55130 2355
rect 55150 2185 55155 2355
rect 55125 2175 55155 2185
rect 55180 2355 55210 2370
rect 55180 2185 55185 2355
rect 55205 2185 55210 2355
rect 55180 2155 55210 2185
rect 55235 2355 55265 2415
rect 55285 2405 55325 2410
rect 55285 2375 55290 2405
rect 55320 2375 55325 2405
rect 55285 2370 55325 2375
rect 55235 2185 55240 2355
rect 55260 2185 55265 2355
rect 55235 2175 55265 2185
rect 55290 2355 55320 2370
rect 55290 2185 55295 2355
rect 55315 2185 55320 2355
rect 55290 2155 55320 2185
rect 55345 2355 55375 2415
rect 55395 2405 55435 2410
rect 55395 2375 55400 2405
rect 55430 2375 55435 2405
rect 55395 2370 55435 2375
rect 55345 2185 55350 2355
rect 55370 2185 55375 2355
rect 55345 2175 55375 2185
rect 55400 2355 55430 2370
rect 55400 2185 55405 2355
rect 55425 2185 55430 2355
rect 55400 2155 55430 2185
rect 55455 2355 55485 2415
rect 55505 2405 55545 2410
rect 55505 2375 55510 2405
rect 55540 2375 55545 2405
rect 55505 2370 55545 2375
rect 55455 2185 55460 2355
rect 55480 2185 55485 2355
rect 55455 2175 55485 2185
rect 55510 2355 55540 2370
rect 55510 2185 55515 2355
rect 55535 2185 55540 2355
rect 55510 2155 55540 2185
rect 55565 2355 55595 2415
rect 55565 2185 55570 2355
rect 55590 2185 55595 2355
rect 55565 2175 55595 2185
rect 55620 2395 55625 2415
rect 55645 2395 55650 2415
rect 55620 2355 55650 2395
rect 55620 2185 55625 2355
rect 55645 2185 55650 2355
rect 55620 2175 55650 2185
rect 54760 2150 54800 2155
rect 54760 2120 54765 2150
rect 54795 2120 54800 2150
rect 54760 2115 54800 2120
rect 55065 2150 55105 2155
rect 55065 2120 55070 2150
rect 55100 2120 55105 2150
rect 55065 2115 55105 2120
rect 55175 2150 55215 2155
rect 55175 2120 55180 2150
rect 55210 2120 55215 2150
rect 55175 2115 55215 2120
rect 55285 2150 55325 2155
rect 55285 2120 55290 2150
rect 55320 2120 55325 2150
rect 55285 2115 55325 2120
rect 55395 2150 55435 2155
rect 55395 2120 55400 2150
rect 55430 2120 55435 2150
rect 55395 2115 55435 2120
rect 55505 2150 55545 2155
rect 55505 2120 55510 2150
rect 55540 2120 55545 2150
rect 55505 2115 55545 2120
rect 54290 1910 54340 1920
rect 54290 1880 54300 1910
rect 54330 1880 54340 1910
rect 54290 1870 54340 1880
rect 54305 1260 54325 1870
rect 54450 1595 54485 1600
rect 54450 1555 54485 1560
rect 54510 1595 54545 1600
rect 54510 1555 54545 1560
rect 54570 1595 54605 1600
rect 54570 1555 54605 1560
rect 54630 1595 54665 1600
rect 54630 1555 54665 1560
rect 54460 1425 54480 1555
rect 54580 1540 54600 1555
rect 54770 1540 54790 2115
rect 55725 2060 55745 2555
rect 55770 2500 55790 2710
rect 55760 2495 55800 2500
rect 55760 2465 55765 2495
rect 55795 2465 55800 2495
rect 55760 2460 55800 2465
rect 55450 2055 55490 2060
rect 55450 2025 55455 2055
rect 55485 2025 55490 2055
rect 55450 2020 55490 2025
rect 55715 2055 55755 2060
rect 55715 2025 55720 2055
rect 55750 2025 55755 2055
rect 55715 2020 55755 2025
rect 54805 1945 54845 1950
rect 54805 1915 54810 1945
rect 54840 1915 54845 1945
rect 54805 1910 54845 1915
rect 55065 1945 55105 1950
rect 55065 1915 55070 1945
rect 55100 1915 55105 1945
rect 55065 1910 55105 1915
rect 55175 1945 55215 1950
rect 55175 1915 55180 1945
rect 55210 1915 55215 1945
rect 55175 1910 55215 1915
rect 55285 1945 55325 1950
rect 55285 1915 55290 1945
rect 55320 1915 55325 1945
rect 55285 1910 55325 1915
rect 55395 1945 55435 1950
rect 55395 1915 55400 1945
rect 55430 1915 55435 1945
rect 55395 1910 55435 1915
rect 55505 1945 55545 1950
rect 55505 1915 55510 1945
rect 55540 1915 55545 1945
rect 55505 1910 55545 1915
rect 54815 1595 54835 1910
rect 54960 1895 54990 1905
rect 54960 1625 54965 1895
rect 54985 1625 54990 1895
rect 54805 1590 54845 1595
rect 54805 1560 54810 1590
rect 54840 1560 54845 1590
rect 54805 1555 54845 1560
rect 54960 1585 54990 1625
rect 54960 1565 54965 1585
rect 54985 1565 54990 1585
rect 55015 1895 55045 1905
rect 55015 1625 55020 1895
rect 55040 1625 55045 1895
rect 55015 1565 55045 1625
rect 55070 1895 55100 1910
rect 55070 1625 55075 1895
rect 55095 1625 55100 1895
rect 55070 1610 55100 1625
rect 55125 1895 55155 1905
rect 55125 1625 55130 1895
rect 55150 1625 55155 1895
rect 55065 1605 55105 1610
rect 55065 1575 55070 1605
rect 55100 1575 55105 1605
rect 55065 1570 55105 1575
rect 55125 1565 55155 1625
rect 55180 1895 55210 1910
rect 55180 1625 55185 1895
rect 55205 1625 55210 1895
rect 55180 1610 55210 1625
rect 55235 1895 55265 1905
rect 55235 1625 55240 1895
rect 55260 1625 55265 1895
rect 55175 1605 55215 1610
rect 55175 1575 55180 1605
rect 55210 1575 55215 1605
rect 55175 1570 55215 1575
rect 55235 1565 55265 1625
rect 55290 1895 55320 1910
rect 55290 1625 55295 1895
rect 55315 1625 55320 1895
rect 55290 1610 55320 1625
rect 55345 1895 55375 1905
rect 55345 1625 55350 1895
rect 55370 1625 55375 1895
rect 55285 1605 55325 1610
rect 55285 1575 55290 1605
rect 55320 1575 55325 1605
rect 55285 1570 55325 1575
rect 55345 1565 55375 1625
rect 55400 1895 55430 1910
rect 55400 1625 55405 1895
rect 55425 1625 55430 1895
rect 55400 1610 55430 1625
rect 55455 1895 55485 1905
rect 55455 1625 55460 1895
rect 55480 1625 55485 1895
rect 55395 1605 55435 1610
rect 55395 1575 55400 1605
rect 55430 1575 55435 1605
rect 55395 1570 55435 1575
rect 55455 1565 55485 1625
rect 55510 1895 55540 1910
rect 55510 1625 55515 1895
rect 55535 1625 55540 1895
rect 55510 1610 55540 1625
rect 55565 1895 55595 1905
rect 55565 1625 55570 1895
rect 55590 1625 55595 1895
rect 55505 1605 55545 1610
rect 55505 1575 55510 1605
rect 55540 1575 55545 1605
rect 55505 1570 55545 1575
rect 55565 1565 55595 1625
rect 55620 1895 55650 1905
rect 55620 1625 55625 1895
rect 55645 1625 55650 1895
rect 55620 1585 55650 1625
rect 55620 1565 55625 1585
rect 55645 1565 55650 1585
rect 55770 1565 55790 2460
rect 55830 2270 55870 2275
rect 55830 2240 55835 2270
rect 55865 2240 55870 2270
rect 55830 2235 55870 2240
rect 54570 1535 54610 1540
rect 54570 1505 54575 1535
rect 54605 1505 54610 1535
rect 54570 1500 54610 1505
rect 54760 1535 54800 1540
rect 54760 1505 54765 1535
rect 54795 1505 54800 1535
rect 54760 1500 54800 1505
rect 54960 1470 54990 1565
rect 55010 1560 55050 1565
rect 55010 1530 55015 1560
rect 55045 1530 55050 1560
rect 55010 1525 55050 1530
rect 55120 1560 55160 1565
rect 55120 1530 55125 1560
rect 55155 1530 55160 1560
rect 55120 1525 55160 1530
rect 55230 1560 55270 1565
rect 55230 1530 55235 1560
rect 55265 1530 55270 1560
rect 55230 1525 55270 1530
rect 55340 1560 55380 1565
rect 55340 1530 55345 1560
rect 55375 1530 55380 1560
rect 55340 1525 55380 1530
rect 55450 1560 55490 1565
rect 55450 1530 55455 1560
rect 55485 1530 55490 1560
rect 55450 1525 55490 1530
rect 55560 1560 55600 1565
rect 55560 1530 55565 1560
rect 55595 1530 55600 1560
rect 55560 1525 55600 1530
rect 55620 1470 55650 1565
rect 55760 1560 55800 1565
rect 55760 1530 55765 1560
rect 55795 1530 55800 1560
rect 55760 1525 55800 1530
rect 54955 1465 54995 1470
rect 54955 1435 54960 1465
rect 54990 1435 54995 1465
rect 54955 1430 54995 1435
rect 55615 1465 55655 1470
rect 55615 1435 55620 1465
rect 55650 1435 55655 1465
rect 55615 1430 55655 1435
rect 55785 1465 55825 1470
rect 55785 1435 55790 1465
rect 55820 1435 55825 1465
rect 55785 1430 55825 1435
rect 54450 1420 54490 1425
rect 54450 1390 54455 1420
rect 54485 1390 54490 1420
rect 54450 1385 54490 1390
rect 54705 1325 54745 1330
rect 54705 1295 54710 1325
rect 54740 1295 54745 1325
rect 54705 1290 54745 1295
rect 55385 1325 55425 1330
rect 55385 1295 55390 1325
rect 55420 1295 55425 1325
rect 54295 1255 54335 1260
rect 54295 1225 54300 1255
rect 54330 1225 54335 1255
rect 54295 1220 54335 1225
rect 54715 1200 54735 1290
rect 55385 1265 55425 1295
rect 54770 1255 54810 1260
rect 54770 1225 54775 1255
rect 54805 1225 54810 1255
rect 54770 1220 54810 1225
rect 55085 1255 55125 1260
rect 55085 1225 55090 1255
rect 55120 1225 55125 1255
rect 55085 1220 55125 1225
rect 55285 1255 55325 1260
rect 55285 1225 55290 1255
rect 55320 1225 55325 1255
rect 55385 1245 55395 1265
rect 55415 1245 55425 1265
rect 55385 1235 55425 1245
rect 55485 1255 55525 1260
rect 55285 1220 55325 1225
rect 55485 1225 55490 1255
rect 55520 1225 55525 1255
rect 55485 1220 55525 1225
rect 54780 1200 54800 1220
rect 54990 1205 55020 1215
rect 54710 1195 54745 1200
rect 54710 1155 54745 1160
rect 54770 1195 54805 1200
rect 54770 1155 54805 1160
rect 54990 535 54995 1205
rect 55015 535 55020 1205
rect 54990 495 55020 535
rect 55090 1205 55120 1220
rect 55090 535 55095 1205
rect 55115 535 55120 1205
rect 55090 520 55120 535
rect 55190 1205 55220 1215
rect 55190 535 55195 1205
rect 55215 535 55220 1205
rect 54990 475 54995 495
rect 55015 475 55020 495
rect 55085 515 55125 520
rect 55085 485 55090 515
rect 55120 485 55125 515
rect 55085 480 55125 485
rect 54990 400 55020 475
rect 55190 400 55220 535
rect 55290 1205 55320 1220
rect 55290 535 55295 1205
rect 55315 535 55320 1205
rect 55290 520 55320 535
rect 55390 1205 55420 1215
rect 55390 535 55395 1205
rect 55415 535 55420 1205
rect 55285 515 55325 520
rect 55285 485 55290 515
rect 55320 485 55325 515
rect 55285 480 55325 485
rect 55390 400 55420 535
rect 55490 1205 55520 1220
rect 55490 535 55495 1205
rect 55515 535 55520 1205
rect 55490 520 55520 535
rect 55590 1205 55620 1215
rect 55590 535 55595 1205
rect 55615 535 55620 1205
rect 55795 895 55815 1430
rect 55785 890 55825 895
rect 55785 860 55790 890
rect 55820 860 55825 890
rect 55785 855 55825 860
rect 55485 515 55525 520
rect 55485 485 55490 515
rect 55520 485 55525 515
rect 55485 480 55525 485
rect 55590 495 55620 535
rect 55590 475 55595 495
rect 55615 475 55620 495
rect 55590 400 55620 475
rect 55795 400 55815 855
rect 55840 750 55860 2235
rect 55950 1425 55970 2985
rect 56085 2980 56125 2985
rect 56085 2950 56090 2980
rect 56120 2950 56125 2980
rect 56085 2945 56125 2950
rect 56035 2930 56065 2940
rect 56035 2910 56040 2930
rect 56060 2910 56065 2930
rect 56035 2870 56065 2910
rect 56035 2850 56040 2870
rect 56060 2850 56065 2870
rect 56090 2930 56120 2945
rect 56090 2910 56095 2930
rect 56115 2910 56120 2930
rect 56090 2850 56120 2910
rect 56145 2930 56175 2990
rect 56195 2980 56235 2985
rect 56195 2950 56200 2980
rect 56230 2950 56235 2980
rect 56195 2945 56235 2950
rect 56145 2910 56150 2930
rect 56170 2910 56175 2930
rect 56145 2895 56175 2910
rect 56200 2930 56230 2945
rect 56200 2910 56205 2930
rect 56225 2910 56230 2930
rect 56140 2890 56180 2895
rect 56140 2860 56145 2890
rect 56175 2860 56180 2890
rect 56140 2855 56180 2860
rect 56200 2850 56230 2910
rect 56255 2930 56285 2990
rect 56305 2980 56345 2985
rect 56305 2950 56310 2980
rect 56340 2950 56345 2980
rect 56305 2945 56345 2950
rect 56255 2910 56260 2930
rect 56280 2910 56285 2930
rect 56255 2895 56285 2910
rect 56310 2930 56340 2945
rect 56310 2910 56315 2930
rect 56335 2910 56340 2930
rect 56250 2890 56290 2895
rect 56250 2860 56255 2890
rect 56285 2860 56290 2890
rect 56250 2855 56290 2860
rect 56310 2850 56340 2910
rect 56365 2930 56395 2990
rect 56415 2980 56455 2985
rect 56415 2950 56420 2980
rect 56450 2950 56455 2980
rect 56415 2945 56455 2950
rect 56365 2910 56370 2930
rect 56390 2910 56395 2930
rect 56365 2895 56395 2910
rect 56420 2930 56450 2945
rect 56420 2910 56425 2930
rect 56445 2910 56450 2930
rect 56360 2890 56400 2895
rect 56360 2860 56365 2890
rect 56395 2860 56400 2890
rect 56360 2855 56400 2860
rect 56420 2850 56450 2910
rect 56475 2930 56505 2990
rect 56525 2980 56565 2985
rect 56525 2950 56530 2980
rect 56560 2950 56565 2980
rect 56525 2945 56565 2950
rect 56475 2910 56480 2930
rect 56500 2910 56505 2930
rect 56475 2895 56505 2910
rect 56530 2930 56560 2945
rect 56530 2910 56535 2930
rect 56555 2910 56560 2930
rect 56470 2890 56510 2895
rect 56470 2860 56475 2890
rect 56505 2860 56510 2890
rect 56470 2855 56510 2860
rect 56530 2850 56560 2910
rect 56585 2930 56615 2990
rect 56690 2985 56720 2990
rect 56635 2980 56675 2985
rect 56635 2950 56640 2980
rect 56670 2950 56675 2980
rect 56635 2945 56675 2950
rect 56585 2910 56590 2930
rect 56610 2910 56615 2930
rect 56585 2895 56615 2910
rect 56640 2930 56670 2945
rect 56640 2910 56645 2930
rect 56665 2910 56670 2930
rect 56580 2890 56620 2895
rect 56580 2860 56585 2890
rect 56615 2860 56620 2890
rect 56580 2855 56620 2860
rect 56640 2850 56670 2910
rect 56695 2930 56725 2940
rect 56695 2910 56700 2930
rect 56720 2910 56725 2930
rect 56695 2870 56725 2910
rect 56695 2850 56700 2870
rect 56720 2850 56725 2870
rect 56835 2850 56855 3150
rect 56885 3135 56915 3220
rect 56940 3240 56970 3345
rect 56990 3335 57030 3340
rect 56990 3305 56995 3335
rect 57025 3305 57030 3335
rect 56990 3300 57030 3305
rect 56940 3220 56945 3240
rect 56965 3220 56970 3240
rect 56940 3210 56970 3220
rect 56995 3240 57025 3300
rect 56995 3220 57000 3240
rect 57020 3220 57025 3240
rect 56995 3205 57025 3220
rect 57050 3240 57080 3345
rect 57100 3290 57140 3295
rect 57100 3260 57105 3290
rect 57135 3260 57140 3290
rect 57100 3255 57140 3260
rect 57050 3220 57055 3240
rect 57075 3220 57080 3240
rect 57050 3210 57080 3220
rect 57105 3240 57135 3255
rect 57105 3220 57110 3240
rect 57130 3220 57135 3240
rect 56990 3200 57030 3205
rect 56990 3170 56995 3200
rect 57025 3170 57030 3200
rect 56990 3165 57030 3170
rect 57105 3135 57135 3220
rect 57160 3240 57190 3345
rect 57210 3335 57250 3340
rect 57210 3305 57215 3335
rect 57245 3305 57250 3335
rect 57210 3300 57250 3305
rect 57160 3220 57165 3240
rect 57185 3220 57190 3240
rect 57160 3210 57190 3220
rect 57215 3240 57245 3300
rect 57215 3220 57220 3240
rect 57240 3220 57245 3240
rect 57215 3205 57245 3220
rect 57270 3240 57300 3345
rect 57320 3290 57360 3295
rect 57320 3260 57325 3290
rect 57355 3260 57360 3290
rect 57320 3255 57360 3260
rect 57270 3220 57275 3240
rect 57295 3220 57300 3240
rect 57270 3210 57300 3220
rect 57325 3240 57355 3255
rect 57325 3220 57330 3240
rect 57350 3220 57355 3240
rect 57210 3200 57250 3205
rect 57210 3170 57215 3200
rect 57245 3170 57250 3200
rect 57210 3165 57250 3170
rect 56880 3130 56920 3135
rect 56880 3100 56885 3130
rect 56915 3100 56920 3130
rect 56880 3095 56920 3100
rect 57100 3130 57140 3135
rect 57100 3100 57105 3130
rect 57135 3100 57140 3130
rect 57100 3095 57140 3100
rect 57220 3030 57240 3165
rect 57325 3135 57355 3220
rect 57380 3240 57410 3345
rect 57430 3335 57470 3340
rect 57430 3305 57435 3335
rect 57465 3305 57470 3335
rect 57430 3300 57470 3305
rect 57380 3220 57385 3240
rect 57405 3220 57410 3240
rect 57380 3210 57410 3220
rect 57435 3240 57465 3300
rect 57435 3220 57440 3240
rect 57460 3220 57465 3240
rect 57435 3205 57465 3220
rect 57490 3240 57520 3345
rect 57705 3330 57725 3650
rect 57760 3645 57765 3665
rect 57785 3645 57790 3665
rect 57850 3685 57890 3690
rect 57850 3655 57855 3685
rect 57885 3655 57890 3685
rect 57850 3650 57890 3655
rect 57760 3635 57790 3645
rect 58015 3385 58035 4165
rect 58490 4125 58510 4165
rect 58120 4120 58160 4125
rect 58120 4090 58125 4120
rect 58155 4090 58160 4120
rect 58120 4085 58160 4090
rect 58240 4120 58280 4125
rect 58240 4090 58245 4120
rect 58275 4090 58280 4120
rect 58240 4085 58280 4090
rect 58360 4120 58400 4125
rect 58360 4090 58365 4120
rect 58395 4090 58400 4120
rect 58360 4085 58400 4090
rect 58480 4120 58520 4125
rect 58480 4090 58485 4120
rect 58515 4090 58520 4120
rect 58480 4085 58520 4090
rect 58600 4120 58640 4125
rect 58600 4090 58605 4120
rect 58635 4090 58640 4120
rect 58600 4085 58640 4090
rect 58720 4120 58760 4125
rect 58720 4090 58725 4120
rect 58755 4090 58760 4120
rect 58720 4085 58760 4090
rect 58840 4120 58880 4125
rect 58840 4090 58845 4120
rect 58875 4090 58880 4120
rect 58840 4085 58880 4090
rect 58125 4025 58155 4085
rect 58180 4075 58220 4080
rect 58180 4045 58185 4075
rect 58215 4045 58220 4075
rect 58180 4040 58220 4045
rect 58125 3705 58130 4025
rect 58150 3705 58155 4025
rect 58125 3665 58155 3705
rect 58185 4025 58215 4040
rect 58185 3705 58190 4025
rect 58210 3705 58215 4025
rect 58185 3690 58215 3705
rect 58245 4025 58275 4085
rect 58300 4075 58340 4080
rect 58300 4045 58305 4075
rect 58335 4045 58340 4075
rect 58300 4040 58340 4045
rect 58245 3705 58250 4025
rect 58270 3705 58275 4025
rect 58245 3695 58275 3705
rect 58305 4025 58335 4040
rect 58305 3705 58310 4025
rect 58330 3705 58335 4025
rect 58305 3690 58335 3705
rect 58365 4025 58395 4085
rect 58420 4075 58460 4080
rect 58420 4045 58425 4075
rect 58455 4045 58460 4075
rect 58420 4040 58460 4045
rect 58365 3705 58370 4025
rect 58390 3705 58395 4025
rect 58365 3695 58395 3705
rect 58425 4025 58455 4040
rect 58425 3705 58430 4025
rect 58450 3705 58455 4025
rect 58425 3690 58455 3705
rect 58485 4025 58515 4085
rect 58540 4075 58580 4080
rect 58540 4045 58545 4075
rect 58575 4045 58580 4075
rect 58540 4040 58580 4045
rect 58485 3705 58490 4025
rect 58510 3705 58515 4025
rect 58485 3695 58515 3705
rect 58545 4025 58575 4040
rect 58545 3705 58550 4025
rect 58570 3705 58575 4025
rect 58545 3690 58575 3705
rect 58605 4025 58635 4085
rect 58660 4075 58700 4080
rect 58660 4045 58665 4075
rect 58695 4045 58700 4075
rect 58660 4040 58700 4045
rect 58605 3705 58610 4025
rect 58630 3705 58635 4025
rect 58605 3695 58635 3705
rect 58665 4025 58695 4040
rect 58665 3705 58670 4025
rect 58690 3705 58695 4025
rect 58665 3690 58695 3705
rect 58725 4025 58755 4085
rect 58780 4075 58820 4080
rect 58780 4045 58785 4075
rect 58815 4045 58820 4075
rect 58780 4040 58820 4045
rect 58725 3705 58730 4025
rect 58750 3705 58755 4025
rect 58725 3695 58755 3705
rect 58785 4025 58815 4040
rect 58785 3705 58790 4025
rect 58810 3705 58815 4025
rect 58785 3690 58815 3705
rect 58845 4025 58875 4085
rect 58845 3705 58850 4025
rect 58870 3705 58875 4025
rect 58125 3645 58130 3665
rect 58150 3645 58155 3665
rect 58180 3685 58220 3690
rect 58180 3655 58185 3685
rect 58215 3655 58220 3685
rect 58180 3650 58220 3655
rect 58300 3685 58340 3690
rect 58300 3655 58305 3685
rect 58335 3655 58340 3685
rect 58300 3650 58340 3655
rect 58420 3685 58460 3690
rect 58420 3655 58425 3685
rect 58455 3655 58460 3685
rect 58420 3650 58460 3655
rect 58540 3685 58580 3690
rect 58540 3655 58545 3685
rect 58575 3655 58580 3685
rect 58540 3650 58580 3655
rect 58660 3685 58700 3690
rect 58660 3655 58665 3685
rect 58695 3655 58700 3685
rect 58660 3650 58700 3655
rect 58780 3685 58820 3690
rect 58780 3655 58785 3685
rect 58815 3655 58820 3685
rect 58780 3650 58820 3655
rect 58845 3665 58875 3705
rect 58125 3635 58155 3645
rect 58845 3645 58850 3665
rect 58870 3645 58875 3665
rect 58845 3635 58875 3645
rect 58480 3560 58520 3565
rect 58480 3530 58485 3560
rect 58515 3530 58520 3560
rect 58480 3525 58520 3530
rect 59155 3400 59195 3405
rect 58005 3380 58045 3385
rect 58005 3350 58010 3380
rect 58040 3350 58045 3380
rect 58005 3345 58045 3350
rect 58150 3380 58190 3385
rect 58150 3350 58155 3380
rect 58185 3350 58190 3380
rect 58150 3345 58190 3350
rect 58260 3380 58300 3385
rect 58260 3350 58265 3380
rect 58295 3350 58300 3380
rect 58260 3345 58300 3350
rect 58370 3380 58410 3385
rect 58370 3350 58375 3380
rect 58405 3350 58410 3380
rect 58370 3345 58410 3350
rect 58480 3380 58520 3385
rect 58480 3350 58485 3380
rect 58515 3350 58520 3380
rect 58480 3345 58520 3350
rect 58590 3380 58630 3385
rect 58590 3350 58595 3380
rect 58625 3350 58630 3380
rect 58590 3345 58630 3350
rect 58700 3380 58740 3385
rect 58700 3350 58705 3380
rect 58735 3350 58740 3380
rect 58700 3345 58740 3350
rect 58810 3380 58850 3385
rect 58810 3350 58815 3380
rect 58845 3350 58850 3380
rect 59155 3370 59160 3400
rect 59190 3370 59195 3400
rect 59155 3365 59195 3370
rect 58810 3345 58850 3350
rect 57695 3325 57735 3330
rect 57695 3295 57700 3325
rect 57730 3295 57735 3325
rect 57695 3290 57735 3295
rect 57490 3220 57495 3240
rect 57515 3220 57520 3240
rect 57430 3200 57470 3205
rect 57430 3170 57435 3200
rect 57465 3170 57470 3200
rect 57430 3165 57470 3170
rect 57490 3180 57520 3220
rect 57490 3160 57495 3180
rect 57515 3160 57520 3180
rect 57490 3150 57520 3160
rect 57320 3130 57360 3135
rect 57320 3100 57325 3130
rect 57355 3100 57360 3130
rect 57320 3095 57360 3100
rect 57180 3025 57240 3030
rect 57080 3020 57110 3025
rect 57180 2995 57185 3025
rect 57215 2995 57240 3025
rect 57180 2990 57240 2995
rect 57290 3025 57330 3030
rect 57290 2995 57295 3025
rect 57325 2995 57330 3025
rect 57290 2990 57330 2995
rect 57400 3025 57440 3030
rect 57400 2995 57405 3025
rect 57435 2995 57440 3025
rect 57400 2990 57440 2995
rect 57510 3025 57550 3030
rect 57510 2995 57515 3025
rect 57545 2995 57550 3025
rect 57510 2990 57550 2995
rect 57620 3025 57660 3030
rect 57620 2995 57625 3025
rect 57655 2995 57660 3025
rect 57620 2990 57660 2995
rect 57730 3020 57760 3025
rect 57080 2985 57110 2990
rect 57125 2980 57165 2985
rect 57125 2950 57130 2980
rect 57160 2950 57165 2980
rect 57125 2945 57165 2950
rect 57075 2930 57105 2940
rect 57075 2910 57080 2930
rect 57100 2910 57105 2930
rect 57075 2870 57105 2910
rect 57075 2850 57080 2870
rect 57100 2850 57105 2870
rect 57130 2930 57160 2945
rect 57130 2910 57135 2930
rect 57155 2910 57160 2930
rect 57130 2850 57160 2910
rect 57185 2930 57215 2990
rect 57185 2910 57190 2930
rect 57210 2910 57215 2930
rect 57185 2895 57215 2910
rect 57240 2930 57270 2940
rect 57240 2910 57245 2930
rect 57265 2910 57270 2930
rect 57180 2890 57220 2895
rect 57180 2860 57185 2890
rect 57215 2860 57220 2890
rect 57180 2855 57220 2860
rect 56035 2750 56065 2850
rect 56085 2845 56125 2850
rect 56085 2815 56090 2845
rect 56120 2815 56125 2845
rect 56085 2810 56125 2815
rect 56195 2845 56235 2850
rect 56195 2815 56200 2845
rect 56230 2815 56235 2845
rect 56195 2810 56235 2815
rect 56305 2845 56345 2850
rect 56305 2815 56310 2845
rect 56340 2815 56345 2845
rect 56305 2810 56345 2815
rect 56415 2845 56455 2850
rect 56415 2815 56420 2845
rect 56450 2815 56455 2845
rect 56415 2810 56455 2815
rect 56525 2845 56565 2850
rect 56525 2815 56530 2845
rect 56560 2815 56565 2845
rect 56525 2810 56565 2815
rect 56635 2845 56675 2850
rect 56635 2815 56640 2845
rect 56670 2815 56675 2845
rect 56635 2810 56675 2815
rect 56095 2790 56125 2795
rect 56095 2755 56125 2760
rect 56580 2790 56610 2795
rect 56580 2755 56610 2760
rect 56695 2750 56725 2850
rect 56825 2845 56865 2850
rect 56825 2815 56830 2845
rect 56860 2815 56865 2845
rect 56825 2810 56865 2815
rect 57075 2750 57105 2850
rect 57125 2845 57165 2850
rect 57125 2815 57130 2845
rect 57160 2815 57165 2845
rect 57125 2810 57165 2815
rect 57190 2790 57220 2795
rect 57190 2755 57220 2760
rect 56030 2745 56070 2750
rect 56030 2715 56035 2745
rect 56065 2715 56070 2745
rect 56030 2710 56070 2715
rect 56690 2745 56730 2750
rect 56690 2715 56695 2745
rect 56725 2715 56730 2745
rect 56690 2710 56730 2715
rect 57070 2745 57110 2750
rect 57070 2715 57075 2745
rect 57105 2715 57110 2745
rect 57070 2710 57110 2715
rect 57240 2695 57270 2910
rect 57295 2930 57325 2990
rect 57345 2980 57385 2985
rect 57345 2950 57350 2980
rect 57380 2950 57385 2980
rect 57345 2945 57385 2950
rect 57295 2910 57300 2930
rect 57320 2910 57325 2930
rect 57295 2895 57325 2910
rect 57350 2930 57380 2945
rect 57350 2910 57355 2930
rect 57375 2910 57380 2930
rect 57290 2890 57330 2895
rect 57290 2860 57295 2890
rect 57325 2860 57330 2890
rect 57290 2855 57330 2860
rect 57350 2850 57380 2910
rect 57405 2930 57435 2990
rect 57405 2910 57410 2930
rect 57430 2910 57435 2930
rect 57405 2895 57435 2910
rect 57460 2930 57490 2940
rect 57460 2910 57465 2930
rect 57485 2910 57490 2930
rect 57400 2890 57440 2895
rect 57400 2860 57405 2890
rect 57435 2860 57440 2890
rect 57400 2855 57440 2860
rect 57345 2845 57385 2850
rect 57345 2815 57350 2845
rect 57380 2815 57385 2845
rect 57345 2810 57385 2815
rect 56605 2690 56645 2695
rect 56605 2660 56610 2690
rect 56640 2660 56645 2690
rect 56605 2655 56645 2660
rect 56825 2690 56865 2695
rect 56825 2660 56830 2690
rect 56860 2660 56865 2690
rect 56825 2655 56865 2660
rect 57045 2690 57085 2695
rect 57045 2660 57050 2690
rect 57080 2660 57085 2690
rect 57045 2655 57085 2660
rect 57235 2690 57275 2695
rect 57235 2660 57240 2690
rect 57270 2660 57275 2690
rect 57235 2655 57275 2660
rect 56305 2590 56345 2595
rect 56305 2560 56310 2590
rect 56340 2560 56345 2590
rect 56305 2555 56345 2560
rect 56555 2570 56585 2580
rect 56095 2270 56125 2275
rect 56095 2235 56125 2240
rect 56140 2260 56180 2265
rect 56140 2230 56145 2260
rect 56175 2230 56180 2260
rect 56140 2225 56180 2230
rect 56250 2260 56290 2265
rect 56250 2230 56255 2260
rect 56285 2230 56290 2260
rect 56250 2225 56290 2230
rect 56085 2215 56125 2220
rect 56085 2185 56090 2215
rect 56120 2185 56125 2215
rect 56085 2180 56125 2185
rect 56030 2165 56065 2175
rect 56030 2045 56040 2165
rect 56060 2045 56065 2165
rect 56030 2035 56065 2045
rect 56035 2030 56065 2035
rect 56090 2165 56120 2180
rect 56090 2045 56095 2165
rect 56115 2045 56120 2165
rect 56035 2005 56065 2015
rect 56035 1985 56040 2005
rect 56060 1985 56065 2005
rect 56090 1985 56120 2045
rect 56145 2165 56175 2225
rect 56195 2215 56235 2220
rect 56195 2185 56200 2215
rect 56230 2185 56235 2215
rect 56195 2180 56235 2185
rect 56145 2045 56150 2165
rect 56170 2045 56175 2165
rect 56145 2030 56175 2045
rect 56200 2165 56230 2180
rect 56200 2045 56205 2165
rect 56225 2045 56230 2165
rect 56140 2025 56180 2030
rect 56140 1995 56145 2025
rect 56175 1995 56180 2025
rect 56140 1990 56180 1995
rect 56200 1985 56230 2045
rect 56255 2165 56285 2225
rect 56315 2220 56335 2555
rect 56555 2550 56560 2570
rect 56580 2550 56585 2570
rect 56555 2520 56585 2550
rect 56610 2570 56640 2655
rect 56715 2635 56755 2640
rect 56715 2605 56720 2635
rect 56750 2605 56755 2635
rect 56715 2600 56755 2605
rect 56610 2550 56615 2570
rect 56635 2550 56640 2570
rect 56550 2515 56590 2520
rect 56550 2485 56555 2515
rect 56585 2485 56590 2515
rect 56550 2480 56590 2485
rect 56610 2465 56640 2550
rect 56665 2570 56695 2580
rect 56665 2550 56670 2570
rect 56690 2550 56695 2570
rect 56665 2520 56695 2550
rect 56720 2570 56750 2600
rect 56720 2550 56725 2570
rect 56745 2550 56750 2570
rect 56660 2515 56700 2520
rect 56660 2485 56665 2515
rect 56695 2485 56700 2515
rect 56660 2480 56700 2485
rect 56605 2460 56645 2465
rect 56605 2430 56610 2460
rect 56640 2430 56645 2460
rect 56605 2425 56645 2430
rect 56720 2420 56750 2550
rect 56775 2570 56805 2580
rect 56775 2550 56780 2570
rect 56800 2550 56805 2570
rect 56775 2520 56805 2550
rect 56830 2570 56860 2655
rect 56935 2635 56975 2640
rect 56935 2605 56940 2635
rect 56970 2605 56975 2635
rect 56935 2600 56975 2605
rect 56830 2550 56835 2570
rect 56855 2550 56860 2570
rect 56770 2515 56810 2520
rect 56770 2485 56775 2515
rect 56805 2485 56810 2515
rect 56770 2480 56810 2485
rect 56830 2465 56860 2550
rect 56885 2570 56915 2580
rect 56885 2550 56890 2570
rect 56910 2550 56915 2570
rect 56885 2520 56915 2550
rect 56940 2570 56970 2600
rect 56940 2550 56945 2570
rect 56965 2550 56970 2570
rect 56880 2515 56920 2520
rect 56880 2485 56885 2515
rect 56915 2485 56920 2515
rect 56880 2480 56920 2485
rect 56825 2460 56865 2465
rect 56825 2430 56830 2460
rect 56860 2430 56865 2460
rect 56825 2425 56865 2430
rect 56940 2420 56970 2550
rect 56995 2570 57025 2580
rect 56995 2550 57000 2570
rect 57020 2550 57025 2570
rect 56995 2520 57025 2550
rect 57050 2570 57080 2655
rect 57350 2640 57380 2810
rect 57460 2695 57490 2910
rect 57515 2930 57545 2990
rect 57565 2980 57605 2985
rect 57565 2950 57570 2980
rect 57600 2950 57605 2980
rect 57565 2945 57605 2950
rect 57515 2910 57520 2930
rect 57540 2910 57545 2930
rect 57515 2895 57545 2910
rect 57570 2930 57600 2945
rect 57570 2910 57575 2930
rect 57595 2910 57600 2930
rect 57510 2890 57550 2895
rect 57510 2860 57515 2890
rect 57545 2860 57550 2890
rect 57510 2855 57550 2860
rect 57570 2850 57600 2910
rect 57625 2930 57655 2990
rect 57730 2985 57760 2990
rect 57820 3020 57860 3025
rect 57820 2990 57825 3020
rect 57855 2990 57860 3020
rect 57820 2985 57860 2990
rect 57625 2910 57630 2930
rect 57650 2910 57655 2930
rect 57625 2895 57655 2910
rect 57680 2930 57710 2940
rect 57680 2910 57685 2930
rect 57705 2910 57710 2930
rect 57620 2890 57660 2895
rect 57620 2860 57625 2890
rect 57655 2860 57660 2890
rect 57620 2855 57660 2860
rect 57565 2845 57605 2850
rect 57565 2815 57570 2845
rect 57600 2815 57605 2845
rect 57565 2810 57605 2815
rect 57680 2695 57710 2910
rect 57735 2930 57765 2940
rect 57735 2910 57740 2930
rect 57760 2910 57765 2930
rect 57735 2870 57765 2910
rect 57735 2850 57740 2870
rect 57760 2850 57765 2870
rect 57735 2750 57765 2850
rect 57730 2745 57770 2750
rect 57730 2715 57735 2745
rect 57765 2715 57770 2745
rect 57730 2710 57770 2715
rect 57455 2690 57495 2695
rect 57455 2660 57460 2690
rect 57490 2660 57495 2690
rect 57455 2655 57495 2660
rect 57675 2690 57715 2695
rect 57675 2660 57680 2690
rect 57710 2660 57715 2690
rect 57675 2655 57715 2660
rect 57155 2635 57195 2640
rect 57155 2605 57160 2635
rect 57190 2605 57195 2635
rect 57155 2600 57195 2605
rect 57345 2635 57385 2640
rect 57345 2605 57350 2635
rect 57380 2605 57385 2635
rect 57345 2600 57385 2605
rect 57050 2550 57055 2570
rect 57075 2550 57080 2570
rect 56990 2515 57030 2520
rect 56990 2485 56995 2515
rect 57025 2485 57030 2515
rect 56990 2480 57030 2485
rect 57050 2465 57080 2550
rect 57105 2570 57135 2580
rect 57105 2550 57110 2570
rect 57130 2550 57135 2570
rect 57105 2520 57135 2550
rect 57160 2570 57190 2600
rect 57455 2590 57495 2595
rect 57160 2550 57165 2570
rect 57185 2550 57190 2570
rect 57100 2515 57140 2520
rect 57100 2485 57105 2515
rect 57135 2485 57140 2515
rect 57100 2480 57140 2485
rect 57045 2460 57085 2465
rect 57045 2430 57050 2460
rect 57080 2430 57085 2460
rect 57045 2425 57085 2430
rect 57160 2420 57190 2550
rect 57215 2570 57245 2580
rect 57215 2550 57220 2570
rect 57240 2550 57245 2570
rect 57455 2560 57460 2590
rect 57490 2560 57495 2590
rect 57455 2555 57495 2560
rect 57215 2520 57245 2550
rect 57210 2515 57250 2520
rect 57210 2485 57215 2515
rect 57245 2485 57250 2515
rect 57210 2480 57250 2485
rect 56715 2415 56755 2420
rect 56715 2385 56720 2415
rect 56750 2385 56755 2415
rect 56715 2380 56755 2385
rect 56935 2415 56975 2420
rect 56935 2385 56940 2415
rect 56970 2385 56975 2415
rect 56935 2380 56975 2385
rect 57155 2415 57195 2420
rect 57155 2385 57160 2415
rect 57190 2385 57195 2415
rect 57155 2380 57195 2385
rect 56635 2270 56665 2275
rect 56360 2260 56400 2265
rect 56360 2230 56365 2260
rect 56395 2230 56400 2260
rect 56360 2225 56400 2230
rect 56470 2260 56510 2265
rect 56470 2230 56475 2260
rect 56505 2230 56510 2260
rect 56470 2225 56510 2230
rect 56580 2260 56620 2265
rect 56580 2230 56585 2260
rect 56615 2230 56620 2260
rect 56635 2235 56665 2240
rect 57135 2270 57165 2275
rect 57135 2235 57165 2240
rect 57180 2260 57220 2265
rect 56580 2225 56620 2230
rect 57180 2230 57185 2260
rect 57215 2230 57220 2260
rect 57180 2225 57220 2230
rect 57290 2260 57330 2265
rect 57290 2230 57295 2260
rect 57325 2230 57330 2260
rect 57290 2225 57330 2230
rect 57400 2260 57440 2265
rect 57400 2230 57405 2260
rect 57435 2230 57440 2260
rect 57400 2225 57440 2230
rect 56305 2215 56345 2220
rect 56305 2185 56310 2215
rect 56340 2185 56345 2215
rect 56305 2180 56345 2185
rect 56255 2045 56260 2165
rect 56280 2045 56285 2165
rect 56255 2030 56285 2045
rect 56310 2165 56340 2180
rect 56310 2045 56315 2165
rect 56335 2045 56340 2165
rect 56250 2025 56290 2030
rect 56250 1995 56255 2025
rect 56285 1995 56290 2025
rect 56250 1990 56290 1995
rect 56310 1985 56340 2045
rect 56365 2165 56395 2225
rect 56415 2215 56455 2220
rect 56415 2185 56420 2215
rect 56450 2185 56455 2215
rect 56415 2180 56455 2185
rect 56365 2045 56370 2165
rect 56390 2045 56395 2165
rect 56365 2030 56395 2045
rect 56420 2165 56450 2180
rect 56420 2045 56425 2165
rect 56445 2045 56450 2165
rect 56360 2025 56400 2030
rect 56360 1995 56365 2025
rect 56395 1995 56400 2025
rect 56360 1990 56400 1995
rect 56035 1940 56065 1985
rect 56085 1980 56125 1985
rect 56085 1950 56090 1980
rect 56120 1950 56125 1980
rect 56085 1945 56125 1950
rect 56195 1980 56235 1985
rect 56195 1950 56200 1980
rect 56230 1950 56235 1980
rect 56195 1945 56235 1950
rect 56305 1980 56345 1985
rect 56305 1950 56310 1980
rect 56340 1950 56345 1980
rect 56305 1945 56345 1950
rect 56030 1935 56070 1940
rect 56030 1905 56035 1935
rect 56065 1905 56070 1935
rect 56030 1900 56070 1905
rect 56370 1810 56390 1990
rect 56420 1985 56450 2045
rect 56475 2165 56505 2225
rect 56525 2215 56565 2220
rect 56525 2185 56530 2215
rect 56560 2185 56565 2215
rect 56525 2180 56565 2185
rect 56475 2045 56480 2165
rect 56500 2045 56505 2165
rect 56475 2030 56505 2045
rect 56530 2165 56560 2180
rect 56530 2045 56535 2165
rect 56555 2045 56560 2165
rect 56470 2025 56510 2030
rect 56470 1995 56475 2025
rect 56505 1995 56510 2025
rect 56470 1990 56510 1995
rect 56530 1985 56560 2045
rect 56585 2165 56615 2225
rect 56635 2215 56675 2220
rect 56635 2185 56640 2215
rect 56670 2185 56675 2215
rect 56635 2180 56675 2185
rect 57125 2215 57165 2220
rect 57125 2185 57130 2215
rect 57160 2185 57165 2215
rect 57125 2180 57165 2185
rect 56585 2045 56590 2165
rect 56610 2045 56615 2165
rect 56585 2030 56615 2045
rect 56640 2165 56670 2180
rect 56640 2045 56645 2165
rect 56665 2045 56670 2165
rect 56580 2025 56620 2030
rect 56580 1995 56585 2025
rect 56615 1995 56620 2025
rect 56580 1990 56620 1995
rect 56640 1985 56670 2045
rect 56695 2165 56765 2175
rect 56695 2045 56700 2165
rect 56720 2045 56765 2165
rect 56695 2035 56765 2045
rect 57035 2165 57105 2175
rect 57035 2045 57080 2165
rect 57100 2045 57105 2165
rect 57035 2035 57105 2045
rect 56695 2005 56725 2035
rect 56695 1985 56700 2005
rect 56720 1985 56725 2005
rect 56415 1980 56455 1985
rect 56415 1950 56420 1980
rect 56450 1950 56455 1980
rect 56415 1945 56455 1950
rect 56525 1980 56565 1985
rect 56525 1950 56530 1980
rect 56560 1950 56565 1980
rect 56525 1945 56565 1950
rect 56635 1980 56675 1985
rect 56635 1950 56640 1980
rect 56670 1950 56675 1980
rect 56635 1945 56675 1950
rect 56695 1940 56725 1985
rect 57075 2005 57105 2035
rect 57075 1985 57080 2005
rect 57100 1985 57105 2005
rect 57130 2165 57160 2180
rect 57130 2045 57135 2165
rect 57155 2045 57160 2165
rect 57130 1985 57160 2045
rect 57185 2165 57215 2225
rect 57235 2215 57275 2220
rect 57235 2185 57240 2215
rect 57270 2185 57275 2215
rect 57235 2180 57275 2185
rect 57185 2045 57190 2165
rect 57210 2045 57215 2165
rect 57185 2030 57215 2045
rect 57240 2165 57270 2180
rect 57240 2045 57245 2165
rect 57265 2045 57270 2165
rect 57180 2025 57220 2030
rect 57180 1995 57185 2025
rect 57215 1995 57220 2025
rect 57180 1990 57220 1995
rect 57240 1985 57270 2045
rect 57295 2165 57325 2225
rect 57345 2215 57385 2220
rect 57345 2185 57350 2215
rect 57380 2185 57385 2215
rect 57345 2180 57385 2185
rect 57295 2045 57300 2165
rect 57320 2045 57325 2165
rect 57295 2030 57325 2045
rect 57350 2165 57380 2180
rect 57350 2045 57355 2165
rect 57375 2045 57380 2165
rect 57290 2025 57330 2030
rect 57290 1995 57295 2025
rect 57325 1995 57330 2025
rect 57290 1990 57330 1995
rect 57350 1985 57380 2045
rect 57405 2165 57435 2225
rect 57465 2220 57485 2555
rect 57510 2260 57550 2265
rect 57510 2230 57515 2260
rect 57545 2230 57550 2260
rect 57510 2225 57550 2230
rect 57620 2260 57660 2265
rect 57620 2230 57625 2260
rect 57655 2230 57660 2260
rect 57620 2225 57660 2230
rect 57455 2215 57495 2220
rect 57455 2185 57460 2215
rect 57490 2185 57495 2215
rect 57455 2180 57495 2185
rect 57405 2045 57410 2165
rect 57430 2045 57435 2165
rect 57405 2030 57435 2045
rect 57460 2165 57490 2180
rect 57460 2045 57465 2165
rect 57485 2045 57490 2165
rect 57400 2025 57440 2030
rect 57400 1995 57405 2025
rect 57435 1995 57440 2025
rect 57400 1990 57440 1995
rect 57075 1940 57105 1985
rect 57125 1980 57165 1985
rect 57125 1950 57130 1980
rect 57160 1950 57165 1980
rect 57125 1945 57165 1950
rect 57235 1980 57275 1985
rect 57235 1950 57240 1980
rect 57270 1950 57275 1980
rect 57235 1945 57275 1950
rect 57345 1980 57385 1985
rect 57345 1950 57350 1980
rect 57380 1950 57385 1980
rect 57345 1945 57385 1950
rect 56690 1935 56730 1940
rect 56690 1905 56695 1935
rect 56725 1905 56730 1935
rect 56690 1900 56730 1905
rect 57070 1935 57110 1940
rect 57070 1905 57075 1935
rect 57105 1905 57110 1935
rect 57070 1900 57110 1905
rect 56365 1805 56395 1810
rect 56085 1795 56125 1800
rect 56040 1785 56070 1790
rect 56085 1765 56090 1795
rect 56120 1765 56125 1795
rect 56085 1760 56125 1765
rect 56195 1795 56235 1800
rect 56195 1765 56200 1795
rect 56230 1765 56235 1795
rect 56195 1760 56235 1765
rect 56305 1795 56345 1800
rect 56305 1765 56310 1795
rect 56340 1765 56345 1795
rect 56365 1770 56395 1775
rect 56415 1795 56455 1800
rect 56305 1760 56345 1765
rect 56415 1765 56420 1795
rect 56450 1765 56455 1795
rect 56415 1760 56455 1765
rect 56525 1795 56565 1800
rect 56525 1765 56530 1795
rect 56560 1765 56565 1795
rect 56525 1760 56565 1765
rect 56635 1795 56675 1800
rect 56635 1765 56640 1795
rect 56670 1765 56675 1795
rect 56635 1760 56675 1765
rect 56690 1785 56720 1790
rect 56040 1750 56070 1755
rect 56035 1695 56065 1705
rect 56035 1575 56040 1695
rect 56060 1575 56065 1695
rect 56035 1565 56065 1575
rect 56090 1695 56120 1760
rect 56140 1750 56180 1755
rect 56140 1720 56145 1750
rect 56175 1720 56180 1750
rect 56140 1715 56180 1720
rect 56090 1575 56095 1695
rect 56115 1575 56120 1695
rect 56090 1560 56120 1575
rect 56145 1695 56175 1715
rect 56145 1575 56150 1695
rect 56170 1575 56175 1695
rect 56085 1555 56125 1560
rect 56035 1535 56065 1545
rect 56035 1515 56040 1535
rect 56060 1515 56065 1535
rect 56085 1525 56090 1555
rect 56120 1525 56125 1555
rect 56085 1520 56125 1525
rect 56145 1515 56175 1575
rect 56200 1695 56230 1760
rect 56250 1750 56290 1755
rect 56250 1720 56255 1750
rect 56285 1720 56290 1750
rect 56250 1715 56290 1720
rect 56200 1575 56205 1695
rect 56225 1575 56230 1695
rect 56200 1560 56230 1575
rect 56255 1695 56285 1715
rect 56255 1575 56260 1695
rect 56280 1575 56285 1695
rect 56195 1555 56235 1560
rect 56195 1525 56200 1555
rect 56230 1525 56235 1555
rect 56195 1520 56235 1525
rect 56255 1515 56285 1575
rect 56310 1695 56340 1760
rect 56360 1750 56400 1755
rect 56360 1720 56365 1750
rect 56395 1720 56400 1750
rect 56360 1715 56400 1720
rect 56310 1575 56315 1695
rect 56335 1575 56340 1695
rect 56310 1560 56340 1575
rect 56365 1695 56395 1715
rect 56365 1575 56370 1695
rect 56390 1575 56395 1695
rect 56305 1555 56345 1560
rect 56305 1525 56310 1555
rect 56340 1525 56345 1555
rect 56305 1520 56345 1525
rect 56365 1515 56395 1575
rect 56420 1695 56450 1760
rect 56470 1750 56510 1755
rect 56470 1720 56475 1750
rect 56505 1720 56510 1750
rect 56470 1715 56510 1720
rect 56420 1575 56425 1695
rect 56445 1575 56450 1695
rect 56420 1560 56450 1575
rect 56475 1695 56505 1715
rect 56475 1575 56480 1695
rect 56500 1575 56505 1695
rect 56415 1555 56455 1560
rect 56415 1525 56420 1555
rect 56450 1525 56455 1555
rect 56415 1520 56455 1525
rect 56475 1515 56505 1575
rect 56530 1695 56560 1760
rect 56580 1750 56620 1755
rect 56580 1720 56585 1750
rect 56615 1720 56620 1750
rect 56580 1715 56620 1720
rect 56530 1575 56535 1695
rect 56555 1575 56560 1695
rect 56530 1560 56560 1575
rect 56585 1695 56615 1715
rect 56585 1575 56590 1695
rect 56610 1575 56615 1695
rect 56525 1555 56565 1560
rect 56525 1525 56530 1555
rect 56560 1525 56565 1555
rect 56525 1520 56565 1525
rect 56585 1515 56615 1575
rect 56640 1695 56670 1760
rect 56690 1750 56720 1755
rect 56850 1785 56880 1790
rect 56850 1750 56880 1755
rect 56903 1785 56933 1790
rect 56903 1750 56933 1755
rect 56950 1705 56970 1855
rect 57410 1810 57430 1990
rect 57460 1985 57490 2045
rect 57515 2165 57545 2225
rect 57565 2215 57605 2220
rect 57565 2185 57570 2215
rect 57600 2185 57605 2215
rect 57565 2180 57605 2185
rect 57515 2045 57520 2165
rect 57540 2045 57545 2165
rect 57515 2030 57545 2045
rect 57570 2165 57600 2180
rect 57570 2045 57575 2165
rect 57595 2045 57600 2165
rect 57510 2025 57550 2030
rect 57510 1995 57515 2025
rect 57545 1995 57550 2025
rect 57510 1990 57550 1995
rect 57570 1985 57600 2045
rect 57625 2165 57655 2225
rect 57675 2215 57715 2220
rect 57675 2185 57680 2215
rect 57710 2185 57715 2215
rect 57675 2180 57715 2185
rect 57625 2045 57630 2165
rect 57650 2045 57655 2165
rect 57625 2030 57655 2045
rect 57680 2165 57710 2180
rect 57680 2045 57685 2165
rect 57705 2045 57710 2165
rect 57620 2025 57660 2030
rect 57620 1995 57625 2025
rect 57655 1995 57660 2025
rect 57620 1990 57660 1995
rect 57680 1985 57710 2045
rect 57735 2165 57765 2175
rect 57735 2045 57740 2165
rect 57760 2045 57765 2165
rect 57735 2035 57765 2045
rect 57735 2005 57765 2015
rect 57735 1985 57740 2005
rect 57760 1985 57765 2005
rect 57455 1980 57495 1985
rect 57455 1950 57460 1980
rect 57490 1950 57495 1980
rect 57455 1945 57495 1950
rect 57565 1980 57605 1985
rect 57565 1950 57570 1980
rect 57600 1950 57605 1980
rect 57565 1945 57605 1950
rect 57675 1980 57715 1985
rect 57675 1950 57680 1980
rect 57710 1950 57715 1980
rect 57675 1945 57715 1950
rect 57735 1940 57765 1985
rect 57730 1935 57770 1940
rect 57730 1905 57735 1935
rect 57765 1905 57770 1935
rect 57730 1900 57770 1905
rect 57405 1805 57435 1810
rect 57125 1795 57165 1800
rect 57080 1785 57110 1790
rect 57125 1765 57130 1795
rect 57160 1765 57165 1795
rect 57125 1760 57165 1765
rect 57235 1795 57275 1800
rect 57235 1765 57240 1795
rect 57270 1765 57275 1795
rect 57235 1760 57275 1765
rect 57345 1795 57385 1800
rect 57345 1765 57350 1795
rect 57380 1765 57385 1795
rect 57405 1770 57435 1775
rect 57455 1795 57495 1800
rect 57345 1760 57385 1765
rect 57455 1765 57460 1795
rect 57490 1765 57495 1795
rect 57455 1760 57495 1765
rect 57565 1795 57605 1800
rect 57565 1765 57570 1795
rect 57600 1765 57605 1795
rect 57565 1760 57605 1765
rect 57675 1795 57715 1800
rect 57675 1765 57680 1795
rect 57710 1765 57715 1795
rect 57675 1760 57715 1765
rect 57730 1785 57760 1790
rect 57080 1750 57110 1755
rect 56640 1575 56645 1695
rect 56665 1575 56670 1695
rect 56640 1560 56670 1575
rect 56695 1695 56805 1705
rect 56695 1575 56700 1695
rect 56720 1575 56780 1695
rect 56800 1575 56805 1695
rect 56695 1565 56805 1575
rect 56830 1695 56860 1705
rect 56830 1575 56835 1695
rect 56855 1575 56860 1695
rect 56830 1565 56860 1575
rect 56885 1695 56915 1705
rect 56885 1575 56890 1695
rect 56910 1575 56915 1695
rect 56885 1565 56915 1575
rect 56940 1695 56970 1705
rect 56940 1575 56945 1695
rect 56965 1575 56970 1695
rect 56940 1565 56970 1575
rect 56995 1695 57105 1705
rect 56995 1575 57000 1695
rect 57020 1575 57080 1695
rect 57100 1575 57105 1695
rect 56995 1565 57105 1575
rect 57130 1695 57160 1760
rect 57180 1750 57220 1755
rect 57180 1720 57185 1750
rect 57215 1720 57220 1750
rect 57180 1715 57220 1720
rect 57130 1575 57135 1695
rect 57155 1575 57160 1695
rect 56635 1555 56675 1560
rect 56635 1525 56640 1555
rect 56670 1525 56675 1555
rect 56740 1545 56760 1565
rect 56635 1520 56675 1525
rect 56735 1535 56765 1545
rect 56735 1515 56740 1535
rect 56760 1515 56765 1535
rect 56035 1505 56065 1515
rect 56140 1510 56180 1515
rect 56040 1470 56060 1505
rect 56140 1480 56145 1510
rect 56175 1480 56180 1510
rect 56140 1475 56180 1480
rect 56250 1510 56290 1515
rect 56250 1480 56255 1510
rect 56285 1480 56290 1510
rect 56250 1475 56290 1480
rect 56360 1510 56400 1515
rect 56360 1480 56365 1510
rect 56395 1480 56400 1510
rect 56360 1475 56400 1480
rect 56470 1510 56510 1515
rect 56470 1480 56475 1510
rect 56505 1480 56510 1510
rect 56470 1475 56510 1480
rect 56580 1510 56620 1515
rect 56580 1480 56585 1510
rect 56615 1480 56620 1510
rect 56735 1505 56765 1515
rect 56580 1475 56620 1480
rect 56740 1470 56760 1505
rect 56030 1465 56070 1470
rect 56030 1435 56035 1465
rect 56065 1435 56070 1465
rect 56030 1430 56070 1435
rect 56730 1465 56770 1470
rect 56730 1435 56735 1465
rect 56765 1435 56770 1465
rect 56730 1430 56770 1435
rect 56835 1425 56855 1565
rect 55940 1420 55980 1425
rect 55940 1390 55945 1420
rect 55975 1390 55980 1420
rect 55940 1385 55980 1390
rect 56825 1420 56865 1425
rect 56825 1390 56830 1420
rect 56860 1390 56865 1420
rect 56825 1385 56865 1390
rect 56330 1265 56370 1270
rect 56330 1235 56335 1265
rect 56365 1235 56370 1265
rect 56330 1230 56370 1235
rect 56185 1145 56255 1155
rect 56185 925 56230 1145
rect 56250 925 56255 1145
rect 56185 915 56255 925
rect 56225 895 56255 915
rect 56280 1145 56310 1155
rect 56280 925 56285 1145
rect 56305 925 56310 1145
rect 56280 895 56310 925
rect 56335 1145 56365 1230
rect 56835 1215 56855 1385
rect 56890 1270 56910 1565
rect 56945 1425 56965 1565
rect 57040 1545 57060 1565
rect 57130 1560 57160 1575
rect 57185 1695 57215 1715
rect 57185 1575 57190 1695
rect 57210 1575 57215 1695
rect 57125 1555 57165 1560
rect 57035 1535 57065 1545
rect 57035 1515 57040 1535
rect 57060 1515 57065 1535
rect 57125 1525 57130 1555
rect 57160 1525 57165 1555
rect 57125 1520 57165 1525
rect 57185 1515 57215 1575
rect 57240 1695 57270 1760
rect 57290 1750 57330 1755
rect 57290 1720 57295 1750
rect 57325 1720 57330 1750
rect 57290 1715 57330 1720
rect 57240 1575 57245 1695
rect 57265 1575 57270 1695
rect 57240 1560 57270 1575
rect 57295 1695 57325 1715
rect 57295 1575 57300 1695
rect 57320 1575 57325 1695
rect 57235 1555 57275 1560
rect 57235 1525 57240 1555
rect 57270 1525 57275 1555
rect 57235 1520 57275 1525
rect 57295 1515 57325 1575
rect 57350 1695 57380 1760
rect 57400 1750 57440 1755
rect 57400 1720 57405 1750
rect 57435 1720 57440 1750
rect 57400 1715 57440 1720
rect 57350 1575 57355 1695
rect 57375 1575 57380 1695
rect 57350 1560 57380 1575
rect 57405 1695 57435 1715
rect 57405 1575 57410 1695
rect 57430 1575 57435 1695
rect 57345 1555 57385 1560
rect 57345 1525 57350 1555
rect 57380 1525 57385 1555
rect 57345 1520 57385 1525
rect 57405 1515 57435 1575
rect 57460 1695 57490 1760
rect 57510 1750 57550 1755
rect 57510 1720 57515 1750
rect 57545 1720 57550 1750
rect 57510 1715 57550 1720
rect 57460 1575 57465 1695
rect 57485 1575 57490 1695
rect 57460 1560 57490 1575
rect 57515 1695 57545 1715
rect 57515 1575 57520 1695
rect 57540 1575 57545 1695
rect 57455 1555 57495 1560
rect 57455 1525 57460 1555
rect 57490 1525 57495 1555
rect 57455 1520 57495 1525
rect 57515 1515 57545 1575
rect 57570 1695 57600 1760
rect 57620 1750 57660 1755
rect 57620 1720 57625 1750
rect 57655 1720 57660 1750
rect 57620 1715 57660 1720
rect 57570 1575 57575 1695
rect 57595 1575 57600 1695
rect 57570 1560 57600 1575
rect 57625 1695 57655 1715
rect 57625 1575 57630 1695
rect 57650 1575 57655 1695
rect 57565 1555 57605 1560
rect 57565 1525 57570 1555
rect 57600 1525 57605 1555
rect 57565 1520 57605 1525
rect 57625 1515 57655 1575
rect 57680 1695 57710 1760
rect 57730 1750 57760 1755
rect 57680 1575 57685 1695
rect 57705 1575 57710 1695
rect 57680 1560 57710 1575
rect 57735 1695 57765 1705
rect 57735 1575 57740 1695
rect 57760 1575 57765 1695
rect 57735 1565 57765 1575
rect 57675 1555 57715 1560
rect 57675 1525 57680 1555
rect 57710 1525 57715 1555
rect 57675 1520 57715 1525
rect 57735 1535 57765 1545
rect 57735 1515 57740 1535
rect 57760 1515 57765 1535
rect 57035 1505 57065 1515
rect 57180 1510 57220 1515
rect 57040 1470 57060 1505
rect 57180 1480 57185 1510
rect 57215 1480 57220 1510
rect 57180 1475 57220 1480
rect 57290 1510 57330 1515
rect 57290 1480 57295 1510
rect 57325 1480 57330 1510
rect 57290 1475 57330 1480
rect 57400 1510 57440 1515
rect 57400 1480 57405 1510
rect 57435 1480 57440 1510
rect 57400 1475 57440 1480
rect 57510 1510 57550 1515
rect 57510 1480 57515 1510
rect 57545 1480 57550 1510
rect 57510 1475 57550 1480
rect 57620 1510 57660 1515
rect 57620 1480 57625 1510
rect 57655 1480 57660 1510
rect 57735 1505 57765 1515
rect 57620 1475 57660 1480
rect 57030 1465 57070 1470
rect 57030 1435 57035 1465
rect 57065 1435 57070 1465
rect 57030 1430 57070 1435
rect 56935 1420 56975 1425
rect 56935 1390 56940 1420
rect 56970 1390 56975 1420
rect 56935 1385 56975 1390
rect 56880 1265 56920 1270
rect 56880 1235 56885 1265
rect 56915 1235 56920 1265
rect 56880 1230 56920 1235
rect 57200 1215 57220 1475
rect 57740 1470 57760 1505
rect 57730 1465 57770 1470
rect 57730 1435 57735 1465
rect 57765 1435 57770 1465
rect 57730 1430 57770 1435
rect 57830 1425 57850 2985
rect 58015 2750 58035 3345
rect 58050 3325 58090 3330
rect 58050 3295 58055 3325
rect 58085 3295 58090 3325
rect 58050 3290 58090 3295
rect 58155 3310 58185 3345
rect 58155 3290 58160 3310
rect 58180 3290 58185 3310
rect 58005 2745 58045 2750
rect 58005 2715 58010 2745
rect 58040 2715 58045 2745
rect 58005 2710 58045 2715
rect 57910 2515 57950 2520
rect 57910 2485 57915 2515
rect 57945 2485 57950 2515
rect 58015 2500 58035 2710
rect 58060 2595 58080 3290
rect 58155 3250 58185 3290
rect 58205 3300 58245 3305
rect 58205 3270 58210 3300
rect 58240 3270 58245 3300
rect 58205 3265 58245 3270
rect 58155 2680 58160 3250
rect 58180 2680 58185 3250
rect 58155 2670 58185 2680
rect 58210 3250 58240 3265
rect 58210 2680 58215 3250
rect 58235 2680 58240 3250
rect 58210 2665 58240 2680
rect 58265 3250 58295 3345
rect 58315 3300 58355 3305
rect 58315 3270 58320 3300
rect 58350 3270 58355 3300
rect 58315 3265 58355 3270
rect 58265 2680 58270 3250
rect 58290 2680 58295 3250
rect 58265 2670 58295 2680
rect 58320 3250 58350 3265
rect 58320 2680 58325 3250
rect 58345 2680 58350 3250
rect 58320 2665 58350 2680
rect 58375 3250 58405 3345
rect 58425 3300 58465 3305
rect 58425 3270 58430 3300
rect 58460 3270 58465 3300
rect 58425 3265 58465 3270
rect 58375 2680 58380 3250
rect 58400 2680 58405 3250
rect 58375 2670 58405 2680
rect 58430 3250 58460 3265
rect 58430 2680 58435 3250
rect 58455 2680 58460 3250
rect 58430 2665 58460 2680
rect 58485 3250 58515 3345
rect 58535 3300 58575 3305
rect 58535 3270 58540 3300
rect 58570 3270 58575 3300
rect 58535 3265 58575 3270
rect 58485 2680 58490 3250
rect 58510 2680 58515 3250
rect 58485 2670 58515 2680
rect 58540 3250 58570 3265
rect 58540 2680 58545 3250
rect 58565 2680 58570 3250
rect 58540 2665 58570 2680
rect 58595 3250 58625 3345
rect 58645 3300 58685 3305
rect 58645 3270 58650 3300
rect 58680 3270 58685 3300
rect 58645 3265 58685 3270
rect 58595 2680 58600 3250
rect 58620 2680 58625 3250
rect 58595 2670 58625 2680
rect 58650 3250 58680 3265
rect 58650 2680 58655 3250
rect 58675 2680 58680 3250
rect 58650 2665 58680 2680
rect 58705 3250 58735 3345
rect 58815 3310 58845 3345
rect 59165 3325 59185 3365
rect 58755 3300 58795 3305
rect 58755 3270 58760 3300
rect 58790 3270 58795 3300
rect 58755 3265 58795 3270
rect 58815 3290 58820 3310
rect 58840 3290 58845 3310
rect 58705 2680 58710 3250
rect 58730 2680 58735 3250
rect 58705 2670 58735 2680
rect 58760 3250 58790 3265
rect 58760 2680 58765 3250
rect 58785 2680 58790 3250
rect 58760 2665 58790 2680
rect 58815 3250 58845 3290
rect 59105 3315 59246 3325
rect 59105 3295 59110 3315
rect 59130 3295 59165 3315
rect 59185 3295 59220 3315
rect 59240 3295 59246 3315
rect 59105 3285 59246 3295
rect 58815 2680 58820 3250
rect 58840 2680 58845 3250
rect 59105 2710 59246 2720
rect 59105 2690 59110 2710
rect 59130 2690 59165 2710
rect 59185 2690 59220 2710
rect 59240 2690 59246 2710
rect 59105 2680 59246 2690
rect 58815 2670 58845 2680
rect 58205 2660 58245 2665
rect 58205 2630 58210 2660
rect 58240 2630 58245 2660
rect 58205 2625 58245 2630
rect 58315 2660 58355 2665
rect 58315 2630 58320 2660
rect 58350 2630 58355 2660
rect 58315 2625 58355 2630
rect 58425 2660 58465 2665
rect 58425 2630 58430 2660
rect 58460 2630 58465 2660
rect 58425 2625 58465 2630
rect 58535 2660 58575 2665
rect 58535 2630 58540 2660
rect 58570 2630 58575 2660
rect 58535 2625 58575 2630
rect 58645 2660 58685 2665
rect 58645 2630 58650 2660
rect 58680 2630 58685 2660
rect 58645 2625 58685 2630
rect 58755 2660 58795 2665
rect 58755 2630 58760 2660
rect 58790 2630 58795 2660
rect 58755 2625 58795 2630
rect 58050 2590 58090 2595
rect 58050 2560 58055 2590
rect 58085 2560 58090 2590
rect 58050 2555 58090 2560
rect 57910 2480 57950 2485
rect 58005 2495 58045 2500
rect 57865 2460 57905 2465
rect 57865 2430 57870 2460
rect 57900 2430 57905 2460
rect 57865 2425 57905 2430
rect 57820 1420 57860 1425
rect 57820 1390 57825 1420
rect 57855 1390 57860 1420
rect 57820 1385 57860 1390
rect 57875 1270 57895 2425
rect 57920 1940 57940 2480
rect 58005 2465 58010 2495
rect 58040 2465 58045 2495
rect 58005 2460 58045 2465
rect 57910 1935 57950 1940
rect 57910 1905 57915 1935
rect 57945 1905 57950 1935
rect 57910 1900 57950 1905
rect 57920 1470 57940 1900
rect 58015 1565 58035 2460
rect 58060 2060 58080 2555
rect 58325 2550 58345 2625
rect 59165 2595 59185 2680
rect 59155 2590 59195 2595
rect 58590 2555 58595 2585
rect 58625 2555 58630 2585
rect 59155 2560 59160 2590
rect 59190 2560 59195 2590
rect 59155 2555 59195 2560
rect 58315 2545 58355 2550
rect 58315 2515 58320 2545
rect 58350 2515 58355 2545
rect 58315 2510 58355 2515
rect 59465 2545 59505 2550
rect 59465 2515 59470 2545
rect 59500 2515 59505 2545
rect 59465 2510 59505 2515
rect 58150 2495 58190 2500
rect 58150 2465 58155 2495
rect 58185 2465 58190 2495
rect 58150 2460 58190 2465
rect 58810 2495 58850 2500
rect 58810 2465 58815 2495
rect 58845 2465 58850 2495
rect 58810 2460 58850 2465
rect 58155 2415 58185 2460
rect 58205 2450 58245 2455
rect 58205 2420 58210 2450
rect 58240 2420 58245 2450
rect 58205 2415 58245 2420
rect 58315 2450 58355 2455
rect 58315 2420 58320 2450
rect 58350 2420 58355 2450
rect 58315 2415 58355 2420
rect 58425 2450 58465 2455
rect 58425 2420 58430 2450
rect 58460 2420 58465 2450
rect 58425 2415 58465 2420
rect 58535 2450 58575 2455
rect 58535 2420 58540 2450
rect 58570 2420 58575 2450
rect 58535 2415 58575 2420
rect 58645 2450 58685 2455
rect 58645 2420 58650 2450
rect 58680 2420 58685 2450
rect 58645 2415 58685 2420
rect 58755 2450 58795 2455
rect 58755 2420 58760 2450
rect 58790 2420 58795 2450
rect 58755 2415 58795 2420
rect 58815 2415 58845 2460
rect 58155 2395 58160 2415
rect 58180 2395 58185 2415
rect 58155 2355 58185 2395
rect 58155 2185 58160 2355
rect 58180 2185 58185 2355
rect 58155 2175 58185 2185
rect 58210 2355 58240 2415
rect 58260 2405 58300 2410
rect 58260 2375 58265 2405
rect 58295 2375 58300 2405
rect 58260 2370 58300 2375
rect 58210 2185 58215 2355
rect 58235 2185 58240 2355
rect 58210 2175 58240 2185
rect 58265 2355 58295 2370
rect 58265 2185 58270 2355
rect 58290 2185 58295 2355
rect 58265 2155 58295 2185
rect 58320 2355 58350 2415
rect 58370 2405 58410 2410
rect 58370 2375 58375 2405
rect 58405 2375 58410 2405
rect 58370 2370 58410 2375
rect 58320 2185 58325 2355
rect 58345 2185 58350 2355
rect 58320 2175 58350 2185
rect 58375 2355 58405 2370
rect 58375 2185 58380 2355
rect 58400 2185 58405 2355
rect 58375 2155 58405 2185
rect 58430 2355 58460 2415
rect 58480 2405 58520 2410
rect 58480 2375 58485 2405
rect 58515 2375 58520 2405
rect 58480 2370 58520 2375
rect 58430 2185 58435 2355
rect 58455 2185 58460 2355
rect 58430 2175 58460 2185
rect 58485 2355 58515 2370
rect 58485 2185 58490 2355
rect 58510 2185 58515 2355
rect 58485 2155 58515 2185
rect 58540 2355 58570 2415
rect 58590 2405 58630 2410
rect 58590 2375 58595 2405
rect 58625 2375 58630 2405
rect 58590 2370 58630 2375
rect 58540 2185 58545 2355
rect 58565 2185 58570 2355
rect 58540 2175 58570 2185
rect 58595 2355 58625 2370
rect 58595 2185 58600 2355
rect 58620 2185 58625 2355
rect 58595 2155 58625 2185
rect 58650 2355 58680 2415
rect 58700 2405 58740 2410
rect 58700 2375 58705 2405
rect 58735 2375 58740 2405
rect 58700 2370 58740 2375
rect 58650 2185 58655 2355
rect 58675 2185 58680 2355
rect 58650 2175 58680 2185
rect 58705 2355 58735 2370
rect 58705 2185 58710 2355
rect 58730 2185 58735 2355
rect 58705 2155 58735 2185
rect 58760 2355 58790 2415
rect 58760 2185 58765 2355
rect 58785 2185 58790 2355
rect 58760 2175 58790 2185
rect 58815 2395 58820 2415
rect 58840 2395 58845 2415
rect 58815 2355 58845 2395
rect 58815 2185 58820 2355
rect 58840 2185 58845 2355
rect 58815 2175 58845 2185
rect 58260 2150 58300 2155
rect 58260 2120 58265 2150
rect 58295 2120 58300 2150
rect 58260 2115 58300 2120
rect 58370 2150 58410 2155
rect 58370 2120 58375 2150
rect 58405 2120 58410 2150
rect 58370 2115 58410 2120
rect 58480 2150 58520 2155
rect 58480 2120 58485 2150
rect 58515 2120 58520 2150
rect 58480 2115 58520 2120
rect 58590 2150 58630 2155
rect 58590 2120 58595 2150
rect 58625 2120 58630 2150
rect 58590 2115 58630 2120
rect 58700 2150 58740 2155
rect 58700 2120 58705 2150
rect 58735 2120 58740 2150
rect 58700 2115 58740 2120
rect 59000 2150 59040 2155
rect 59000 2120 59005 2150
rect 59035 2120 59040 2150
rect 59000 2115 59040 2120
rect 58050 2055 58090 2060
rect 58050 2025 58055 2055
rect 58085 2025 58090 2055
rect 58050 2020 58090 2025
rect 58315 2055 58355 2060
rect 58315 2025 58320 2055
rect 58350 2025 58355 2055
rect 58315 2020 58355 2025
rect 58260 1945 58300 1950
rect 58260 1915 58265 1945
rect 58295 1915 58300 1945
rect 58260 1910 58300 1915
rect 58370 1945 58410 1950
rect 58370 1915 58375 1945
rect 58405 1915 58410 1945
rect 58370 1910 58410 1915
rect 58480 1945 58520 1950
rect 58480 1915 58485 1945
rect 58515 1915 58520 1945
rect 58480 1910 58520 1915
rect 58590 1945 58630 1950
rect 58590 1915 58595 1945
rect 58625 1915 58630 1945
rect 58590 1910 58630 1915
rect 58700 1945 58740 1950
rect 58700 1915 58705 1945
rect 58735 1915 58740 1945
rect 58700 1910 58740 1915
rect 58955 1945 58995 1950
rect 58955 1915 58960 1945
rect 58990 1915 58995 1945
rect 58955 1910 58995 1915
rect 58155 1895 58185 1905
rect 58155 1625 58160 1895
rect 58180 1625 58185 1895
rect 58155 1585 58185 1625
rect 58155 1565 58160 1585
rect 58180 1565 58185 1585
rect 58210 1895 58240 1905
rect 58210 1625 58215 1895
rect 58235 1625 58240 1895
rect 58210 1565 58240 1625
rect 58265 1895 58295 1910
rect 58265 1625 58270 1895
rect 58290 1625 58295 1895
rect 58265 1610 58295 1625
rect 58320 1895 58350 1905
rect 58320 1625 58325 1895
rect 58345 1625 58350 1895
rect 58260 1605 58300 1610
rect 58260 1575 58265 1605
rect 58295 1575 58300 1605
rect 58260 1570 58300 1575
rect 58320 1565 58350 1625
rect 58375 1895 58405 1910
rect 58375 1625 58380 1895
rect 58400 1625 58405 1895
rect 58375 1610 58405 1625
rect 58430 1895 58460 1905
rect 58430 1625 58435 1895
rect 58455 1625 58460 1895
rect 58370 1605 58410 1610
rect 58370 1575 58375 1605
rect 58405 1575 58410 1605
rect 58370 1570 58410 1575
rect 58430 1565 58460 1625
rect 58485 1895 58515 1910
rect 58485 1625 58490 1895
rect 58510 1625 58515 1895
rect 58485 1610 58515 1625
rect 58540 1895 58570 1905
rect 58540 1625 58545 1895
rect 58565 1625 58570 1895
rect 58480 1605 58520 1610
rect 58480 1575 58485 1605
rect 58515 1575 58520 1605
rect 58480 1570 58520 1575
rect 58540 1565 58570 1625
rect 58595 1895 58625 1910
rect 58595 1625 58600 1895
rect 58620 1625 58625 1895
rect 58595 1610 58625 1625
rect 58650 1895 58680 1905
rect 58650 1625 58655 1895
rect 58675 1625 58680 1895
rect 58590 1605 58630 1610
rect 58590 1575 58595 1605
rect 58625 1575 58630 1605
rect 58590 1570 58630 1575
rect 58650 1565 58680 1625
rect 58705 1895 58735 1910
rect 58705 1625 58710 1895
rect 58730 1625 58735 1895
rect 58705 1610 58735 1625
rect 58760 1895 58790 1905
rect 58760 1625 58765 1895
rect 58785 1625 58790 1895
rect 58700 1605 58740 1610
rect 58700 1575 58705 1605
rect 58735 1575 58740 1605
rect 58700 1570 58740 1575
rect 58760 1565 58790 1625
rect 58815 1895 58845 1905
rect 58815 1625 58820 1895
rect 58840 1625 58845 1895
rect 58815 1585 58845 1625
rect 58815 1565 58820 1585
rect 58840 1565 58845 1585
rect 58005 1560 58045 1565
rect 58005 1530 58010 1560
rect 58040 1530 58045 1560
rect 58005 1525 58045 1530
rect 58155 1470 58185 1565
rect 58205 1560 58245 1565
rect 58205 1530 58210 1560
rect 58240 1530 58245 1560
rect 58205 1525 58245 1530
rect 58315 1560 58355 1565
rect 58315 1530 58320 1560
rect 58350 1530 58355 1560
rect 58315 1525 58355 1530
rect 58425 1560 58465 1565
rect 58425 1530 58430 1560
rect 58460 1530 58465 1560
rect 58425 1525 58465 1530
rect 58535 1560 58575 1565
rect 58535 1530 58540 1560
rect 58570 1530 58575 1560
rect 58535 1525 58575 1530
rect 58645 1560 58685 1565
rect 58645 1530 58650 1560
rect 58680 1530 58685 1560
rect 58645 1525 58685 1530
rect 58755 1560 58795 1565
rect 58755 1530 58760 1560
rect 58790 1530 58795 1560
rect 58755 1525 58795 1530
rect 58815 1470 58845 1565
rect 58965 1545 58985 1910
rect 58955 1540 58995 1545
rect 58955 1510 58960 1540
rect 58990 1510 58995 1540
rect 58955 1505 58995 1510
rect 59010 1490 59030 2115
rect 59475 1920 59495 2510
rect 59515 2450 59555 2455
rect 59515 2420 59520 2450
rect 59550 2420 59555 2450
rect 59515 2415 59555 2420
rect 59460 1910 59510 1920
rect 59460 1880 59470 1910
rect 59500 1880 59510 1910
rect 59460 1870 59510 1880
rect 59135 1545 59170 1550
rect 59135 1505 59170 1510
rect 59195 1545 59230 1550
rect 59195 1505 59230 1510
rect 59255 1545 59290 1550
rect 59255 1505 59290 1510
rect 59315 1545 59350 1551
rect 59315 1505 59350 1510
rect 59200 1490 59220 1505
rect 59000 1485 59040 1490
rect 57910 1465 57950 1470
rect 57910 1435 57915 1465
rect 57945 1435 57950 1465
rect 57910 1430 57950 1435
rect 58150 1465 58190 1470
rect 58150 1435 58155 1465
rect 58185 1435 58190 1465
rect 58150 1430 58190 1435
rect 58810 1465 58850 1470
rect 58810 1435 58815 1465
rect 58845 1435 58850 1465
rect 59000 1455 59005 1485
rect 59035 1455 59040 1485
rect 59000 1450 59040 1455
rect 59190 1485 59230 1490
rect 59190 1455 59195 1485
rect 59225 1455 59230 1485
rect 59190 1450 59230 1455
rect 58810 1430 58850 1435
rect 57405 1265 57445 1270
rect 57405 1235 57410 1265
rect 57440 1235 57445 1265
rect 57405 1230 57445 1235
rect 57865 1265 57905 1270
rect 57865 1235 57870 1265
rect 57900 1235 57905 1265
rect 57865 1230 57905 1235
rect 56440 1210 56480 1215
rect 56440 1180 56445 1210
rect 56475 1180 56480 1210
rect 56440 1175 56480 1180
rect 56550 1210 56590 1215
rect 56550 1180 56555 1210
rect 56585 1180 56590 1210
rect 56550 1175 56590 1180
rect 56660 1210 56700 1215
rect 56660 1180 56665 1210
rect 56695 1180 56700 1210
rect 56660 1175 56700 1180
rect 56770 1210 56810 1215
rect 56770 1180 56775 1210
rect 56805 1180 56810 1210
rect 56770 1175 56810 1180
rect 56830 1205 56860 1215
rect 56830 1185 56835 1205
rect 56855 1185 56860 1205
rect 56830 1175 56860 1185
rect 56880 1210 56920 1215
rect 56880 1180 56885 1210
rect 56915 1180 56920 1210
rect 56880 1175 56920 1180
rect 56990 1210 57030 1215
rect 56990 1180 56995 1210
rect 57025 1180 57030 1210
rect 56990 1175 57030 1180
rect 57100 1210 57140 1215
rect 57100 1180 57105 1210
rect 57135 1180 57140 1210
rect 57100 1175 57140 1180
rect 57200 1210 57250 1215
rect 57200 1180 57215 1210
rect 57245 1180 57250 1210
rect 57200 1175 57250 1180
rect 57320 1210 57360 1215
rect 57320 1180 57325 1210
rect 57355 1180 57360 1210
rect 57320 1175 57360 1180
rect 57430 1210 57470 1215
rect 57430 1180 57435 1210
rect 57465 1180 57470 1210
rect 57430 1175 57470 1180
rect 56335 925 56340 1145
rect 56360 925 56365 1145
rect 56335 915 56365 925
rect 56390 1145 56420 1155
rect 56390 925 56395 1145
rect 56415 925 56420 1145
rect 56390 895 56420 925
rect 56445 1145 56475 1175
rect 56445 925 56450 1145
rect 56470 925 56475 1145
rect 56220 890 56260 895
rect 56220 860 56225 890
rect 56255 860 56260 890
rect 56220 855 56260 860
rect 56275 890 56315 895
rect 56275 860 56280 890
rect 56310 860 56315 890
rect 56275 855 56315 860
rect 56385 890 56425 895
rect 56385 860 56390 890
rect 56420 860 56425 890
rect 56385 855 56425 860
rect 56445 850 56475 925
rect 56500 1145 56530 1155
rect 56500 925 56505 1145
rect 56525 925 56530 1145
rect 56500 895 56530 925
rect 56555 1145 56585 1175
rect 56555 925 56560 1145
rect 56580 925 56585 1145
rect 56495 890 56535 895
rect 56495 860 56500 890
rect 56530 860 56535 890
rect 56495 855 56535 860
rect 56555 850 56585 925
rect 56610 1145 56640 1155
rect 56610 925 56615 1145
rect 56635 925 56640 1145
rect 56610 895 56640 925
rect 56665 1145 56695 1175
rect 56665 925 56670 1145
rect 56690 925 56695 1145
rect 56605 890 56645 895
rect 56605 860 56610 890
rect 56640 860 56645 890
rect 56605 855 56645 860
rect 56665 850 56695 925
rect 56720 1145 56750 1155
rect 56720 925 56725 1145
rect 56745 925 56750 1145
rect 56720 895 56750 925
rect 56775 1145 56805 1175
rect 56775 925 56780 1145
rect 56800 925 56805 1145
rect 56715 890 56755 895
rect 56715 860 56720 890
rect 56750 860 56755 890
rect 56715 855 56755 860
rect 56775 850 56805 925
rect 56830 1145 56860 1155
rect 56830 925 56835 1145
rect 56855 925 56860 1145
rect 56830 895 56860 925
rect 56885 1145 56915 1175
rect 56885 925 56890 1145
rect 56910 925 56915 1145
rect 56825 890 56865 895
rect 56825 860 56830 890
rect 56860 860 56865 890
rect 56825 855 56865 860
rect 56885 850 56915 925
rect 56940 1145 56970 1155
rect 56940 925 56945 1145
rect 56965 925 56970 1145
rect 56940 895 56970 925
rect 56995 1145 57025 1175
rect 56995 925 57000 1145
rect 57020 925 57025 1145
rect 56935 890 56975 895
rect 56935 860 56940 890
rect 56970 860 56975 890
rect 56935 855 56975 860
rect 56995 850 57025 925
rect 57050 1145 57080 1155
rect 57050 925 57055 1145
rect 57075 925 57080 1145
rect 57050 895 57080 925
rect 57105 1145 57135 1175
rect 57105 925 57110 1145
rect 57130 925 57135 1145
rect 57045 890 57085 895
rect 57045 860 57050 890
rect 57080 860 57085 890
rect 57045 855 57085 860
rect 57105 850 57135 925
rect 57160 1145 57190 1155
rect 57160 925 57165 1145
rect 57185 925 57190 1145
rect 57160 895 57190 925
rect 57215 1145 57245 1175
rect 57215 925 57220 1145
rect 57240 925 57245 1145
rect 57155 890 57195 895
rect 57155 860 57160 890
rect 57190 860 57195 890
rect 57155 855 57195 860
rect 57215 850 57245 925
rect 57270 1145 57300 1155
rect 57270 925 57275 1145
rect 57295 925 57300 1145
rect 57270 895 57300 925
rect 57325 1145 57355 1175
rect 57325 925 57330 1145
rect 57350 925 57355 1145
rect 57265 890 57305 895
rect 57265 860 57270 890
rect 57300 860 57305 890
rect 57265 855 57305 860
rect 57325 850 57355 925
rect 57380 1145 57410 1155
rect 57380 925 57385 1145
rect 57405 925 57410 1145
rect 57380 895 57410 925
rect 57435 1145 57465 1175
rect 57435 925 57440 1145
rect 57460 925 57465 1145
rect 57375 890 57415 895
rect 57375 860 57380 890
rect 57410 860 57415 890
rect 57375 855 57415 860
rect 57435 850 57465 925
rect 57490 1145 57520 1155
rect 57490 925 57495 1145
rect 57515 925 57520 1145
rect 57490 895 57520 925
rect 57485 890 57525 895
rect 57485 860 57490 890
rect 57520 860 57525 890
rect 57920 885 57940 1430
rect 59320 1425 59340 1505
rect 59310 1420 59350 1425
rect 59310 1390 59315 1420
rect 59345 1390 59350 1420
rect 59310 1385 59350 1390
rect 58430 1325 58470 1330
rect 58430 1295 58435 1325
rect 58465 1295 58470 1325
rect 58430 1290 58470 1295
rect 59035 1325 59075 1330
rect 59035 1295 59040 1325
rect 59070 1295 59075 1325
rect 59035 1290 59075 1295
rect 58435 1265 58465 1290
rect 58280 1255 58320 1260
rect 58280 1225 58285 1255
rect 58315 1225 58320 1255
rect 58435 1245 58440 1265
rect 58460 1245 58465 1265
rect 58435 1235 58465 1245
rect 58480 1255 58520 1260
rect 58970 1255 59010 1260
rect 58280 1220 58320 1225
rect 58480 1225 58485 1255
rect 58515 1225 58520 1255
rect 58480 1220 58520 1225
rect 58680 1225 58685 1255
rect 58715 1225 58720 1255
rect 58680 1220 58720 1225
rect 58970 1225 58975 1255
rect 59005 1225 59010 1255
rect 58970 1220 59010 1225
rect 58185 1205 58215 1215
rect 57485 855 57525 860
rect 57910 880 57950 885
rect 57910 850 57915 880
rect 57945 850 57950 880
rect 56440 845 56480 850
rect 56440 815 56445 845
rect 56475 815 56480 845
rect 56440 810 56480 815
rect 56550 845 56590 850
rect 56550 815 56555 845
rect 56585 815 56590 845
rect 56550 810 56590 815
rect 56660 845 56700 850
rect 56660 815 56665 845
rect 56695 815 56700 845
rect 56660 810 56700 815
rect 56770 845 56810 850
rect 56770 815 56775 845
rect 56805 815 56810 845
rect 56770 810 56810 815
rect 56880 845 56920 850
rect 56880 815 56885 845
rect 56915 815 56920 845
rect 56880 810 56920 815
rect 56990 845 57030 850
rect 56990 815 56995 845
rect 57025 815 57030 845
rect 56990 810 57030 815
rect 57100 845 57140 850
rect 57100 815 57105 845
rect 57135 815 57140 845
rect 57100 810 57140 815
rect 57210 845 57250 850
rect 57210 815 57215 845
rect 57245 815 57250 845
rect 57210 810 57250 815
rect 57320 845 57360 850
rect 57320 815 57325 845
rect 57355 815 57360 845
rect 57320 810 57360 815
rect 57430 845 57470 850
rect 57910 845 57950 850
rect 57430 815 57435 845
rect 57465 815 57470 845
rect 57430 810 57470 815
rect 56540 790 56580 795
rect 56540 760 56545 790
rect 56575 760 56580 790
rect 56540 755 56580 760
rect 56650 790 56690 795
rect 56650 760 56655 790
rect 56685 760 56690 790
rect 56650 755 56690 760
rect 56870 790 56910 795
rect 56870 760 56875 790
rect 56905 760 56910 790
rect 56870 755 56910 760
rect 55830 745 55870 750
rect 55830 715 55835 745
rect 55865 715 55870 745
rect 55830 710 55870 715
rect 56485 745 56525 750
rect 56485 715 56490 745
rect 56520 715 56525 745
rect 56485 710 56525 715
rect 56395 680 56465 690
rect 56395 560 56440 680
rect 56460 560 56465 680
rect 56395 550 56465 560
rect 56435 520 56465 550
rect 56435 500 56440 520
rect 56460 500 56465 520
rect 56490 680 56520 710
rect 56490 560 56495 680
rect 56515 560 56520 680
rect 56490 500 56520 560
rect 56545 680 56575 755
rect 56595 745 56635 750
rect 56595 715 56600 745
rect 56630 715 56635 745
rect 56595 710 56635 715
rect 56545 560 56550 680
rect 56570 560 56575 680
rect 56545 545 56575 560
rect 56600 680 56630 710
rect 56600 560 56605 680
rect 56625 560 56630 680
rect 56540 540 56580 545
rect 56540 510 56545 540
rect 56575 510 56580 540
rect 56540 505 56580 510
rect 56600 500 56630 560
rect 56655 680 56685 755
rect 56705 745 56745 750
rect 56705 715 56710 745
rect 56740 715 56745 745
rect 56705 710 56745 715
rect 56655 560 56660 680
rect 56680 560 56685 680
rect 56655 545 56685 560
rect 56710 680 56740 710
rect 56710 560 56715 680
rect 56735 560 56740 680
rect 56650 540 56690 545
rect 56650 510 56655 540
rect 56685 510 56690 540
rect 56650 505 56690 510
rect 56710 500 56740 560
rect 56765 680 56835 690
rect 56765 560 56770 680
rect 56790 560 56835 680
rect 56765 550 56835 560
rect 56875 680 56905 755
rect 57040 745 57080 750
rect 57040 715 57045 745
rect 57075 715 57080 745
rect 57040 710 57080 715
rect 56875 560 56880 680
rect 56900 560 56905 680
rect 56765 520 56795 550
rect 56875 545 56905 560
rect 57215 680 57245 810
rect 57215 560 57220 680
rect 57240 560 57245 680
rect 57215 550 57245 560
rect 56765 500 56770 520
rect 56790 500 56795 520
rect 56870 540 56910 545
rect 56870 510 56875 540
rect 56905 510 56910 540
rect 56870 505 56910 510
rect 56435 400 56465 500
rect 56485 495 56525 500
rect 56485 465 56490 495
rect 56520 465 56525 495
rect 56485 460 56525 465
rect 56595 495 56635 500
rect 56595 465 56600 495
rect 56630 465 56635 495
rect 56595 460 56635 465
rect 56705 495 56745 500
rect 56705 465 56710 495
rect 56740 465 56745 495
rect 56705 460 56745 465
rect 56765 400 56795 500
rect 57920 400 57940 845
rect 58185 535 58190 1205
rect 58210 535 58215 1205
rect 58185 495 58215 535
rect 58285 1205 58315 1220
rect 58285 535 58290 1205
rect 58310 535 58315 1205
rect 58285 520 58315 535
rect 58385 1205 58415 1215
rect 58385 535 58390 1205
rect 58410 535 58415 1205
rect 58185 475 58190 495
rect 58210 475 58215 495
rect 58280 515 58320 520
rect 58280 485 58285 515
rect 58315 485 58320 515
rect 58280 480 58320 485
rect 58185 400 58215 475
rect 58385 400 58415 535
rect 58485 1205 58515 1220
rect 58485 535 58490 1205
rect 58510 535 58515 1205
rect 58485 520 58515 535
rect 58585 1205 58615 1215
rect 58585 535 58590 1205
rect 58610 535 58615 1205
rect 58480 515 58520 520
rect 58480 485 58485 515
rect 58515 485 58520 515
rect 58480 480 58520 485
rect 58585 400 58615 535
rect 58685 1205 58715 1220
rect 58685 535 58690 1205
rect 58710 535 58715 1205
rect 58685 520 58715 535
rect 58785 1205 58815 1215
rect 58980 1205 59000 1220
rect 59045 1205 59065 1290
rect 59475 1260 59495 1870
rect 59465 1255 59505 1260
rect 59465 1225 59470 1255
rect 59500 1225 59505 1255
rect 59465 1220 59505 1225
rect 58785 535 58790 1205
rect 58810 535 58815 1205
rect 58975 1200 59010 1205
rect 58975 1160 59010 1165
rect 59035 1200 59070 1205
rect 59035 1160 59070 1165
rect 58680 515 58720 520
rect 58680 485 58685 515
rect 58715 485 58720 515
rect 58680 480 58720 485
rect 58785 495 58815 535
rect 58785 475 58790 495
rect 58810 475 58815 495
rect 58785 400 58815 475
rect 59525 400 59545 2415
rect 54245 395 54285 400
rect 54245 365 54250 395
rect 54280 365 54285 395
rect 54245 360 54285 365
rect 54985 395 55025 400
rect 54985 365 54990 395
rect 55020 365 55025 395
rect 54985 360 55025 365
rect 55185 395 55225 400
rect 55185 365 55190 395
rect 55220 365 55225 395
rect 55185 360 55225 365
rect 55385 395 55425 400
rect 55385 365 55390 395
rect 55420 365 55425 395
rect 55385 360 55425 365
rect 55585 395 55625 400
rect 55585 365 55590 395
rect 55620 365 55625 395
rect 55585 360 55625 365
rect 55785 395 55825 400
rect 55785 365 55790 395
rect 55820 365 55825 395
rect 55785 360 55825 365
rect 56430 395 56470 400
rect 56430 365 56435 395
rect 56465 365 56470 395
rect 56430 360 56470 365
rect 56760 395 56800 400
rect 56760 365 56765 395
rect 56795 365 56800 395
rect 56760 360 56800 365
rect 56880 395 56920 400
rect 56880 365 56885 395
rect 56915 365 56920 395
rect 56880 360 56920 365
rect 57910 395 57950 400
rect 57910 365 57915 395
rect 57945 365 57950 395
rect 57910 360 57950 365
rect 58180 395 58220 400
rect 58180 365 58185 395
rect 58215 365 58220 395
rect 58180 360 58220 365
rect 58380 395 58420 400
rect 58380 365 58385 395
rect 58415 365 58420 395
rect 58380 360 58420 365
rect 58580 395 58620 400
rect 58580 365 58585 395
rect 58615 365 58620 395
rect 58580 360 58620 365
rect 58780 395 58820 400
rect 58780 365 58785 395
rect 58815 365 58820 395
rect 58780 360 58820 365
rect 59515 395 59555 400
rect 59515 365 59520 395
rect 59550 365 59555 395
rect 59515 360 59555 365
rect 56890 -455 56910 360
<< via1 >>
rect 56210 4785 56240 4815
rect 56090 4755 56120 4760
rect 56090 4735 56095 4755
rect 56095 4735 56115 4755
rect 56115 4735 56120 4755
rect 56090 4730 56120 4735
rect 56680 4785 56710 4815
rect 56210 4730 56240 4760
rect 56270 4755 56300 4760
rect 56270 4735 56275 4755
rect 56275 4735 56295 4755
rect 56295 4735 56300 4755
rect 56270 4730 56300 4735
rect 56560 4585 56590 4590
rect 56560 4565 56565 4585
rect 56565 4565 56585 4585
rect 56585 4565 56590 4585
rect 56560 4560 56590 4565
rect 56620 4560 56650 4590
rect 57090 4785 57120 4815
rect 57560 4785 57590 4815
rect 56885 4730 56915 4760
rect 57030 4755 57060 4760
rect 57030 4735 57035 4755
rect 57035 4735 57055 4755
rect 57055 4735 57060 4755
rect 57030 4730 57060 4735
rect 56740 4585 56770 4590
rect 56740 4565 56745 4585
rect 56745 4565 56765 4585
rect 56765 4565 56770 4585
rect 56740 4560 56770 4565
rect 56885 4560 56915 4590
rect 56210 4325 56240 4355
rect 56680 4325 56710 4355
rect 56155 4305 56185 4310
rect 56155 4285 56160 4305
rect 56160 4285 56180 4305
rect 56180 4285 56185 4305
rect 56155 4280 56185 4285
rect 56630 4305 56660 4310
rect 56630 4285 56635 4305
rect 56635 4285 56655 4305
rect 56655 4285 56660 4305
rect 56630 4280 56660 4285
rect 56830 4280 56860 4310
rect 55290 4170 55320 4200
rect 55765 4170 55795 4200
rect 54930 4090 54960 4120
rect 55050 4090 55080 4120
rect 55170 4090 55200 4120
rect 55290 4090 55320 4120
rect 55410 4090 55440 4120
rect 55530 4090 55560 4120
rect 55650 4090 55680 4120
rect 54990 4045 55020 4075
rect 55110 4045 55140 4075
rect 55230 4045 55260 4075
rect 55350 4045 55380 4075
rect 55470 4045 55500 4075
rect 55590 4045 55620 4075
rect 54990 3655 55020 3685
rect 55110 3655 55140 3685
rect 55230 3655 55260 3685
rect 55350 3655 55380 3685
rect 55470 3655 55500 3685
rect 55590 3655 55620 3685
rect 55290 3555 55320 3560
rect 55290 3535 55295 3555
rect 55295 3535 55315 3555
rect 55315 3535 55320 3555
rect 55290 3530 55320 3535
rect 54610 3370 54640 3400
rect 55915 4090 55945 4120
rect 56010 4090 56040 4120
rect 56130 4090 56160 4120
rect 56250 4090 56280 4120
rect 56370 4090 56400 4120
rect 56490 4090 56520 4120
rect 56610 4090 56640 4120
rect 56730 4090 56760 4120
rect 56070 4045 56100 4075
rect 55915 3655 55945 3685
rect 56190 4045 56220 4075
rect 56310 4045 56340 4075
rect 56430 4045 56460 4075
rect 56550 4045 56580 4075
rect 56670 4045 56700 4075
rect 56070 3655 56100 3685
rect 56190 3655 56220 3685
rect 56310 3655 56340 3685
rect 56430 3655 56460 3685
rect 56550 3655 56580 3685
rect 56670 3655 56700 3685
rect 54960 3350 54990 3380
rect 55070 3350 55100 3380
rect 55180 3350 55210 3380
rect 55290 3350 55320 3380
rect 55400 3350 55430 3380
rect 55510 3350 55540 3380
rect 55620 3350 55650 3380
rect 55765 3350 55795 3380
rect 55015 3270 55045 3300
rect 55125 3270 55155 3300
rect 55235 3270 55265 3300
rect 55345 3270 55375 3300
rect 55455 3270 55485 3300
rect 55565 3270 55595 3300
rect 55720 3295 55750 3325
rect 55015 2630 55045 2660
rect 55125 2630 55155 2660
rect 55235 2630 55265 2660
rect 55345 2630 55375 2660
rect 55455 2630 55485 2660
rect 55565 2630 55595 2660
rect 54610 2560 54640 2590
rect 55180 2580 55210 2585
rect 55180 2560 55185 2580
rect 55185 2560 55205 2580
rect 55205 2560 55210 2580
rect 55180 2555 55210 2560
rect 57150 4730 57180 4760
rect 57210 4755 57240 4760
rect 57210 4735 57215 4755
rect 57215 4735 57235 4755
rect 57235 4735 57240 4755
rect 57210 4730 57240 4735
rect 57500 4755 57530 4760
rect 57500 4735 57505 4755
rect 57505 4735 57525 4755
rect 57525 4735 57530 4755
rect 57500 4730 57530 4735
rect 57560 4730 57590 4760
rect 57680 4755 57710 4760
rect 57680 4735 57685 4755
rect 57685 4735 57705 4755
rect 57705 4735 57710 4755
rect 57680 4730 57710 4735
rect 57090 4325 57120 4355
rect 57560 4325 57590 4355
rect 56940 4225 56970 4255
rect 57576 4295 57606 4300
rect 57576 4275 57581 4295
rect 57581 4275 57601 4295
rect 57601 4275 57606 4295
rect 57576 4270 57606 4275
rect 56885 4170 56915 4200
rect 56370 3600 56400 3605
rect 56370 3580 56375 3600
rect 56375 3580 56395 3600
rect 56395 3580 56400 3600
rect 56370 3575 56400 3580
rect 56840 3575 56870 3605
rect 57140 4215 57170 4245
rect 57620 4215 57650 4245
rect 58010 4170 58040 4200
rect 58485 4170 58515 4200
rect 57040 4090 57070 4120
rect 57160 4090 57190 4120
rect 57280 4090 57310 4120
rect 57400 4090 57430 4120
rect 57520 4090 57550 4120
rect 57640 4090 57670 4120
rect 57760 4090 57790 4120
rect 57855 4090 57885 4120
rect 57100 4045 57130 4075
rect 57220 4045 57250 4075
rect 57340 4045 57370 4075
rect 57460 4045 57490 4075
rect 57580 4045 57610 4075
rect 57700 4045 57730 4075
rect 57100 3655 57130 3685
rect 57220 3655 57250 3685
rect 57340 3655 57370 3685
rect 57460 3655 57490 3685
rect 57580 3655 57610 3685
rect 57700 3655 57730 3685
rect 57400 3600 57430 3605
rect 57400 3580 57405 3600
rect 57405 3580 57425 3600
rect 57425 3580 57430 3600
rect 57400 3575 57430 3580
rect 56930 3530 56960 3560
rect 56280 3350 56310 3380
rect 56390 3350 56420 3380
rect 56500 3350 56530 3380
rect 56610 3350 56640 3380
rect 56720 3350 56750 3380
rect 56830 3350 56860 3380
rect 56940 3350 56970 3380
rect 57050 3350 57080 3380
rect 57160 3350 57190 3380
rect 57270 3350 57300 3380
rect 57380 3350 57410 3380
rect 57490 3350 57520 3380
rect 56070 3295 56100 3325
rect 56335 3305 56365 3335
rect 56445 3260 56475 3290
rect 56335 3170 56365 3200
rect 56555 3305 56585 3335
rect 56665 3260 56695 3290
rect 56555 3170 56585 3200
rect 56775 3305 56805 3335
rect 56885 3260 56915 3290
rect 56775 3170 56805 3200
rect 56445 3100 56475 3130
rect 56665 3100 56695 3130
rect 55945 2990 55975 3020
rect 56040 3015 56070 3020
rect 56040 2995 56045 3015
rect 56045 2995 56065 3015
rect 56065 2995 56070 3015
rect 56040 2990 56070 2995
rect 56145 2995 56175 3025
rect 56255 2995 56285 3025
rect 56365 2995 56395 3025
rect 56475 2995 56505 3025
rect 56585 2995 56615 3025
rect 56690 3015 56720 3020
rect 56690 2995 56695 3015
rect 56695 2995 56715 3015
rect 56715 2995 56720 3015
rect 56690 2990 56720 2995
rect 55765 2715 55795 2745
rect 55720 2560 55750 2590
rect 54300 2515 54330 2545
rect 55455 2515 55485 2545
rect 54250 2420 54280 2450
rect 54960 2465 54990 2495
rect 55620 2465 55650 2495
rect 55015 2420 55045 2450
rect 55125 2420 55155 2450
rect 55235 2420 55265 2450
rect 55345 2420 55375 2450
rect 55455 2420 55485 2450
rect 55565 2420 55595 2450
rect 55070 2375 55100 2405
rect 55180 2375 55210 2405
rect 55290 2375 55320 2405
rect 55400 2375 55430 2405
rect 55510 2375 55540 2405
rect 54765 2120 54795 2150
rect 55070 2145 55100 2150
rect 55070 2125 55075 2145
rect 55075 2125 55095 2145
rect 55095 2125 55100 2145
rect 55070 2120 55100 2125
rect 55180 2145 55210 2150
rect 55180 2125 55185 2145
rect 55185 2125 55205 2145
rect 55205 2125 55210 2145
rect 55180 2120 55210 2125
rect 55290 2145 55320 2150
rect 55290 2125 55295 2145
rect 55295 2125 55315 2145
rect 55315 2125 55320 2145
rect 55290 2120 55320 2125
rect 55400 2145 55430 2150
rect 55400 2125 55405 2145
rect 55405 2125 55425 2145
rect 55425 2125 55430 2145
rect 55400 2120 55430 2125
rect 55510 2145 55540 2150
rect 55510 2125 55515 2145
rect 55515 2125 55535 2145
rect 55535 2125 55540 2145
rect 55510 2120 55540 2125
rect 54300 1880 54330 1910
rect 54450 1590 54485 1595
rect 54450 1565 54455 1590
rect 54455 1565 54480 1590
rect 54480 1565 54485 1590
rect 54450 1560 54485 1565
rect 54510 1590 54545 1595
rect 54510 1565 54515 1590
rect 54515 1565 54540 1590
rect 54540 1565 54545 1590
rect 54510 1560 54545 1565
rect 54570 1590 54605 1595
rect 54570 1565 54575 1590
rect 54575 1565 54600 1590
rect 54600 1565 54605 1590
rect 54570 1560 54605 1565
rect 54630 1590 54665 1595
rect 54630 1565 54635 1590
rect 54635 1565 54660 1590
rect 54660 1565 54665 1590
rect 54630 1560 54665 1565
rect 55765 2465 55795 2495
rect 55455 2050 55485 2055
rect 55455 2030 55460 2050
rect 55460 2030 55480 2050
rect 55480 2030 55485 2050
rect 55455 2025 55485 2030
rect 55720 2025 55750 2055
rect 54810 1915 54840 1945
rect 55070 1915 55100 1945
rect 55180 1915 55210 1945
rect 55290 1915 55320 1945
rect 55400 1915 55430 1945
rect 55510 1915 55540 1945
rect 54810 1560 54840 1590
rect 55070 1575 55100 1605
rect 55180 1575 55210 1605
rect 55290 1575 55320 1605
rect 55400 1575 55430 1605
rect 55510 1575 55540 1605
rect 55835 2240 55865 2270
rect 54575 1505 54605 1535
rect 54765 1505 54795 1535
rect 55015 1530 55045 1560
rect 55125 1530 55155 1560
rect 55235 1530 55265 1560
rect 55345 1530 55375 1560
rect 55455 1530 55485 1560
rect 55565 1530 55595 1560
rect 55765 1530 55795 1560
rect 54960 1435 54990 1465
rect 55620 1435 55650 1465
rect 55790 1435 55820 1465
rect 54455 1390 54485 1420
rect 54710 1295 54740 1325
rect 55390 1295 55420 1325
rect 54300 1225 54330 1255
rect 54775 1225 54805 1255
rect 55090 1225 55120 1255
rect 55290 1225 55320 1255
rect 55490 1225 55520 1255
rect 54710 1190 54745 1195
rect 54710 1165 54715 1190
rect 54715 1165 54740 1190
rect 54740 1165 54745 1190
rect 54710 1160 54745 1165
rect 54770 1190 54805 1195
rect 54770 1165 54775 1190
rect 54775 1165 54800 1190
rect 54800 1165 54805 1190
rect 54770 1160 54805 1165
rect 55090 485 55120 515
rect 55290 485 55320 515
rect 55790 860 55820 890
rect 55490 485 55520 515
rect 56090 2950 56120 2980
rect 56200 2950 56230 2980
rect 56145 2860 56175 2890
rect 56310 2950 56340 2980
rect 56255 2860 56285 2890
rect 56420 2950 56450 2980
rect 56365 2860 56395 2890
rect 56530 2950 56560 2980
rect 56475 2860 56505 2890
rect 56640 2950 56670 2980
rect 56585 2860 56615 2890
rect 56995 3305 57025 3335
rect 57105 3260 57135 3290
rect 56995 3170 57025 3200
rect 57215 3305 57245 3335
rect 57325 3260 57355 3290
rect 57215 3170 57245 3200
rect 56885 3100 56915 3130
rect 57105 3100 57135 3130
rect 57435 3305 57465 3335
rect 57855 3655 57885 3685
rect 58125 4090 58155 4120
rect 58245 4090 58275 4120
rect 58365 4090 58395 4120
rect 58485 4090 58515 4120
rect 58605 4090 58635 4120
rect 58725 4090 58755 4120
rect 58845 4090 58875 4120
rect 58185 4045 58215 4075
rect 58305 4045 58335 4075
rect 58425 4045 58455 4075
rect 58545 4045 58575 4075
rect 58665 4045 58695 4075
rect 58785 4045 58815 4075
rect 58185 3655 58215 3685
rect 58305 3655 58335 3685
rect 58425 3655 58455 3685
rect 58545 3655 58575 3685
rect 58665 3655 58695 3685
rect 58785 3655 58815 3685
rect 58485 3555 58515 3560
rect 58485 3535 58490 3555
rect 58490 3535 58510 3555
rect 58510 3535 58515 3555
rect 58485 3530 58515 3535
rect 58010 3350 58040 3380
rect 58155 3350 58185 3380
rect 58265 3350 58295 3380
rect 58375 3350 58405 3380
rect 58485 3350 58515 3380
rect 58595 3350 58625 3380
rect 58705 3350 58735 3380
rect 58815 3350 58845 3380
rect 59160 3370 59190 3400
rect 57700 3295 57730 3325
rect 57435 3170 57465 3200
rect 57325 3100 57355 3130
rect 57080 3015 57110 3020
rect 57080 2995 57085 3015
rect 57085 2995 57105 3015
rect 57105 2995 57110 3015
rect 57080 2990 57110 2995
rect 57185 2995 57215 3025
rect 57295 2995 57325 3025
rect 57405 2995 57435 3025
rect 57515 2995 57545 3025
rect 57625 2995 57655 3025
rect 57730 3015 57760 3020
rect 57730 2995 57735 3015
rect 57735 2995 57755 3015
rect 57755 2995 57760 3015
rect 57730 2990 57760 2995
rect 57130 2950 57160 2980
rect 57185 2860 57215 2890
rect 56090 2815 56120 2845
rect 56200 2815 56230 2845
rect 56310 2815 56340 2845
rect 56420 2815 56450 2845
rect 56530 2815 56560 2845
rect 56640 2815 56670 2845
rect 56095 2785 56125 2790
rect 56095 2765 56100 2785
rect 56100 2765 56120 2785
rect 56120 2765 56125 2785
rect 56095 2760 56125 2765
rect 56580 2785 56610 2790
rect 56580 2765 56585 2785
rect 56585 2765 56605 2785
rect 56605 2765 56610 2785
rect 56580 2760 56610 2765
rect 56830 2815 56860 2845
rect 57130 2815 57160 2845
rect 57190 2785 57220 2790
rect 57190 2765 57195 2785
rect 57195 2765 57215 2785
rect 57215 2765 57220 2785
rect 57190 2760 57220 2765
rect 56035 2715 56065 2745
rect 56695 2715 56725 2745
rect 57075 2715 57105 2745
rect 57350 2950 57380 2980
rect 57295 2860 57325 2890
rect 57405 2860 57435 2890
rect 57350 2815 57380 2845
rect 56610 2660 56640 2690
rect 56830 2660 56860 2690
rect 57050 2660 57080 2690
rect 57240 2660 57270 2690
rect 56310 2560 56340 2590
rect 56095 2265 56125 2270
rect 56095 2245 56100 2265
rect 56100 2245 56120 2265
rect 56120 2245 56125 2265
rect 56095 2240 56125 2245
rect 56145 2230 56175 2260
rect 56255 2230 56285 2260
rect 56090 2185 56120 2215
rect 56200 2185 56230 2215
rect 56145 1995 56175 2025
rect 56720 2630 56750 2635
rect 56720 2610 56725 2630
rect 56725 2610 56745 2630
rect 56745 2610 56750 2630
rect 56720 2605 56750 2610
rect 56555 2510 56585 2515
rect 56555 2490 56560 2510
rect 56560 2490 56580 2510
rect 56580 2490 56585 2510
rect 56555 2485 56585 2490
rect 56665 2485 56695 2515
rect 56610 2430 56640 2460
rect 56940 2630 56970 2635
rect 56940 2610 56945 2630
rect 56945 2610 56965 2630
rect 56965 2610 56970 2630
rect 56940 2605 56970 2610
rect 56775 2485 56805 2515
rect 56885 2485 56915 2515
rect 56830 2430 56860 2460
rect 57570 2950 57600 2980
rect 57515 2860 57545 2890
rect 57825 2990 57855 3020
rect 57625 2860 57655 2890
rect 57570 2815 57600 2845
rect 57735 2715 57765 2745
rect 57460 2660 57490 2690
rect 57680 2660 57710 2690
rect 57160 2605 57190 2635
rect 57350 2605 57380 2635
rect 56995 2485 57025 2515
rect 57105 2485 57135 2515
rect 57050 2430 57080 2460
rect 57460 2560 57490 2590
rect 57215 2510 57245 2515
rect 57215 2490 57220 2510
rect 57220 2490 57240 2510
rect 57240 2490 57245 2510
rect 57215 2485 57245 2490
rect 56720 2385 56750 2415
rect 56940 2385 56970 2415
rect 57160 2385 57190 2415
rect 56635 2265 56665 2270
rect 56365 2230 56395 2260
rect 56475 2230 56505 2260
rect 56585 2230 56615 2260
rect 56635 2245 56640 2265
rect 56640 2245 56660 2265
rect 56660 2245 56665 2265
rect 56635 2240 56665 2245
rect 57135 2265 57165 2270
rect 57135 2245 57140 2265
rect 57140 2245 57160 2265
rect 57160 2245 57165 2265
rect 57135 2240 57165 2245
rect 57185 2230 57215 2260
rect 57295 2230 57325 2260
rect 57405 2230 57435 2260
rect 56310 2185 56340 2215
rect 56255 1995 56285 2025
rect 56420 2185 56450 2215
rect 56365 1995 56395 2025
rect 56090 1950 56120 1980
rect 56200 1950 56230 1980
rect 56310 1950 56340 1980
rect 56035 1905 56065 1935
rect 56530 2185 56560 2215
rect 56475 1995 56505 2025
rect 56640 2185 56670 2215
rect 57130 2185 57160 2215
rect 56585 1995 56615 2025
rect 56420 1950 56450 1980
rect 56530 1950 56560 1980
rect 56640 1950 56670 1980
rect 57240 2185 57270 2215
rect 57185 1995 57215 2025
rect 57350 2185 57380 2215
rect 57295 1995 57325 2025
rect 57515 2230 57545 2260
rect 57625 2230 57655 2260
rect 57460 2185 57490 2215
rect 57405 1995 57435 2025
rect 57130 1950 57160 1980
rect 57240 1950 57270 1980
rect 57350 1950 57380 1980
rect 56695 1905 56725 1935
rect 57075 1905 57105 1935
rect 56040 1780 56070 1785
rect 56040 1760 56045 1780
rect 56045 1760 56065 1780
rect 56065 1760 56070 1780
rect 56090 1765 56120 1795
rect 56200 1765 56230 1795
rect 56310 1765 56340 1795
rect 56365 1775 56395 1805
rect 56420 1765 56450 1795
rect 56530 1765 56560 1795
rect 56640 1765 56670 1795
rect 56690 1780 56720 1785
rect 56690 1760 56695 1780
rect 56695 1760 56715 1780
rect 56715 1760 56720 1780
rect 56040 1755 56070 1760
rect 56145 1720 56175 1750
rect 56090 1525 56120 1555
rect 56255 1720 56285 1750
rect 56200 1525 56230 1555
rect 56365 1720 56395 1750
rect 56310 1525 56340 1555
rect 56475 1720 56505 1750
rect 56420 1525 56450 1555
rect 56585 1720 56615 1750
rect 56530 1525 56560 1555
rect 56690 1755 56720 1760
rect 56850 1780 56880 1785
rect 56850 1760 56855 1780
rect 56855 1760 56875 1780
rect 56875 1760 56880 1780
rect 56850 1755 56880 1760
rect 56903 1780 56933 1785
rect 56903 1760 56908 1780
rect 56908 1760 56928 1780
rect 56928 1760 56933 1780
rect 56903 1755 56933 1760
rect 57570 2185 57600 2215
rect 57515 1995 57545 2025
rect 57680 2185 57710 2215
rect 57625 1995 57655 2025
rect 57460 1950 57490 1980
rect 57570 1950 57600 1980
rect 57680 1950 57710 1980
rect 57735 1905 57765 1935
rect 57080 1780 57110 1785
rect 57080 1760 57085 1780
rect 57085 1760 57105 1780
rect 57105 1760 57110 1780
rect 57130 1765 57160 1795
rect 57240 1765 57270 1795
rect 57350 1765 57380 1795
rect 57405 1775 57435 1805
rect 57460 1765 57490 1795
rect 57570 1765 57600 1795
rect 57680 1765 57710 1795
rect 57730 1780 57760 1785
rect 57730 1760 57735 1780
rect 57735 1760 57755 1780
rect 57755 1760 57760 1780
rect 57080 1755 57110 1760
rect 57185 1720 57215 1750
rect 56640 1525 56670 1555
rect 56145 1480 56175 1510
rect 56255 1480 56285 1510
rect 56365 1480 56395 1510
rect 56475 1480 56505 1510
rect 56585 1480 56615 1510
rect 56035 1435 56065 1465
rect 56735 1435 56765 1465
rect 55945 1390 55975 1420
rect 56830 1390 56860 1420
rect 56335 1235 56365 1265
rect 57130 1525 57160 1555
rect 57295 1720 57325 1750
rect 57240 1525 57270 1555
rect 57405 1720 57435 1750
rect 57350 1525 57380 1555
rect 57515 1720 57545 1750
rect 57460 1525 57490 1555
rect 57625 1720 57655 1750
rect 57570 1525 57600 1555
rect 57730 1755 57760 1760
rect 57680 1525 57710 1555
rect 57185 1480 57215 1510
rect 57295 1480 57325 1510
rect 57405 1480 57435 1510
rect 57515 1480 57545 1510
rect 57625 1480 57655 1510
rect 57035 1435 57065 1465
rect 56940 1390 56970 1420
rect 56885 1235 56915 1265
rect 57735 1435 57765 1465
rect 58055 3295 58085 3325
rect 58010 2715 58040 2745
rect 57915 2485 57945 2515
rect 58210 3270 58240 3300
rect 58320 3270 58350 3300
rect 58430 3270 58460 3300
rect 58540 3270 58570 3300
rect 58650 3270 58680 3300
rect 58760 3270 58790 3300
rect 58210 2630 58240 2660
rect 58320 2630 58350 2660
rect 58430 2630 58460 2660
rect 58540 2630 58570 2660
rect 58650 2630 58680 2660
rect 58760 2630 58790 2660
rect 58055 2560 58085 2590
rect 57870 2430 57900 2460
rect 57825 1390 57855 1420
rect 58010 2465 58040 2495
rect 57915 1905 57945 1935
rect 58595 2580 58625 2585
rect 58595 2560 58600 2580
rect 58600 2560 58620 2580
rect 58620 2560 58625 2580
rect 58595 2555 58625 2560
rect 59160 2560 59190 2590
rect 58320 2515 58350 2545
rect 59470 2515 59500 2545
rect 58155 2465 58185 2495
rect 58815 2465 58845 2495
rect 58210 2420 58240 2450
rect 58320 2420 58350 2450
rect 58430 2420 58460 2450
rect 58540 2420 58570 2450
rect 58650 2420 58680 2450
rect 58760 2420 58790 2450
rect 58265 2375 58295 2405
rect 58375 2375 58405 2405
rect 58485 2375 58515 2405
rect 58595 2375 58625 2405
rect 58705 2375 58735 2405
rect 58265 2145 58295 2150
rect 58265 2125 58270 2145
rect 58270 2125 58290 2145
rect 58290 2125 58295 2145
rect 58265 2120 58295 2125
rect 58375 2145 58405 2150
rect 58375 2125 58380 2145
rect 58380 2125 58400 2145
rect 58400 2125 58405 2145
rect 58375 2120 58405 2125
rect 58485 2145 58515 2150
rect 58485 2125 58490 2145
rect 58490 2125 58510 2145
rect 58510 2125 58515 2145
rect 58485 2120 58515 2125
rect 58595 2145 58625 2150
rect 58595 2125 58600 2145
rect 58600 2125 58620 2145
rect 58620 2125 58625 2145
rect 58595 2120 58625 2125
rect 58705 2145 58735 2150
rect 58705 2125 58710 2145
rect 58710 2125 58730 2145
rect 58730 2125 58735 2145
rect 58705 2120 58735 2125
rect 59005 2120 59035 2150
rect 58055 2025 58085 2055
rect 58320 2050 58350 2055
rect 58320 2030 58325 2050
rect 58325 2030 58345 2050
rect 58345 2030 58350 2050
rect 58320 2025 58350 2030
rect 58265 1915 58295 1945
rect 58375 1915 58405 1945
rect 58485 1915 58515 1945
rect 58595 1915 58625 1945
rect 58705 1915 58735 1945
rect 58960 1915 58990 1945
rect 58265 1575 58295 1605
rect 58375 1575 58405 1605
rect 58485 1575 58515 1605
rect 58595 1575 58625 1605
rect 58705 1575 58735 1605
rect 58010 1530 58040 1560
rect 58210 1530 58240 1560
rect 58320 1530 58350 1560
rect 58430 1530 58460 1560
rect 58540 1530 58570 1560
rect 58650 1530 58680 1560
rect 58760 1530 58790 1560
rect 58960 1510 58990 1540
rect 59520 2420 59550 2450
rect 59470 1880 59500 1910
rect 59135 1540 59170 1545
rect 59135 1515 59140 1540
rect 59140 1515 59165 1540
rect 59165 1515 59170 1540
rect 59135 1510 59170 1515
rect 59195 1540 59230 1545
rect 59195 1515 59200 1540
rect 59200 1515 59225 1540
rect 59225 1515 59230 1540
rect 59195 1510 59230 1515
rect 59255 1540 59290 1545
rect 59255 1515 59260 1540
rect 59260 1515 59285 1540
rect 59285 1515 59290 1540
rect 59255 1510 59290 1515
rect 59315 1540 59350 1545
rect 59315 1515 59320 1540
rect 59320 1515 59345 1540
rect 59345 1515 59350 1540
rect 59315 1510 59350 1515
rect 57915 1435 57945 1465
rect 58155 1435 58185 1465
rect 58815 1435 58845 1465
rect 59005 1455 59035 1485
rect 59195 1455 59225 1485
rect 57410 1260 57440 1265
rect 57410 1240 57415 1260
rect 57415 1240 57435 1260
rect 57435 1240 57440 1260
rect 57410 1235 57440 1240
rect 57870 1235 57900 1265
rect 56445 1180 56475 1210
rect 56555 1180 56585 1210
rect 56665 1180 56695 1210
rect 56775 1180 56805 1210
rect 56885 1180 56915 1210
rect 56995 1180 57025 1210
rect 57105 1180 57135 1210
rect 57215 1180 57245 1210
rect 57325 1180 57355 1210
rect 57435 1180 57465 1210
rect 56225 885 56255 890
rect 56225 865 56230 885
rect 56230 865 56250 885
rect 56250 865 56255 885
rect 56225 860 56255 865
rect 56280 860 56310 890
rect 56390 860 56420 890
rect 56500 860 56530 890
rect 56610 860 56640 890
rect 56720 860 56750 890
rect 56830 860 56860 890
rect 56940 860 56970 890
rect 57050 860 57080 890
rect 57160 860 57190 890
rect 57270 860 57300 890
rect 57380 860 57410 890
rect 57490 885 57520 890
rect 57490 865 57495 885
rect 57495 865 57515 885
rect 57515 865 57520 885
rect 57490 860 57520 865
rect 59315 1390 59345 1420
rect 58435 1295 58465 1325
rect 59040 1295 59070 1325
rect 58285 1225 58315 1255
rect 58485 1225 58515 1255
rect 58685 1225 58715 1255
rect 58975 1225 59005 1255
rect 57915 850 57945 880
rect 56445 815 56475 845
rect 56555 815 56585 845
rect 56665 815 56695 845
rect 56775 815 56805 845
rect 56885 815 56915 845
rect 56995 815 57025 845
rect 57105 815 57135 845
rect 57215 815 57245 845
rect 57325 815 57355 845
rect 57435 815 57465 845
rect 56545 760 56575 790
rect 56655 760 56685 790
rect 56875 760 56905 790
rect 55835 715 55865 745
rect 56490 715 56520 745
rect 56600 740 56630 745
rect 56600 720 56605 740
rect 56605 720 56625 740
rect 56625 720 56630 740
rect 56600 715 56630 720
rect 56545 510 56575 540
rect 56710 715 56740 745
rect 56655 510 56685 540
rect 57045 740 57075 745
rect 57045 720 57050 740
rect 57050 720 57070 740
rect 57070 720 57075 740
rect 57045 715 57075 720
rect 56875 510 56905 540
rect 56490 465 56520 495
rect 56600 465 56630 495
rect 56710 465 56740 495
rect 58285 485 58315 515
rect 58485 485 58515 515
rect 59470 1225 59500 1255
rect 58975 1195 59010 1200
rect 58975 1170 58980 1195
rect 58980 1170 59005 1195
rect 59005 1170 59010 1195
rect 58975 1165 59010 1170
rect 59035 1195 59070 1200
rect 59035 1170 59040 1195
rect 59040 1170 59065 1195
rect 59065 1170 59070 1195
rect 59035 1165 59070 1170
rect 58685 485 58715 515
rect 54250 365 54280 395
rect 54990 365 55020 395
rect 55190 365 55220 395
rect 55390 365 55420 395
rect 55590 365 55620 395
rect 55790 365 55820 395
rect 56435 365 56465 395
rect 56765 365 56795 395
rect 56885 365 56915 395
rect 57915 365 57945 395
rect 58185 365 58215 395
rect 58385 365 58415 395
rect 58585 365 58615 395
rect 58785 365 58815 395
rect 59520 365 59550 395
<< metal2 >>
rect 56205 4815 56245 4820
rect 56205 4785 56210 4815
rect 56240 4810 56245 4815
rect 56675 4815 56715 4820
rect 56675 4810 56680 4815
rect 56240 4790 56680 4810
rect 56240 4785 56245 4790
rect 56205 4780 56245 4785
rect 56675 4785 56680 4790
rect 56710 4785 56715 4815
rect 56675 4780 56715 4785
rect 57085 4815 57125 4820
rect 57085 4785 57090 4815
rect 57120 4810 57125 4815
rect 57555 4815 57595 4820
rect 57555 4810 57560 4815
rect 57120 4790 57560 4810
rect 57120 4785 57125 4790
rect 57085 4780 57125 4785
rect 57555 4785 57560 4790
rect 57590 4785 57595 4815
rect 57555 4780 57595 4785
rect 56085 4760 56125 4765
rect 56085 4730 56090 4760
rect 56120 4755 56125 4760
rect 56205 4760 56245 4765
rect 56205 4755 56210 4760
rect 56120 4735 56210 4755
rect 56120 4730 56125 4735
rect 56085 4725 56125 4730
rect 56205 4730 56210 4735
rect 56240 4755 56245 4760
rect 56265 4760 56305 4765
rect 56265 4755 56270 4760
rect 56240 4735 56270 4755
rect 56240 4730 56245 4735
rect 56205 4725 56245 4730
rect 56265 4730 56270 4735
rect 56300 4730 56305 4760
rect 56265 4725 56305 4730
rect 56880 4760 56920 4765
rect 56880 4730 56885 4760
rect 56915 4755 56920 4760
rect 57025 4760 57065 4765
rect 57025 4755 57030 4760
rect 56915 4735 57030 4755
rect 56915 4730 56920 4735
rect 56880 4725 56920 4730
rect 57025 4730 57030 4735
rect 57060 4755 57065 4760
rect 57145 4760 57185 4765
rect 57145 4755 57150 4760
rect 57060 4735 57150 4755
rect 57060 4730 57065 4735
rect 57025 4725 57065 4730
rect 57145 4730 57150 4735
rect 57180 4755 57185 4760
rect 57205 4760 57245 4765
rect 57205 4755 57210 4760
rect 57180 4735 57210 4755
rect 57180 4730 57185 4735
rect 57145 4725 57185 4730
rect 57205 4730 57210 4735
rect 57240 4730 57245 4760
rect 57205 4725 57245 4730
rect 57495 4760 57535 4765
rect 57495 4730 57500 4760
rect 57530 4755 57535 4760
rect 57555 4760 57595 4765
rect 57555 4755 57560 4760
rect 57530 4735 57560 4755
rect 57530 4730 57535 4735
rect 57495 4725 57535 4730
rect 57555 4730 57560 4735
rect 57590 4755 57595 4760
rect 57675 4760 57715 4765
rect 57675 4755 57680 4760
rect 57590 4735 57680 4755
rect 57590 4730 57595 4735
rect 57555 4725 57595 4730
rect 57675 4730 57680 4735
rect 57710 4730 57715 4760
rect 57675 4725 57715 4730
rect 56555 4590 56595 4595
rect 56555 4560 56560 4590
rect 56590 4585 56595 4590
rect 56615 4590 56655 4595
rect 56615 4585 56620 4590
rect 56590 4565 56620 4585
rect 56590 4560 56595 4565
rect 56555 4555 56595 4560
rect 56615 4560 56620 4565
rect 56650 4585 56655 4590
rect 56735 4590 56775 4595
rect 56735 4585 56740 4590
rect 56650 4565 56740 4585
rect 56650 4560 56655 4565
rect 56615 4555 56655 4560
rect 56735 4560 56740 4565
rect 56770 4585 56775 4590
rect 56880 4590 56920 4595
rect 56880 4585 56885 4590
rect 56770 4565 56885 4585
rect 56770 4560 56775 4565
rect 56735 4555 56775 4560
rect 56880 4560 56885 4565
rect 56915 4560 56920 4590
rect 56880 4555 56920 4560
rect 56205 4355 56245 4360
rect 56205 4325 56210 4355
rect 56240 4350 56245 4355
rect 56675 4355 56715 4360
rect 56675 4350 56680 4355
rect 56240 4330 56680 4350
rect 56240 4325 56245 4330
rect 56205 4320 56245 4325
rect 56675 4325 56680 4330
rect 56710 4325 56715 4355
rect 56675 4320 56715 4325
rect 57085 4355 57125 4360
rect 57085 4325 57090 4355
rect 57120 4350 57125 4355
rect 57555 4355 57595 4360
rect 57555 4350 57560 4355
rect 57120 4330 57560 4350
rect 57120 4325 57125 4330
rect 57085 4320 57125 4325
rect 57555 4325 57560 4330
rect 57590 4325 57595 4355
rect 57555 4320 57595 4325
rect 56150 4310 56190 4315
rect 56150 4280 56155 4310
rect 56185 4305 56190 4310
rect 56630 4310 56660 4315
rect 56185 4285 56630 4305
rect 56185 4280 56190 4285
rect 56150 4275 56190 4280
rect 56825 4310 56865 4315
rect 56825 4305 56830 4310
rect 56660 4285 56830 4305
rect 56630 4275 56660 4280
rect 56825 4280 56830 4285
rect 56860 4305 56865 4310
rect 56860 4300 57606 4305
rect 56860 4285 57576 4300
rect 56860 4280 56865 4285
rect 56825 4275 56865 4280
rect 57576 4265 57606 4270
rect 56935 4255 56975 4260
rect 56935 4225 56940 4255
rect 56970 4240 56975 4255
rect 57135 4245 57175 4250
rect 57135 4240 57140 4245
rect 56970 4225 57140 4240
rect 56935 4220 57140 4225
rect 57135 4215 57140 4220
rect 57170 4240 57175 4245
rect 57615 4245 57655 4250
rect 57615 4240 57620 4245
rect 57170 4220 57620 4240
rect 57170 4215 57175 4220
rect 57135 4210 57175 4215
rect 57615 4215 57620 4220
rect 57650 4215 57655 4245
rect 57615 4210 57655 4215
rect 55285 4200 55325 4205
rect 55285 4170 55290 4200
rect 55320 4195 55325 4200
rect 55760 4200 55800 4205
rect 55760 4195 55765 4200
rect 55320 4175 55765 4195
rect 55320 4170 55325 4175
rect 55285 4165 55325 4170
rect 55760 4170 55765 4175
rect 55795 4195 55800 4200
rect 56880 4200 56920 4205
rect 56880 4195 56885 4200
rect 55795 4175 56885 4195
rect 55795 4170 55800 4175
rect 55760 4165 55800 4170
rect 56880 4170 56885 4175
rect 56915 4195 56920 4200
rect 58005 4200 58045 4205
rect 58005 4195 58010 4200
rect 56915 4175 58010 4195
rect 56915 4170 56920 4175
rect 56880 4165 56920 4170
rect 58005 4170 58010 4175
rect 58040 4195 58045 4200
rect 58480 4200 58520 4205
rect 58480 4195 58485 4200
rect 58040 4175 58485 4195
rect 58040 4170 58045 4175
rect 58005 4165 58045 4170
rect 58480 4170 58485 4175
rect 58515 4170 58520 4200
rect 58480 4165 58520 4170
rect 54925 4120 54965 4125
rect 54925 4090 54930 4120
rect 54960 4115 54965 4120
rect 55045 4120 55085 4125
rect 55045 4115 55050 4120
rect 54960 4095 55050 4115
rect 54960 4090 54965 4095
rect 54925 4085 54965 4090
rect 55045 4090 55050 4095
rect 55080 4115 55085 4120
rect 55165 4120 55205 4125
rect 55165 4115 55170 4120
rect 55080 4095 55170 4115
rect 55080 4090 55085 4095
rect 55045 4085 55085 4090
rect 55165 4090 55170 4095
rect 55200 4115 55205 4120
rect 55285 4120 55325 4125
rect 55285 4115 55290 4120
rect 55200 4095 55290 4115
rect 55200 4090 55205 4095
rect 55165 4085 55205 4090
rect 55285 4090 55290 4095
rect 55320 4115 55325 4120
rect 55405 4120 55445 4125
rect 55405 4115 55410 4120
rect 55320 4095 55410 4115
rect 55320 4090 55325 4095
rect 55285 4085 55325 4090
rect 55405 4090 55410 4095
rect 55440 4115 55445 4120
rect 55525 4120 55565 4125
rect 55525 4115 55530 4120
rect 55440 4095 55530 4115
rect 55440 4090 55445 4095
rect 55405 4085 55445 4090
rect 55525 4090 55530 4095
rect 55560 4115 55565 4120
rect 55645 4120 55685 4125
rect 55645 4115 55650 4120
rect 55560 4095 55650 4115
rect 55560 4090 55565 4095
rect 55525 4085 55565 4090
rect 55645 4090 55650 4095
rect 55680 4090 55685 4120
rect 55645 4085 55685 4090
rect 55910 4120 55950 4125
rect 55910 4090 55915 4120
rect 55945 4115 55950 4120
rect 56005 4120 56045 4125
rect 56005 4115 56010 4120
rect 55945 4095 56010 4115
rect 55945 4090 55950 4095
rect 55910 4085 55950 4090
rect 56005 4090 56010 4095
rect 56040 4115 56045 4120
rect 56125 4120 56165 4125
rect 56125 4115 56130 4120
rect 56040 4095 56130 4115
rect 56040 4090 56045 4095
rect 56005 4085 56045 4090
rect 56125 4090 56130 4095
rect 56160 4115 56165 4120
rect 56245 4120 56285 4125
rect 56245 4115 56250 4120
rect 56160 4095 56250 4115
rect 56160 4090 56165 4095
rect 56125 4085 56165 4090
rect 56245 4090 56250 4095
rect 56280 4115 56285 4120
rect 56365 4120 56405 4125
rect 56365 4115 56370 4120
rect 56280 4095 56370 4115
rect 56280 4090 56285 4095
rect 56245 4085 56285 4090
rect 56365 4090 56370 4095
rect 56400 4115 56405 4120
rect 56485 4120 56525 4125
rect 56485 4115 56490 4120
rect 56400 4095 56490 4115
rect 56400 4090 56405 4095
rect 56365 4085 56405 4090
rect 56485 4090 56490 4095
rect 56520 4115 56525 4120
rect 56605 4120 56645 4125
rect 56605 4115 56610 4120
rect 56520 4095 56610 4115
rect 56520 4090 56525 4095
rect 56485 4085 56525 4090
rect 56605 4090 56610 4095
rect 56640 4115 56645 4120
rect 56725 4120 56765 4125
rect 56725 4115 56730 4120
rect 56640 4095 56730 4115
rect 56640 4090 56645 4095
rect 56605 4085 56645 4090
rect 56725 4090 56730 4095
rect 56760 4090 56765 4120
rect 56725 4085 56765 4090
rect 57035 4120 57075 4125
rect 57035 4090 57040 4120
rect 57070 4115 57075 4120
rect 57155 4120 57195 4125
rect 57155 4115 57160 4120
rect 57070 4095 57160 4115
rect 57070 4090 57075 4095
rect 57035 4085 57075 4090
rect 57155 4090 57160 4095
rect 57190 4115 57195 4120
rect 57275 4120 57315 4125
rect 57275 4115 57280 4120
rect 57190 4095 57280 4115
rect 57190 4090 57195 4095
rect 57155 4085 57195 4090
rect 57275 4090 57280 4095
rect 57310 4115 57315 4120
rect 57395 4120 57435 4125
rect 57395 4115 57400 4120
rect 57310 4095 57400 4115
rect 57310 4090 57315 4095
rect 57275 4085 57315 4090
rect 57395 4090 57400 4095
rect 57430 4115 57435 4120
rect 57515 4120 57555 4125
rect 57515 4115 57520 4120
rect 57430 4095 57520 4115
rect 57430 4090 57435 4095
rect 57395 4085 57435 4090
rect 57515 4090 57520 4095
rect 57550 4115 57555 4120
rect 57635 4120 57675 4125
rect 57635 4115 57640 4120
rect 57550 4095 57640 4115
rect 57550 4090 57555 4095
rect 57515 4085 57555 4090
rect 57635 4090 57640 4095
rect 57670 4115 57675 4120
rect 57755 4120 57795 4125
rect 57755 4115 57760 4120
rect 57670 4095 57760 4115
rect 57670 4090 57675 4095
rect 57635 4085 57675 4090
rect 57755 4090 57760 4095
rect 57790 4115 57795 4120
rect 57850 4120 57890 4125
rect 57850 4115 57855 4120
rect 57790 4095 57855 4115
rect 57790 4090 57795 4095
rect 57755 4085 57795 4090
rect 57850 4090 57855 4095
rect 57885 4090 57890 4120
rect 57850 4085 57890 4090
rect 58120 4120 58160 4125
rect 58120 4090 58125 4120
rect 58155 4115 58160 4120
rect 58240 4120 58280 4125
rect 58240 4115 58245 4120
rect 58155 4095 58245 4115
rect 58155 4090 58160 4095
rect 58120 4085 58160 4090
rect 58240 4090 58245 4095
rect 58275 4115 58280 4120
rect 58360 4120 58400 4125
rect 58360 4115 58365 4120
rect 58275 4095 58365 4115
rect 58275 4090 58280 4095
rect 58240 4085 58280 4090
rect 58360 4090 58365 4095
rect 58395 4115 58400 4120
rect 58480 4120 58520 4125
rect 58480 4115 58485 4120
rect 58395 4095 58485 4115
rect 58395 4090 58400 4095
rect 58360 4085 58400 4090
rect 58480 4090 58485 4095
rect 58515 4115 58520 4120
rect 58600 4120 58640 4125
rect 58600 4115 58605 4120
rect 58515 4095 58605 4115
rect 58515 4090 58520 4095
rect 58480 4085 58520 4090
rect 58600 4090 58605 4095
rect 58635 4115 58640 4120
rect 58720 4120 58760 4125
rect 58720 4115 58725 4120
rect 58635 4095 58725 4115
rect 58635 4090 58640 4095
rect 58600 4085 58640 4090
rect 58720 4090 58725 4095
rect 58755 4115 58760 4120
rect 58840 4120 58880 4125
rect 58840 4115 58845 4120
rect 58755 4095 58845 4115
rect 58755 4090 58760 4095
rect 58720 4085 58760 4090
rect 58840 4090 58845 4095
rect 58875 4090 58880 4120
rect 58840 4085 58880 4090
rect 54985 4075 55025 4080
rect 54985 4045 54990 4075
rect 55020 4070 55025 4075
rect 55105 4075 55145 4080
rect 55105 4070 55110 4075
rect 55020 4050 55110 4070
rect 55020 4045 55025 4050
rect 54985 4040 55025 4045
rect 55105 4045 55110 4050
rect 55140 4070 55145 4075
rect 55225 4075 55265 4080
rect 55225 4070 55230 4075
rect 55140 4050 55230 4070
rect 55140 4045 55145 4050
rect 55105 4040 55145 4045
rect 55225 4045 55230 4050
rect 55260 4070 55265 4075
rect 55345 4075 55385 4080
rect 55345 4070 55350 4075
rect 55260 4050 55350 4070
rect 55260 4045 55265 4050
rect 55225 4040 55265 4045
rect 55345 4045 55350 4050
rect 55380 4070 55385 4075
rect 55465 4075 55505 4080
rect 55465 4070 55470 4075
rect 55380 4050 55470 4070
rect 55380 4045 55385 4050
rect 55345 4040 55385 4045
rect 55465 4045 55470 4050
rect 55500 4070 55505 4075
rect 55585 4075 55625 4080
rect 55585 4070 55590 4075
rect 55500 4050 55590 4070
rect 55500 4045 55505 4050
rect 55465 4040 55505 4045
rect 55585 4045 55590 4050
rect 55620 4045 55625 4075
rect 55585 4040 55625 4045
rect 56065 4075 56105 4080
rect 56065 4045 56070 4075
rect 56100 4070 56105 4075
rect 56185 4075 56225 4080
rect 56185 4070 56190 4075
rect 56100 4050 56190 4070
rect 56100 4045 56105 4050
rect 56065 4040 56105 4045
rect 56185 4045 56190 4050
rect 56220 4070 56225 4075
rect 56305 4075 56345 4080
rect 56305 4070 56310 4075
rect 56220 4050 56310 4070
rect 56220 4045 56225 4050
rect 56185 4040 56225 4045
rect 56305 4045 56310 4050
rect 56340 4070 56345 4075
rect 56425 4075 56465 4080
rect 56425 4070 56430 4075
rect 56340 4050 56430 4070
rect 56340 4045 56345 4050
rect 56305 4040 56345 4045
rect 56425 4045 56430 4050
rect 56460 4070 56465 4075
rect 56545 4075 56585 4080
rect 56545 4070 56550 4075
rect 56460 4050 56550 4070
rect 56460 4045 56465 4050
rect 56425 4040 56465 4045
rect 56545 4045 56550 4050
rect 56580 4070 56585 4075
rect 56665 4075 56705 4080
rect 56665 4070 56670 4075
rect 56580 4050 56670 4070
rect 56580 4045 56585 4050
rect 56545 4040 56585 4045
rect 56665 4045 56670 4050
rect 56700 4045 56705 4075
rect 56665 4040 56705 4045
rect 57095 4075 57135 4080
rect 57095 4045 57100 4075
rect 57130 4070 57135 4075
rect 57215 4075 57255 4080
rect 57215 4070 57220 4075
rect 57130 4050 57220 4070
rect 57130 4045 57135 4050
rect 57095 4040 57135 4045
rect 57215 4045 57220 4050
rect 57250 4070 57255 4075
rect 57335 4075 57375 4080
rect 57335 4070 57340 4075
rect 57250 4050 57340 4070
rect 57250 4045 57255 4050
rect 57215 4040 57255 4045
rect 57335 4045 57340 4050
rect 57370 4070 57375 4075
rect 57455 4075 57495 4080
rect 57455 4070 57460 4075
rect 57370 4050 57460 4070
rect 57370 4045 57375 4050
rect 57335 4040 57375 4045
rect 57455 4045 57460 4050
rect 57490 4070 57495 4075
rect 57575 4075 57615 4080
rect 57575 4070 57580 4075
rect 57490 4050 57580 4070
rect 57490 4045 57495 4050
rect 57455 4040 57495 4045
rect 57575 4045 57580 4050
rect 57610 4070 57615 4075
rect 57695 4075 57735 4080
rect 57695 4070 57700 4075
rect 57610 4050 57700 4070
rect 57610 4045 57615 4050
rect 57575 4040 57615 4045
rect 57695 4045 57700 4050
rect 57730 4045 57735 4075
rect 57695 4040 57735 4045
rect 58180 4075 58220 4080
rect 58180 4045 58185 4075
rect 58215 4070 58220 4075
rect 58300 4075 58340 4080
rect 58300 4070 58305 4075
rect 58215 4050 58305 4070
rect 58215 4045 58220 4050
rect 58180 4040 58220 4045
rect 58300 4045 58305 4050
rect 58335 4070 58340 4075
rect 58420 4075 58460 4080
rect 58420 4070 58425 4075
rect 58335 4050 58425 4070
rect 58335 4045 58340 4050
rect 58300 4040 58340 4045
rect 58420 4045 58425 4050
rect 58455 4070 58460 4075
rect 58540 4075 58580 4080
rect 58540 4070 58545 4075
rect 58455 4050 58545 4070
rect 58455 4045 58460 4050
rect 58420 4040 58460 4045
rect 58540 4045 58545 4050
rect 58575 4070 58580 4075
rect 58660 4075 58700 4080
rect 58660 4070 58665 4075
rect 58575 4050 58665 4070
rect 58575 4045 58580 4050
rect 58540 4040 58580 4045
rect 58660 4045 58665 4050
rect 58695 4070 58700 4075
rect 58780 4075 58820 4080
rect 58780 4070 58785 4075
rect 58695 4050 58785 4070
rect 58695 4045 58700 4050
rect 58660 4040 58700 4045
rect 58780 4045 58785 4050
rect 58815 4045 58820 4075
rect 58780 4040 58820 4045
rect 54985 3685 55025 3690
rect 54985 3655 54990 3685
rect 55020 3680 55025 3685
rect 55105 3685 55145 3690
rect 55105 3680 55110 3685
rect 55020 3660 55110 3680
rect 55020 3655 55025 3660
rect 54985 3650 55025 3655
rect 55105 3655 55110 3660
rect 55140 3680 55145 3685
rect 55225 3685 55265 3690
rect 55225 3680 55230 3685
rect 55140 3660 55230 3680
rect 55140 3655 55145 3660
rect 55105 3650 55145 3655
rect 55225 3655 55230 3660
rect 55260 3680 55265 3685
rect 55345 3685 55385 3690
rect 55345 3680 55350 3685
rect 55260 3660 55350 3680
rect 55260 3655 55265 3660
rect 55225 3650 55265 3655
rect 55345 3655 55350 3660
rect 55380 3680 55385 3685
rect 55465 3685 55505 3690
rect 55465 3680 55470 3685
rect 55380 3660 55470 3680
rect 55380 3655 55385 3660
rect 55345 3650 55385 3655
rect 55465 3655 55470 3660
rect 55500 3680 55505 3685
rect 55585 3685 55625 3690
rect 55585 3680 55590 3685
rect 55500 3660 55590 3680
rect 55500 3655 55505 3660
rect 55465 3650 55505 3655
rect 55585 3655 55590 3660
rect 55620 3680 55625 3685
rect 55910 3685 55950 3690
rect 55910 3680 55915 3685
rect 55620 3660 55915 3680
rect 55620 3655 55625 3660
rect 55585 3650 55625 3655
rect 55910 3655 55915 3660
rect 55945 3655 55950 3685
rect 55910 3650 55950 3655
rect 56065 3685 56105 3690
rect 56065 3655 56070 3685
rect 56100 3680 56105 3685
rect 56185 3685 56225 3690
rect 56185 3680 56190 3685
rect 56100 3660 56190 3680
rect 56100 3655 56105 3660
rect 56065 3650 56105 3655
rect 56185 3655 56190 3660
rect 56220 3680 56225 3685
rect 56305 3685 56345 3690
rect 56305 3680 56310 3685
rect 56220 3660 56310 3680
rect 56220 3655 56225 3660
rect 56185 3650 56225 3655
rect 56305 3655 56310 3660
rect 56340 3680 56345 3685
rect 56425 3685 56465 3690
rect 56425 3680 56430 3685
rect 56340 3660 56430 3680
rect 56340 3655 56345 3660
rect 56305 3650 56345 3655
rect 56425 3655 56430 3660
rect 56460 3680 56465 3685
rect 56545 3685 56585 3690
rect 56545 3680 56550 3685
rect 56460 3660 56550 3680
rect 56460 3655 56465 3660
rect 56425 3650 56465 3655
rect 56545 3655 56550 3660
rect 56580 3680 56585 3685
rect 56665 3685 56705 3690
rect 56665 3680 56670 3685
rect 56580 3660 56670 3680
rect 56580 3655 56585 3660
rect 56545 3650 56585 3655
rect 56665 3655 56670 3660
rect 56700 3655 56705 3685
rect 56665 3650 56705 3655
rect 57095 3685 57135 3690
rect 57095 3655 57100 3685
rect 57130 3680 57135 3685
rect 57215 3685 57255 3690
rect 57215 3680 57220 3685
rect 57130 3660 57220 3680
rect 57130 3655 57135 3660
rect 57095 3650 57135 3655
rect 57215 3655 57220 3660
rect 57250 3680 57255 3685
rect 57335 3685 57375 3690
rect 57335 3680 57340 3685
rect 57250 3660 57340 3680
rect 57250 3655 57255 3660
rect 57215 3650 57255 3655
rect 57335 3655 57340 3660
rect 57370 3680 57375 3685
rect 57455 3685 57495 3690
rect 57455 3680 57460 3685
rect 57370 3660 57460 3680
rect 57370 3655 57375 3660
rect 57335 3650 57375 3655
rect 57455 3655 57460 3660
rect 57490 3680 57495 3685
rect 57575 3685 57615 3690
rect 57575 3680 57580 3685
rect 57490 3660 57580 3680
rect 57490 3655 57495 3660
rect 57455 3650 57495 3655
rect 57575 3655 57580 3660
rect 57610 3680 57615 3685
rect 57695 3685 57735 3690
rect 57695 3680 57700 3685
rect 57610 3660 57700 3680
rect 57610 3655 57615 3660
rect 57575 3650 57615 3655
rect 57695 3655 57700 3660
rect 57730 3655 57735 3685
rect 57695 3650 57735 3655
rect 57850 3685 57890 3690
rect 57850 3655 57855 3685
rect 57885 3680 57890 3685
rect 58180 3685 58220 3690
rect 58180 3680 58185 3685
rect 57885 3660 58185 3680
rect 57885 3655 57890 3660
rect 57850 3650 57890 3655
rect 58180 3655 58185 3660
rect 58215 3680 58220 3685
rect 58300 3685 58340 3690
rect 58300 3680 58305 3685
rect 58215 3660 58305 3680
rect 58215 3655 58220 3660
rect 58180 3650 58220 3655
rect 58300 3655 58305 3660
rect 58335 3680 58340 3685
rect 58420 3685 58460 3690
rect 58420 3680 58425 3685
rect 58335 3660 58425 3680
rect 58335 3655 58340 3660
rect 58300 3650 58340 3655
rect 58420 3655 58425 3660
rect 58455 3680 58460 3685
rect 58540 3685 58580 3690
rect 58540 3680 58545 3685
rect 58455 3660 58545 3680
rect 58455 3655 58460 3660
rect 58420 3650 58460 3655
rect 58540 3655 58545 3660
rect 58575 3680 58580 3685
rect 58660 3685 58700 3690
rect 58660 3680 58665 3685
rect 58575 3660 58665 3680
rect 58575 3655 58580 3660
rect 58540 3650 58580 3655
rect 58660 3655 58665 3660
rect 58695 3680 58700 3685
rect 58780 3685 58820 3690
rect 58780 3680 58785 3685
rect 58695 3660 58785 3680
rect 58695 3655 58700 3660
rect 58660 3650 58700 3655
rect 58780 3655 58785 3660
rect 58815 3655 58820 3685
rect 58780 3650 58820 3655
rect 56365 3605 56405 3610
rect 56365 3575 56370 3605
rect 56400 3600 56405 3605
rect 56835 3605 56875 3610
rect 56835 3600 56840 3605
rect 56400 3580 56840 3600
rect 56400 3575 56405 3580
rect 56365 3570 56405 3575
rect 56835 3575 56840 3580
rect 56870 3600 56875 3605
rect 57395 3605 57435 3610
rect 57395 3600 57400 3605
rect 56870 3580 57400 3600
rect 56870 3575 56875 3580
rect 56835 3570 56875 3575
rect 57395 3575 57400 3580
rect 57430 3575 57435 3605
rect 57395 3570 57435 3575
rect 55285 3560 55325 3565
rect 55285 3530 55290 3560
rect 55320 3555 55325 3560
rect 56925 3560 56965 3565
rect 56925 3555 56930 3560
rect 55320 3535 56930 3555
rect 55320 3530 55325 3535
rect 55285 3525 55325 3530
rect 56925 3530 56930 3535
rect 56960 3555 56965 3560
rect 58480 3560 58520 3565
rect 58480 3555 58485 3560
rect 56960 3535 58485 3555
rect 56960 3530 56965 3535
rect 56925 3525 56965 3530
rect 58480 3530 58485 3535
rect 58515 3530 58520 3560
rect 58480 3525 58520 3530
rect 54605 3400 54645 3405
rect 54605 3370 54610 3400
rect 54640 3370 54645 3400
rect 59155 3400 59195 3405
rect 54605 3365 54645 3370
rect 54955 3380 54995 3385
rect 54955 3350 54960 3380
rect 54990 3375 54995 3380
rect 55065 3380 55105 3385
rect 55065 3375 55070 3380
rect 54990 3355 55070 3375
rect 54990 3350 54995 3355
rect 54955 3345 54995 3350
rect 55065 3350 55070 3355
rect 55100 3375 55105 3380
rect 55175 3380 55215 3385
rect 55175 3375 55180 3380
rect 55100 3355 55180 3375
rect 55100 3350 55105 3355
rect 55065 3345 55105 3350
rect 55175 3350 55180 3355
rect 55210 3375 55215 3380
rect 55285 3380 55325 3385
rect 55285 3375 55290 3380
rect 55210 3355 55290 3375
rect 55210 3350 55215 3355
rect 55175 3345 55215 3350
rect 55285 3350 55290 3355
rect 55320 3375 55325 3380
rect 55395 3380 55435 3385
rect 55395 3375 55400 3380
rect 55320 3355 55400 3375
rect 55320 3350 55325 3355
rect 55285 3345 55325 3350
rect 55395 3350 55400 3355
rect 55430 3375 55435 3380
rect 55505 3380 55545 3385
rect 55505 3375 55510 3380
rect 55430 3355 55510 3375
rect 55430 3350 55435 3355
rect 55395 3345 55435 3350
rect 55505 3350 55510 3355
rect 55540 3375 55545 3380
rect 55615 3380 55655 3385
rect 55615 3375 55620 3380
rect 55540 3355 55620 3375
rect 55540 3350 55545 3355
rect 55505 3345 55545 3350
rect 55615 3350 55620 3355
rect 55650 3375 55655 3380
rect 55760 3380 55800 3385
rect 55760 3375 55765 3380
rect 55650 3355 55765 3375
rect 55650 3350 55655 3355
rect 55615 3345 55655 3350
rect 55760 3350 55765 3355
rect 55795 3350 55800 3380
rect 55760 3345 55800 3350
rect 56275 3380 56315 3385
rect 56275 3350 56280 3380
rect 56310 3375 56315 3380
rect 56385 3380 56425 3385
rect 56385 3375 56390 3380
rect 56310 3355 56390 3375
rect 56310 3350 56315 3355
rect 56275 3345 56315 3350
rect 56385 3350 56390 3355
rect 56420 3375 56425 3380
rect 56495 3380 56535 3385
rect 56495 3375 56500 3380
rect 56420 3355 56500 3375
rect 56420 3350 56425 3355
rect 56385 3345 56425 3350
rect 56495 3350 56500 3355
rect 56530 3375 56535 3380
rect 56605 3380 56645 3385
rect 56605 3375 56610 3380
rect 56530 3355 56610 3375
rect 56530 3350 56535 3355
rect 56495 3345 56535 3350
rect 56605 3350 56610 3355
rect 56640 3375 56645 3380
rect 56715 3380 56755 3385
rect 56715 3375 56720 3380
rect 56640 3355 56720 3375
rect 56640 3350 56645 3355
rect 56605 3345 56645 3350
rect 56715 3350 56720 3355
rect 56750 3375 56755 3380
rect 56825 3380 56865 3385
rect 56825 3375 56830 3380
rect 56750 3355 56830 3375
rect 56750 3350 56755 3355
rect 56715 3345 56755 3350
rect 56825 3350 56830 3355
rect 56860 3375 56865 3380
rect 56935 3380 56975 3385
rect 56935 3375 56940 3380
rect 56860 3355 56940 3375
rect 56860 3350 56865 3355
rect 56825 3345 56865 3350
rect 56935 3350 56940 3355
rect 56970 3375 56975 3380
rect 57045 3380 57085 3385
rect 57045 3375 57050 3380
rect 56970 3355 57050 3375
rect 56970 3350 56975 3355
rect 56935 3345 56975 3350
rect 57045 3350 57050 3355
rect 57080 3375 57085 3380
rect 57155 3380 57195 3385
rect 57155 3375 57160 3380
rect 57080 3355 57160 3375
rect 57080 3350 57085 3355
rect 57045 3345 57085 3350
rect 57155 3350 57160 3355
rect 57190 3375 57195 3380
rect 57265 3380 57305 3385
rect 57265 3375 57270 3380
rect 57190 3355 57270 3375
rect 57190 3350 57195 3355
rect 57155 3345 57195 3350
rect 57265 3350 57270 3355
rect 57300 3375 57305 3380
rect 57375 3380 57415 3385
rect 57375 3375 57380 3380
rect 57300 3355 57380 3375
rect 57300 3350 57305 3355
rect 57265 3345 57305 3350
rect 57375 3350 57380 3355
rect 57410 3375 57415 3380
rect 57485 3380 57525 3385
rect 57485 3375 57490 3380
rect 57410 3355 57490 3375
rect 57410 3350 57415 3355
rect 57375 3345 57415 3350
rect 57485 3350 57490 3355
rect 57520 3375 57525 3380
rect 58005 3380 58045 3385
rect 58005 3375 58010 3380
rect 57520 3355 58010 3375
rect 57520 3350 57525 3355
rect 57485 3345 57525 3350
rect 58005 3350 58010 3355
rect 58040 3375 58045 3380
rect 58150 3380 58190 3385
rect 58150 3375 58155 3380
rect 58040 3355 58155 3375
rect 58040 3350 58045 3355
rect 58005 3345 58045 3350
rect 58150 3350 58155 3355
rect 58185 3375 58190 3380
rect 58260 3380 58300 3385
rect 58260 3375 58265 3380
rect 58185 3355 58265 3375
rect 58185 3350 58190 3355
rect 58150 3345 58190 3350
rect 58260 3350 58265 3355
rect 58295 3375 58300 3380
rect 58370 3380 58410 3385
rect 58370 3375 58375 3380
rect 58295 3355 58375 3375
rect 58295 3350 58300 3355
rect 58260 3345 58300 3350
rect 58370 3350 58375 3355
rect 58405 3375 58410 3380
rect 58480 3380 58520 3385
rect 58480 3375 58485 3380
rect 58405 3355 58485 3375
rect 58405 3350 58410 3355
rect 58370 3345 58410 3350
rect 58480 3350 58485 3355
rect 58515 3375 58520 3380
rect 58590 3380 58630 3385
rect 58590 3375 58595 3380
rect 58515 3355 58595 3375
rect 58515 3350 58520 3355
rect 58480 3345 58520 3350
rect 58590 3350 58595 3355
rect 58625 3375 58630 3380
rect 58700 3380 58740 3385
rect 58700 3375 58705 3380
rect 58625 3355 58705 3375
rect 58625 3350 58630 3355
rect 58590 3345 58630 3350
rect 58700 3350 58705 3355
rect 58735 3375 58740 3380
rect 58810 3380 58850 3385
rect 58810 3375 58815 3380
rect 58735 3355 58815 3375
rect 58735 3350 58740 3355
rect 58700 3345 58740 3350
rect 58810 3350 58815 3355
rect 58845 3350 58850 3380
rect 59155 3370 59160 3400
rect 59190 3370 59195 3400
rect 59155 3365 59195 3370
rect 58810 3345 58850 3350
rect 56330 3335 56370 3340
rect 55715 3325 55755 3330
rect 55010 3300 55050 3305
rect 55010 3270 55015 3300
rect 55045 3295 55050 3300
rect 55120 3300 55160 3305
rect 55120 3295 55125 3300
rect 55045 3275 55125 3295
rect 55045 3270 55050 3275
rect 55010 3265 55050 3270
rect 55120 3270 55125 3275
rect 55155 3295 55160 3300
rect 55230 3300 55270 3305
rect 55230 3295 55235 3300
rect 55155 3275 55235 3295
rect 55155 3270 55160 3275
rect 55120 3265 55160 3270
rect 55230 3270 55235 3275
rect 55265 3295 55270 3300
rect 55340 3300 55380 3305
rect 55340 3295 55345 3300
rect 55265 3275 55345 3295
rect 55265 3270 55270 3275
rect 55230 3265 55270 3270
rect 55340 3270 55345 3275
rect 55375 3295 55380 3300
rect 55450 3300 55490 3305
rect 55450 3295 55455 3300
rect 55375 3275 55455 3295
rect 55375 3270 55380 3275
rect 55340 3265 55380 3270
rect 55450 3270 55455 3275
rect 55485 3295 55490 3300
rect 55560 3300 55600 3305
rect 55560 3295 55565 3300
rect 55485 3275 55565 3295
rect 55485 3270 55490 3275
rect 55450 3265 55490 3270
rect 55560 3270 55565 3275
rect 55595 3270 55600 3300
rect 55715 3295 55720 3325
rect 55750 3320 55755 3325
rect 56065 3325 56105 3330
rect 56065 3320 56070 3325
rect 55750 3300 56070 3320
rect 55750 3295 55755 3300
rect 55715 3290 55755 3295
rect 56065 3295 56070 3300
rect 56100 3295 56105 3325
rect 56330 3305 56335 3335
rect 56365 3330 56370 3335
rect 56550 3335 56590 3340
rect 56550 3330 56555 3335
rect 56365 3310 56555 3330
rect 56365 3305 56370 3310
rect 56330 3300 56370 3305
rect 56550 3305 56555 3310
rect 56585 3330 56590 3335
rect 56770 3335 56810 3340
rect 56770 3330 56775 3335
rect 56585 3310 56775 3330
rect 56585 3305 56590 3310
rect 56550 3300 56590 3305
rect 56770 3305 56775 3310
rect 56805 3330 56810 3335
rect 56990 3335 57030 3340
rect 56990 3330 56995 3335
rect 56805 3310 56995 3330
rect 56805 3305 56810 3310
rect 56770 3300 56810 3305
rect 56990 3305 56995 3310
rect 57025 3330 57030 3335
rect 57210 3335 57250 3340
rect 57210 3330 57215 3335
rect 57025 3310 57215 3330
rect 57025 3305 57030 3310
rect 56990 3300 57030 3305
rect 57210 3305 57215 3310
rect 57245 3330 57250 3335
rect 57430 3335 57470 3340
rect 57430 3330 57435 3335
rect 57245 3310 57435 3330
rect 57245 3305 57250 3310
rect 57210 3300 57250 3305
rect 57430 3305 57435 3310
rect 57465 3305 57470 3335
rect 57430 3300 57470 3305
rect 57695 3325 57735 3330
rect 57695 3295 57700 3325
rect 57730 3320 57735 3325
rect 58050 3325 58090 3330
rect 58050 3320 58055 3325
rect 57730 3300 58055 3320
rect 57730 3295 57735 3300
rect 56065 3290 56105 3295
rect 56440 3290 56480 3295
rect 55560 3265 55600 3270
rect 56440 3260 56445 3290
rect 56475 3285 56480 3290
rect 56660 3290 56700 3295
rect 56660 3285 56665 3290
rect 56475 3265 56665 3285
rect 56475 3260 56480 3265
rect 56440 3255 56480 3260
rect 56660 3260 56665 3265
rect 56695 3285 56700 3290
rect 56880 3290 56920 3295
rect 56880 3285 56885 3290
rect 56695 3265 56885 3285
rect 56695 3260 56700 3265
rect 56660 3255 56700 3260
rect 56880 3260 56885 3265
rect 56915 3285 56920 3290
rect 57100 3290 57140 3295
rect 57100 3285 57105 3290
rect 56915 3265 57105 3285
rect 56915 3260 56920 3265
rect 56880 3255 56920 3260
rect 57100 3260 57105 3265
rect 57135 3285 57140 3290
rect 57320 3290 57360 3295
rect 57695 3290 57735 3295
rect 58050 3295 58055 3300
rect 58085 3295 58090 3325
rect 58050 3290 58090 3295
rect 58205 3300 58245 3305
rect 57320 3285 57325 3290
rect 57135 3265 57325 3285
rect 57135 3260 57140 3265
rect 57100 3255 57140 3260
rect 57320 3260 57325 3265
rect 57355 3260 57360 3290
rect 58205 3270 58210 3300
rect 58240 3295 58245 3300
rect 58315 3300 58355 3305
rect 58315 3295 58320 3300
rect 58240 3275 58320 3295
rect 58240 3270 58245 3275
rect 58205 3265 58245 3270
rect 58315 3270 58320 3275
rect 58350 3295 58355 3300
rect 58425 3300 58465 3305
rect 58425 3295 58430 3300
rect 58350 3275 58430 3295
rect 58350 3270 58355 3275
rect 58315 3265 58355 3270
rect 58425 3270 58430 3275
rect 58460 3295 58465 3300
rect 58535 3300 58575 3305
rect 58535 3295 58540 3300
rect 58460 3275 58540 3295
rect 58460 3270 58465 3275
rect 58425 3265 58465 3270
rect 58535 3270 58540 3275
rect 58570 3295 58575 3300
rect 58645 3300 58685 3305
rect 58645 3295 58650 3300
rect 58570 3275 58650 3295
rect 58570 3270 58575 3275
rect 58535 3265 58575 3270
rect 58645 3270 58650 3275
rect 58680 3295 58685 3300
rect 58755 3300 58795 3305
rect 58755 3295 58760 3300
rect 58680 3275 58760 3295
rect 58680 3270 58685 3275
rect 58645 3265 58685 3270
rect 58755 3270 58760 3275
rect 58790 3270 58795 3300
rect 58755 3265 58795 3270
rect 57320 3255 57360 3260
rect 56330 3200 56370 3205
rect 56330 3170 56335 3200
rect 56365 3195 56370 3200
rect 56550 3200 56590 3205
rect 56550 3195 56555 3200
rect 56365 3175 56555 3195
rect 56365 3170 56370 3175
rect 56330 3165 56370 3170
rect 56550 3170 56555 3175
rect 56585 3195 56590 3200
rect 56770 3200 56810 3205
rect 56770 3195 56775 3200
rect 56585 3175 56775 3195
rect 56585 3170 56590 3175
rect 56550 3165 56590 3170
rect 56770 3170 56775 3175
rect 56805 3195 56810 3200
rect 56990 3200 57030 3205
rect 56990 3195 56995 3200
rect 56805 3175 56995 3195
rect 56805 3170 56810 3175
rect 56770 3165 56810 3170
rect 56990 3170 56995 3175
rect 57025 3195 57030 3200
rect 57210 3200 57250 3205
rect 57210 3195 57215 3200
rect 57025 3175 57215 3195
rect 57025 3170 57030 3175
rect 56990 3165 57030 3170
rect 57210 3170 57215 3175
rect 57245 3195 57250 3200
rect 57430 3200 57470 3205
rect 57430 3195 57435 3200
rect 57245 3175 57435 3195
rect 57245 3170 57250 3175
rect 57210 3165 57250 3170
rect 57430 3170 57435 3175
rect 57465 3170 57470 3200
rect 57430 3165 57470 3170
rect 56440 3130 56480 3135
rect 56440 3100 56445 3130
rect 56475 3125 56480 3130
rect 56660 3130 56700 3135
rect 56660 3125 56665 3130
rect 56475 3105 56665 3125
rect 56475 3100 56480 3105
rect 56440 3095 56480 3100
rect 56660 3100 56665 3105
rect 56695 3125 56700 3130
rect 56880 3130 56920 3135
rect 56880 3125 56885 3130
rect 56695 3105 56885 3125
rect 56695 3100 56700 3105
rect 56660 3095 56700 3100
rect 56880 3100 56885 3105
rect 56915 3125 56920 3130
rect 57100 3130 57140 3135
rect 57100 3125 57105 3130
rect 56915 3105 57105 3125
rect 56915 3100 56920 3105
rect 56880 3095 56920 3100
rect 57100 3100 57105 3105
rect 57135 3125 57140 3130
rect 57320 3130 57360 3135
rect 57320 3125 57325 3130
rect 57135 3105 57325 3125
rect 57135 3100 57140 3105
rect 57100 3095 57140 3100
rect 57320 3100 57325 3105
rect 57355 3100 57360 3130
rect 57320 3095 57360 3100
rect 56140 3025 56180 3030
rect 55940 3020 55980 3025
rect 55940 2990 55945 3020
rect 55975 3015 55980 3020
rect 56040 3020 56070 3025
rect 55975 2995 56040 3015
rect 55975 2990 55980 2995
rect 55940 2985 55980 2990
rect 56140 2995 56145 3025
rect 56175 3020 56180 3025
rect 56250 3025 56290 3030
rect 56250 3020 56255 3025
rect 56175 3000 56255 3020
rect 56175 2995 56180 3000
rect 56140 2990 56180 2995
rect 56250 2995 56255 3000
rect 56285 3020 56290 3025
rect 56360 3025 56400 3030
rect 56360 3020 56365 3025
rect 56285 3000 56365 3020
rect 56285 2995 56290 3000
rect 56250 2990 56290 2995
rect 56360 2995 56365 3000
rect 56395 3020 56400 3025
rect 56470 3025 56510 3030
rect 56470 3020 56475 3025
rect 56395 3000 56475 3020
rect 56395 2995 56400 3000
rect 56360 2990 56400 2995
rect 56470 2995 56475 3000
rect 56505 3020 56510 3025
rect 56580 3025 56620 3030
rect 57180 3025 57220 3030
rect 56580 3020 56585 3025
rect 56505 3000 56585 3020
rect 56505 2995 56510 3000
rect 56470 2990 56510 2995
rect 56580 2995 56585 3000
rect 56615 2995 56620 3025
rect 56580 2990 56620 2995
rect 56690 3020 56720 3025
rect 57080 3020 57110 3025
rect 56720 2995 57080 3015
rect 56040 2985 56070 2990
rect 56690 2985 56720 2990
rect 57180 2995 57185 3025
rect 57215 3020 57220 3025
rect 57290 3025 57330 3030
rect 57290 3020 57295 3025
rect 57215 3000 57295 3020
rect 57215 2995 57220 3000
rect 57180 2990 57220 2995
rect 57290 2995 57295 3000
rect 57325 3020 57330 3025
rect 57400 3025 57440 3030
rect 57400 3020 57405 3025
rect 57325 3000 57405 3020
rect 57325 2995 57330 3000
rect 57290 2990 57330 2995
rect 57400 2995 57405 3000
rect 57435 3020 57440 3025
rect 57510 3025 57550 3030
rect 57510 3020 57515 3025
rect 57435 3000 57515 3020
rect 57435 2995 57440 3000
rect 57400 2990 57440 2995
rect 57510 2995 57515 3000
rect 57545 3020 57550 3025
rect 57620 3025 57660 3030
rect 57620 3020 57625 3025
rect 57545 3000 57625 3020
rect 57545 2995 57550 3000
rect 57510 2990 57550 2995
rect 57620 2995 57625 3000
rect 57655 2995 57660 3025
rect 57620 2990 57660 2995
rect 57730 3020 57760 3025
rect 57820 3020 57860 3025
rect 57820 3015 57825 3020
rect 57760 2995 57825 3015
rect 57080 2985 57110 2990
rect 57730 2985 57760 2990
rect 57820 2990 57825 2995
rect 57855 2990 57860 3020
rect 57820 2985 57860 2990
rect 56085 2980 56125 2985
rect 56085 2950 56090 2980
rect 56120 2975 56125 2980
rect 56195 2980 56235 2985
rect 56195 2975 56200 2980
rect 56120 2955 56200 2975
rect 56120 2950 56125 2955
rect 56085 2945 56125 2950
rect 56195 2950 56200 2955
rect 56230 2975 56235 2980
rect 56305 2980 56345 2985
rect 56305 2975 56310 2980
rect 56230 2955 56310 2975
rect 56230 2950 56235 2955
rect 56195 2945 56235 2950
rect 56305 2950 56310 2955
rect 56340 2975 56345 2980
rect 56415 2980 56455 2985
rect 56415 2975 56420 2980
rect 56340 2955 56420 2975
rect 56340 2950 56345 2955
rect 56305 2945 56345 2950
rect 56415 2950 56420 2955
rect 56450 2975 56455 2980
rect 56525 2980 56565 2985
rect 56525 2975 56530 2980
rect 56450 2955 56530 2975
rect 56450 2950 56455 2955
rect 56415 2945 56455 2950
rect 56525 2950 56530 2955
rect 56560 2975 56565 2980
rect 56635 2980 56675 2985
rect 56635 2975 56640 2980
rect 56560 2955 56640 2975
rect 56560 2950 56565 2955
rect 56525 2945 56565 2950
rect 56635 2950 56640 2955
rect 56670 2950 56675 2980
rect 56635 2945 56675 2950
rect 57125 2980 57165 2985
rect 57125 2950 57130 2980
rect 57160 2975 57165 2980
rect 57345 2980 57385 2985
rect 57345 2975 57350 2980
rect 57160 2955 57350 2975
rect 57160 2950 57165 2955
rect 57125 2945 57165 2950
rect 57345 2950 57350 2955
rect 57380 2975 57385 2980
rect 57565 2980 57605 2985
rect 57565 2975 57570 2980
rect 57380 2955 57570 2975
rect 57380 2950 57385 2955
rect 57345 2945 57385 2950
rect 57565 2950 57570 2955
rect 57600 2950 57605 2980
rect 57565 2945 57605 2950
rect 56140 2890 56180 2895
rect 56140 2860 56145 2890
rect 56175 2885 56180 2890
rect 56250 2890 56290 2895
rect 56250 2885 56255 2890
rect 56175 2865 56255 2885
rect 56175 2860 56180 2865
rect 56140 2855 56180 2860
rect 56250 2860 56255 2865
rect 56285 2885 56290 2890
rect 56360 2890 56400 2895
rect 56360 2885 56365 2890
rect 56285 2865 56365 2885
rect 56285 2860 56290 2865
rect 56250 2855 56290 2860
rect 56360 2860 56365 2865
rect 56395 2885 56400 2890
rect 56470 2890 56510 2895
rect 56470 2885 56475 2890
rect 56395 2865 56475 2885
rect 56395 2860 56400 2865
rect 56360 2855 56400 2860
rect 56470 2860 56475 2865
rect 56505 2885 56510 2890
rect 56580 2890 56620 2895
rect 56580 2885 56585 2890
rect 56505 2865 56585 2885
rect 56505 2860 56510 2865
rect 56470 2855 56510 2860
rect 56580 2860 56585 2865
rect 56615 2860 56620 2890
rect 56580 2855 56620 2860
rect 57180 2890 57220 2895
rect 57180 2860 57185 2890
rect 57215 2885 57220 2890
rect 57290 2890 57330 2895
rect 57290 2885 57295 2890
rect 57215 2865 57295 2885
rect 57215 2860 57220 2865
rect 57180 2855 57220 2860
rect 57290 2860 57295 2865
rect 57325 2885 57330 2890
rect 57400 2890 57440 2895
rect 57400 2885 57405 2890
rect 57325 2865 57405 2885
rect 57325 2860 57330 2865
rect 57290 2855 57330 2860
rect 57400 2860 57405 2865
rect 57435 2885 57440 2890
rect 57510 2890 57550 2895
rect 57510 2885 57515 2890
rect 57435 2865 57515 2885
rect 57435 2860 57440 2865
rect 57400 2855 57440 2860
rect 57510 2860 57515 2865
rect 57545 2885 57550 2890
rect 57620 2890 57660 2895
rect 57620 2885 57625 2890
rect 57545 2865 57625 2885
rect 57545 2860 57550 2865
rect 57510 2855 57550 2860
rect 57620 2860 57625 2865
rect 57655 2860 57660 2890
rect 57620 2855 57660 2860
rect 56085 2845 56125 2850
rect 56085 2815 56090 2845
rect 56120 2840 56125 2845
rect 56195 2845 56235 2850
rect 56195 2840 56200 2845
rect 56120 2820 56200 2840
rect 56120 2815 56125 2820
rect 56085 2810 56125 2815
rect 56195 2815 56200 2820
rect 56230 2840 56235 2845
rect 56305 2845 56345 2850
rect 56305 2840 56310 2845
rect 56230 2820 56310 2840
rect 56230 2815 56235 2820
rect 56195 2810 56235 2815
rect 56305 2815 56310 2820
rect 56340 2840 56345 2845
rect 56415 2845 56455 2850
rect 56415 2840 56420 2845
rect 56340 2820 56420 2840
rect 56340 2815 56345 2820
rect 56305 2810 56345 2815
rect 56415 2815 56420 2820
rect 56450 2840 56455 2845
rect 56525 2845 56565 2850
rect 56525 2840 56530 2845
rect 56450 2820 56530 2840
rect 56450 2815 56455 2820
rect 56415 2810 56455 2815
rect 56525 2815 56530 2820
rect 56560 2840 56565 2845
rect 56635 2845 56675 2850
rect 56635 2840 56640 2845
rect 56560 2820 56640 2840
rect 56560 2815 56565 2820
rect 56525 2810 56565 2815
rect 56635 2815 56640 2820
rect 56670 2840 56675 2845
rect 56825 2845 56865 2850
rect 56825 2840 56830 2845
rect 56670 2820 56830 2840
rect 56670 2815 56675 2820
rect 56635 2810 56675 2815
rect 56825 2815 56830 2820
rect 56860 2815 56865 2845
rect 56825 2810 56865 2815
rect 57125 2845 57165 2850
rect 57125 2815 57130 2845
rect 57160 2840 57165 2845
rect 57345 2845 57385 2850
rect 57345 2840 57350 2845
rect 57160 2820 57350 2840
rect 57160 2815 57165 2820
rect 57125 2810 57165 2815
rect 57345 2815 57350 2820
rect 57380 2840 57385 2845
rect 57565 2845 57605 2850
rect 57565 2840 57570 2845
rect 57380 2820 57570 2840
rect 57380 2815 57385 2820
rect 57345 2810 57385 2815
rect 57565 2815 57570 2820
rect 57600 2815 57605 2845
rect 57565 2810 57605 2815
rect 56095 2790 56125 2795
rect 55955 2765 56095 2785
rect 56095 2755 56125 2760
rect 56580 2790 56610 2795
rect 57190 2790 57220 2795
rect 56610 2765 57190 2785
rect 56580 2755 56610 2760
rect 57190 2755 57220 2760
rect 55760 2745 55800 2750
rect 55760 2715 55765 2745
rect 55795 2740 55800 2745
rect 56030 2745 56070 2750
rect 56030 2740 56035 2745
rect 55795 2720 56035 2740
rect 55795 2715 55800 2720
rect 55760 2710 55800 2715
rect 56030 2715 56035 2720
rect 56065 2740 56070 2745
rect 56690 2745 56730 2750
rect 56690 2740 56695 2745
rect 56065 2720 56695 2740
rect 56065 2715 56070 2720
rect 56030 2710 56070 2715
rect 56690 2715 56695 2720
rect 56725 2715 56730 2745
rect 56690 2710 56730 2715
rect 57070 2745 57110 2750
rect 57070 2715 57075 2745
rect 57105 2740 57110 2745
rect 57730 2745 57770 2750
rect 57730 2740 57735 2745
rect 57105 2720 57735 2740
rect 57105 2715 57110 2720
rect 57070 2710 57110 2715
rect 57730 2715 57735 2720
rect 57765 2740 57770 2745
rect 58005 2745 58045 2750
rect 58005 2740 58010 2745
rect 57765 2720 58010 2740
rect 57765 2715 57770 2720
rect 57730 2710 57770 2715
rect 58005 2715 58010 2720
rect 58040 2715 58045 2745
rect 58005 2710 58045 2715
rect 56605 2690 56645 2695
rect 55010 2660 55050 2665
rect 55010 2630 55015 2660
rect 55045 2655 55050 2660
rect 55120 2660 55160 2665
rect 55120 2655 55125 2660
rect 55045 2635 55125 2655
rect 55045 2630 55050 2635
rect 55010 2625 55050 2630
rect 55120 2630 55125 2635
rect 55155 2655 55160 2660
rect 55230 2660 55270 2665
rect 55230 2655 55235 2660
rect 55155 2635 55235 2655
rect 55155 2630 55160 2635
rect 55120 2625 55160 2630
rect 55230 2630 55235 2635
rect 55265 2655 55270 2660
rect 55340 2660 55380 2665
rect 55340 2655 55345 2660
rect 55265 2635 55345 2655
rect 55265 2630 55270 2635
rect 55230 2625 55270 2630
rect 55340 2630 55345 2635
rect 55375 2655 55380 2660
rect 55450 2660 55490 2665
rect 55450 2655 55455 2660
rect 55375 2635 55455 2655
rect 55375 2630 55380 2635
rect 55340 2625 55380 2630
rect 55450 2630 55455 2635
rect 55485 2655 55490 2660
rect 55560 2660 55600 2665
rect 55560 2655 55565 2660
rect 55485 2635 55565 2655
rect 55485 2630 55490 2635
rect 55450 2625 55490 2630
rect 55560 2630 55565 2635
rect 55595 2630 55600 2660
rect 56605 2660 56610 2690
rect 56640 2685 56645 2690
rect 56825 2690 56865 2695
rect 56825 2685 56830 2690
rect 56640 2665 56830 2685
rect 56640 2660 56645 2665
rect 56605 2655 56645 2660
rect 56825 2660 56830 2665
rect 56860 2685 56865 2690
rect 57045 2690 57085 2695
rect 57045 2685 57050 2690
rect 56860 2665 57050 2685
rect 56860 2660 56865 2665
rect 56825 2655 56865 2660
rect 57045 2660 57050 2665
rect 57080 2685 57085 2690
rect 57235 2690 57275 2695
rect 57235 2685 57240 2690
rect 57080 2665 57240 2685
rect 57080 2660 57085 2665
rect 57045 2655 57085 2660
rect 57235 2660 57240 2665
rect 57270 2685 57275 2690
rect 57455 2690 57495 2695
rect 57455 2685 57460 2690
rect 57270 2665 57460 2685
rect 57270 2660 57275 2665
rect 57235 2655 57275 2660
rect 57455 2660 57460 2665
rect 57490 2685 57495 2690
rect 57675 2690 57715 2695
rect 57675 2685 57680 2690
rect 57490 2665 57680 2685
rect 57490 2660 57495 2665
rect 57455 2655 57495 2660
rect 57675 2660 57680 2665
rect 57710 2660 57715 2690
rect 57675 2655 57715 2660
rect 58205 2660 58245 2665
rect 55560 2625 55600 2630
rect 56715 2635 56755 2640
rect 56715 2605 56720 2635
rect 56750 2630 56755 2635
rect 56935 2635 56975 2640
rect 56935 2630 56940 2635
rect 56750 2610 56940 2630
rect 56750 2605 56755 2610
rect 56715 2600 56755 2605
rect 56935 2605 56940 2610
rect 56970 2630 56975 2635
rect 57155 2635 57195 2640
rect 57155 2630 57160 2635
rect 56970 2610 57160 2630
rect 56970 2605 56975 2610
rect 56935 2600 56975 2605
rect 57155 2605 57160 2610
rect 57190 2630 57195 2635
rect 57345 2635 57385 2640
rect 57345 2630 57350 2635
rect 57190 2610 57350 2630
rect 57190 2605 57195 2610
rect 57155 2600 57195 2605
rect 57345 2605 57350 2610
rect 57380 2605 57385 2635
rect 58205 2630 58210 2660
rect 58240 2655 58245 2660
rect 58315 2660 58355 2665
rect 58315 2655 58320 2660
rect 58240 2635 58320 2655
rect 58240 2630 58245 2635
rect 58205 2625 58245 2630
rect 58315 2630 58320 2635
rect 58350 2655 58355 2660
rect 58425 2660 58465 2665
rect 58425 2655 58430 2660
rect 58350 2635 58430 2655
rect 58350 2630 58355 2635
rect 58315 2625 58355 2630
rect 58425 2630 58430 2635
rect 58460 2655 58465 2660
rect 58535 2660 58575 2665
rect 58535 2655 58540 2660
rect 58460 2635 58540 2655
rect 58460 2630 58465 2635
rect 58425 2625 58465 2630
rect 58535 2630 58540 2635
rect 58570 2655 58575 2660
rect 58645 2660 58685 2665
rect 58645 2655 58650 2660
rect 58570 2635 58650 2655
rect 58570 2630 58575 2635
rect 58535 2625 58575 2630
rect 58645 2630 58650 2635
rect 58680 2655 58685 2660
rect 58755 2660 58795 2665
rect 58755 2655 58760 2660
rect 58680 2635 58760 2655
rect 58680 2630 58685 2635
rect 58645 2625 58685 2630
rect 58755 2630 58760 2635
rect 58790 2630 58795 2660
rect 58755 2625 58795 2630
rect 57345 2600 57385 2605
rect 54605 2590 54645 2595
rect 54605 2560 54610 2590
rect 54640 2585 54645 2590
rect 55715 2590 55755 2595
rect 55715 2585 55720 2590
rect 54640 2565 55180 2585
rect 54640 2560 54645 2565
rect 54605 2555 54645 2560
rect 55175 2555 55180 2565
rect 55210 2565 55720 2585
rect 55210 2555 55215 2565
rect 55715 2560 55720 2565
rect 55750 2585 55755 2590
rect 56305 2590 56345 2595
rect 56305 2585 56310 2590
rect 55750 2565 56310 2585
rect 55750 2560 55755 2565
rect 55715 2555 55755 2560
rect 56305 2560 56310 2565
rect 56340 2560 56345 2590
rect 56305 2555 56345 2560
rect 57455 2590 57495 2595
rect 57455 2560 57460 2590
rect 57490 2585 57495 2590
rect 58050 2590 58090 2595
rect 58050 2585 58055 2590
rect 57490 2565 58055 2585
rect 57490 2560 57495 2565
rect 57455 2555 57495 2560
rect 58050 2560 58055 2565
rect 58085 2585 58090 2590
rect 59155 2590 59195 2595
rect 59155 2585 59160 2590
rect 58085 2565 58595 2585
rect 58085 2560 58090 2565
rect 58050 2555 58090 2560
rect 58590 2555 58595 2565
rect 58625 2565 59160 2585
rect 58625 2555 58630 2565
rect 59155 2560 59160 2565
rect 59190 2560 59195 2590
rect 59155 2555 59195 2560
rect 54295 2545 54335 2550
rect 54295 2515 54300 2545
rect 54330 2540 54335 2545
rect 55450 2545 55490 2550
rect 55450 2540 55455 2545
rect 54330 2520 55455 2540
rect 54330 2515 54335 2520
rect 54295 2510 54335 2515
rect 55450 2515 55455 2520
rect 55485 2515 55490 2545
rect 58315 2545 58355 2550
rect 55450 2510 55490 2515
rect 56550 2515 56590 2520
rect 54955 2495 54995 2500
rect 54955 2465 54960 2495
rect 54990 2490 54995 2495
rect 55615 2495 55655 2500
rect 55615 2490 55620 2495
rect 54990 2470 55620 2490
rect 54990 2465 54995 2470
rect 54955 2460 54995 2465
rect 55615 2465 55620 2470
rect 55650 2490 55655 2495
rect 55760 2495 55800 2500
rect 55760 2490 55765 2495
rect 55650 2470 55765 2490
rect 55650 2465 55655 2470
rect 55615 2460 55655 2465
rect 55760 2465 55765 2470
rect 55795 2465 55800 2495
rect 56550 2485 56555 2515
rect 56585 2510 56590 2515
rect 56660 2515 56700 2520
rect 56660 2510 56665 2515
rect 56585 2490 56665 2510
rect 56585 2485 56590 2490
rect 56550 2480 56590 2485
rect 56660 2485 56665 2490
rect 56695 2510 56700 2515
rect 56770 2515 56810 2520
rect 56770 2510 56775 2515
rect 56695 2490 56775 2510
rect 56695 2485 56700 2490
rect 56660 2480 56700 2485
rect 56770 2485 56775 2490
rect 56805 2510 56810 2515
rect 56880 2515 56920 2520
rect 56880 2510 56885 2515
rect 56805 2490 56885 2510
rect 56805 2485 56810 2490
rect 56770 2480 56810 2485
rect 56880 2485 56885 2490
rect 56915 2510 56920 2515
rect 56990 2515 57030 2520
rect 56990 2510 56995 2515
rect 56915 2490 56995 2510
rect 56915 2485 56920 2490
rect 56880 2480 56920 2485
rect 56990 2485 56995 2490
rect 57025 2510 57030 2515
rect 57100 2515 57140 2520
rect 57100 2510 57105 2515
rect 57025 2490 57105 2510
rect 57025 2485 57030 2490
rect 56990 2480 57030 2485
rect 57100 2485 57105 2490
rect 57135 2510 57140 2515
rect 57210 2515 57250 2520
rect 57210 2510 57215 2515
rect 57135 2490 57215 2510
rect 57135 2485 57140 2490
rect 57100 2480 57140 2485
rect 57210 2485 57215 2490
rect 57245 2510 57250 2515
rect 57910 2515 57950 2520
rect 57910 2510 57915 2515
rect 57245 2490 57915 2510
rect 57245 2485 57250 2490
rect 57210 2480 57250 2485
rect 57910 2485 57915 2490
rect 57945 2485 57950 2515
rect 58315 2515 58320 2545
rect 58350 2540 58355 2545
rect 59465 2545 59505 2550
rect 59465 2540 59470 2545
rect 58350 2520 59470 2540
rect 58350 2515 58355 2520
rect 58315 2510 58355 2515
rect 59465 2515 59470 2520
rect 59500 2515 59505 2545
rect 59465 2510 59505 2515
rect 57910 2480 57950 2485
rect 58005 2495 58045 2500
rect 58005 2465 58010 2495
rect 58040 2490 58045 2495
rect 58150 2495 58190 2500
rect 58150 2490 58155 2495
rect 58040 2470 58155 2490
rect 58040 2465 58045 2470
rect 55760 2460 55800 2465
rect 56605 2460 56645 2465
rect 54245 2450 54285 2455
rect 54245 2420 54250 2450
rect 54280 2445 54285 2450
rect 55010 2450 55050 2455
rect 55010 2445 55015 2450
rect 54280 2425 55015 2445
rect 54280 2420 54285 2425
rect 54245 2415 54285 2420
rect 55010 2420 55015 2425
rect 55045 2445 55050 2450
rect 55120 2450 55160 2455
rect 55120 2445 55125 2450
rect 55045 2425 55125 2445
rect 55045 2420 55050 2425
rect 55010 2415 55050 2420
rect 55120 2420 55125 2425
rect 55155 2445 55160 2450
rect 55230 2450 55270 2455
rect 55230 2445 55235 2450
rect 55155 2425 55235 2445
rect 55155 2420 55160 2425
rect 55120 2415 55160 2420
rect 55230 2420 55235 2425
rect 55265 2445 55270 2450
rect 55340 2450 55380 2455
rect 55340 2445 55345 2450
rect 55265 2425 55345 2445
rect 55265 2420 55270 2425
rect 55230 2415 55270 2420
rect 55340 2420 55345 2425
rect 55375 2445 55380 2450
rect 55450 2450 55490 2455
rect 55450 2445 55455 2450
rect 55375 2425 55455 2445
rect 55375 2420 55380 2425
rect 55340 2415 55380 2420
rect 55450 2420 55455 2425
rect 55485 2445 55490 2450
rect 55560 2450 55600 2455
rect 55560 2445 55565 2450
rect 55485 2425 55565 2445
rect 55485 2420 55490 2425
rect 55450 2415 55490 2420
rect 55560 2420 55565 2425
rect 55595 2420 55600 2450
rect 56605 2430 56610 2460
rect 56640 2455 56645 2460
rect 56825 2460 56865 2465
rect 56825 2455 56830 2460
rect 56640 2435 56830 2455
rect 56640 2430 56645 2435
rect 56605 2425 56645 2430
rect 56825 2430 56830 2435
rect 56860 2455 56865 2460
rect 57045 2460 57085 2465
rect 57045 2455 57050 2460
rect 56860 2435 57050 2455
rect 56860 2430 56865 2435
rect 56825 2425 56865 2430
rect 57045 2430 57050 2435
rect 57080 2455 57085 2460
rect 57865 2460 57905 2465
rect 58005 2460 58045 2465
rect 58150 2465 58155 2470
rect 58185 2490 58190 2495
rect 58810 2495 58850 2500
rect 58810 2490 58815 2495
rect 58185 2470 58815 2490
rect 58185 2465 58190 2470
rect 58150 2460 58190 2465
rect 58810 2465 58815 2470
rect 58845 2465 58850 2495
rect 58810 2460 58850 2465
rect 57865 2455 57870 2460
rect 57080 2435 57870 2455
rect 57080 2430 57085 2435
rect 57045 2425 57085 2430
rect 57865 2430 57870 2435
rect 57900 2430 57905 2460
rect 57865 2425 57905 2430
rect 58205 2450 58245 2455
rect 58205 2420 58210 2450
rect 58240 2445 58245 2450
rect 58315 2450 58355 2455
rect 58315 2445 58320 2450
rect 58240 2425 58320 2445
rect 58240 2420 58245 2425
rect 55560 2415 55600 2420
rect 56715 2415 56755 2420
rect 55065 2405 55105 2410
rect 55065 2375 55070 2405
rect 55100 2400 55105 2405
rect 55175 2405 55215 2410
rect 55175 2400 55180 2405
rect 55100 2380 55180 2400
rect 55100 2375 55105 2380
rect 55065 2370 55105 2375
rect 55175 2375 55180 2380
rect 55210 2400 55215 2405
rect 55285 2405 55325 2410
rect 55285 2400 55290 2405
rect 55210 2380 55290 2400
rect 55210 2375 55215 2380
rect 55175 2370 55215 2375
rect 55285 2375 55290 2380
rect 55320 2400 55325 2405
rect 55395 2405 55435 2410
rect 55395 2400 55400 2405
rect 55320 2380 55400 2400
rect 55320 2375 55325 2380
rect 55285 2370 55325 2375
rect 55395 2375 55400 2380
rect 55430 2400 55435 2405
rect 55505 2405 55545 2410
rect 55505 2400 55510 2405
rect 55430 2380 55510 2400
rect 55430 2375 55435 2380
rect 55395 2370 55435 2375
rect 55505 2375 55510 2380
rect 55540 2375 55545 2405
rect 56715 2385 56720 2415
rect 56750 2410 56755 2415
rect 56935 2415 56975 2420
rect 56935 2410 56940 2415
rect 56750 2390 56940 2410
rect 56750 2385 56755 2390
rect 56715 2380 56755 2385
rect 56935 2385 56940 2390
rect 56970 2410 56975 2415
rect 57155 2415 57195 2420
rect 58205 2415 58245 2420
rect 58315 2420 58320 2425
rect 58350 2445 58355 2450
rect 58425 2450 58465 2455
rect 58425 2445 58430 2450
rect 58350 2425 58430 2445
rect 58350 2420 58355 2425
rect 58315 2415 58355 2420
rect 58425 2420 58430 2425
rect 58460 2445 58465 2450
rect 58535 2450 58575 2455
rect 58535 2445 58540 2450
rect 58460 2425 58540 2445
rect 58460 2420 58465 2425
rect 58425 2415 58465 2420
rect 58535 2420 58540 2425
rect 58570 2445 58575 2450
rect 58645 2450 58685 2455
rect 58645 2445 58650 2450
rect 58570 2425 58650 2445
rect 58570 2420 58575 2425
rect 58535 2415 58575 2420
rect 58645 2420 58650 2425
rect 58680 2445 58685 2450
rect 58755 2450 58795 2455
rect 58755 2445 58760 2450
rect 58680 2425 58760 2445
rect 58680 2420 58685 2425
rect 58645 2415 58685 2420
rect 58755 2420 58760 2425
rect 58790 2445 58795 2450
rect 59515 2450 59555 2455
rect 59515 2445 59520 2450
rect 58790 2425 59520 2445
rect 58790 2420 58795 2425
rect 58755 2415 58795 2420
rect 59515 2420 59520 2425
rect 59550 2420 59555 2450
rect 59515 2415 59555 2420
rect 57155 2410 57160 2415
rect 56970 2390 57160 2410
rect 56970 2385 56975 2390
rect 56935 2380 56975 2385
rect 57155 2385 57160 2390
rect 57190 2385 57195 2415
rect 57155 2380 57195 2385
rect 58260 2405 58300 2410
rect 55505 2370 55545 2375
rect 58260 2375 58265 2405
rect 58295 2400 58300 2405
rect 58370 2405 58410 2410
rect 58370 2400 58375 2405
rect 58295 2380 58375 2400
rect 58295 2375 58300 2380
rect 58260 2370 58300 2375
rect 58370 2375 58375 2380
rect 58405 2400 58410 2405
rect 58480 2405 58520 2410
rect 58480 2400 58485 2405
rect 58405 2380 58485 2400
rect 58405 2375 58410 2380
rect 58370 2370 58410 2375
rect 58480 2375 58485 2380
rect 58515 2400 58520 2405
rect 58590 2405 58630 2410
rect 58590 2400 58595 2405
rect 58515 2380 58595 2400
rect 58515 2375 58520 2380
rect 58480 2370 58520 2375
rect 58590 2375 58595 2380
rect 58625 2400 58630 2405
rect 58700 2405 58740 2410
rect 58700 2400 58705 2405
rect 58625 2380 58705 2400
rect 58625 2375 58630 2380
rect 58590 2370 58630 2375
rect 58700 2375 58705 2380
rect 58735 2375 58740 2405
rect 58700 2370 58740 2375
rect 55830 2270 55870 2275
rect 55830 2240 55835 2270
rect 55865 2265 55870 2270
rect 56095 2270 56125 2275
rect 55865 2245 56095 2265
rect 55865 2240 55870 2245
rect 55830 2235 55870 2240
rect 56635 2270 56665 2275
rect 56095 2235 56125 2240
rect 56140 2260 56180 2265
rect 56140 2230 56145 2260
rect 56175 2255 56180 2260
rect 56250 2260 56290 2265
rect 56250 2255 56255 2260
rect 56175 2235 56255 2255
rect 56175 2230 56180 2235
rect 56140 2225 56180 2230
rect 56250 2230 56255 2235
rect 56285 2255 56290 2260
rect 56360 2260 56400 2265
rect 56360 2255 56365 2260
rect 56285 2235 56365 2255
rect 56285 2230 56290 2235
rect 56250 2225 56290 2230
rect 56360 2230 56365 2235
rect 56395 2255 56400 2260
rect 56470 2260 56510 2265
rect 56470 2255 56475 2260
rect 56395 2235 56475 2255
rect 56395 2230 56400 2235
rect 56360 2225 56400 2230
rect 56470 2230 56475 2235
rect 56505 2255 56510 2260
rect 56580 2260 56620 2265
rect 56580 2255 56585 2260
rect 56505 2235 56585 2255
rect 56505 2230 56510 2235
rect 56470 2225 56510 2230
rect 56580 2230 56585 2235
rect 56615 2230 56620 2260
rect 57135 2270 57165 2275
rect 56665 2245 57135 2265
rect 56635 2235 56665 2240
rect 57135 2235 57165 2240
rect 57180 2260 57220 2265
rect 56580 2225 56620 2230
rect 57180 2230 57185 2260
rect 57215 2255 57220 2260
rect 57290 2260 57330 2265
rect 57290 2255 57295 2260
rect 57215 2235 57295 2255
rect 57215 2230 57220 2235
rect 57180 2225 57220 2230
rect 57290 2230 57295 2235
rect 57325 2255 57330 2260
rect 57400 2260 57440 2265
rect 57400 2255 57405 2260
rect 57325 2235 57405 2255
rect 57325 2230 57330 2235
rect 57290 2225 57330 2230
rect 57400 2230 57405 2235
rect 57435 2255 57440 2260
rect 57510 2260 57550 2265
rect 57510 2255 57515 2260
rect 57435 2235 57515 2255
rect 57435 2230 57440 2235
rect 57400 2225 57440 2230
rect 57510 2230 57515 2235
rect 57545 2255 57550 2260
rect 57620 2260 57660 2265
rect 57620 2255 57625 2260
rect 57545 2235 57625 2255
rect 57545 2230 57550 2235
rect 57510 2225 57550 2230
rect 57620 2230 57625 2235
rect 57655 2230 57660 2260
rect 57620 2225 57660 2230
rect 56085 2215 56125 2220
rect 56085 2185 56090 2215
rect 56120 2210 56125 2215
rect 56195 2215 56235 2220
rect 56195 2210 56200 2215
rect 56120 2190 56200 2210
rect 56120 2185 56125 2190
rect 56085 2180 56125 2185
rect 56195 2185 56200 2190
rect 56230 2210 56235 2215
rect 56305 2215 56345 2220
rect 56305 2210 56310 2215
rect 56230 2190 56310 2210
rect 56230 2185 56235 2190
rect 56195 2180 56235 2185
rect 56305 2185 56310 2190
rect 56340 2210 56345 2215
rect 56415 2215 56455 2220
rect 56415 2210 56420 2215
rect 56340 2190 56420 2210
rect 56340 2185 56345 2190
rect 56305 2180 56345 2185
rect 56415 2185 56420 2190
rect 56450 2210 56455 2215
rect 56525 2215 56565 2220
rect 56525 2210 56530 2215
rect 56450 2190 56530 2210
rect 56450 2185 56455 2190
rect 56415 2180 56455 2185
rect 56525 2185 56530 2190
rect 56560 2210 56565 2215
rect 56635 2215 56675 2220
rect 56635 2210 56640 2215
rect 56560 2190 56640 2210
rect 56560 2185 56565 2190
rect 56525 2180 56565 2185
rect 56635 2185 56640 2190
rect 56670 2185 56675 2215
rect 56635 2180 56675 2185
rect 57125 2215 57165 2220
rect 57125 2185 57130 2215
rect 57160 2210 57165 2215
rect 57235 2215 57275 2220
rect 57235 2210 57240 2215
rect 57160 2190 57240 2210
rect 57160 2185 57165 2190
rect 57125 2180 57165 2185
rect 57235 2185 57240 2190
rect 57270 2210 57275 2215
rect 57345 2215 57385 2220
rect 57345 2210 57350 2215
rect 57270 2190 57350 2210
rect 57270 2185 57275 2190
rect 57235 2180 57275 2185
rect 57345 2185 57350 2190
rect 57380 2210 57385 2215
rect 57455 2215 57495 2220
rect 57455 2210 57460 2215
rect 57380 2190 57460 2210
rect 57380 2185 57385 2190
rect 57345 2180 57385 2185
rect 57455 2185 57460 2190
rect 57490 2210 57495 2215
rect 57565 2215 57605 2220
rect 57565 2210 57570 2215
rect 57490 2190 57570 2210
rect 57490 2185 57495 2190
rect 57455 2180 57495 2185
rect 57565 2185 57570 2190
rect 57600 2210 57605 2215
rect 57675 2215 57715 2220
rect 57675 2210 57680 2215
rect 57600 2190 57680 2210
rect 57600 2185 57605 2190
rect 57565 2180 57605 2185
rect 57675 2185 57680 2190
rect 57710 2185 57715 2215
rect 57675 2180 57715 2185
rect 54760 2150 54800 2155
rect 54760 2120 54765 2150
rect 54795 2145 54800 2150
rect 55065 2150 55105 2155
rect 55065 2145 55070 2150
rect 54795 2125 55070 2145
rect 54795 2120 54800 2125
rect 54760 2115 54800 2120
rect 55065 2120 55070 2125
rect 55100 2145 55105 2150
rect 55175 2150 55215 2155
rect 55175 2145 55180 2150
rect 55100 2125 55180 2145
rect 55100 2120 55105 2125
rect 55065 2115 55105 2120
rect 55175 2120 55180 2125
rect 55210 2145 55215 2150
rect 55285 2150 55325 2155
rect 55285 2145 55290 2150
rect 55210 2125 55290 2145
rect 55210 2120 55215 2125
rect 55175 2115 55215 2120
rect 55285 2120 55290 2125
rect 55320 2145 55325 2150
rect 55395 2150 55435 2155
rect 55395 2145 55400 2150
rect 55320 2125 55400 2145
rect 55320 2120 55325 2125
rect 55285 2115 55325 2120
rect 55395 2120 55400 2125
rect 55430 2145 55435 2150
rect 55505 2150 55545 2155
rect 55505 2145 55510 2150
rect 55430 2125 55510 2145
rect 55430 2120 55435 2125
rect 55395 2115 55435 2120
rect 55505 2120 55510 2125
rect 55540 2120 55545 2150
rect 55505 2115 55545 2120
rect 58260 2150 58300 2155
rect 58260 2120 58265 2150
rect 58295 2145 58300 2150
rect 58370 2150 58410 2155
rect 58370 2145 58375 2150
rect 58295 2125 58375 2145
rect 58295 2120 58300 2125
rect 58260 2115 58300 2120
rect 58370 2120 58375 2125
rect 58405 2145 58410 2150
rect 58480 2150 58520 2155
rect 58480 2145 58485 2150
rect 58405 2125 58485 2145
rect 58405 2120 58410 2125
rect 58370 2115 58410 2120
rect 58480 2120 58485 2125
rect 58515 2145 58520 2150
rect 58590 2150 58630 2155
rect 58590 2145 58595 2150
rect 58515 2125 58595 2145
rect 58515 2120 58520 2125
rect 58480 2115 58520 2120
rect 58590 2120 58595 2125
rect 58625 2145 58630 2150
rect 58700 2150 58740 2155
rect 58700 2145 58705 2150
rect 58625 2125 58705 2145
rect 58625 2120 58630 2125
rect 58590 2115 58630 2120
rect 58700 2120 58705 2125
rect 58735 2145 58740 2150
rect 59000 2150 59040 2155
rect 59000 2145 59005 2150
rect 58735 2125 59005 2145
rect 58735 2120 58740 2125
rect 58700 2115 58740 2120
rect 59000 2120 59005 2125
rect 59035 2120 59040 2150
rect 59000 2115 59040 2120
rect 55450 2055 55490 2060
rect 55450 2025 55455 2055
rect 55485 2050 55490 2055
rect 55715 2055 55755 2060
rect 55715 2050 55720 2055
rect 55485 2030 55720 2050
rect 55485 2025 55490 2030
rect 55450 2020 55490 2025
rect 55715 2025 55720 2030
rect 55750 2025 55755 2055
rect 58050 2055 58090 2060
rect 55715 2020 55755 2025
rect 56140 2025 56180 2030
rect 56140 1995 56145 2025
rect 56175 2020 56180 2025
rect 56250 2025 56290 2030
rect 56250 2020 56255 2025
rect 56175 2000 56255 2020
rect 56175 1995 56180 2000
rect 56140 1990 56180 1995
rect 56250 1995 56255 2000
rect 56285 2020 56290 2025
rect 56360 2025 56400 2030
rect 56360 2020 56365 2025
rect 56285 2000 56365 2020
rect 56285 1995 56290 2000
rect 56250 1990 56290 1995
rect 56360 1995 56365 2000
rect 56395 2020 56400 2025
rect 56470 2025 56510 2030
rect 56470 2020 56475 2025
rect 56395 2000 56475 2020
rect 56395 1995 56400 2000
rect 56360 1990 56400 1995
rect 56470 1995 56475 2000
rect 56505 2020 56510 2025
rect 56580 2025 56620 2030
rect 56580 2020 56585 2025
rect 56505 2000 56585 2020
rect 56505 1995 56510 2000
rect 56470 1990 56510 1995
rect 56580 1995 56585 2000
rect 56615 1995 56620 2025
rect 56580 1990 56620 1995
rect 57180 2025 57220 2030
rect 57180 1995 57185 2025
rect 57215 2020 57220 2025
rect 57290 2025 57330 2030
rect 57290 2020 57295 2025
rect 57215 2000 57295 2020
rect 57215 1995 57220 2000
rect 57180 1990 57220 1995
rect 57290 1995 57295 2000
rect 57325 2020 57330 2025
rect 57400 2025 57440 2030
rect 57400 2020 57405 2025
rect 57325 2000 57405 2020
rect 57325 1995 57330 2000
rect 57290 1990 57330 1995
rect 57400 1995 57405 2000
rect 57435 2020 57440 2025
rect 57510 2025 57550 2030
rect 57510 2020 57515 2025
rect 57435 2000 57515 2020
rect 57435 1995 57440 2000
rect 57400 1990 57440 1995
rect 57510 1995 57515 2000
rect 57545 2020 57550 2025
rect 57620 2025 57660 2030
rect 57620 2020 57625 2025
rect 57545 2000 57625 2020
rect 57545 1995 57550 2000
rect 57510 1990 57550 1995
rect 57620 1995 57625 2000
rect 57655 1995 57660 2025
rect 58050 2025 58055 2055
rect 58085 2050 58090 2055
rect 58315 2055 58355 2060
rect 58315 2050 58320 2055
rect 58085 2030 58320 2050
rect 58085 2025 58090 2030
rect 58050 2020 58090 2025
rect 58315 2025 58320 2030
rect 58350 2025 58355 2055
rect 58315 2020 58355 2025
rect 57620 1990 57660 1995
rect 56085 1980 56125 1985
rect 56085 1950 56090 1980
rect 56120 1975 56125 1980
rect 56195 1980 56235 1985
rect 56195 1975 56200 1980
rect 56120 1955 56200 1975
rect 56120 1950 56125 1955
rect 54805 1945 54845 1950
rect 54290 1910 54340 1920
rect 54805 1915 54810 1945
rect 54840 1940 54845 1945
rect 55065 1945 55105 1950
rect 55065 1940 55070 1945
rect 54840 1920 55070 1940
rect 54840 1915 54845 1920
rect 54805 1910 54845 1915
rect 55065 1915 55070 1920
rect 55100 1940 55105 1945
rect 55175 1945 55215 1950
rect 55175 1940 55180 1945
rect 55100 1920 55180 1940
rect 55100 1915 55105 1920
rect 55065 1910 55105 1915
rect 55175 1915 55180 1920
rect 55210 1940 55215 1945
rect 55285 1945 55325 1950
rect 55285 1940 55290 1945
rect 55210 1920 55290 1940
rect 55210 1915 55215 1920
rect 55175 1910 55215 1915
rect 55285 1915 55290 1920
rect 55320 1940 55325 1945
rect 55395 1945 55435 1950
rect 55395 1940 55400 1945
rect 55320 1920 55400 1940
rect 55320 1915 55325 1920
rect 55285 1910 55325 1915
rect 55395 1915 55400 1920
rect 55430 1940 55435 1945
rect 55505 1945 55545 1950
rect 56085 1945 56125 1950
rect 56195 1950 56200 1955
rect 56230 1975 56235 1980
rect 56305 1980 56345 1985
rect 56305 1975 56310 1980
rect 56230 1955 56310 1975
rect 56230 1950 56235 1955
rect 56195 1945 56235 1950
rect 56305 1950 56310 1955
rect 56340 1975 56345 1980
rect 56415 1980 56455 1985
rect 56415 1975 56420 1980
rect 56340 1955 56420 1975
rect 56340 1950 56345 1955
rect 56305 1945 56345 1950
rect 56415 1950 56420 1955
rect 56450 1975 56455 1980
rect 56525 1980 56565 1985
rect 56525 1975 56530 1980
rect 56450 1955 56530 1975
rect 56450 1950 56455 1955
rect 56415 1945 56455 1950
rect 56525 1950 56530 1955
rect 56560 1975 56565 1980
rect 56635 1980 56675 1985
rect 56635 1975 56640 1980
rect 56560 1955 56640 1975
rect 56560 1950 56565 1955
rect 56525 1945 56565 1950
rect 56635 1950 56640 1955
rect 56670 1950 56675 1980
rect 56635 1945 56675 1950
rect 57125 1980 57165 1985
rect 57125 1950 57130 1980
rect 57160 1975 57165 1980
rect 57235 1980 57275 1985
rect 57235 1975 57240 1980
rect 57160 1955 57240 1975
rect 57160 1950 57165 1955
rect 57125 1945 57165 1950
rect 57235 1950 57240 1955
rect 57270 1975 57275 1980
rect 57345 1980 57385 1985
rect 57345 1975 57350 1980
rect 57270 1955 57350 1975
rect 57270 1950 57275 1955
rect 57235 1945 57275 1950
rect 57345 1950 57350 1955
rect 57380 1975 57385 1980
rect 57455 1980 57495 1985
rect 57455 1975 57460 1980
rect 57380 1955 57460 1975
rect 57380 1950 57385 1955
rect 57345 1945 57385 1950
rect 57455 1950 57460 1955
rect 57490 1975 57495 1980
rect 57565 1980 57605 1985
rect 57565 1975 57570 1980
rect 57490 1955 57570 1975
rect 57490 1950 57495 1955
rect 57455 1945 57495 1950
rect 57565 1950 57570 1955
rect 57600 1975 57605 1980
rect 57675 1980 57715 1985
rect 57675 1975 57680 1980
rect 57600 1955 57680 1975
rect 57600 1950 57605 1955
rect 57565 1945 57605 1950
rect 57675 1950 57680 1955
rect 57710 1950 57715 1980
rect 57675 1945 57715 1950
rect 58260 1945 58300 1950
rect 55505 1940 55510 1945
rect 55430 1920 55510 1940
rect 55430 1915 55435 1920
rect 55395 1910 55435 1915
rect 55505 1915 55510 1920
rect 55540 1915 55545 1945
rect 55505 1910 55545 1915
rect 56030 1935 56070 1940
rect 54290 1880 54300 1910
rect 54330 1880 54340 1910
rect 56030 1905 56035 1935
rect 56065 1930 56070 1935
rect 56690 1935 56730 1940
rect 56690 1930 56695 1935
rect 56065 1910 56695 1930
rect 56065 1905 56070 1910
rect 56030 1900 56070 1905
rect 56690 1905 56695 1910
rect 56725 1930 56730 1935
rect 57070 1935 57110 1940
rect 57070 1930 57075 1935
rect 56725 1910 57075 1930
rect 56725 1905 56730 1910
rect 56690 1900 56730 1905
rect 57070 1905 57075 1910
rect 57105 1930 57110 1935
rect 57730 1935 57770 1940
rect 57730 1930 57735 1935
rect 57105 1910 57735 1930
rect 57105 1905 57110 1910
rect 57070 1900 57110 1905
rect 57730 1905 57735 1910
rect 57765 1930 57770 1935
rect 57910 1935 57950 1940
rect 57910 1930 57915 1935
rect 57765 1910 57915 1930
rect 57765 1905 57770 1910
rect 57730 1900 57770 1905
rect 57910 1905 57915 1910
rect 57945 1905 57950 1935
rect 58260 1915 58265 1945
rect 58295 1940 58300 1945
rect 58370 1945 58410 1950
rect 58370 1940 58375 1945
rect 58295 1920 58375 1940
rect 58295 1915 58300 1920
rect 58260 1910 58300 1915
rect 58370 1915 58375 1920
rect 58405 1940 58410 1945
rect 58480 1945 58520 1950
rect 58480 1940 58485 1945
rect 58405 1920 58485 1940
rect 58405 1915 58410 1920
rect 58370 1910 58410 1915
rect 58480 1915 58485 1920
rect 58515 1940 58520 1945
rect 58590 1945 58630 1950
rect 58590 1940 58595 1945
rect 58515 1920 58595 1940
rect 58515 1915 58520 1920
rect 58480 1910 58520 1915
rect 58590 1915 58595 1920
rect 58625 1940 58630 1945
rect 58700 1945 58740 1950
rect 58700 1940 58705 1945
rect 58625 1920 58705 1940
rect 58625 1915 58630 1920
rect 58590 1910 58630 1915
rect 58700 1915 58705 1920
rect 58735 1940 58740 1945
rect 58955 1945 58995 1950
rect 58955 1940 58960 1945
rect 58735 1920 58960 1940
rect 58735 1915 58740 1920
rect 58700 1910 58740 1915
rect 58955 1915 58960 1920
rect 58990 1915 58995 1945
rect 58955 1910 58995 1915
rect 59460 1910 59510 1920
rect 57910 1900 57950 1905
rect 54290 1870 54340 1880
rect 59460 1880 59470 1910
rect 59500 1880 59510 1910
rect 59460 1870 59510 1880
rect 56365 1805 56395 1810
rect 56085 1795 56125 1800
rect 56040 1785 56070 1790
rect 56030 1760 56040 1780
rect 56085 1765 56090 1795
rect 56120 1790 56125 1795
rect 56195 1795 56235 1800
rect 56195 1790 56200 1795
rect 56120 1770 56200 1790
rect 56120 1765 56125 1770
rect 56085 1760 56125 1765
rect 56195 1765 56200 1770
rect 56230 1790 56235 1795
rect 56305 1795 56345 1800
rect 56305 1790 56310 1795
rect 56230 1770 56310 1790
rect 56230 1765 56235 1770
rect 56195 1760 56235 1765
rect 56305 1765 56310 1770
rect 56340 1790 56345 1795
rect 56340 1775 56365 1790
rect 57405 1805 57435 1810
rect 56415 1795 56455 1800
rect 56415 1790 56420 1795
rect 56395 1775 56420 1790
rect 56340 1770 56420 1775
rect 56340 1765 56345 1770
rect 56305 1760 56345 1765
rect 56415 1765 56420 1770
rect 56450 1790 56455 1795
rect 56525 1795 56565 1800
rect 56525 1790 56530 1795
rect 56450 1770 56530 1790
rect 56450 1765 56455 1770
rect 56415 1760 56455 1765
rect 56525 1765 56530 1770
rect 56560 1790 56565 1795
rect 56635 1795 56675 1800
rect 56635 1790 56640 1795
rect 56560 1770 56640 1790
rect 56560 1765 56565 1770
rect 56525 1760 56565 1765
rect 56635 1765 56640 1770
rect 56670 1765 56675 1795
rect 57125 1795 57165 1800
rect 56635 1760 56675 1765
rect 56690 1785 56720 1790
rect 56850 1785 56880 1790
rect 56720 1760 56850 1780
rect 56040 1750 56070 1755
rect 56140 1750 56180 1755
rect 56140 1720 56145 1750
rect 56175 1745 56180 1750
rect 56250 1750 56290 1755
rect 56250 1745 56255 1750
rect 56175 1725 56255 1745
rect 56175 1720 56180 1725
rect 56140 1715 56180 1720
rect 56250 1720 56255 1725
rect 56285 1745 56290 1750
rect 56360 1750 56400 1755
rect 56360 1745 56365 1750
rect 56285 1725 56365 1745
rect 56285 1720 56290 1725
rect 56250 1715 56290 1720
rect 56360 1720 56365 1725
rect 56395 1745 56400 1750
rect 56470 1750 56510 1755
rect 56470 1745 56475 1750
rect 56395 1725 56475 1745
rect 56395 1720 56400 1725
rect 56360 1715 56400 1720
rect 56470 1720 56475 1725
rect 56505 1745 56510 1750
rect 56580 1750 56620 1755
rect 56690 1750 56720 1755
rect 56850 1750 56880 1755
rect 56903 1785 56933 1790
rect 57080 1785 57110 1790
rect 56933 1760 57080 1780
rect 56903 1750 56933 1755
rect 57125 1765 57130 1795
rect 57160 1790 57165 1795
rect 57235 1795 57275 1800
rect 57235 1790 57240 1795
rect 57160 1770 57240 1790
rect 57160 1765 57165 1770
rect 57125 1760 57165 1765
rect 57235 1765 57240 1770
rect 57270 1790 57275 1795
rect 57345 1795 57385 1800
rect 57345 1790 57350 1795
rect 57270 1770 57350 1790
rect 57270 1765 57275 1770
rect 57235 1760 57275 1765
rect 57345 1765 57350 1770
rect 57380 1790 57385 1795
rect 57380 1775 57405 1790
rect 57455 1795 57495 1800
rect 57455 1790 57460 1795
rect 57435 1775 57460 1790
rect 57380 1770 57460 1775
rect 57380 1765 57385 1770
rect 57345 1760 57385 1765
rect 57455 1765 57460 1770
rect 57490 1790 57495 1795
rect 57565 1795 57605 1800
rect 57565 1790 57570 1795
rect 57490 1770 57570 1790
rect 57490 1765 57495 1770
rect 57455 1760 57495 1765
rect 57565 1765 57570 1770
rect 57600 1790 57605 1795
rect 57675 1795 57715 1800
rect 57675 1790 57680 1795
rect 57600 1770 57680 1790
rect 57600 1765 57605 1770
rect 57565 1760 57605 1765
rect 57675 1765 57680 1770
rect 57710 1765 57715 1795
rect 57675 1760 57715 1765
rect 57730 1785 57760 1790
rect 57760 1760 57770 1780
rect 57080 1750 57110 1755
rect 57180 1750 57220 1755
rect 56580 1745 56585 1750
rect 56505 1725 56585 1745
rect 56505 1720 56510 1725
rect 56470 1715 56510 1720
rect 56580 1720 56585 1725
rect 56615 1720 56620 1750
rect 56580 1715 56620 1720
rect 57180 1720 57185 1750
rect 57215 1745 57220 1750
rect 57290 1750 57330 1755
rect 57290 1745 57295 1750
rect 57215 1725 57295 1745
rect 57215 1720 57220 1725
rect 57180 1715 57220 1720
rect 57290 1720 57295 1725
rect 57325 1745 57330 1750
rect 57400 1750 57440 1755
rect 57400 1745 57405 1750
rect 57325 1725 57405 1745
rect 57325 1720 57330 1725
rect 57290 1715 57330 1720
rect 57400 1720 57405 1725
rect 57435 1745 57440 1750
rect 57510 1750 57550 1755
rect 57510 1745 57515 1750
rect 57435 1725 57515 1745
rect 57435 1720 57440 1725
rect 57400 1715 57440 1720
rect 57510 1720 57515 1725
rect 57545 1745 57550 1750
rect 57620 1750 57660 1755
rect 57730 1750 57760 1755
rect 57620 1745 57625 1750
rect 57545 1725 57625 1745
rect 57545 1720 57550 1725
rect 57510 1715 57550 1720
rect 57620 1720 57625 1725
rect 57655 1720 57660 1750
rect 57620 1715 57660 1720
rect 55065 1605 55105 1610
rect 54450 1595 54545 1600
rect 54485 1560 54510 1595
rect 54450 1555 54545 1560
rect 54570 1595 54605 1600
rect 54570 1555 54605 1560
rect 54630 1595 54665 1600
rect 54805 1590 54845 1595
rect 54805 1585 54810 1590
rect 54665 1565 54810 1585
rect 54630 1555 54665 1560
rect 54805 1560 54810 1565
rect 54840 1560 54845 1590
rect 55065 1575 55070 1605
rect 55100 1600 55105 1605
rect 55175 1605 55215 1610
rect 55175 1600 55180 1605
rect 55100 1580 55180 1600
rect 55100 1575 55105 1580
rect 55065 1570 55105 1575
rect 55175 1575 55180 1580
rect 55210 1600 55215 1605
rect 55285 1605 55325 1610
rect 55285 1600 55290 1605
rect 55210 1580 55290 1600
rect 55210 1575 55215 1580
rect 55175 1570 55215 1575
rect 55285 1575 55290 1580
rect 55320 1600 55325 1605
rect 55395 1605 55435 1610
rect 55395 1600 55400 1605
rect 55320 1580 55400 1600
rect 55320 1575 55325 1580
rect 55285 1570 55325 1575
rect 55395 1575 55400 1580
rect 55430 1600 55435 1605
rect 55505 1605 55545 1610
rect 55505 1600 55510 1605
rect 55430 1580 55510 1600
rect 55430 1575 55435 1580
rect 55395 1570 55435 1575
rect 55505 1575 55510 1580
rect 55540 1575 55545 1605
rect 55505 1570 55545 1575
rect 58260 1605 58300 1610
rect 58260 1575 58265 1605
rect 58295 1600 58300 1605
rect 58370 1605 58410 1610
rect 58370 1600 58375 1605
rect 58295 1580 58375 1600
rect 58295 1575 58300 1580
rect 58260 1570 58300 1575
rect 58370 1575 58375 1580
rect 58405 1600 58410 1605
rect 58480 1605 58520 1610
rect 58480 1600 58485 1605
rect 58405 1580 58485 1600
rect 58405 1575 58410 1580
rect 58370 1570 58410 1575
rect 58480 1575 58485 1580
rect 58515 1600 58520 1605
rect 58590 1605 58630 1610
rect 58590 1600 58595 1605
rect 58515 1580 58595 1600
rect 58515 1575 58520 1580
rect 58480 1570 58520 1575
rect 58590 1575 58595 1580
rect 58625 1600 58630 1605
rect 58700 1605 58740 1610
rect 58700 1600 58705 1605
rect 58625 1580 58705 1600
rect 58625 1575 58630 1580
rect 58590 1570 58630 1575
rect 58700 1575 58705 1580
rect 58735 1575 58740 1605
rect 58700 1570 58740 1575
rect 54805 1555 54845 1560
rect 55010 1560 55050 1565
rect 54570 1535 54610 1540
rect 54570 1505 54575 1535
rect 54605 1530 54610 1535
rect 54760 1535 54800 1540
rect 54760 1530 54765 1535
rect 54605 1510 54765 1530
rect 54605 1505 54610 1510
rect 54570 1500 54610 1505
rect 54760 1505 54765 1510
rect 54795 1505 54800 1535
rect 55010 1530 55015 1560
rect 55045 1555 55050 1560
rect 55120 1560 55160 1565
rect 55120 1555 55125 1560
rect 55045 1535 55125 1555
rect 55045 1530 55050 1535
rect 55010 1525 55050 1530
rect 55120 1530 55125 1535
rect 55155 1555 55160 1560
rect 55230 1560 55270 1565
rect 55230 1555 55235 1560
rect 55155 1535 55235 1555
rect 55155 1530 55160 1535
rect 55120 1525 55160 1530
rect 55230 1530 55235 1535
rect 55265 1555 55270 1560
rect 55340 1560 55380 1565
rect 55340 1555 55345 1560
rect 55265 1535 55345 1555
rect 55265 1530 55270 1535
rect 55230 1525 55270 1530
rect 55340 1530 55345 1535
rect 55375 1555 55380 1560
rect 55450 1560 55490 1565
rect 55450 1555 55455 1560
rect 55375 1535 55455 1555
rect 55375 1530 55380 1535
rect 55340 1525 55380 1530
rect 55450 1530 55455 1535
rect 55485 1555 55490 1560
rect 55560 1560 55600 1565
rect 55560 1555 55565 1560
rect 55485 1535 55565 1555
rect 55485 1530 55490 1535
rect 55450 1525 55490 1530
rect 55560 1530 55565 1535
rect 55595 1555 55600 1560
rect 55760 1560 55800 1565
rect 58005 1560 58045 1565
rect 55760 1555 55765 1560
rect 55595 1535 55765 1555
rect 55595 1530 55600 1535
rect 55560 1525 55600 1530
rect 55760 1530 55765 1535
rect 55795 1530 55800 1560
rect 55760 1525 55800 1530
rect 56085 1555 56125 1560
rect 56085 1525 56090 1555
rect 56120 1550 56125 1555
rect 56195 1555 56235 1560
rect 56195 1550 56200 1555
rect 56120 1530 56200 1550
rect 56120 1525 56125 1530
rect 56085 1520 56125 1525
rect 56195 1525 56200 1530
rect 56230 1550 56235 1555
rect 56305 1555 56345 1560
rect 56305 1550 56310 1555
rect 56230 1530 56310 1550
rect 56230 1525 56235 1530
rect 56195 1520 56235 1525
rect 56305 1525 56310 1530
rect 56340 1550 56345 1555
rect 56415 1555 56455 1560
rect 56415 1550 56420 1555
rect 56340 1530 56420 1550
rect 56340 1525 56345 1530
rect 56305 1520 56345 1525
rect 56415 1525 56420 1530
rect 56450 1550 56455 1555
rect 56525 1555 56565 1560
rect 56525 1550 56530 1555
rect 56450 1530 56530 1550
rect 56450 1525 56455 1530
rect 56415 1520 56455 1525
rect 56525 1525 56530 1530
rect 56560 1550 56565 1555
rect 56635 1555 56675 1560
rect 56635 1550 56640 1555
rect 56560 1530 56640 1550
rect 56560 1525 56565 1530
rect 56525 1520 56565 1525
rect 56635 1525 56640 1530
rect 56670 1525 56675 1555
rect 56635 1520 56675 1525
rect 57125 1555 57165 1560
rect 57125 1525 57130 1555
rect 57160 1550 57165 1555
rect 57235 1555 57275 1560
rect 57235 1550 57240 1555
rect 57160 1530 57240 1550
rect 57160 1525 57165 1530
rect 57125 1520 57165 1525
rect 57235 1525 57240 1530
rect 57270 1550 57275 1555
rect 57345 1555 57385 1560
rect 57345 1550 57350 1555
rect 57270 1530 57350 1550
rect 57270 1525 57275 1530
rect 57235 1520 57275 1525
rect 57345 1525 57350 1530
rect 57380 1550 57385 1555
rect 57455 1555 57495 1560
rect 57455 1550 57460 1555
rect 57380 1530 57460 1550
rect 57380 1525 57385 1530
rect 57345 1520 57385 1525
rect 57455 1525 57460 1530
rect 57490 1550 57495 1555
rect 57565 1555 57605 1560
rect 57565 1550 57570 1555
rect 57490 1530 57570 1550
rect 57490 1525 57495 1530
rect 57455 1520 57495 1525
rect 57565 1525 57570 1530
rect 57600 1550 57605 1555
rect 57675 1555 57715 1560
rect 57675 1550 57680 1555
rect 57600 1530 57680 1550
rect 57600 1525 57605 1530
rect 57565 1520 57605 1525
rect 57675 1525 57680 1530
rect 57710 1525 57715 1555
rect 58005 1530 58010 1560
rect 58040 1555 58045 1560
rect 58205 1560 58245 1565
rect 58205 1555 58210 1560
rect 58040 1535 58210 1555
rect 58040 1530 58045 1535
rect 58005 1525 58045 1530
rect 58205 1530 58210 1535
rect 58240 1555 58245 1560
rect 58315 1560 58355 1565
rect 58315 1555 58320 1560
rect 58240 1535 58320 1555
rect 58240 1530 58245 1535
rect 58205 1525 58245 1530
rect 58315 1530 58320 1535
rect 58350 1555 58355 1560
rect 58425 1560 58465 1565
rect 58425 1555 58430 1560
rect 58350 1535 58430 1555
rect 58350 1530 58355 1535
rect 58315 1525 58355 1530
rect 58425 1530 58430 1535
rect 58460 1555 58465 1560
rect 58535 1560 58575 1565
rect 58535 1555 58540 1560
rect 58460 1535 58540 1555
rect 58460 1530 58465 1535
rect 58425 1525 58465 1530
rect 58535 1530 58540 1535
rect 58570 1555 58575 1560
rect 58645 1560 58685 1565
rect 58645 1555 58650 1560
rect 58570 1535 58650 1555
rect 58570 1530 58575 1535
rect 58535 1525 58575 1530
rect 58645 1530 58650 1535
rect 58680 1555 58685 1560
rect 58755 1560 58795 1565
rect 58755 1555 58760 1560
rect 58680 1535 58760 1555
rect 58680 1530 58685 1535
rect 58645 1525 58685 1530
rect 58755 1530 58760 1535
rect 58790 1530 58795 1560
rect 59315 1550 59350 1551
rect 59135 1545 59170 1550
rect 58755 1525 58795 1530
rect 58955 1540 58995 1545
rect 57675 1520 57715 1525
rect 54760 1500 54800 1505
rect 56140 1510 56180 1515
rect 56140 1480 56145 1510
rect 56175 1505 56180 1510
rect 56250 1510 56290 1515
rect 56250 1505 56255 1510
rect 56175 1485 56255 1505
rect 56175 1480 56180 1485
rect 56140 1475 56180 1480
rect 56250 1480 56255 1485
rect 56285 1505 56290 1510
rect 56360 1510 56400 1515
rect 56360 1505 56365 1510
rect 56285 1485 56365 1505
rect 56285 1480 56290 1485
rect 56250 1475 56290 1480
rect 56360 1480 56365 1485
rect 56395 1505 56400 1510
rect 56470 1510 56510 1515
rect 56470 1505 56475 1510
rect 56395 1485 56475 1505
rect 56395 1480 56400 1485
rect 56360 1475 56400 1480
rect 56470 1480 56475 1485
rect 56505 1505 56510 1510
rect 56580 1510 56620 1515
rect 56580 1505 56585 1510
rect 56505 1485 56585 1505
rect 56505 1480 56510 1485
rect 56470 1475 56510 1480
rect 56580 1480 56585 1485
rect 56615 1505 56620 1510
rect 57180 1510 57220 1515
rect 57180 1505 57185 1510
rect 56615 1485 57185 1505
rect 56615 1480 56620 1485
rect 56580 1475 56620 1480
rect 57180 1480 57185 1485
rect 57215 1505 57220 1510
rect 57290 1510 57330 1515
rect 57290 1505 57295 1510
rect 57215 1485 57295 1505
rect 57215 1480 57220 1485
rect 57180 1475 57220 1480
rect 57290 1480 57295 1485
rect 57325 1505 57330 1510
rect 57400 1510 57440 1515
rect 57400 1505 57405 1510
rect 57325 1485 57405 1505
rect 57325 1480 57330 1485
rect 57290 1475 57330 1480
rect 57400 1480 57405 1485
rect 57435 1505 57440 1510
rect 57510 1510 57550 1515
rect 57510 1505 57515 1510
rect 57435 1485 57515 1505
rect 57435 1480 57440 1485
rect 57400 1475 57440 1480
rect 57510 1480 57515 1485
rect 57545 1505 57550 1510
rect 57620 1510 57660 1515
rect 57620 1505 57625 1510
rect 57545 1485 57625 1505
rect 57545 1480 57550 1485
rect 57510 1475 57550 1480
rect 57620 1480 57625 1485
rect 57655 1480 57660 1510
rect 58955 1510 58960 1540
rect 58990 1535 58995 1540
rect 58990 1515 59135 1535
rect 58990 1510 58995 1515
rect 58955 1505 58995 1510
rect 59135 1505 59170 1510
rect 59195 1545 59230 1550
rect 59195 1505 59230 1510
rect 59255 1545 59350 1550
rect 59290 1510 59315 1545
rect 59255 1505 59350 1510
rect 57620 1475 57660 1480
rect 59000 1485 59040 1490
rect 54955 1465 54995 1470
rect 54955 1435 54960 1465
rect 54990 1460 54995 1465
rect 55615 1465 55655 1470
rect 55615 1460 55620 1465
rect 54990 1440 55620 1460
rect 54990 1435 54995 1440
rect 54955 1430 54995 1435
rect 55615 1435 55620 1440
rect 55650 1460 55655 1465
rect 55785 1465 55825 1470
rect 55785 1460 55790 1465
rect 55650 1440 55790 1460
rect 55650 1435 55655 1440
rect 55615 1430 55655 1435
rect 55785 1435 55790 1440
rect 55820 1435 55825 1465
rect 55785 1430 55825 1435
rect 56030 1465 56070 1470
rect 56030 1435 56035 1465
rect 56065 1460 56070 1465
rect 56730 1465 56770 1470
rect 56730 1460 56735 1465
rect 56065 1440 56735 1460
rect 56065 1435 56070 1440
rect 56030 1430 56070 1435
rect 56730 1435 56735 1440
rect 56765 1460 56770 1465
rect 57030 1465 57070 1470
rect 57030 1460 57035 1465
rect 56765 1440 57035 1460
rect 56765 1435 56770 1440
rect 56730 1430 56770 1435
rect 57030 1435 57035 1440
rect 57065 1460 57070 1465
rect 57730 1465 57770 1470
rect 57730 1460 57735 1465
rect 57065 1440 57735 1460
rect 57065 1435 57070 1440
rect 57030 1430 57070 1435
rect 57730 1435 57735 1440
rect 57765 1460 57770 1465
rect 57910 1465 57950 1470
rect 57910 1460 57915 1465
rect 57765 1440 57915 1460
rect 57765 1435 57770 1440
rect 57730 1430 57770 1435
rect 57910 1435 57915 1440
rect 57945 1460 57950 1465
rect 58150 1465 58190 1470
rect 58150 1460 58155 1465
rect 57945 1440 58155 1460
rect 57945 1435 57950 1440
rect 57910 1430 57950 1435
rect 58150 1435 58155 1440
rect 58185 1460 58190 1465
rect 58810 1465 58850 1470
rect 58810 1460 58815 1465
rect 58185 1440 58815 1460
rect 58185 1435 58190 1440
rect 58150 1430 58190 1435
rect 58810 1435 58815 1440
rect 58845 1435 58850 1465
rect 59000 1455 59005 1485
rect 59035 1480 59040 1485
rect 59190 1485 59230 1490
rect 59190 1480 59195 1485
rect 59035 1460 59195 1480
rect 59035 1455 59040 1460
rect 59000 1450 59040 1455
rect 59190 1455 59195 1460
rect 59225 1455 59230 1485
rect 59190 1450 59230 1455
rect 58810 1430 58850 1435
rect 54450 1420 54490 1425
rect 54450 1390 54455 1420
rect 54485 1415 54490 1420
rect 55940 1420 55980 1425
rect 55940 1415 55945 1420
rect 54485 1395 55945 1415
rect 54485 1390 54490 1395
rect 54450 1385 54490 1390
rect 55940 1390 55945 1395
rect 55975 1390 55980 1420
rect 55940 1385 55980 1390
rect 56825 1420 56865 1425
rect 56825 1390 56830 1420
rect 56860 1415 56865 1420
rect 56935 1420 56975 1425
rect 56935 1415 56940 1420
rect 56860 1395 56940 1415
rect 56860 1390 56865 1395
rect 56825 1385 56865 1390
rect 56935 1390 56940 1395
rect 56970 1390 56975 1420
rect 56935 1385 56975 1390
rect 57820 1420 57860 1425
rect 57820 1390 57825 1420
rect 57855 1415 57860 1420
rect 59310 1420 59350 1425
rect 59310 1415 59315 1420
rect 57855 1395 59315 1415
rect 57855 1390 57860 1395
rect 57820 1385 57860 1390
rect 59310 1390 59315 1395
rect 59345 1390 59350 1420
rect 59310 1385 59350 1390
rect 54705 1325 54745 1330
rect 54705 1295 54710 1325
rect 54740 1320 54745 1325
rect 55385 1325 55425 1330
rect 55385 1320 55390 1325
rect 54740 1300 55390 1320
rect 54740 1295 54745 1300
rect 54705 1290 54745 1295
rect 55385 1295 55390 1300
rect 55420 1320 55425 1325
rect 58430 1325 58470 1330
rect 58430 1320 58435 1325
rect 55420 1300 58435 1320
rect 55420 1295 55425 1300
rect 55385 1290 55425 1295
rect 58430 1295 58435 1300
rect 58465 1320 58470 1325
rect 59035 1325 59075 1330
rect 59035 1320 59040 1325
rect 58465 1300 59040 1320
rect 58465 1295 58470 1300
rect 58430 1290 58470 1295
rect 59035 1295 59040 1300
rect 59070 1295 59075 1325
rect 59035 1290 59075 1295
rect 56330 1265 56370 1270
rect 54295 1255 54335 1260
rect 54295 1225 54300 1255
rect 54330 1250 54335 1255
rect 54770 1255 54810 1260
rect 54770 1250 54775 1255
rect 54330 1230 54775 1250
rect 54330 1225 54335 1230
rect 54295 1220 54335 1225
rect 54770 1225 54775 1230
rect 54805 1250 54810 1255
rect 55085 1255 55125 1260
rect 55085 1250 55090 1255
rect 54805 1230 55090 1250
rect 54805 1225 54810 1230
rect 54770 1220 54810 1225
rect 55085 1225 55090 1230
rect 55120 1250 55125 1255
rect 55285 1255 55325 1260
rect 55285 1250 55290 1255
rect 55120 1230 55290 1250
rect 55120 1225 55125 1230
rect 55085 1220 55125 1225
rect 55285 1225 55290 1230
rect 55320 1250 55325 1255
rect 55485 1255 55525 1260
rect 55485 1250 55490 1255
rect 55320 1230 55490 1250
rect 55320 1225 55325 1230
rect 55285 1220 55325 1225
rect 55485 1225 55490 1230
rect 55520 1225 55525 1255
rect 56330 1235 56335 1265
rect 56365 1260 56370 1265
rect 56880 1265 56920 1270
rect 56880 1260 56885 1265
rect 56365 1240 56885 1260
rect 56365 1235 56370 1240
rect 56330 1230 56370 1235
rect 56880 1235 56885 1240
rect 56915 1235 56920 1265
rect 56880 1230 56920 1235
rect 57405 1265 57445 1270
rect 57405 1235 57410 1265
rect 57440 1260 57445 1265
rect 57865 1265 57905 1270
rect 57865 1260 57870 1265
rect 57440 1240 57870 1260
rect 57440 1235 57445 1240
rect 57405 1230 57445 1235
rect 57865 1235 57870 1240
rect 57900 1235 57905 1265
rect 57865 1230 57905 1235
rect 58280 1255 58320 1260
rect 55485 1220 55525 1225
rect 58280 1225 58285 1255
rect 58315 1250 58320 1255
rect 58480 1255 58520 1260
rect 58970 1255 59010 1260
rect 58480 1250 58485 1255
rect 58315 1230 58485 1250
rect 58315 1225 58320 1230
rect 58280 1220 58320 1225
rect 58480 1225 58485 1230
rect 58515 1250 58520 1255
rect 58680 1250 58685 1255
rect 58515 1230 58685 1250
rect 58515 1225 58520 1230
rect 58480 1220 58520 1225
rect 58680 1225 58685 1230
rect 58715 1250 58720 1255
rect 58970 1250 58975 1255
rect 58715 1230 58975 1250
rect 58715 1225 58720 1230
rect 58680 1220 58720 1225
rect 58970 1225 58975 1230
rect 59005 1250 59010 1255
rect 59465 1255 59505 1260
rect 59465 1250 59470 1255
rect 59005 1230 59470 1250
rect 59005 1225 59010 1230
rect 58970 1220 59010 1225
rect 59465 1225 59470 1230
rect 59500 1225 59505 1255
rect 59465 1220 59505 1225
rect 56440 1210 56480 1215
rect 54710 1195 54745 1200
rect 54710 1155 54745 1160
rect 54770 1195 54805 1200
rect 56440 1180 56445 1210
rect 56475 1205 56480 1210
rect 56550 1210 56590 1215
rect 56550 1205 56555 1210
rect 56475 1185 56555 1205
rect 56475 1180 56480 1185
rect 56440 1175 56480 1180
rect 56550 1180 56555 1185
rect 56585 1205 56590 1210
rect 56660 1210 56700 1215
rect 56660 1205 56665 1210
rect 56585 1185 56665 1205
rect 56585 1180 56590 1185
rect 56550 1175 56590 1180
rect 56660 1180 56665 1185
rect 56695 1205 56700 1210
rect 56770 1210 56810 1215
rect 56770 1205 56775 1210
rect 56695 1185 56775 1205
rect 56695 1180 56700 1185
rect 56660 1175 56700 1180
rect 56770 1180 56775 1185
rect 56805 1205 56810 1210
rect 56880 1210 56920 1215
rect 56880 1205 56885 1210
rect 56805 1185 56885 1205
rect 56805 1180 56810 1185
rect 56770 1175 56810 1180
rect 56880 1180 56885 1185
rect 56915 1205 56920 1210
rect 56990 1210 57030 1215
rect 56990 1205 56995 1210
rect 56915 1185 56995 1205
rect 56915 1180 56920 1185
rect 56880 1175 56920 1180
rect 56990 1180 56995 1185
rect 57025 1205 57030 1210
rect 57100 1210 57140 1215
rect 57100 1205 57105 1210
rect 57025 1185 57105 1205
rect 57025 1180 57030 1185
rect 56990 1175 57030 1180
rect 57100 1180 57105 1185
rect 57135 1205 57140 1210
rect 57210 1210 57250 1215
rect 57210 1205 57215 1210
rect 57135 1185 57215 1205
rect 57135 1180 57140 1185
rect 57100 1175 57140 1180
rect 57210 1180 57215 1185
rect 57245 1205 57250 1210
rect 57320 1210 57360 1215
rect 57320 1205 57325 1210
rect 57245 1185 57325 1205
rect 57245 1180 57250 1185
rect 57210 1175 57250 1180
rect 57320 1180 57325 1185
rect 57355 1205 57360 1210
rect 57430 1210 57470 1215
rect 57430 1205 57435 1210
rect 57355 1185 57435 1205
rect 57355 1180 57360 1185
rect 57320 1175 57360 1180
rect 57430 1180 57435 1185
rect 57465 1180 57470 1210
rect 57430 1175 57470 1180
rect 58975 1200 59010 1205
rect 58975 1160 59010 1165
rect 59035 1200 59070 1205
rect 59035 1160 59070 1165
rect 54770 1155 54805 1160
rect 55785 890 55825 895
rect 55785 860 55790 890
rect 55820 885 55825 890
rect 56220 890 56260 895
rect 56220 885 56225 890
rect 55820 865 56225 885
rect 55820 860 55825 865
rect 55785 855 55825 860
rect 56220 860 56225 865
rect 56255 885 56260 890
rect 56275 890 56315 895
rect 56275 885 56280 890
rect 56255 865 56280 885
rect 56255 860 56260 865
rect 56220 855 56260 860
rect 56275 860 56280 865
rect 56310 885 56315 890
rect 56385 890 56425 895
rect 56385 885 56390 890
rect 56310 865 56390 885
rect 56310 860 56315 865
rect 56275 855 56315 860
rect 56385 860 56390 865
rect 56420 885 56425 890
rect 56495 890 56535 895
rect 56495 885 56500 890
rect 56420 865 56500 885
rect 56420 860 56425 865
rect 56385 855 56425 860
rect 56495 860 56500 865
rect 56530 885 56535 890
rect 56605 890 56645 895
rect 56605 885 56610 890
rect 56530 865 56610 885
rect 56530 860 56535 865
rect 56495 855 56535 860
rect 56605 860 56610 865
rect 56640 885 56645 890
rect 56715 890 56755 895
rect 56715 885 56720 890
rect 56640 865 56720 885
rect 56640 860 56645 865
rect 56605 855 56645 860
rect 56715 860 56720 865
rect 56750 885 56755 890
rect 56825 890 56865 895
rect 56825 885 56830 890
rect 56750 865 56830 885
rect 56750 860 56755 865
rect 56715 855 56755 860
rect 56825 860 56830 865
rect 56860 885 56865 890
rect 56935 890 56975 895
rect 56935 885 56940 890
rect 56860 865 56940 885
rect 56860 860 56865 865
rect 56825 855 56865 860
rect 56935 860 56940 865
rect 56970 885 56975 890
rect 57045 890 57085 895
rect 57045 885 57050 890
rect 56970 865 57050 885
rect 56970 860 56975 865
rect 56935 855 56975 860
rect 57045 860 57050 865
rect 57080 885 57085 890
rect 57155 890 57195 895
rect 57155 885 57160 890
rect 57080 865 57160 885
rect 57080 860 57085 865
rect 57045 855 57085 860
rect 57155 860 57160 865
rect 57190 885 57195 890
rect 57265 890 57305 895
rect 57265 885 57270 890
rect 57190 865 57270 885
rect 57190 860 57195 865
rect 57155 855 57195 860
rect 57265 860 57270 865
rect 57300 885 57305 890
rect 57375 890 57415 895
rect 57375 885 57380 890
rect 57300 865 57380 885
rect 57300 860 57305 865
rect 57265 855 57305 860
rect 57375 860 57380 865
rect 57410 885 57415 890
rect 57485 890 57525 895
rect 57485 885 57490 890
rect 57410 865 57490 885
rect 57410 860 57415 865
rect 57375 855 57415 860
rect 57485 860 57490 865
rect 57520 885 57525 890
rect 57520 880 57950 885
rect 57520 865 57915 880
rect 57520 860 57525 865
rect 57485 855 57525 860
rect 57910 850 57915 865
rect 57945 850 57950 880
rect 56440 845 56480 850
rect 56440 815 56445 845
rect 56475 840 56480 845
rect 56550 845 56590 850
rect 56550 840 56555 845
rect 56475 820 56555 840
rect 56475 815 56480 820
rect 56440 810 56480 815
rect 56550 815 56555 820
rect 56585 840 56590 845
rect 56660 845 56700 850
rect 56660 840 56665 845
rect 56585 820 56665 840
rect 56585 815 56590 820
rect 56550 810 56590 815
rect 56660 815 56665 820
rect 56695 840 56700 845
rect 56770 845 56810 850
rect 56770 840 56775 845
rect 56695 820 56775 840
rect 56695 815 56700 820
rect 56660 810 56700 815
rect 56770 815 56775 820
rect 56805 840 56810 845
rect 56880 845 56920 850
rect 56880 840 56885 845
rect 56805 820 56885 840
rect 56805 815 56810 820
rect 56770 810 56810 815
rect 56880 815 56885 820
rect 56915 840 56920 845
rect 56990 845 57030 850
rect 56990 840 56995 845
rect 56915 820 56995 840
rect 56915 815 56920 820
rect 56880 810 56920 815
rect 56990 815 56995 820
rect 57025 840 57030 845
rect 57100 845 57140 850
rect 57100 840 57105 845
rect 57025 820 57105 840
rect 57025 815 57030 820
rect 56990 810 57030 815
rect 57100 815 57105 820
rect 57135 840 57140 845
rect 57210 845 57250 850
rect 57210 840 57215 845
rect 57135 820 57215 840
rect 57135 815 57140 820
rect 57100 810 57140 815
rect 57210 815 57215 820
rect 57245 840 57250 845
rect 57320 845 57360 850
rect 57320 840 57325 845
rect 57245 820 57325 840
rect 57245 815 57250 820
rect 57210 810 57250 815
rect 57320 815 57325 820
rect 57355 840 57360 845
rect 57430 845 57470 850
rect 57910 845 57950 850
rect 57430 840 57435 845
rect 57355 820 57435 840
rect 57355 815 57360 820
rect 57320 810 57360 815
rect 57430 815 57435 820
rect 57465 815 57470 845
rect 57430 810 57470 815
rect 56540 790 56580 795
rect 56540 760 56545 790
rect 56575 785 56580 790
rect 56650 790 56690 795
rect 56650 785 56655 790
rect 56575 765 56655 785
rect 56575 760 56580 765
rect 56540 755 56580 760
rect 56650 760 56655 765
rect 56685 785 56690 790
rect 56870 790 56910 795
rect 56870 785 56875 790
rect 56685 765 56875 785
rect 56685 760 56690 765
rect 56650 755 56690 760
rect 56870 760 56875 765
rect 56905 760 56910 790
rect 56870 755 56910 760
rect 55830 745 55870 750
rect 55830 715 55835 745
rect 55865 740 55870 745
rect 56485 745 56525 750
rect 56485 740 56490 745
rect 55865 720 56490 740
rect 55865 715 55870 720
rect 55830 710 55870 715
rect 56485 715 56490 720
rect 56520 740 56525 745
rect 56595 745 56635 750
rect 56595 740 56600 745
rect 56520 720 56600 740
rect 56520 715 56525 720
rect 56485 710 56525 715
rect 56595 715 56600 720
rect 56630 740 56635 745
rect 56705 745 56745 750
rect 56705 740 56710 745
rect 56630 720 56710 740
rect 56630 715 56635 720
rect 56595 710 56635 715
rect 56705 715 56710 720
rect 56740 740 56745 745
rect 57040 745 57080 750
rect 57040 740 57045 745
rect 56740 720 57045 740
rect 56740 715 56745 720
rect 56705 710 56745 715
rect 57040 715 57045 720
rect 57075 715 57080 745
rect 57040 710 57080 715
rect 56540 540 56580 545
rect 55085 515 55125 520
rect 55085 485 55090 515
rect 55120 510 55125 515
rect 55285 515 55325 520
rect 55285 510 55290 515
rect 55120 490 55290 510
rect 55120 485 55125 490
rect 55085 480 55125 485
rect 55285 485 55290 490
rect 55320 510 55325 515
rect 55485 515 55525 520
rect 55485 510 55490 515
rect 55320 490 55490 510
rect 55320 485 55325 490
rect 55285 480 55325 485
rect 55485 485 55490 490
rect 55520 485 55525 515
rect 56540 510 56545 540
rect 56575 535 56580 540
rect 56650 540 56690 545
rect 56650 535 56655 540
rect 56575 515 56655 535
rect 56575 510 56580 515
rect 56540 505 56580 510
rect 56650 510 56655 515
rect 56685 535 56690 540
rect 56870 540 56910 545
rect 56870 535 56875 540
rect 56685 515 56875 535
rect 56685 510 56690 515
rect 56650 505 56690 510
rect 56870 510 56875 515
rect 56905 510 56910 540
rect 56870 505 56910 510
rect 58280 515 58320 520
rect 55485 480 55525 485
rect 56485 495 56525 500
rect 56485 465 56490 495
rect 56520 490 56525 495
rect 56595 495 56635 500
rect 56595 490 56600 495
rect 56520 470 56600 490
rect 56520 465 56525 470
rect 56485 460 56525 465
rect 56595 465 56600 470
rect 56630 490 56635 495
rect 56705 495 56745 500
rect 56705 490 56710 495
rect 56630 470 56710 490
rect 56630 465 56635 470
rect 56595 460 56635 465
rect 56705 465 56710 470
rect 56740 465 56745 495
rect 58280 485 58285 515
rect 58315 510 58320 515
rect 58480 515 58520 520
rect 58480 510 58485 515
rect 58315 490 58485 510
rect 58315 485 58320 490
rect 58280 480 58320 485
rect 58480 485 58485 490
rect 58515 510 58520 515
rect 58680 515 58720 520
rect 58680 510 58685 515
rect 58515 490 58685 510
rect 58515 485 58520 490
rect 58480 480 58520 485
rect 58680 485 58685 490
rect 58715 485 58720 515
rect 58680 480 58720 485
rect 56705 460 56745 465
rect 54245 395 54285 400
rect 54245 365 54250 395
rect 54280 390 54285 395
rect 54985 395 55025 400
rect 54985 390 54990 395
rect 54280 370 54990 390
rect 54280 365 54285 370
rect 54245 360 54285 365
rect 54985 365 54990 370
rect 55020 390 55025 395
rect 55185 395 55225 400
rect 55185 390 55190 395
rect 55020 370 55190 390
rect 55020 365 55025 370
rect 54985 360 55025 365
rect 55185 365 55190 370
rect 55220 390 55225 395
rect 55385 395 55425 400
rect 55385 390 55390 395
rect 55220 370 55390 390
rect 55220 365 55225 370
rect 55185 360 55225 365
rect 55385 365 55390 370
rect 55420 390 55425 395
rect 55585 395 55625 400
rect 55585 390 55590 395
rect 55420 370 55590 390
rect 55420 365 55425 370
rect 55385 360 55425 365
rect 55585 365 55590 370
rect 55620 390 55625 395
rect 55785 395 55825 400
rect 55785 390 55790 395
rect 55620 370 55790 390
rect 55620 365 55625 370
rect 55585 360 55625 365
rect 55785 365 55790 370
rect 55820 390 55825 395
rect 56430 395 56470 400
rect 56430 390 56435 395
rect 55820 370 56435 390
rect 55820 365 55825 370
rect 55785 360 55825 365
rect 56430 365 56435 370
rect 56465 390 56470 395
rect 56760 395 56800 400
rect 56760 390 56765 395
rect 56465 370 56765 390
rect 56465 365 56470 370
rect 56430 360 56470 365
rect 56760 365 56765 370
rect 56795 390 56800 395
rect 56880 395 56920 400
rect 56880 390 56885 395
rect 56795 370 56885 390
rect 56795 365 56800 370
rect 56760 360 56800 365
rect 56880 365 56885 370
rect 56915 390 56920 395
rect 57910 395 57950 400
rect 57910 390 57915 395
rect 56915 370 57915 390
rect 56915 365 56920 370
rect 56880 360 56920 365
rect 57910 365 57915 370
rect 57945 390 57950 395
rect 58180 395 58220 400
rect 58180 390 58185 395
rect 57945 370 58185 390
rect 57945 365 57950 370
rect 57910 360 57950 365
rect 58180 365 58185 370
rect 58215 390 58220 395
rect 58380 395 58420 400
rect 58380 390 58385 395
rect 58215 370 58385 390
rect 58215 365 58220 370
rect 58180 360 58220 365
rect 58380 365 58385 370
rect 58415 390 58420 395
rect 58580 395 58620 400
rect 58580 390 58585 395
rect 58415 370 58585 390
rect 58415 365 58420 370
rect 58380 360 58420 365
rect 58580 365 58585 370
rect 58615 390 58620 395
rect 58780 395 58820 400
rect 58780 390 58785 395
rect 58615 370 58785 390
rect 58615 365 58620 370
rect 58580 360 58620 365
rect 58780 365 58785 370
rect 58815 390 58820 395
rect 59515 395 59555 400
rect 59515 390 59520 395
rect 58815 370 59520 390
rect 58815 365 58820 370
rect 58780 360 58820 365
rect 59515 365 59520 370
rect 59550 365 59555 395
rect 59515 360 59555 365
<< via2 >>
rect 54610 3370 54640 3400
rect 59160 3370 59190 3400
rect 54300 1880 54330 1910
rect 59470 1880 59500 1910
<< metal3 >>
rect 52410 5770 52640 5855
rect 52760 5770 52990 5855
rect 53110 5770 53340 5855
rect 52410 5720 53340 5770
rect 52410 5625 52640 5720
rect 52760 5625 52990 5720
rect 53110 5625 53340 5720
rect 53460 5625 53690 5855
rect 53810 5625 54040 5855
rect 54160 5625 54390 5855
rect 54510 5625 54740 5855
rect 54860 5625 55090 5855
rect 55210 5625 55440 5855
rect 55560 5625 55790 5855
rect 55910 5625 56140 5855
rect 56260 5625 56490 5855
rect 56610 5625 56840 5855
rect 56960 5625 57190 5855
rect 57310 5625 57540 5855
rect 57660 5625 57890 5855
rect 58010 5625 58240 5855
rect 58360 5625 58590 5855
rect 58710 5625 58940 5855
rect 59060 5625 59290 5855
rect 59410 5625 59640 5855
rect 59760 5625 59990 5855
rect 60110 5625 60340 5855
rect 60460 5770 60690 5855
rect 60810 5770 61040 5855
rect 61160 5770 61390 5855
rect 60460 5720 61390 5770
rect 60460 5625 60690 5720
rect 60810 5625 61040 5720
rect 61160 5625 61390 5720
rect 53200 5505 53250 5625
rect 53550 5505 53600 5625
rect 53900 5505 53950 5625
rect 54250 5505 54300 5625
rect 54600 5505 54650 5625
rect 54950 5505 55000 5625
rect 55300 5505 55350 5625
rect 55650 5505 55700 5625
rect 56000 5505 56050 5625
rect 56350 5505 56400 5625
rect 56700 5505 56750 5625
rect 57050 5505 57100 5625
rect 57400 5505 57450 5625
rect 57750 5505 57800 5625
rect 58100 5505 58150 5625
rect 58450 5505 58500 5625
rect 58800 5505 58850 5625
rect 59150 5505 59200 5625
rect 59500 5505 59550 5625
rect 59850 5505 59900 5625
rect 60200 5505 60250 5625
rect 60550 5505 60600 5625
rect 52410 5420 52640 5505
rect 52760 5420 52990 5505
rect 53110 5420 53340 5505
rect 53460 5420 53690 5505
rect 53810 5420 54040 5505
rect 54160 5420 54390 5505
rect 54510 5420 54740 5505
rect 54860 5420 55090 5505
rect 55210 5420 55440 5505
rect 55560 5420 55790 5505
rect 55910 5420 56140 5505
rect 56260 5420 56490 5505
rect 56610 5420 56840 5505
rect 52410 5370 56840 5420
rect 52410 5275 52640 5370
rect 52760 5275 52990 5370
rect 53110 5275 53340 5370
rect 53460 5275 53690 5370
rect 53810 5275 54040 5370
rect 54160 5275 54390 5370
rect 54510 5275 54740 5370
rect 54860 5275 55090 5370
rect 55210 5275 55440 5370
rect 55560 5275 55790 5370
rect 55910 5275 56140 5370
rect 56260 5275 56490 5370
rect 56610 5275 56840 5370
rect 56960 5420 57190 5505
rect 57310 5420 57540 5505
rect 57660 5420 57890 5505
rect 58010 5420 58240 5505
rect 58360 5420 58590 5505
rect 58710 5420 58940 5505
rect 59060 5420 59290 5505
rect 59410 5420 59640 5505
rect 59760 5420 59990 5505
rect 60110 5420 60340 5505
rect 60460 5420 60690 5505
rect 60810 5420 61040 5505
rect 61160 5420 61390 5505
rect 56960 5370 61390 5420
rect 56960 5275 57190 5370
rect 57310 5275 57540 5370
rect 57660 5275 57890 5370
rect 58010 5275 58240 5370
rect 58360 5275 58590 5370
rect 58710 5275 58940 5370
rect 59060 5275 59290 5370
rect 59410 5275 59640 5370
rect 59760 5275 59990 5370
rect 60110 5275 60340 5370
rect 60460 5275 60690 5370
rect 60810 5275 61040 5370
rect 61160 5275 61390 5370
rect 53200 5155 53250 5275
rect 54250 5155 54300 5275
rect 54600 5155 54650 5275
rect 54950 5155 55000 5275
rect 55300 5155 55350 5275
rect 55650 5155 55700 5275
rect 56000 5155 56050 5275
rect 56350 5155 56400 5275
rect 56700 5155 56750 5275
rect 57050 5155 57100 5275
rect 57400 5155 57450 5275
rect 57750 5155 57800 5275
rect 58100 5155 58150 5275
rect 58450 5155 58500 5275
rect 58800 5155 58850 5275
rect 59150 5155 59200 5275
rect 59500 5155 59550 5275
rect 60550 5155 60600 5275
rect 52410 5070 52640 5155
rect 52760 5070 52990 5155
rect 53110 5070 53340 5155
rect 53460 5070 53690 5155
rect 53810 5070 54040 5155
rect 52410 5020 54040 5070
rect 52410 4925 52640 5020
rect 52760 4925 52990 5020
rect 53110 4925 53340 5020
rect 53460 4925 53690 5020
rect 53810 4925 54040 5020
rect 54160 4925 54390 5155
rect 54510 4925 54740 5155
rect 54860 4925 55090 5155
rect 55210 4925 55440 5155
rect 55560 4925 55790 5155
rect 55910 4925 56140 5155
rect 56260 4925 56490 5155
rect 56610 4925 56840 5155
rect 56960 4925 57190 5155
rect 57310 4925 57540 5155
rect 57660 4925 57890 5155
rect 58010 4925 58240 5155
rect 58360 4925 58590 5155
rect 58710 4925 58940 5155
rect 59060 4925 59290 5155
rect 59410 4925 59640 5155
rect 59760 5070 59990 5155
rect 60110 5070 60340 5155
rect 60460 5070 60690 5155
rect 60810 5070 61040 5155
rect 61160 5070 61390 5155
rect 59760 5020 61390 5070
rect 59760 4925 59990 5020
rect 60110 4925 60340 5020
rect 60460 4925 60690 5020
rect 60810 4925 61040 5020
rect 61160 4925 61390 5020
rect 53200 4805 53250 4925
rect 54250 4805 54300 4925
rect 54600 4805 54650 4925
rect 54950 4805 55000 4925
rect 55300 4805 55350 4925
rect 58450 4805 58500 4925
rect 58800 4805 58850 4925
rect 59150 4805 59200 4925
rect 59500 4805 59550 4925
rect 60550 4805 60600 4925
rect 52410 4720 52640 4805
rect 52760 4720 52990 4805
rect 53110 4720 53340 4805
rect 53460 4720 53690 4805
rect 53810 4720 54040 4805
rect 52410 4670 54040 4720
rect 52410 4575 52640 4670
rect 52760 4575 52990 4670
rect 53110 4575 53340 4670
rect 53460 4575 53690 4670
rect 53810 4575 54040 4670
rect 54160 4575 54390 4805
rect 54510 4575 54740 4805
rect 54860 4575 55090 4805
rect 55210 4575 55440 4805
rect 58360 4575 58590 4805
rect 58710 4575 58940 4805
rect 59060 4575 59290 4805
rect 59410 4575 59640 4805
rect 59760 4720 59990 4805
rect 60110 4720 60340 4805
rect 60460 4720 60690 4805
rect 60810 4720 61040 4805
rect 61160 4720 61390 4805
rect 59760 4670 61390 4720
rect 59760 4575 59990 4670
rect 60110 4575 60340 4670
rect 60460 4575 60690 4670
rect 60810 4575 61040 4670
rect 61160 4575 61390 4670
rect 53200 4455 53250 4575
rect 54250 4455 54300 4575
rect 54600 4455 54650 4575
rect 54950 4455 55000 4575
rect 55300 4455 55350 4575
rect 58450 4455 58500 4575
rect 58800 4455 58850 4575
rect 59150 4455 59200 4575
rect 59500 4455 59550 4575
rect 60550 4455 60600 4575
rect 52410 4370 52640 4455
rect 52760 4370 52990 4455
rect 53110 4370 53340 4455
rect 53460 4370 53690 4455
rect 53810 4370 54040 4455
rect 52410 4320 54040 4370
rect 52410 4225 52640 4320
rect 52760 4225 52990 4320
rect 53110 4225 53340 4320
rect 53460 4225 53690 4320
rect 53810 4225 54040 4320
rect 54160 4225 54390 4455
rect 54510 4225 54740 4455
rect 54860 4225 55090 4455
rect 55210 4225 55440 4455
rect 58360 4225 58590 4455
rect 58710 4225 58940 4455
rect 59060 4225 59290 4455
rect 59410 4225 59640 4455
rect 59760 4370 59990 4455
rect 60110 4370 60340 4455
rect 60460 4370 60690 4455
rect 60810 4370 61040 4455
rect 61160 4370 61390 4455
rect 59760 4320 61390 4370
rect 59760 4225 59990 4320
rect 60110 4225 60340 4320
rect 60460 4225 60690 4320
rect 60810 4225 61040 4320
rect 61160 4225 61390 4320
rect 53200 4105 53250 4225
rect 52410 4020 52640 4105
rect 52760 4020 52990 4105
rect 53110 4020 53340 4105
rect 53460 4020 53690 4105
rect 53810 4020 54040 4105
rect 52410 3970 54040 4020
rect 52410 3875 52640 3970
rect 52760 3875 52990 3970
rect 53110 3875 53340 3970
rect 53460 3875 53690 3970
rect 53810 3875 54040 3970
rect 53200 3755 53250 3875
rect 52410 3670 52640 3755
rect 52760 3670 52990 3755
rect 53110 3670 53340 3755
rect 53460 3670 53690 3755
rect 53810 3670 54040 3755
rect 52410 3620 54040 3670
rect 52410 3525 52640 3620
rect 52760 3525 52990 3620
rect 53110 3525 53340 3620
rect 53460 3525 53690 3620
rect 53810 3525 54040 3620
rect 53200 3405 53250 3525
rect 52410 3320 52640 3405
rect 52760 3320 52990 3405
rect 53110 3320 53340 3405
rect 53460 3320 53690 3405
rect 53810 3320 54040 3405
rect 54605 3400 54645 4225
rect 54605 3370 54610 3400
rect 54640 3370 54645 3400
rect 54605 3365 54645 3370
rect 59155 3400 59195 4225
rect 60550 4105 60600 4225
rect 59760 4020 59990 4105
rect 60110 4020 60340 4105
rect 60460 4020 60690 4105
rect 60810 4020 61040 4105
rect 61160 4020 61390 4105
rect 59760 3970 61390 4020
rect 59760 3875 59990 3970
rect 60110 3875 60340 3970
rect 60460 3875 60690 3970
rect 60810 3875 61040 3970
rect 61160 3875 61390 3970
rect 60550 3755 60600 3875
rect 59760 3670 59990 3755
rect 60110 3670 60340 3755
rect 60460 3670 60690 3755
rect 60810 3670 61040 3755
rect 61160 3670 61390 3755
rect 59760 3620 61390 3670
rect 59760 3525 59990 3620
rect 60110 3525 60340 3620
rect 60460 3525 60690 3620
rect 60810 3525 61040 3620
rect 61160 3525 61390 3620
rect 60550 3405 60600 3525
rect 59155 3370 59160 3400
rect 59190 3370 59195 3400
rect 59155 3365 59195 3370
rect 52410 3270 54040 3320
rect 52410 3175 52640 3270
rect 52760 3175 52990 3270
rect 53110 3175 53340 3270
rect 53460 3175 53690 3270
rect 53810 3175 54040 3270
rect 59760 3320 59990 3405
rect 60110 3320 60340 3405
rect 60460 3320 60690 3405
rect 60810 3320 61040 3405
rect 61160 3320 61390 3405
rect 59760 3270 61390 3320
rect 59760 3175 59990 3270
rect 60110 3175 60340 3270
rect 60460 3175 60690 3270
rect 60810 3175 61040 3270
rect 61160 3175 61390 3270
rect 53200 3055 53250 3175
rect 60550 3055 60600 3175
rect 52410 2970 52640 3055
rect 52760 2970 52990 3055
rect 53110 2970 53340 3055
rect 53460 2970 53690 3055
rect 53810 2970 54040 3055
rect 52410 2920 54040 2970
rect 52410 2825 52640 2920
rect 52760 2825 52990 2920
rect 53110 2825 53340 2920
rect 53460 2825 53690 2920
rect 53810 2825 54040 2920
rect 59760 2970 59990 3055
rect 60110 2970 60340 3055
rect 60460 2970 60690 3055
rect 60810 2970 61040 3055
rect 61160 2970 61390 3055
rect 59760 2920 61390 2970
rect 59760 2825 59990 2920
rect 60110 2825 60340 2920
rect 60460 2825 60690 2920
rect 60810 2825 61040 2920
rect 61160 2825 61390 2920
rect 53200 2705 53250 2825
rect 60550 2705 60600 2825
rect 52410 2620 52640 2705
rect 52760 2620 52990 2705
rect 53110 2620 53340 2705
rect 53460 2620 53690 2705
rect 53810 2620 54040 2705
rect 52410 2570 54040 2620
rect 52410 2475 52640 2570
rect 52760 2475 52990 2570
rect 53110 2475 53340 2570
rect 53460 2475 53690 2570
rect 53810 2475 54040 2570
rect 59760 2620 59990 2705
rect 60110 2620 60340 2705
rect 60460 2620 60690 2705
rect 60810 2620 61040 2705
rect 61160 2620 61390 2705
rect 59760 2570 61390 2620
rect 59760 2475 59990 2570
rect 60110 2475 60340 2570
rect 60460 2475 60690 2570
rect 60810 2475 61040 2570
rect 61160 2475 61390 2570
rect 53200 2355 53250 2475
rect 60550 2355 60600 2475
rect 52410 2270 52640 2355
rect 52760 2270 52990 2355
rect 53110 2270 53340 2355
rect 53460 2270 53690 2355
rect 53810 2270 54040 2355
rect 52410 2220 54040 2270
rect 52410 2125 52640 2220
rect 52760 2125 52990 2220
rect 53110 2125 53340 2220
rect 53460 2125 53690 2220
rect 53810 2125 54040 2220
rect 59760 2270 59990 2355
rect 60110 2270 60340 2355
rect 60460 2270 60690 2355
rect 60810 2270 61040 2355
rect 61160 2270 61390 2355
rect 59760 2220 61390 2270
rect 59760 2125 59990 2220
rect 60110 2125 60340 2220
rect 60460 2125 60690 2220
rect 60810 2125 61040 2220
rect 61160 2125 61390 2220
rect 53200 2005 53250 2125
rect 60550 2005 60600 2125
rect 52410 1920 52640 2005
rect 52760 1920 52990 2005
rect 53110 1920 53340 2005
rect 53460 1920 53690 2005
rect 53810 1920 54040 2005
rect 59760 1920 59990 2005
rect 60110 1920 60340 2005
rect 60460 1920 60690 2005
rect 60810 1920 61040 2005
rect 61160 1920 61390 2005
rect 52410 1870 54040 1920
rect 54290 1915 54340 1920
rect 54290 1875 54295 1915
rect 54335 1875 54340 1915
rect 54290 1870 54340 1875
rect 59460 1915 59510 1920
rect 59460 1875 59465 1915
rect 59505 1875 59510 1915
rect 59460 1870 59510 1875
rect 59760 1870 61390 1920
rect 52410 1775 52640 1870
rect 52760 1775 52990 1870
rect 53110 1775 53340 1870
rect 53460 1775 53690 1870
rect 53810 1775 54040 1870
rect 59760 1775 59990 1870
rect 60110 1775 60340 1870
rect 60460 1775 60690 1870
rect 60810 1775 61040 1870
rect 61160 1775 61390 1870
rect 53200 1655 53250 1775
rect 60550 1655 60600 1775
rect 52410 1570 52640 1655
rect 52760 1570 52990 1655
rect 53110 1570 53340 1655
rect 53460 1570 53690 1655
rect 53810 1570 54040 1655
rect 52410 1520 54040 1570
rect 52410 1425 52640 1520
rect 52760 1425 52990 1520
rect 53110 1425 53340 1520
rect 53460 1425 53690 1520
rect 53810 1425 54040 1520
rect 59760 1570 59990 1655
rect 60110 1570 60340 1655
rect 60460 1570 60690 1655
rect 60810 1570 61040 1655
rect 61160 1570 61390 1655
rect 59760 1520 61390 1570
rect 59760 1425 59990 1520
rect 60110 1425 60340 1520
rect 60460 1425 60690 1520
rect 60810 1425 61040 1520
rect 61160 1425 61390 1520
rect 53200 1305 53250 1425
rect 60550 1305 60600 1425
rect 52410 1220 52640 1305
rect 52760 1220 52990 1305
rect 53110 1220 53340 1305
rect 53460 1220 53690 1305
rect 53810 1220 54040 1305
rect 52410 1170 54040 1220
rect 52410 1075 52640 1170
rect 52760 1075 52990 1170
rect 53110 1075 53340 1170
rect 53460 1075 53690 1170
rect 53810 1075 54040 1170
rect 59760 1220 59990 1305
rect 60110 1220 60340 1305
rect 60460 1220 60690 1305
rect 60810 1220 61040 1305
rect 61160 1220 61390 1305
rect 59760 1170 61390 1220
rect 59760 1075 59990 1170
rect 60110 1075 60340 1170
rect 60460 1075 60690 1170
rect 60810 1075 61040 1170
rect 61160 1075 61390 1170
rect 53200 955 53250 1075
rect 60550 955 60600 1075
rect 52410 870 52640 955
rect 52760 870 52990 955
rect 53110 870 53340 955
rect 53460 870 53690 955
rect 53810 870 54040 955
rect 52410 820 54040 870
rect 52410 725 52640 820
rect 52760 725 52990 820
rect 53110 725 53340 820
rect 53460 725 53690 820
rect 53810 725 54040 820
rect 59760 870 59990 955
rect 60110 870 60340 955
rect 60460 870 60690 955
rect 60810 870 61040 955
rect 61160 870 61390 955
rect 59760 820 61390 870
rect 59760 725 59990 820
rect 60110 725 60340 820
rect 60460 725 60690 820
rect 60810 725 61040 820
rect 61160 725 61390 820
rect 53200 605 53250 725
rect 60550 605 60600 725
rect 52410 520 52640 605
rect 52760 520 52990 605
rect 53110 520 53340 605
rect 53460 520 53690 605
rect 53810 520 54040 605
rect 52410 470 54040 520
rect 52410 375 52640 470
rect 52760 375 52990 470
rect 53110 375 53340 470
rect 53460 375 53690 470
rect 53810 375 54040 470
rect 59760 520 59990 605
rect 60110 520 60340 605
rect 60460 520 60690 605
rect 60810 520 61040 605
rect 61160 520 61390 605
rect 59760 470 61390 520
rect 59760 375 59990 470
rect 60110 375 60340 470
rect 60460 375 60690 470
rect 60810 375 61040 470
rect 61160 375 61390 470
rect 53200 255 53250 375
rect 60550 255 60600 375
rect 52410 170 52640 255
rect 52760 170 52990 255
rect 53110 170 53340 255
rect 53460 170 53690 255
rect 53810 170 54040 255
rect 54160 170 54390 255
rect 54510 170 54740 255
rect 54860 170 55090 255
rect 55210 170 55440 255
rect 55560 170 55790 255
rect 55910 170 56140 255
rect 56260 170 56490 255
rect 56610 170 56840 255
rect 52410 120 56840 170
rect 52410 25 52640 120
rect 52760 25 52990 120
rect 53110 25 53340 120
rect 53460 25 53690 120
rect 53810 25 54040 120
rect 54160 25 54390 120
rect 54510 25 54740 120
rect 54860 25 55090 120
rect 55210 25 55440 120
rect 55560 25 55790 120
rect 55910 25 56140 120
rect 56260 25 56490 120
rect 56610 25 56840 120
rect 56960 170 57190 255
rect 57310 170 57540 255
rect 57660 170 57890 255
rect 58010 170 58240 255
rect 58360 170 58590 255
rect 58710 170 58940 255
rect 59060 170 59290 255
rect 59410 170 59640 255
rect 59760 170 59990 255
rect 60110 170 60340 255
rect 60460 170 60690 255
rect 60810 170 61040 255
rect 61160 170 61390 255
rect 56960 120 61390 170
rect 56960 25 57190 120
rect 57310 25 57540 120
rect 57660 25 57890 120
rect 58010 25 58240 120
rect 58360 25 58590 120
rect 58710 25 58940 120
rect 59060 25 59290 120
rect 59410 25 59640 120
rect 59760 25 59990 120
rect 60110 25 60340 120
rect 60460 25 60690 120
rect 60810 25 61040 120
rect 61160 25 61390 120
rect 53200 -95 53250 25
rect 53550 -95 53600 25
rect 53900 -95 53950 25
rect 54250 -95 54300 25
rect 54600 -95 54650 25
rect 54950 -95 55000 25
rect 55300 -95 55350 25
rect 55650 -95 55700 25
rect 56000 -95 56050 25
rect 56350 -95 56400 25
rect 56700 -95 56750 25
rect 57050 -95 57100 25
rect 57400 -95 57450 25
rect 57750 -95 57800 25
rect 58100 -95 58150 25
rect 58450 -95 58500 25
rect 58800 -95 58850 25
rect 59150 -95 59200 25
rect 59500 -95 59550 25
rect 59850 -95 59900 25
rect 60200 -95 60250 25
rect 60550 -95 60600 25
rect 52410 -180 52640 -95
rect 52760 -180 52990 -95
rect 53110 -180 53340 -95
rect 52410 -230 53340 -180
rect 52410 -325 52640 -230
rect 52760 -325 52990 -230
rect 53110 -325 53340 -230
rect 53460 -325 53690 -95
rect 53810 -325 54040 -95
rect 54160 -325 54390 -95
rect 54510 -325 54740 -95
rect 54860 -325 55090 -95
rect 55210 -325 55440 -95
rect 55560 -325 55790 -95
rect 55910 -325 56140 -95
rect 56260 -325 56490 -95
rect 56610 -325 56840 -95
rect 56960 -325 57190 -95
rect 57310 -325 57540 -95
rect 57660 -325 57890 -95
rect 58010 -325 58240 -95
rect 58360 -325 58590 -95
rect 58710 -325 58940 -95
rect 59060 -325 59290 -95
rect 59410 -325 59640 -95
rect 59760 -325 59990 -95
rect 60110 -325 60340 -95
rect 60460 -180 60690 -95
rect 60810 -180 61040 -95
rect 61160 -180 61390 -95
rect 60460 -230 61390 -180
rect 60460 -325 60690 -230
rect 60810 -325 61040 -230
rect 61160 -325 61390 -230
<< via3 >>
rect 54295 1910 54335 1915
rect 54295 1880 54300 1910
rect 54300 1880 54330 1910
rect 54330 1880 54335 1910
rect 54295 1875 54335 1880
rect 59465 1910 59505 1915
rect 59465 1880 59470 1910
rect 59470 1880 59500 1910
rect 59500 1880 59505 1910
rect 59465 1875 59505 1880
<< mimcap >>
rect 52425 5765 52625 5840
rect 52425 5725 52505 5765
rect 52545 5725 52625 5765
rect 52425 5640 52625 5725
rect 52775 5765 52975 5840
rect 52775 5725 52855 5765
rect 52895 5725 52975 5765
rect 52775 5640 52975 5725
rect 53125 5765 53325 5840
rect 53125 5725 53205 5765
rect 53245 5725 53325 5765
rect 53125 5640 53325 5725
rect 53475 5765 53675 5840
rect 53475 5725 53555 5765
rect 53595 5725 53675 5765
rect 53475 5640 53675 5725
rect 53825 5765 54025 5840
rect 53825 5725 53905 5765
rect 53945 5725 54025 5765
rect 53825 5640 54025 5725
rect 54175 5765 54375 5840
rect 54175 5725 54255 5765
rect 54295 5725 54375 5765
rect 54175 5640 54375 5725
rect 54525 5765 54725 5840
rect 54525 5725 54605 5765
rect 54645 5725 54725 5765
rect 54525 5640 54725 5725
rect 54875 5765 55075 5840
rect 54875 5725 54955 5765
rect 54995 5725 55075 5765
rect 54875 5640 55075 5725
rect 55225 5765 55425 5840
rect 55225 5725 55305 5765
rect 55345 5725 55425 5765
rect 55225 5640 55425 5725
rect 55575 5765 55775 5840
rect 55575 5725 55655 5765
rect 55695 5725 55775 5765
rect 55575 5640 55775 5725
rect 55925 5765 56125 5840
rect 55925 5725 56005 5765
rect 56045 5725 56125 5765
rect 55925 5640 56125 5725
rect 56275 5765 56475 5840
rect 56275 5725 56355 5765
rect 56395 5725 56475 5765
rect 56275 5640 56475 5725
rect 56625 5765 56825 5840
rect 56625 5725 56705 5765
rect 56745 5725 56825 5765
rect 56625 5640 56825 5725
rect 56975 5765 57175 5840
rect 56975 5725 57055 5765
rect 57095 5725 57175 5765
rect 56975 5640 57175 5725
rect 57325 5765 57525 5840
rect 57325 5725 57405 5765
rect 57445 5725 57525 5765
rect 57325 5640 57525 5725
rect 57675 5765 57875 5840
rect 57675 5725 57755 5765
rect 57795 5725 57875 5765
rect 57675 5640 57875 5725
rect 58025 5765 58225 5840
rect 58025 5725 58105 5765
rect 58145 5725 58225 5765
rect 58025 5640 58225 5725
rect 58375 5765 58575 5840
rect 58375 5725 58455 5765
rect 58495 5725 58575 5765
rect 58375 5640 58575 5725
rect 58725 5765 58925 5840
rect 58725 5725 58805 5765
rect 58845 5725 58925 5765
rect 58725 5640 58925 5725
rect 59075 5765 59275 5840
rect 59075 5725 59155 5765
rect 59195 5725 59275 5765
rect 59075 5640 59275 5725
rect 59425 5765 59625 5840
rect 59425 5725 59505 5765
rect 59545 5725 59625 5765
rect 59425 5640 59625 5725
rect 59775 5765 59975 5840
rect 59775 5725 59855 5765
rect 59895 5725 59975 5765
rect 59775 5640 59975 5725
rect 60125 5765 60325 5840
rect 60125 5725 60205 5765
rect 60245 5725 60325 5765
rect 60125 5640 60325 5725
rect 60475 5765 60675 5840
rect 60475 5725 60555 5765
rect 60595 5725 60675 5765
rect 60475 5640 60675 5725
rect 60825 5765 61025 5840
rect 60825 5725 60905 5765
rect 60945 5725 61025 5765
rect 60825 5640 61025 5725
rect 61175 5765 61375 5840
rect 61175 5725 61255 5765
rect 61295 5725 61375 5765
rect 61175 5640 61375 5725
rect 52425 5415 52625 5490
rect 52425 5375 52505 5415
rect 52545 5375 52625 5415
rect 52425 5290 52625 5375
rect 52775 5415 52975 5490
rect 52775 5375 52855 5415
rect 52895 5375 52975 5415
rect 52775 5290 52975 5375
rect 53125 5415 53325 5490
rect 53125 5375 53205 5415
rect 53245 5375 53325 5415
rect 53125 5290 53325 5375
rect 53475 5415 53675 5490
rect 53475 5375 53555 5415
rect 53595 5375 53675 5415
rect 53475 5290 53675 5375
rect 53825 5415 54025 5490
rect 53825 5375 53905 5415
rect 53945 5375 54025 5415
rect 53825 5290 54025 5375
rect 54175 5415 54375 5490
rect 54175 5375 54255 5415
rect 54295 5375 54375 5415
rect 54175 5290 54375 5375
rect 54525 5415 54725 5490
rect 54525 5375 54605 5415
rect 54645 5375 54725 5415
rect 54525 5290 54725 5375
rect 54875 5415 55075 5490
rect 54875 5375 54955 5415
rect 54995 5375 55075 5415
rect 54875 5290 55075 5375
rect 55225 5415 55425 5490
rect 55225 5375 55305 5415
rect 55345 5375 55425 5415
rect 55225 5290 55425 5375
rect 55575 5415 55775 5490
rect 55575 5375 55655 5415
rect 55695 5375 55775 5415
rect 55575 5290 55775 5375
rect 55925 5415 56125 5490
rect 55925 5375 56005 5415
rect 56045 5375 56125 5415
rect 55925 5290 56125 5375
rect 56275 5415 56475 5490
rect 56275 5375 56355 5415
rect 56395 5375 56475 5415
rect 56275 5290 56475 5375
rect 56625 5415 56825 5490
rect 56625 5375 56705 5415
rect 56745 5375 56825 5415
rect 56625 5290 56825 5375
rect 56975 5415 57175 5490
rect 56975 5375 57055 5415
rect 57095 5375 57175 5415
rect 56975 5290 57175 5375
rect 57325 5415 57525 5490
rect 57325 5375 57405 5415
rect 57445 5375 57525 5415
rect 57325 5290 57525 5375
rect 57675 5415 57875 5490
rect 57675 5375 57755 5415
rect 57795 5375 57875 5415
rect 57675 5290 57875 5375
rect 58025 5415 58225 5490
rect 58025 5375 58105 5415
rect 58145 5375 58225 5415
rect 58025 5290 58225 5375
rect 58375 5415 58575 5490
rect 58375 5375 58455 5415
rect 58495 5375 58575 5415
rect 58375 5290 58575 5375
rect 58725 5415 58925 5490
rect 58725 5375 58805 5415
rect 58845 5375 58925 5415
rect 58725 5290 58925 5375
rect 59075 5415 59275 5490
rect 59075 5375 59155 5415
rect 59195 5375 59275 5415
rect 59075 5290 59275 5375
rect 59425 5415 59625 5490
rect 59425 5375 59505 5415
rect 59545 5375 59625 5415
rect 59425 5290 59625 5375
rect 59775 5415 59975 5490
rect 59775 5375 59855 5415
rect 59895 5375 59975 5415
rect 59775 5290 59975 5375
rect 60125 5415 60325 5490
rect 60125 5375 60205 5415
rect 60245 5375 60325 5415
rect 60125 5290 60325 5375
rect 60475 5415 60675 5490
rect 60475 5375 60555 5415
rect 60595 5375 60675 5415
rect 60475 5290 60675 5375
rect 60825 5415 61025 5490
rect 60825 5375 60905 5415
rect 60945 5375 61025 5415
rect 60825 5290 61025 5375
rect 61175 5415 61375 5490
rect 61175 5375 61255 5415
rect 61295 5375 61375 5415
rect 61175 5290 61375 5375
rect 52425 5065 52625 5140
rect 52425 5025 52505 5065
rect 52545 5025 52625 5065
rect 52425 4940 52625 5025
rect 52775 5065 52975 5140
rect 52775 5025 52855 5065
rect 52895 5025 52975 5065
rect 52775 4940 52975 5025
rect 53125 5065 53325 5140
rect 53125 5025 53205 5065
rect 53245 5025 53325 5065
rect 53125 4940 53325 5025
rect 53475 5065 53675 5140
rect 53475 5025 53555 5065
rect 53595 5025 53675 5065
rect 53475 4940 53675 5025
rect 53825 5065 54025 5140
rect 53825 5025 53905 5065
rect 53945 5025 54025 5065
rect 53825 4940 54025 5025
rect 54175 5065 54375 5140
rect 54175 5025 54255 5065
rect 54295 5025 54375 5065
rect 54175 4940 54375 5025
rect 54525 5065 54725 5140
rect 54525 5025 54605 5065
rect 54645 5025 54725 5065
rect 54525 4940 54725 5025
rect 54875 5065 55075 5140
rect 54875 5025 54955 5065
rect 54995 5025 55075 5065
rect 54875 4940 55075 5025
rect 55225 5065 55425 5140
rect 55225 5025 55305 5065
rect 55345 5025 55425 5065
rect 55225 4940 55425 5025
rect 55575 5055 55775 5140
rect 55575 5015 55655 5055
rect 55695 5015 55775 5055
rect 55575 4940 55775 5015
rect 55925 5055 56125 5140
rect 55925 5015 56005 5055
rect 56045 5015 56125 5055
rect 55925 4940 56125 5015
rect 56275 5055 56475 5140
rect 56275 5015 56355 5055
rect 56395 5015 56475 5055
rect 56275 4940 56475 5015
rect 56625 5055 56825 5140
rect 56625 5015 56705 5055
rect 56745 5015 56825 5055
rect 56625 4940 56825 5015
rect 56975 5055 57175 5140
rect 56975 5015 57055 5055
rect 57095 5015 57175 5055
rect 56975 4940 57175 5015
rect 57325 5055 57525 5140
rect 57325 5015 57405 5055
rect 57445 5015 57525 5055
rect 57325 4940 57525 5015
rect 57675 5055 57875 5140
rect 57675 5015 57755 5055
rect 57795 5015 57875 5055
rect 57675 4940 57875 5015
rect 58025 5055 58225 5140
rect 58025 5015 58105 5055
rect 58145 5015 58225 5055
rect 58025 4940 58225 5015
rect 58375 5065 58575 5140
rect 58375 5025 58455 5065
rect 58495 5025 58575 5065
rect 58375 4940 58575 5025
rect 58725 5065 58925 5140
rect 58725 5025 58805 5065
rect 58845 5025 58925 5065
rect 58725 4940 58925 5025
rect 59075 5065 59275 5140
rect 59075 5025 59155 5065
rect 59195 5025 59275 5065
rect 59075 4940 59275 5025
rect 59425 5065 59625 5140
rect 59425 5025 59505 5065
rect 59545 5025 59625 5065
rect 59425 4940 59625 5025
rect 59775 5065 59975 5140
rect 59775 5025 59855 5065
rect 59895 5025 59975 5065
rect 59775 4940 59975 5025
rect 60125 5065 60325 5140
rect 60125 5025 60205 5065
rect 60245 5025 60325 5065
rect 60125 4940 60325 5025
rect 60475 5065 60675 5140
rect 60475 5025 60555 5065
rect 60595 5025 60675 5065
rect 60475 4940 60675 5025
rect 60825 5065 61025 5140
rect 60825 5025 60905 5065
rect 60945 5025 61025 5065
rect 60825 4940 61025 5025
rect 61175 5065 61375 5140
rect 61175 5025 61255 5065
rect 61295 5025 61375 5065
rect 61175 4940 61375 5025
rect 52425 4715 52625 4790
rect 52425 4675 52505 4715
rect 52545 4675 52625 4715
rect 52425 4590 52625 4675
rect 52775 4715 52975 4790
rect 52775 4675 52855 4715
rect 52895 4675 52975 4715
rect 52775 4590 52975 4675
rect 53125 4715 53325 4790
rect 53125 4675 53205 4715
rect 53245 4675 53325 4715
rect 53125 4590 53325 4675
rect 53475 4715 53675 4790
rect 53475 4675 53555 4715
rect 53595 4675 53675 4715
rect 53475 4590 53675 4675
rect 53825 4715 54025 4790
rect 53825 4675 53905 4715
rect 53945 4675 54025 4715
rect 53825 4590 54025 4675
rect 54175 4715 54375 4790
rect 54175 4675 54255 4715
rect 54295 4675 54375 4715
rect 54175 4590 54375 4675
rect 54525 4715 54725 4790
rect 54525 4675 54605 4715
rect 54645 4675 54725 4715
rect 54525 4590 54725 4675
rect 54875 4715 55075 4790
rect 54875 4675 54955 4715
rect 54995 4675 55075 4715
rect 54875 4590 55075 4675
rect 55225 4715 55425 4790
rect 55225 4675 55305 4715
rect 55345 4675 55425 4715
rect 55225 4590 55425 4675
rect 58375 4715 58575 4790
rect 58375 4675 58455 4715
rect 58495 4675 58575 4715
rect 58375 4590 58575 4675
rect 58725 4715 58925 4790
rect 58725 4675 58805 4715
rect 58845 4675 58925 4715
rect 58725 4590 58925 4675
rect 59075 4715 59275 4790
rect 59075 4675 59155 4715
rect 59195 4675 59275 4715
rect 59075 4590 59275 4675
rect 59425 4715 59625 4790
rect 59425 4675 59505 4715
rect 59545 4675 59625 4715
rect 59425 4590 59625 4675
rect 59775 4715 59975 4790
rect 59775 4675 59855 4715
rect 59895 4675 59975 4715
rect 59775 4590 59975 4675
rect 60125 4715 60325 4790
rect 60125 4675 60205 4715
rect 60245 4675 60325 4715
rect 60125 4590 60325 4675
rect 60475 4715 60675 4790
rect 60475 4675 60555 4715
rect 60595 4675 60675 4715
rect 60475 4590 60675 4675
rect 60825 4715 61025 4790
rect 60825 4675 60905 4715
rect 60945 4675 61025 4715
rect 60825 4590 61025 4675
rect 61175 4715 61375 4790
rect 61175 4675 61255 4715
rect 61295 4675 61375 4715
rect 61175 4590 61375 4675
rect 52425 4365 52625 4440
rect 52425 4325 52505 4365
rect 52545 4325 52625 4365
rect 52425 4240 52625 4325
rect 52775 4365 52975 4440
rect 52775 4325 52855 4365
rect 52895 4325 52975 4365
rect 52775 4240 52975 4325
rect 53125 4365 53325 4440
rect 53125 4325 53205 4365
rect 53245 4325 53325 4365
rect 53125 4240 53325 4325
rect 53475 4365 53675 4440
rect 53475 4325 53555 4365
rect 53595 4325 53675 4365
rect 53475 4240 53675 4325
rect 53825 4365 54025 4440
rect 53825 4325 53905 4365
rect 53945 4325 54025 4365
rect 53825 4240 54025 4325
rect 54175 4365 54375 4440
rect 54175 4325 54255 4365
rect 54295 4325 54375 4365
rect 54175 4240 54375 4325
rect 54525 4365 54725 4440
rect 54525 4325 54605 4365
rect 54645 4325 54725 4365
rect 54525 4240 54725 4325
rect 54875 4365 55075 4440
rect 54875 4325 54955 4365
rect 54995 4325 55075 4365
rect 54875 4240 55075 4325
rect 55225 4365 55425 4440
rect 55225 4325 55305 4365
rect 55345 4325 55425 4365
rect 55225 4240 55425 4325
rect 58375 4365 58575 4440
rect 58375 4325 58455 4365
rect 58495 4325 58575 4365
rect 58375 4240 58575 4325
rect 58725 4365 58925 4440
rect 58725 4325 58805 4365
rect 58845 4325 58925 4365
rect 58725 4240 58925 4325
rect 59075 4365 59275 4440
rect 59075 4325 59155 4365
rect 59195 4325 59275 4365
rect 59075 4240 59275 4325
rect 59425 4365 59625 4440
rect 59425 4325 59505 4365
rect 59545 4325 59625 4365
rect 59425 4240 59625 4325
rect 59775 4365 59975 4440
rect 59775 4325 59855 4365
rect 59895 4325 59975 4365
rect 59775 4240 59975 4325
rect 60125 4365 60325 4440
rect 60125 4325 60205 4365
rect 60245 4325 60325 4365
rect 60125 4240 60325 4325
rect 60475 4365 60675 4440
rect 60475 4325 60555 4365
rect 60595 4325 60675 4365
rect 60475 4240 60675 4325
rect 60825 4365 61025 4440
rect 60825 4325 60905 4365
rect 60945 4325 61025 4365
rect 60825 4240 61025 4325
rect 61175 4365 61375 4440
rect 61175 4325 61255 4365
rect 61295 4325 61375 4365
rect 61175 4240 61375 4325
rect 52425 4015 52625 4090
rect 52425 3975 52505 4015
rect 52545 3975 52625 4015
rect 52425 3890 52625 3975
rect 52775 4015 52975 4090
rect 52775 3975 52855 4015
rect 52895 3975 52975 4015
rect 52775 3890 52975 3975
rect 53125 4015 53325 4090
rect 53125 3975 53205 4015
rect 53245 3975 53325 4015
rect 53125 3890 53325 3975
rect 53475 4015 53675 4090
rect 53475 3975 53555 4015
rect 53595 3975 53675 4015
rect 53475 3890 53675 3975
rect 53825 4015 54025 4090
rect 53825 3975 53905 4015
rect 53945 3975 54025 4015
rect 53825 3890 54025 3975
rect 59775 4015 59975 4090
rect 59775 3975 59855 4015
rect 59895 3975 59975 4015
rect 59775 3890 59975 3975
rect 60125 4015 60325 4090
rect 60125 3975 60205 4015
rect 60245 3975 60325 4015
rect 60125 3890 60325 3975
rect 60475 4015 60675 4090
rect 60475 3975 60555 4015
rect 60595 3975 60675 4015
rect 60475 3890 60675 3975
rect 60825 4015 61025 4090
rect 60825 3975 60905 4015
rect 60945 3975 61025 4015
rect 60825 3890 61025 3975
rect 61175 4015 61375 4090
rect 61175 3975 61255 4015
rect 61295 3975 61375 4015
rect 61175 3890 61375 3975
rect 52425 3665 52625 3740
rect 52425 3625 52505 3665
rect 52545 3625 52625 3665
rect 52425 3540 52625 3625
rect 52775 3665 52975 3740
rect 52775 3625 52855 3665
rect 52895 3625 52975 3665
rect 52775 3540 52975 3625
rect 53125 3665 53325 3740
rect 53125 3625 53205 3665
rect 53245 3625 53325 3665
rect 53125 3540 53325 3625
rect 53475 3665 53675 3740
rect 53475 3625 53555 3665
rect 53595 3625 53675 3665
rect 53475 3540 53675 3625
rect 53825 3665 54025 3740
rect 53825 3625 53905 3665
rect 53945 3625 54025 3665
rect 53825 3540 54025 3625
rect 59775 3665 59975 3740
rect 59775 3625 59855 3665
rect 59895 3625 59975 3665
rect 59775 3540 59975 3625
rect 60125 3665 60325 3740
rect 60125 3625 60205 3665
rect 60245 3625 60325 3665
rect 60125 3540 60325 3625
rect 60475 3665 60675 3740
rect 60475 3625 60555 3665
rect 60595 3625 60675 3665
rect 60475 3540 60675 3625
rect 60825 3665 61025 3740
rect 60825 3625 60905 3665
rect 60945 3625 61025 3665
rect 60825 3540 61025 3625
rect 61175 3665 61375 3740
rect 61175 3625 61255 3665
rect 61295 3625 61375 3665
rect 61175 3540 61375 3625
rect 52425 3315 52625 3390
rect 52425 3275 52505 3315
rect 52545 3275 52625 3315
rect 52425 3190 52625 3275
rect 52775 3315 52975 3390
rect 52775 3275 52855 3315
rect 52895 3275 52975 3315
rect 52775 3190 52975 3275
rect 53125 3315 53325 3390
rect 53125 3275 53205 3315
rect 53245 3275 53325 3315
rect 53125 3190 53325 3275
rect 53475 3315 53675 3390
rect 53475 3275 53555 3315
rect 53595 3275 53675 3315
rect 53475 3190 53675 3275
rect 53825 3315 54025 3390
rect 53825 3275 53905 3315
rect 53945 3275 54025 3315
rect 53825 3190 54025 3275
rect 59775 3315 59975 3390
rect 59775 3275 59855 3315
rect 59895 3275 59975 3315
rect 59775 3190 59975 3275
rect 60125 3315 60325 3390
rect 60125 3275 60205 3315
rect 60245 3275 60325 3315
rect 60125 3190 60325 3275
rect 60475 3315 60675 3390
rect 60475 3275 60555 3315
rect 60595 3275 60675 3315
rect 60475 3190 60675 3275
rect 60825 3315 61025 3390
rect 60825 3275 60905 3315
rect 60945 3275 61025 3315
rect 60825 3190 61025 3275
rect 61175 3315 61375 3390
rect 61175 3275 61255 3315
rect 61295 3275 61375 3315
rect 61175 3190 61375 3275
rect 52425 2965 52625 3040
rect 52425 2925 52505 2965
rect 52545 2925 52625 2965
rect 52425 2840 52625 2925
rect 52775 2965 52975 3040
rect 52775 2925 52855 2965
rect 52895 2925 52975 2965
rect 52775 2840 52975 2925
rect 53125 2965 53325 3040
rect 53125 2925 53205 2965
rect 53245 2925 53325 2965
rect 53125 2840 53325 2925
rect 53475 2965 53675 3040
rect 53475 2925 53555 2965
rect 53595 2925 53675 2965
rect 53475 2840 53675 2925
rect 53825 2965 54025 3040
rect 53825 2925 53905 2965
rect 53945 2925 54025 2965
rect 53825 2840 54025 2925
rect 59775 2965 59975 3040
rect 59775 2925 59855 2965
rect 59895 2925 59975 2965
rect 59775 2840 59975 2925
rect 60125 2965 60325 3040
rect 60125 2925 60205 2965
rect 60245 2925 60325 2965
rect 60125 2840 60325 2925
rect 60475 2965 60675 3040
rect 60475 2925 60555 2965
rect 60595 2925 60675 2965
rect 60475 2840 60675 2925
rect 60825 2965 61025 3040
rect 60825 2925 60905 2965
rect 60945 2925 61025 2965
rect 60825 2840 61025 2925
rect 61175 2965 61375 3040
rect 61175 2925 61255 2965
rect 61295 2925 61375 2965
rect 61175 2840 61375 2925
rect 52425 2615 52625 2690
rect 52425 2575 52505 2615
rect 52545 2575 52625 2615
rect 52425 2490 52625 2575
rect 52775 2615 52975 2690
rect 52775 2575 52855 2615
rect 52895 2575 52975 2615
rect 52775 2490 52975 2575
rect 53125 2615 53325 2690
rect 53125 2575 53205 2615
rect 53245 2575 53325 2615
rect 53125 2490 53325 2575
rect 53475 2615 53675 2690
rect 53475 2575 53555 2615
rect 53595 2575 53675 2615
rect 53475 2490 53675 2575
rect 53825 2615 54025 2690
rect 53825 2575 53905 2615
rect 53945 2575 54025 2615
rect 53825 2490 54025 2575
rect 59775 2615 59975 2690
rect 59775 2575 59855 2615
rect 59895 2575 59975 2615
rect 59775 2490 59975 2575
rect 60125 2615 60325 2690
rect 60125 2575 60205 2615
rect 60245 2575 60325 2615
rect 60125 2490 60325 2575
rect 60475 2615 60675 2690
rect 60475 2575 60555 2615
rect 60595 2575 60675 2615
rect 60475 2490 60675 2575
rect 60825 2615 61025 2690
rect 60825 2575 60905 2615
rect 60945 2575 61025 2615
rect 60825 2490 61025 2575
rect 61175 2615 61375 2690
rect 61175 2575 61255 2615
rect 61295 2575 61375 2615
rect 61175 2490 61375 2575
rect 52425 2265 52625 2340
rect 52425 2225 52505 2265
rect 52545 2225 52625 2265
rect 52425 2140 52625 2225
rect 52775 2265 52975 2340
rect 52775 2225 52855 2265
rect 52895 2225 52975 2265
rect 52775 2140 52975 2225
rect 53125 2265 53325 2340
rect 53125 2225 53205 2265
rect 53245 2225 53325 2265
rect 53125 2140 53325 2225
rect 53475 2265 53675 2340
rect 53475 2225 53555 2265
rect 53595 2225 53675 2265
rect 53475 2140 53675 2225
rect 53825 2265 54025 2340
rect 53825 2225 53905 2265
rect 53945 2225 54025 2265
rect 53825 2140 54025 2225
rect 59775 2265 59975 2340
rect 59775 2225 59855 2265
rect 59895 2225 59975 2265
rect 59775 2140 59975 2225
rect 60125 2265 60325 2340
rect 60125 2225 60205 2265
rect 60245 2225 60325 2265
rect 60125 2140 60325 2225
rect 60475 2265 60675 2340
rect 60475 2225 60555 2265
rect 60595 2225 60675 2265
rect 60475 2140 60675 2225
rect 60825 2265 61025 2340
rect 60825 2225 60905 2265
rect 60945 2225 61025 2265
rect 60825 2140 61025 2225
rect 61175 2265 61375 2340
rect 61175 2225 61255 2265
rect 61295 2225 61375 2265
rect 61175 2140 61375 2225
rect 52425 1915 52625 1990
rect 52425 1875 52505 1915
rect 52545 1875 52625 1915
rect 52425 1790 52625 1875
rect 52775 1915 52975 1990
rect 52775 1875 52855 1915
rect 52895 1875 52975 1915
rect 52775 1790 52975 1875
rect 53125 1915 53325 1990
rect 53125 1875 53205 1915
rect 53245 1875 53325 1915
rect 53125 1790 53325 1875
rect 53475 1915 53675 1990
rect 53475 1875 53555 1915
rect 53595 1875 53675 1915
rect 53475 1790 53675 1875
rect 53825 1915 54025 1990
rect 53825 1875 53905 1915
rect 53945 1875 54025 1915
rect 53825 1790 54025 1875
rect 59775 1915 59975 1990
rect 59775 1875 59855 1915
rect 59895 1875 59975 1915
rect 59775 1790 59975 1875
rect 60125 1915 60325 1990
rect 60125 1875 60205 1915
rect 60245 1875 60325 1915
rect 60125 1790 60325 1875
rect 60475 1915 60675 1990
rect 60475 1875 60555 1915
rect 60595 1875 60675 1915
rect 60475 1790 60675 1875
rect 60825 1915 61025 1990
rect 60825 1875 60905 1915
rect 60945 1875 61025 1915
rect 60825 1790 61025 1875
rect 61175 1915 61375 1990
rect 61175 1875 61255 1915
rect 61295 1875 61375 1915
rect 61175 1790 61375 1875
rect 52425 1565 52625 1640
rect 52425 1525 52505 1565
rect 52545 1525 52625 1565
rect 52425 1440 52625 1525
rect 52775 1565 52975 1640
rect 52775 1525 52855 1565
rect 52895 1525 52975 1565
rect 52775 1440 52975 1525
rect 53125 1565 53325 1640
rect 53125 1525 53205 1565
rect 53245 1525 53325 1565
rect 53125 1440 53325 1525
rect 53475 1565 53675 1640
rect 53475 1525 53555 1565
rect 53595 1525 53675 1565
rect 53475 1440 53675 1525
rect 53825 1565 54025 1640
rect 53825 1525 53905 1565
rect 53945 1525 54025 1565
rect 53825 1440 54025 1525
rect 59775 1565 59975 1640
rect 59775 1525 59855 1565
rect 59895 1525 59975 1565
rect 59775 1440 59975 1525
rect 60125 1565 60325 1640
rect 60125 1525 60205 1565
rect 60245 1525 60325 1565
rect 60125 1440 60325 1525
rect 60475 1565 60675 1640
rect 60475 1525 60555 1565
rect 60595 1525 60675 1565
rect 60475 1440 60675 1525
rect 60825 1565 61025 1640
rect 60825 1525 60905 1565
rect 60945 1525 61025 1565
rect 60825 1440 61025 1525
rect 61175 1565 61375 1640
rect 61175 1525 61255 1565
rect 61295 1525 61375 1565
rect 61175 1440 61375 1525
rect 52425 1215 52625 1290
rect 52425 1175 52505 1215
rect 52545 1175 52625 1215
rect 52425 1090 52625 1175
rect 52775 1215 52975 1290
rect 52775 1175 52855 1215
rect 52895 1175 52975 1215
rect 52775 1090 52975 1175
rect 53125 1215 53325 1290
rect 53125 1175 53205 1215
rect 53245 1175 53325 1215
rect 53125 1090 53325 1175
rect 53475 1215 53675 1290
rect 53475 1175 53555 1215
rect 53595 1175 53675 1215
rect 53475 1090 53675 1175
rect 53825 1215 54025 1290
rect 53825 1175 53905 1215
rect 53945 1175 54025 1215
rect 53825 1090 54025 1175
rect 59775 1215 59975 1290
rect 59775 1175 59855 1215
rect 59895 1175 59975 1215
rect 59775 1090 59975 1175
rect 60125 1215 60325 1290
rect 60125 1175 60205 1215
rect 60245 1175 60325 1215
rect 60125 1090 60325 1175
rect 60475 1215 60675 1290
rect 60475 1175 60555 1215
rect 60595 1175 60675 1215
rect 60475 1090 60675 1175
rect 60825 1215 61025 1290
rect 60825 1175 60905 1215
rect 60945 1175 61025 1215
rect 60825 1090 61025 1175
rect 61175 1215 61375 1290
rect 61175 1175 61255 1215
rect 61295 1175 61375 1215
rect 61175 1090 61375 1175
rect 52425 865 52625 940
rect 52425 825 52505 865
rect 52545 825 52625 865
rect 52425 740 52625 825
rect 52775 865 52975 940
rect 52775 825 52855 865
rect 52895 825 52975 865
rect 52775 740 52975 825
rect 53125 865 53325 940
rect 53125 825 53205 865
rect 53245 825 53325 865
rect 53125 740 53325 825
rect 53475 865 53675 940
rect 53475 825 53555 865
rect 53595 825 53675 865
rect 53475 740 53675 825
rect 53825 865 54025 940
rect 53825 825 53905 865
rect 53945 825 54025 865
rect 53825 740 54025 825
rect 59775 865 59975 940
rect 59775 825 59855 865
rect 59895 825 59975 865
rect 59775 740 59975 825
rect 60125 865 60325 940
rect 60125 825 60205 865
rect 60245 825 60325 865
rect 60125 740 60325 825
rect 60475 865 60675 940
rect 60475 825 60555 865
rect 60595 825 60675 865
rect 60475 740 60675 825
rect 60825 865 61025 940
rect 60825 825 60905 865
rect 60945 825 61025 865
rect 60825 740 61025 825
rect 61175 865 61375 940
rect 61175 825 61255 865
rect 61295 825 61375 865
rect 61175 740 61375 825
rect 52425 515 52625 590
rect 52425 475 52505 515
rect 52545 475 52625 515
rect 52425 390 52625 475
rect 52775 515 52975 590
rect 52775 475 52855 515
rect 52895 475 52975 515
rect 52775 390 52975 475
rect 53125 515 53325 590
rect 53125 475 53205 515
rect 53245 475 53325 515
rect 53125 390 53325 475
rect 53475 515 53675 590
rect 53475 475 53555 515
rect 53595 475 53675 515
rect 53475 390 53675 475
rect 53825 515 54025 590
rect 53825 475 53905 515
rect 53945 475 54025 515
rect 53825 390 54025 475
rect 59775 515 59975 590
rect 59775 475 59855 515
rect 59895 475 59975 515
rect 59775 390 59975 475
rect 60125 515 60325 590
rect 60125 475 60205 515
rect 60245 475 60325 515
rect 60125 390 60325 475
rect 60475 515 60675 590
rect 60475 475 60555 515
rect 60595 475 60675 515
rect 60475 390 60675 475
rect 60825 515 61025 590
rect 60825 475 60905 515
rect 60945 475 61025 515
rect 60825 390 61025 475
rect 61175 515 61375 590
rect 61175 475 61255 515
rect 61295 475 61375 515
rect 61175 390 61375 475
rect 52425 165 52625 240
rect 52425 125 52505 165
rect 52545 125 52625 165
rect 52425 40 52625 125
rect 52775 165 52975 240
rect 52775 125 52855 165
rect 52895 125 52975 165
rect 52775 40 52975 125
rect 53125 165 53325 240
rect 53125 125 53205 165
rect 53245 125 53325 165
rect 53125 40 53325 125
rect 53475 165 53675 240
rect 53475 125 53555 165
rect 53595 125 53675 165
rect 53475 40 53675 125
rect 53825 165 54025 240
rect 53825 125 53905 165
rect 53945 125 54025 165
rect 53825 40 54025 125
rect 54175 165 54375 240
rect 54175 125 54255 165
rect 54295 125 54375 165
rect 54175 40 54375 125
rect 54525 165 54725 240
rect 54525 125 54605 165
rect 54645 125 54725 165
rect 54525 40 54725 125
rect 54875 165 55075 240
rect 54875 125 54955 165
rect 54995 125 55075 165
rect 54875 40 55075 125
rect 55225 165 55425 240
rect 55225 125 55305 165
rect 55345 125 55425 165
rect 55225 40 55425 125
rect 55575 165 55775 240
rect 55575 125 55655 165
rect 55695 125 55775 165
rect 55575 40 55775 125
rect 55925 165 56125 240
rect 55925 125 56005 165
rect 56045 125 56125 165
rect 55925 40 56125 125
rect 56275 165 56475 240
rect 56275 125 56355 165
rect 56395 125 56475 165
rect 56275 40 56475 125
rect 56625 165 56825 240
rect 56625 125 56705 165
rect 56745 125 56825 165
rect 56625 40 56825 125
rect 56975 165 57175 240
rect 56975 125 57055 165
rect 57095 125 57175 165
rect 56975 40 57175 125
rect 57325 165 57525 240
rect 57325 125 57405 165
rect 57445 125 57525 165
rect 57325 40 57525 125
rect 57675 165 57875 240
rect 57675 125 57755 165
rect 57795 125 57875 165
rect 57675 40 57875 125
rect 58025 165 58225 240
rect 58025 125 58105 165
rect 58145 125 58225 165
rect 58025 40 58225 125
rect 58375 165 58575 240
rect 58375 125 58455 165
rect 58495 125 58575 165
rect 58375 40 58575 125
rect 58725 165 58925 240
rect 58725 125 58805 165
rect 58845 125 58925 165
rect 58725 40 58925 125
rect 59075 165 59275 240
rect 59075 125 59155 165
rect 59195 125 59275 165
rect 59075 40 59275 125
rect 59425 165 59625 240
rect 59425 125 59505 165
rect 59545 125 59625 165
rect 59425 40 59625 125
rect 59775 165 59975 240
rect 59775 125 59855 165
rect 59895 125 59975 165
rect 59775 40 59975 125
rect 60125 165 60325 240
rect 60125 125 60205 165
rect 60245 125 60325 165
rect 60125 40 60325 125
rect 60475 165 60675 240
rect 60475 125 60555 165
rect 60595 125 60675 165
rect 60475 40 60675 125
rect 60825 165 61025 240
rect 60825 125 60905 165
rect 60945 125 61025 165
rect 60825 40 61025 125
rect 61175 165 61375 240
rect 61175 125 61255 165
rect 61295 125 61375 165
rect 61175 40 61375 125
rect 52425 -185 52625 -110
rect 52425 -225 52505 -185
rect 52545 -225 52625 -185
rect 52425 -310 52625 -225
rect 52775 -185 52975 -110
rect 52775 -225 52855 -185
rect 52895 -225 52975 -185
rect 52775 -310 52975 -225
rect 53125 -185 53325 -110
rect 53125 -225 53205 -185
rect 53245 -225 53325 -185
rect 53125 -310 53325 -225
rect 53475 -185 53675 -110
rect 53475 -225 53555 -185
rect 53595 -225 53675 -185
rect 53475 -310 53675 -225
rect 53825 -185 54025 -110
rect 53825 -225 53905 -185
rect 53945 -225 54025 -185
rect 53825 -310 54025 -225
rect 54175 -185 54375 -110
rect 54175 -225 54255 -185
rect 54295 -225 54375 -185
rect 54175 -310 54375 -225
rect 54525 -185 54725 -110
rect 54525 -225 54605 -185
rect 54645 -225 54725 -185
rect 54525 -310 54725 -225
rect 54875 -185 55075 -110
rect 54875 -225 54955 -185
rect 54995 -225 55075 -185
rect 54875 -310 55075 -225
rect 55225 -185 55425 -110
rect 55225 -225 55305 -185
rect 55345 -225 55425 -185
rect 55225 -310 55425 -225
rect 55575 -185 55775 -110
rect 55575 -225 55655 -185
rect 55695 -225 55775 -185
rect 55575 -310 55775 -225
rect 55925 -185 56125 -110
rect 55925 -225 56005 -185
rect 56045 -225 56125 -185
rect 55925 -310 56125 -225
rect 56275 -185 56475 -110
rect 56275 -225 56355 -185
rect 56395 -225 56475 -185
rect 56275 -310 56475 -225
rect 56625 -185 56825 -110
rect 56625 -225 56705 -185
rect 56745 -225 56825 -185
rect 56625 -310 56825 -225
rect 56975 -185 57175 -110
rect 56975 -225 57055 -185
rect 57095 -225 57175 -185
rect 56975 -310 57175 -225
rect 57325 -185 57525 -110
rect 57325 -225 57405 -185
rect 57445 -225 57525 -185
rect 57325 -310 57525 -225
rect 57675 -185 57875 -110
rect 57675 -225 57755 -185
rect 57795 -225 57875 -185
rect 57675 -310 57875 -225
rect 58025 -185 58225 -110
rect 58025 -225 58105 -185
rect 58145 -225 58225 -185
rect 58025 -310 58225 -225
rect 58375 -185 58575 -110
rect 58375 -225 58455 -185
rect 58495 -225 58575 -185
rect 58375 -310 58575 -225
rect 58725 -185 58925 -110
rect 58725 -225 58805 -185
rect 58845 -225 58925 -185
rect 58725 -310 58925 -225
rect 59075 -185 59275 -110
rect 59075 -225 59155 -185
rect 59195 -225 59275 -185
rect 59075 -310 59275 -225
rect 59425 -185 59625 -110
rect 59425 -225 59505 -185
rect 59545 -225 59625 -185
rect 59425 -310 59625 -225
rect 59775 -185 59975 -110
rect 59775 -225 59855 -185
rect 59895 -225 59975 -185
rect 59775 -310 59975 -225
rect 60125 -185 60325 -110
rect 60125 -225 60205 -185
rect 60245 -225 60325 -185
rect 60125 -310 60325 -225
rect 60475 -185 60675 -110
rect 60475 -225 60555 -185
rect 60595 -225 60675 -185
rect 60475 -310 60675 -225
rect 60825 -185 61025 -110
rect 60825 -225 60905 -185
rect 60945 -225 61025 -185
rect 60825 -310 61025 -225
rect 61175 -185 61375 -110
rect 61175 -225 61255 -185
rect 61295 -225 61375 -185
rect 61175 -310 61375 -225
<< mimcapcontact >>
rect 52505 5725 52545 5765
rect 52855 5725 52895 5765
rect 53205 5725 53245 5765
rect 53555 5725 53595 5765
rect 53905 5725 53945 5765
rect 54255 5725 54295 5765
rect 54605 5725 54645 5765
rect 54955 5725 54995 5765
rect 55305 5725 55345 5765
rect 55655 5725 55695 5765
rect 56005 5725 56045 5765
rect 56355 5725 56395 5765
rect 56705 5725 56745 5765
rect 57055 5725 57095 5765
rect 57405 5725 57445 5765
rect 57755 5725 57795 5765
rect 58105 5725 58145 5765
rect 58455 5725 58495 5765
rect 58805 5725 58845 5765
rect 59155 5725 59195 5765
rect 59505 5725 59545 5765
rect 59855 5725 59895 5765
rect 60205 5725 60245 5765
rect 60555 5725 60595 5765
rect 60905 5725 60945 5765
rect 61255 5725 61295 5765
rect 52505 5375 52545 5415
rect 52855 5375 52895 5415
rect 53205 5375 53245 5415
rect 53555 5375 53595 5415
rect 53905 5375 53945 5415
rect 54255 5375 54295 5415
rect 54605 5375 54645 5415
rect 54955 5375 54995 5415
rect 55305 5375 55345 5415
rect 55655 5375 55695 5415
rect 56005 5375 56045 5415
rect 56355 5375 56395 5415
rect 56705 5375 56745 5415
rect 57055 5375 57095 5415
rect 57405 5375 57445 5415
rect 57755 5375 57795 5415
rect 58105 5375 58145 5415
rect 58455 5375 58495 5415
rect 58805 5375 58845 5415
rect 59155 5375 59195 5415
rect 59505 5375 59545 5415
rect 59855 5375 59895 5415
rect 60205 5375 60245 5415
rect 60555 5375 60595 5415
rect 60905 5375 60945 5415
rect 61255 5375 61295 5415
rect 52505 5025 52545 5065
rect 52855 5025 52895 5065
rect 53205 5025 53245 5065
rect 53555 5025 53595 5065
rect 53905 5025 53945 5065
rect 54255 5025 54295 5065
rect 54605 5025 54645 5065
rect 54955 5025 54995 5065
rect 55305 5025 55345 5065
rect 55655 5015 55695 5055
rect 56005 5015 56045 5055
rect 56355 5015 56395 5055
rect 56705 5015 56745 5055
rect 57055 5015 57095 5055
rect 57405 5015 57445 5055
rect 57755 5015 57795 5055
rect 58105 5015 58145 5055
rect 58455 5025 58495 5065
rect 58805 5025 58845 5065
rect 59155 5025 59195 5065
rect 59505 5025 59545 5065
rect 59855 5025 59895 5065
rect 60205 5025 60245 5065
rect 60555 5025 60595 5065
rect 60905 5025 60945 5065
rect 61255 5025 61295 5065
rect 52505 4675 52545 4715
rect 52855 4675 52895 4715
rect 53205 4675 53245 4715
rect 53555 4675 53595 4715
rect 53905 4675 53945 4715
rect 54255 4675 54295 4715
rect 54605 4675 54645 4715
rect 54955 4675 54995 4715
rect 55305 4675 55345 4715
rect 58455 4675 58495 4715
rect 58805 4675 58845 4715
rect 59155 4675 59195 4715
rect 59505 4675 59545 4715
rect 59855 4675 59895 4715
rect 60205 4675 60245 4715
rect 60555 4675 60595 4715
rect 60905 4675 60945 4715
rect 61255 4675 61295 4715
rect 52505 4325 52545 4365
rect 52855 4325 52895 4365
rect 53205 4325 53245 4365
rect 53555 4325 53595 4365
rect 53905 4325 53945 4365
rect 54255 4325 54295 4365
rect 54605 4325 54645 4365
rect 54955 4325 54995 4365
rect 55305 4325 55345 4365
rect 58455 4325 58495 4365
rect 58805 4325 58845 4365
rect 59155 4325 59195 4365
rect 59505 4325 59545 4365
rect 59855 4325 59895 4365
rect 60205 4325 60245 4365
rect 60555 4325 60595 4365
rect 60905 4325 60945 4365
rect 61255 4325 61295 4365
rect 52505 3975 52545 4015
rect 52855 3975 52895 4015
rect 53205 3975 53245 4015
rect 53555 3975 53595 4015
rect 53905 3975 53945 4015
rect 59855 3975 59895 4015
rect 60205 3975 60245 4015
rect 60555 3975 60595 4015
rect 60905 3975 60945 4015
rect 61255 3975 61295 4015
rect 52505 3625 52545 3665
rect 52855 3625 52895 3665
rect 53205 3625 53245 3665
rect 53555 3625 53595 3665
rect 53905 3625 53945 3665
rect 59855 3625 59895 3665
rect 60205 3625 60245 3665
rect 60555 3625 60595 3665
rect 60905 3625 60945 3665
rect 61255 3625 61295 3665
rect 52505 3275 52545 3315
rect 52855 3275 52895 3315
rect 53205 3275 53245 3315
rect 53555 3275 53595 3315
rect 53905 3275 53945 3315
rect 59855 3275 59895 3315
rect 60205 3275 60245 3315
rect 60555 3275 60595 3315
rect 60905 3275 60945 3315
rect 61255 3275 61295 3315
rect 52505 2925 52545 2965
rect 52855 2925 52895 2965
rect 53205 2925 53245 2965
rect 53555 2925 53595 2965
rect 53905 2925 53945 2965
rect 59855 2925 59895 2965
rect 60205 2925 60245 2965
rect 60555 2925 60595 2965
rect 60905 2925 60945 2965
rect 61255 2925 61295 2965
rect 52505 2575 52545 2615
rect 52855 2575 52895 2615
rect 53205 2575 53245 2615
rect 53555 2575 53595 2615
rect 53905 2575 53945 2615
rect 59855 2575 59895 2615
rect 60205 2575 60245 2615
rect 60555 2575 60595 2615
rect 60905 2575 60945 2615
rect 61255 2575 61295 2615
rect 52505 2225 52545 2265
rect 52855 2225 52895 2265
rect 53205 2225 53245 2265
rect 53555 2225 53595 2265
rect 53905 2225 53945 2265
rect 59855 2225 59895 2265
rect 60205 2225 60245 2265
rect 60555 2225 60595 2265
rect 60905 2225 60945 2265
rect 61255 2225 61295 2265
rect 52505 1875 52545 1915
rect 52855 1875 52895 1915
rect 53205 1875 53245 1915
rect 53555 1875 53595 1915
rect 53905 1875 53945 1915
rect 59855 1875 59895 1915
rect 60205 1875 60245 1915
rect 60555 1875 60595 1915
rect 60905 1875 60945 1915
rect 61255 1875 61295 1915
rect 52505 1525 52545 1565
rect 52855 1525 52895 1565
rect 53205 1525 53245 1565
rect 53555 1525 53595 1565
rect 53905 1525 53945 1565
rect 59855 1525 59895 1565
rect 60205 1525 60245 1565
rect 60555 1525 60595 1565
rect 60905 1525 60945 1565
rect 61255 1525 61295 1565
rect 52505 1175 52545 1215
rect 52855 1175 52895 1215
rect 53205 1175 53245 1215
rect 53555 1175 53595 1215
rect 53905 1175 53945 1215
rect 59855 1175 59895 1215
rect 60205 1175 60245 1215
rect 60555 1175 60595 1215
rect 60905 1175 60945 1215
rect 61255 1175 61295 1215
rect 52505 825 52545 865
rect 52855 825 52895 865
rect 53205 825 53245 865
rect 53555 825 53595 865
rect 53905 825 53945 865
rect 59855 825 59895 865
rect 60205 825 60245 865
rect 60555 825 60595 865
rect 60905 825 60945 865
rect 61255 825 61295 865
rect 52505 475 52545 515
rect 52855 475 52895 515
rect 53205 475 53245 515
rect 53555 475 53595 515
rect 53905 475 53945 515
rect 59855 475 59895 515
rect 60205 475 60245 515
rect 60555 475 60595 515
rect 60905 475 60945 515
rect 61255 475 61295 515
rect 52505 125 52545 165
rect 52855 125 52895 165
rect 53205 125 53245 165
rect 53555 125 53595 165
rect 53905 125 53945 165
rect 54255 125 54295 165
rect 54605 125 54645 165
rect 54955 125 54995 165
rect 55305 125 55345 165
rect 55655 125 55695 165
rect 56005 125 56045 165
rect 56355 125 56395 165
rect 56705 125 56745 165
rect 57055 125 57095 165
rect 57405 125 57445 165
rect 57755 125 57795 165
rect 58105 125 58145 165
rect 58455 125 58495 165
rect 58805 125 58845 165
rect 59155 125 59195 165
rect 59505 125 59545 165
rect 59855 125 59895 165
rect 60205 125 60245 165
rect 60555 125 60595 165
rect 60905 125 60945 165
rect 61255 125 61295 165
rect 52505 -225 52545 -185
rect 52855 -225 52895 -185
rect 53205 -225 53245 -185
rect 53555 -225 53595 -185
rect 53905 -225 53945 -185
rect 54255 -225 54295 -185
rect 54605 -225 54645 -185
rect 54955 -225 54995 -185
rect 55305 -225 55345 -185
rect 55655 -225 55695 -185
rect 56005 -225 56045 -185
rect 56355 -225 56395 -185
rect 56705 -225 56745 -185
rect 57055 -225 57095 -185
rect 57405 -225 57445 -185
rect 57755 -225 57795 -185
rect 58105 -225 58145 -185
rect 58455 -225 58495 -185
rect 58805 -225 58845 -185
rect 59155 -225 59195 -185
rect 59505 -225 59545 -185
rect 59855 -225 59895 -185
rect 60205 -225 60245 -185
rect 60555 -225 60595 -185
rect 60905 -225 60945 -185
rect 61255 -225 61295 -185
<< metal4 >>
rect 52500 5765 53250 5770
rect 52500 5725 52505 5765
rect 52545 5725 52855 5765
rect 52895 5725 53205 5765
rect 53245 5725 53250 5765
rect 52500 5720 53250 5725
rect 53200 5420 53250 5720
rect 53550 5765 53600 5770
rect 53550 5725 53555 5765
rect 53595 5725 53600 5765
rect 53550 5420 53600 5725
rect 53900 5765 53950 5770
rect 53900 5725 53905 5765
rect 53945 5725 53950 5765
rect 53900 5420 53950 5725
rect 54250 5765 54300 5770
rect 54250 5725 54255 5765
rect 54295 5725 54300 5765
rect 54250 5420 54300 5725
rect 54600 5765 54650 5770
rect 54600 5725 54605 5765
rect 54645 5725 54650 5765
rect 54600 5420 54650 5725
rect 54950 5765 55000 5770
rect 54950 5725 54955 5765
rect 54995 5725 55000 5765
rect 54950 5420 55000 5725
rect 55300 5765 55350 5770
rect 55300 5725 55305 5765
rect 55345 5725 55350 5765
rect 55300 5420 55350 5725
rect 55650 5765 55700 5770
rect 55650 5725 55655 5765
rect 55695 5725 55700 5765
rect 55650 5420 55700 5725
rect 56000 5765 56050 5770
rect 56000 5725 56005 5765
rect 56045 5725 56050 5765
rect 56000 5420 56050 5725
rect 56350 5765 56400 5770
rect 56350 5725 56355 5765
rect 56395 5725 56400 5765
rect 56350 5420 56400 5725
rect 56700 5765 56750 5770
rect 56700 5725 56705 5765
rect 56745 5725 56750 5765
rect 56700 5420 56750 5725
rect 52500 5415 56750 5420
rect 52500 5375 52505 5415
rect 52545 5375 52855 5415
rect 52895 5375 53205 5415
rect 53245 5375 53555 5415
rect 53595 5375 53905 5415
rect 53945 5375 54255 5415
rect 54295 5375 54605 5415
rect 54645 5375 54955 5415
rect 54995 5375 55305 5415
rect 55345 5375 55655 5415
rect 55695 5375 56005 5415
rect 56045 5375 56355 5415
rect 56395 5375 56705 5415
rect 56745 5375 56750 5415
rect 52500 5370 56750 5375
rect 53200 5070 53250 5370
rect 52500 5065 53950 5070
rect 52500 5025 52505 5065
rect 52545 5025 52855 5065
rect 52895 5025 53205 5065
rect 53245 5025 53555 5065
rect 53595 5025 53905 5065
rect 53945 5025 53950 5065
rect 52500 5020 53950 5025
rect 54250 5065 54300 5370
rect 54250 5025 54255 5065
rect 54295 5025 54300 5065
rect 53200 4720 53250 5020
rect 52500 4715 53950 4720
rect 52500 4675 52505 4715
rect 52545 4675 52855 4715
rect 52895 4675 53205 4715
rect 53245 4675 53555 4715
rect 53595 4675 53905 4715
rect 53945 4675 53950 4715
rect 52500 4670 53950 4675
rect 54250 4715 54300 5025
rect 54250 4675 54255 4715
rect 54295 4675 54300 4715
rect 53200 4370 53250 4670
rect 52500 4365 53950 4370
rect 52500 4325 52505 4365
rect 52545 4325 52855 4365
rect 52895 4325 53205 4365
rect 53245 4325 53555 4365
rect 53595 4325 53905 4365
rect 53945 4325 53950 4365
rect 52500 4320 53950 4325
rect 54250 4365 54300 4675
rect 54250 4325 54255 4365
rect 54295 4325 54300 4365
rect 54250 4320 54300 4325
rect 54600 5065 54650 5370
rect 54600 5025 54605 5065
rect 54645 5025 54650 5065
rect 54600 4715 54650 5025
rect 54600 4675 54605 4715
rect 54645 4675 54650 4715
rect 54600 4365 54650 4675
rect 54600 4325 54605 4365
rect 54645 4325 54650 4365
rect 54600 4320 54650 4325
rect 54950 5065 55000 5370
rect 54950 5025 54955 5065
rect 54995 5025 55000 5065
rect 54950 4715 55000 5025
rect 54950 4675 54955 4715
rect 54995 4675 55000 4715
rect 54950 4365 55000 4675
rect 54950 4325 54955 4365
rect 54995 4325 55000 4365
rect 54950 4320 55000 4325
rect 55300 5065 55350 5370
rect 55300 5025 55305 5065
rect 55345 5025 55350 5065
rect 55300 4715 55350 5025
rect 55650 5055 55700 5370
rect 55650 5015 55655 5055
rect 55695 5015 55700 5055
rect 55650 5010 55700 5015
rect 56000 5055 56050 5370
rect 56000 5015 56005 5055
rect 56045 5015 56050 5055
rect 56000 5010 56050 5015
rect 56350 5055 56400 5370
rect 56350 5015 56355 5055
rect 56395 5015 56400 5055
rect 56350 5010 56400 5015
rect 56700 5055 56750 5370
rect 56700 5015 56705 5055
rect 56745 5015 56750 5055
rect 56700 5010 56750 5015
rect 57050 5765 57100 5770
rect 57050 5725 57055 5765
rect 57095 5725 57100 5765
rect 57050 5420 57100 5725
rect 57400 5765 57450 5770
rect 57400 5725 57405 5765
rect 57445 5725 57450 5765
rect 57400 5420 57450 5725
rect 57750 5765 57800 5770
rect 57750 5725 57755 5765
rect 57795 5725 57800 5765
rect 57750 5420 57800 5725
rect 58100 5765 58150 5770
rect 58100 5725 58105 5765
rect 58145 5725 58150 5765
rect 58100 5420 58150 5725
rect 58450 5765 58500 5770
rect 58450 5725 58455 5765
rect 58495 5725 58500 5765
rect 58450 5420 58500 5725
rect 58800 5765 58850 5770
rect 58800 5725 58805 5765
rect 58845 5725 58850 5765
rect 58800 5420 58850 5725
rect 59150 5765 59200 5770
rect 59150 5725 59155 5765
rect 59195 5725 59200 5765
rect 59150 5420 59200 5725
rect 59500 5765 59550 5770
rect 59500 5725 59505 5765
rect 59545 5725 59550 5765
rect 59500 5420 59550 5725
rect 59850 5765 59900 5770
rect 59850 5725 59855 5765
rect 59895 5725 59900 5765
rect 59850 5420 59900 5725
rect 60200 5765 60250 5770
rect 60200 5725 60205 5765
rect 60245 5725 60250 5765
rect 60200 5420 60250 5725
rect 60550 5765 61300 5770
rect 60550 5725 60555 5765
rect 60595 5725 60905 5765
rect 60945 5725 61255 5765
rect 61295 5725 61300 5765
rect 60550 5720 61300 5725
rect 60550 5420 60600 5720
rect 57050 5415 61300 5420
rect 57050 5375 57055 5415
rect 57095 5375 57405 5415
rect 57445 5375 57755 5415
rect 57795 5375 58105 5415
rect 58145 5375 58455 5415
rect 58495 5375 58805 5415
rect 58845 5375 59155 5415
rect 59195 5375 59505 5415
rect 59545 5375 59855 5415
rect 59895 5375 60205 5415
rect 60245 5375 60555 5415
rect 60595 5375 60905 5415
rect 60945 5375 61255 5415
rect 61295 5375 61300 5415
rect 57050 5370 61300 5375
rect 57050 5055 57100 5370
rect 57050 5015 57055 5055
rect 57095 5015 57100 5055
rect 57050 5010 57100 5015
rect 57400 5055 57450 5370
rect 57400 5015 57405 5055
rect 57445 5015 57450 5055
rect 57400 5010 57450 5015
rect 57750 5055 57800 5370
rect 57750 5015 57755 5055
rect 57795 5015 57800 5055
rect 57750 5010 57800 5015
rect 58100 5055 58150 5370
rect 58100 5015 58105 5055
rect 58145 5015 58150 5055
rect 58100 5010 58150 5015
rect 58450 5065 58500 5370
rect 58450 5025 58455 5065
rect 58495 5025 58500 5065
rect 55300 4675 55305 4715
rect 55345 4675 55350 4715
rect 55300 4365 55350 4675
rect 55300 4325 55305 4365
rect 55345 4325 55350 4365
rect 55300 4320 55350 4325
rect 58450 4715 58500 5025
rect 58450 4675 58455 4715
rect 58495 4675 58500 4715
rect 58450 4365 58500 4675
rect 58450 4325 58455 4365
rect 58495 4325 58500 4365
rect 58450 4320 58500 4325
rect 58800 5065 58850 5370
rect 58800 5025 58805 5065
rect 58845 5025 58850 5065
rect 58800 4715 58850 5025
rect 58800 4675 58805 4715
rect 58845 4675 58850 4715
rect 58800 4365 58850 4675
rect 58800 4325 58805 4365
rect 58845 4325 58850 4365
rect 58800 4320 58850 4325
rect 59150 5065 59200 5370
rect 59150 5025 59155 5065
rect 59195 5025 59200 5065
rect 59150 4715 59200 5025
rect 59150 4675 59155 4715
rect 59195 4675 59200 4715
rect 59150 4365 59200 4675
rect 59150 4325 59155 4365
rect 59195 4325 59200 4365
rect 59150 4320 59200 4325
rect 59500 5065 59550 5370
rect 60550 5070 60600 5370
rect 59500 5025 59505 5065
rect 59545 5025 59550 5065
rect 59500 4715 59550 5025
rect 59850 5065 61300 5070
rect 59850 5025 59855 5065
rect 59895 5025 60205 5065
rect 60245 5025 60555 5065
rect 60595 5025 60905 5065
rect 60945 5025 61255 5065
rect 61295 5025 61300 5065
rect 59850 5020 61300 5025
rect 60550 4720 60600 5020
rect 59500 4675 59505 4715
rect 59545 4675 59550 4715
rect 59500 4365 59550 4675
rect 59850 4715 61300 4720
rect 59850 4675 59855 4715
rect 59895 4675 60205 4715
rect 60245 4675 60555 4715
rect 60595 4675 60905 4715
rect 60945 4675 61255 4715
rect 61295 4675 61300 4715
rect 59850 4670 61300 4675
rect 60550 4370 60600 4670
rect 59500 4325 59505 4365
rect 59545 4325 59550 4365
rect 59500 4320 59550 4325
rect 59850 4365 61300 4370
rect 59850 4325 59855 4365
rect 59895 4325 60205 4365
rect 60245 4325 60555 4365
rect 60595 4325 60905 4365
rect 60945 4325 61255 4365
rect 61295 4325 61300 4365
rect 59850 4320 61300 4325
rect 53200 4020 53250 4320
rect 60550 4020 60600 4320
rect 52500 4015 53950 4020
rect 52500 3975 52505 4015
rect 52545 3975 52855 4015
rect 52895 3975 53205 4015
rect 53245 3975 53555 4015
rect 53595 3975 53905 4015
rect 53945 3975 53950 4015
rect 52500 3970 53950 3975
rect 59850 4015 61300 4020
rect 59850 3975 59855 4015
rect 59895 3975 60205 4015
rect 60245 3975 60555 4015
rect 60595 3975 60905 4015
rect 60945 3975 61255 4015
rect 61295 3975 61300 4015
rect 59850 3970 61300 3975
rect 53200 3670 53250 3970
rect 60550 3670 60600 3970
rect 52500 3665 53950 3670
rect 52500 3625 52505 3665
rect 52545 3625 52855 3665
rect 52895 3625 53205 3665
rect 53245 3625 53555 3665
rect 53595 3625 53905 3665
rect 53945 3625 53950 3665
rect 52500 3620 53950 3625
rect 59850 3665 61300 3670
rect 59850 3625 59855 3665
rect 59895 3625 60205 3665
rect 60245 3625 60555 3665
rect 60595 3625 60905 3665
rect 60945 3625 61255 3665
rect 61295 3625 61300 3665
rect 59850 3620 61300 3625
rect 53200 3320 53250 3620
rect 60550 3320 60600 3620
rect 52500 3315 53950 3320
rect 52500 3275 52505 3315
rect 52545 3275 52855 3315
rect 52895 3275 53205 3315
rect 53245 3275 53555 3315
rect 53595 3275 53905 3315
rect 53945 3275 53950 3315
rect 52500 3270 53950 3275
rect 59850 3315 61300 3320
rect 59850 3275 59855 3315
rect 59895 3275 60205 3315
rect 60245 3275 60555 3315
rect 60595 3275 60905 3315
rect 60945 3275 61255 3315
rect 61295 3275 61300 3315
rect 59850 3270 61300 3275
rect 53200 2970 53250 3270
rect 60550 2970 60600 3270
rect 52500 2965 53950 2970
rect 52500 2925 52505 2965
rect 52545 2925 52855 2965
rect 52895 2925 53205 2965
rect 53245 2925 53555 2965
rect 53595 2925 53905 2965
rect 53945 2925 53950 2965
rect 52500 2920 53950 2925
rect 59850 2965 61300 2970
rect 59850 2925 59855 2965
rect 59895 2925 60205 2965
rect 60245 2925 60555 2965
rect 60595 2925 60905 2965
rect 60945 2925 61255 2965
rect 61295 2925 61300 2965
rect 59850 2920 61300 2925
rect 53200 2620 53250 2920
rect 60550 2620 60600 2920
rect 52500 2615 53950 2620
rect 52500 2575 52505 2615
rect 52545 2575 52855 2615
rect 52895 2575 53205 2615
rect 53245 2575 53555 2615
rect 53595 2575 53905 2615
rect 53945 2575 53950 2615
rect 52500 2570 53950 2575
rect 59850 2615 61300 2620
rect 59850 2575 59855 2615
rect 59895 2575 60205 2615
rect 60245 2575 60555 2615
rect 60595 2575 60905 2615
rect 60945 2575 61255 2615
rect 61295 2575 61300 2615
rect 59850 2570 61300 2575
rect 53200 2270 53250 2570
rect 60550 2270 60600 2570
rect 52500 2265 53950 2270
rect 52500 2225 52505 2265
rect 52545 2225 52855 2265
rect 52895 2225 53205 2265
rect 53245 2225 53555 2265
rect 53595 2225 53905 2265
rect 53945 2225 53950 2265
rect 52500 2220 53950 2225
rect 59850 2265 61300 2270
rect 59850 2225 59855 2265
rect 59895 2225 60205 2265
rect 60245 2225 60555 2265
rect 60595 2225 60905 2265
rect 60945 2225 61255 2265
rect 61295 2225 61300 2265
rect 59850 2220 61300 2225
rect 53200 1920 53250 2220
rect 60550 1920 60600 2220
rect 52500 1915 54340 1920
rect 52500 1875 52505 1915
rect 52545 1875 52855 1915
rect 52895 1875 53205 1915
rect 53245 1875 53555 1915
rect 53595 1875 53905 1915
rect 53945 1875 54295 1915
rect 54335 1875 54340 1915
rect 52500 1870 54340 1875
rect 59460 1915 61300 1920
rect 59460 1875 59465 1915
rect 59505 1875 59855 1915
rect 59895 1875 60205 1915
rect 60245 1875 60555 1915
rect 60595 1875 60905 1915
rect 60945 1875 61255 1915
rect 61295 1875 61300 1915
rect 59460 1870 61300 1875
rect 53200 1570 53250 1870
rect 60550 1570 60600 1870
rect 52500 1565 53950 1570
rect 52500 1525 52505 1565
rect 52545 1525 52855 1565
rect 52895 1525 53205 1565
rect 53245 1525 53555 1565
rect 53595 1525 53905 1565
rect 53945 1525 53950 1565
rect 52500 1520 53950 1525
rect 59850 1565 61300 1570
rect 59850 1525 59855 1565
rect 59895 1525 60205 1565
rect 60245 1525 60555 1565
rect 60595 1525 60905 1565
rect 60945 1525 61255 1565
rect 61295 1525 61300 1565
rect 59850 1520 61300 1525
rect 53200 1220 53250 1520
rect 60550 1220 60600 1520
rect 52500 1215 53950 1220
rect 52500 1175 52505 1215
rect 52545 1175 52855 1215
rect 52895 1175 53205 1215
rect 53245 1175 53555 1215
rect 53595 1175 53905 1215
rect 53945 1175 53950 1215
rect 52500 1170 53950 1175
rect 59850 1215 61300 1220
rect 59850 1175 59855 1215
rect 59895 1175 60205 1215
rect 60245 1175 60555 1215
rect 60595 1175 60905 1215
rect 60945 1175 61255 1215
rect 61295 1175 61300 1215
rect 59850 1170 61300 1175
rect 53200 870 53250 1170
rect 60550 870 60600 1170
rect 52500 865 53950 870
rect 52500 825 52505 865
rect 52545 825 52855 865
rect 52895 825 53205 865
rect 53245 825 53555 865
rect 53595 825 53905 865
rect 53945 825 53950 865
rect 52500 820 53950 825
rect 59850 865 61300 870
rect 59850 825 59855 865
rect 59895 825 60205 865
rect 60245 825 60555 865
rect 60595 825 60905 865
rect 60945 825 61255 865
rect 61295 825 61300 865
rect 59850 820 61300 825
rect 53200 520 53250 820
rect 60550 520 60600 820
rect 52500 515 53950 520
rect 52500 475 52505 515
rect 52545 475 52855 515
rect 52895 475 53205 515
rect 53245 475 53555 515
rect 53595 475 53905 515
rect 53945 475 53950 515
rect 52500 470 53950 475
rect 59850 515 61300 520
rect 59850 475 59855 515
rect 59895 475 60205 515
rect 60245 475 60555 515
rect 60595 475 60905 515
rect 60945 475 61255 515
rect 61295 475 61300 515
rect 59850 470 61300 475
rect 53200 170 53250 470
rect 60550 170 60600 470
rect 52500 165 56750 170
rect 52500 125 52505 165
rect 52545 125 52855 165
rect 52895 125 53205 165
rect 53245 125 53555 165
rect 53595 125 53905 165
rect 53945 125 54255 165
rect 54295 125 54605 165
rect 54645 125 54955 165
rect 54995 125 55305 165
rect 55345 125 55655 165
rect 55695 125 56005 165
rect 56045 125 56355 165
rect 56395 125 56705 165
rect 56745 125 56750 165
rect 52500 120 56750 125
rect 53200 -180 53250 120
rect 52500 -185 53250 -180
rect 52500 -225 52505 -185
rect 52545 -225 52855 -185
rect 52895 -225 53205 -185
rect 53245 -225 53250 -185
rect 52500 -230 53250 -225
rect 53550 -185 53600 120
rect 53550 -225 53555 -185
rect 53595 -225 53600 -185
rect 53550 -230 53600 -225
rect 53900 -185 53950 120
rect 53900 -225 53905 -185
rect 53945 -225 53950 -185
rect 53900 -230 53950 -225
rect 54250 -185 54300 120
rect 54250 -225 54255 -185
rect 54295 -225 54300 -185
rect 54250 -230 54300 -225
rect 54600 -185 54650 120
rect 54600 -225 54605 -185
rect 54645 -225 54650 -185
rect 54600 -230 54650 -225
rect 54950 -185 55000 120
rect 54950 -225 54955 -185
rect 54995 -225 55000 -185
rect 54950 -230 55000 -225
rect 55300 -185 55350 120
rect 55300 -225 55305 -185
rect 55345 -225 55350 -185
rect 55300 -230 55350 -225
rect 55650 -185 55700 120
rect 55650 -225 55655 -185
rect 55695 -225 55700 -185
rect 55650 -230 55700 -225
rect 56000 -185 56050 120
rect 56000 -225 56005 -185
rect 56045 -225 56050 -185
rect 56000 -230 56050 -225
rect 56350 -185 56400 120
rect 56350 -225 56355 -185
rect 56395 -225 56400 -185
rect 56350 -230 56400 -225
rect 56700 -185 56750 120
rect 56700 -225 56705 -185
rect 56745 -225 56750 -185
rect 56700 -230 56750 -225
rect 57050 165 61300 170
rect 57050 125 57055 165
rect 57095 125 57405 165
rect 57445 125 57755 165
rect 57795 125 58105 165
rect 58145 125 58455 165
rect 58495 125 58805 165
rect 58845 125 59155 165
rect 59195 125 59505 165
rect 59545 125 59855 165
rect 59895 125 60205 165
rect 60245 125 60555 165
rect 60595 125 60905 165
rect 60945 125 61255 165
rect 61295 125 61300 165
rect 57050 120 61300 125
rect 57050 -185 57100 120
rect 57050 -225 57055 -185
rect 57095 -225 57100 -185
rect 57050 -230 57100 -225
rect 57400 -185 57450 120
rect 57400 -225 57405 -185
rect 57445 -225 57450 -185
rect 57400 -230 57450 -225
rect 57750 -185 57800 120
rect 57750 -225 57755 -185
rect 57795 -225 57800 -185
rect 57750 -230 57800 -225
rect 58100 -185 58150 120
rect 58100 -225 58105 -185
rect 58145 -225 58150 -185
rect 58100 -230 58150 -225
rect 58450 -185 58500 120
rect 58450 -225 58455 -185
rect 58495 -225 58500 -185
rect 58450 -230 58500 -225
rect 58800 -185 58850 120
rect 58800 -225 58805 -185
rect 58845 -225 58850 -185
rect 58800 -230 58850 -225
rect 59150 -185 59200 120
rect 59150 -225 59155 -185
rect 59195 -225 59200 -185
rect 59150 -230 59200 -225
rect 59500 -185 59550 120
rect 59500 -225 59505 -185
rect 59545 -225 59550 -185
rect 59500 -230 59550 -225
rect 59850 -185 59900 120
rect 59850 -225 59855 -185
rect 59895 -225 59900 -185
rect 59850 -230 59900 -225
rect 60200 -185 60250 120
rect 60200 -225 60205 -185
rect 60245 -225 60250 -185
rect 60200 -230 60250 -225
rect 60550 -180 60600 120
rect 60550 -185 61300 -180
rect 60550 -225 60555 -185
rect 60595 -225 60905 -185
rect 60945 -225 61255 -185
rect 61295 -225 61300 -185
rect 60550 -230 61300 -225
<< labels >>
flabel metal3 59195 3460 59195 3460 3 FreeSans 240 0 80 0 cap_res_X
flabel metal3 54605 3460 54605 3460 7 FreeSans 240 0 -80 0 cap_res_Y
flabel metal1 55920 4030 55920 4030 7 FreeSans 240 0 -80 0 VD4
flabel metal1 57880 4015 57880 4015 3 FreeSans 240 0 80 0 VD3
flabel metal1 56910 1290 56910 1290 3 FreeSans 200 0 80 0 V_p_mir
flabel metal1 56370 1880 56370 1880 7 FreeSans 240 0 -80 0 VD2
flabel metal1 57430 1875 57430 1875 3 FreeSans 240 0 80 0 VD1
flabel metal1 56950 1825 56950 1825 7 FreeSans 240 0 -80 0 V_tail_gate
flabel metal1 55850 2275 55850 2275 1 FreeSans 200 0 0 80 Vb1
port 6 n
flabel metal1 56345 2575 56345 2575 3 FreeSans 240 0 80 0 Y
flabel metal1 57455 2575 57455 2575 7 FreeSans 240 0 -80 0 X
flabel metal2 57720 1300 57720 1300 5 FreeSans 200 0 0 -80 V_b_2nd_stage
flabel metal2 57235 2675 57235 2675 7 FreeSans 200 0 -80 0 err_amp_out
flabel metal2 57605 2830 57605 2830 3 FreeSans 200 0 80 0 err_amp_mir
flabel metal2 56900 3015 56900 3015 1 FreeSans 240 0 0 80 V_tot
flabel metal1 57240 3065 57240 3065 3 FreeSans 200 0 80 0 V_err_p
flabel metal1 54315 1220 54315 1220 5 FreeSans 240 0 0 -80 VOUT+
port 10 s
flabel metal2 57365 4810 57365 4810 1 FreeSans 240 0 0 80 Vb2_Vb3
flabel metal2 56455 4810 56455 4810 1 FreeSans 240 0 0 80 Vb2_2
flabel metal2 57770 1770 57770 1770 3 FreeSans 240 0 80 0 VIN-
flabel metal2 56030 1770 56030 1770 7 FreeSans 240 0 -80 0 VIN+
flabel metal1 57220 1285 57220 1285 3 FreeSans 240 0 80 0 V_source
flabel metal1 56835 3065 56835 3065 7 FreeSans 200 0 -80 0 V_err_gate
port 13 w
flabel metal2 55960 2775 55960 2775 7 FreeSans 200 0 -80 0 V_err_amp_ref
port 12 w
flabel metal1 59020 2155 59020 2155 1 FreeSans 240 0 0 80 V_CMFB_S1
port 2 n
flabel metal1 58975 1950 58975 1950 1 FreeSans 240 0 0 80 V_CMFB_S2
port 7 n
flabel metal1 54780 2155 54780 2155 1 FreeSans 240 0 0 80 V_CMFB_S3
port 3 n
flabel metal1 54825 1950 54825 1950 1 FreeSans 240 0 0 80 V_CMFB_S4
port 8 n
flabel metal1 59485 1220 59485 1220 5 FreeSans 240 0 0 -80 VOUT-
port 9 s
flabel metal2 57000 3535 57000 3535 5 FreeSans 200 0 0 -80 Vb3
port 4 s
flabel metal1 56855 3570 56855 3570 5 FreeSans 200 0 0 -80 Vb2
port 5 s
<< end >>
