magic
tech sky130A
magscale 1 2
timestamp 1755645661
<< nwell >>
rect 112050 9020 112730 9800
rect 112990 9020 113670 9460
rect 113930 9020 114610 9800
rect 114870 9020 115550 9800
rect 109060 7020 110820 7800
rect 111890 7020 113650 7800
rect 113950 7020 115710 7800
rect 116780 7020 118540 7800
rect 109120 5070 110760 6350
rect 112900 5800 114700 6380
rect 116840 5070 118480 6350
rect 117830 5060 118110 5070
rect 109120 3320 110760 3800
rect 116840 3320 118480 3800
<< nmos >>
rect 113620 4630 113650 5130
rect 113730 4630 113760 5130
rect 113840 4630 113870 5130
rect 113950 4630 113980 5130
rect 112140 3510 112170 3810
rect 112250 3510 112280 3810
rect 112360 3510 112390 3810
rect 112470 3510 112500 3810
rect 112580 3510 112610 3810
rect 112690 3510 112720 3810
rect 112800 3510 112830 3810
rect 112910 3510 112940 3810
rect 113020 3510 113050 3810
rect 113130 3510 113160 3810
rect 113240 3510 113270 3810
rect 113350 3510 113380 3810
rect 114220 3510 114250 3810
rect 114330 3510 114360 3810
rect 114440 3510 114470 3810
rect 114550 3510 114580 3810
rect 114660 3510 114690 3810
rect 114770 3510 114800 3810
rect 114880 3510 114910 3810
rect 114990 3510 115020 3810
rect 115100 3510 115130 3810
rect 115210 3510 115240 3810
rect 115320 3510 115350 3810
rect 115430 3510 115460 3810
rect 109320 2280 109350 2880
rect 109430 2280 109460 2880
rect 109540 2280 109570 2880
rect 109650 2280 109680 2880
rect 109760 2280 109790 2880
rect 109870 2280 109900 2880
rect 109980 2280 110010 2880
rect 110090 2280 110120 2880
rect 110200 2280 110230 2880
rect 110310 2280 110340 2880
rect 110420 2280 110450 2880
rect 110530 2280 110560 2880
rect 112140 2140 112170 2440
rect 112250 2140 112280 2440
rect 112360 2140 112390 2440
rect 112470 2140 112500 2440
rect 112580 2140 112610 2440
rect 112690 2140 112720 2440
rect 112800 2140 112830 2440
rect 112910 2140 112940 2440
rect 113020 2140 113050 2440
rect 113130 2140 113160 2440
rect 113240 2140 113270 2440
rect 113350 2140 113380 2440
rect 113620 2140 113650 2440
rect 113730 2140 113760 2440
rect 113840 2140 113870 2440
rect 113950 2140 113980 2440
rect 114220 2140 114250 2440
rect 114330 2140 114360 2440
rect 114440 2140 114470 2440
rect 114550 2140 114580 2440
rect 114660 2140 114690 2440
rect 114770 2140 114800 2440
rect 114880 2140 114910 2440
rect 114990 2140 115020 2440
rect 115100 2140 115130 2440
rect 115210 2140 115240 2440
rect 115320 2140 115350 2440
rect 115430 2140 115460 2440
rect 117040 2280 117070 2880
rect 117150 2280 117180 2880
rect 117260 2280 117290 2880
rect 117370 2280 117400 2880
rect 117480 2280 117510 2880
rect 117590 2280 117620 2880
rect 117700 2280 117730 2880
rect 117810 2280 117840 2880
rect 117920 2280 117950 2880
rect 118030 2280 118060 2880
rect 118140 2280 118170 2880
rect 118250 2280 118280 2880
rect 109380 -720 109500 680
rect 109580 -720 109700 680
rect 109780 -720 109900 680
rect 109980 -720 110100 680
rect 110180 -720 110300 680
rect 110380 -720 110500 680
rect 112520 410 112550 910
rect 112630 410 112660 910
rect 112740 410 112770 910
rect 112850 410 112880 910
rect 112960 410 112990 910
rect 113070 410 113100 910
rect 113180 410 113210 910
rect 113290 410 113320 910
rect 113400 410 113430 910
rect 113510 410 113540 910
rect 113620 410 113650 910
rect 113730 410 113760 910
rect 113840 410 113870 910
rect 113950 410 113980 910
rect 114060 410 114090 910
rect 114170 410 114200 910
rect 114280 410 114310 910
rect 114390 410 114420 910
rect 114500 410 114530 910
rect 114610 410 114640 910
rect 114720 410 114750 910
rect 114830 410 114860 910
rect 114940 410 114970 910
rect 112940 -900 112970 -600
rect 113050 -900 113080 -600
rect 113160 -900 113190 -600
rect 113270 -900 113300 -600
rect 113380 -900 113410 -600
rect 113490 -900 113520 -600
rect 113820 -900 114420 -600
rect 117100 -720 117220 680
rect 117300 -720 117420 680
rect 117500 -720 117620 680
rect 117700 -720 117820 680
rect 117900 -720 118020 680
rect 118100 -720 118220 680
<< pmos >>
rect 112250 9060 112290 9760
rect 112370 9060 112410 9760
rect 112490 9060 112530 9760
rect 113190 9060 113230 9420
rect 113310 9060 113350 9420
rect 113430 9060 113470 9420
rect 114130 9060 114170 9760
rect 114250 9060 114290 9760
rect 114370 9060 114410 9760
rect 115070 9060 115110 9760
rect 115190 9060 115230 9760
rect 115310 9060 115350 9760
rect 109260 7060 109300 7760
rect 109380 7060 109420 7760
rect 109500 7060 109540 7760
rect 109620 7060 109660 7760
rect 109740 7060 109780 7760
rect 109860 7060 109900 7760
rect 109980 7060 110020 7760
rect 110100 7060 110140 7760
rect 110220 7060 110260 7760
rect 110340 7060 110380 7760
rect 110460 7060 110500 7760
rect 110580 7060 110620 7760
rect 112090 7060 112130 7760
rect 112210 7060 112250 7760
rect 112330 7060 112370 7760
rect 112450 7060 112490 7760
rect 112570 7060 112610 7760
rect 112690 7060 112730 7760
rect 112810 7060 112850 7760
rect 112930 7060 112970 7760
rect 113050 7060 113090 7760
rect 113170 7060 113210 7760
rect 113290 7060 113330 7760
rect 113410 7060 113450 7760
rect 114150 7060 114190 7760
rect 114270 7060 114310 7760
rect 114390 7060 114430 7760
rect 114510 7060 114550 7760
rect 114630 7060 114670 7760
rect 114750 7060 114790 7760
rect 114870 7060 114910 7760
rect 114990 7060 115030 7760
rect 115110 7060 115150 7760
rect 115230 7060 115270 7760
rect 115350 7060 115390 7760
rect 115470 7060 115510 7760
rect 116980 7060 117020 7760
rect 117100 7060 117140 7760
rect 117220 7060 117260 7760
rect 117340 7060 117380 7760
rect 117460 7060 117500 7760
rect 117580 7060 117620 7760
rect 117700 7060 117740 7760
rect 117820 7060 117860 7760
rect 117940 7060 117980 7760
rect 118060 7060 118100 7760
rect 118180 7060 118220 7760
rect 118300 7060 118340 7760
rect 109320 5110 109350 6310
rect 109430 5110 109460 6310
rect 109540 5110 109570 6310
rect 109650 5110 109680 6310
rect 109760 5110 109790 6310
rect 109870 5110 109900 6310
rect 109980 5110 110010 6310
rect 110090 5110 110120 6310
rect 110200 5110 110230 6310
rect 110310 5110 110340 6310
rect 110420 5110 110450 6310
rect 110530 5110 110560 6310
rect 113100 5840 113130 6340
rect 113210 5840 113240 6340
rect 113320 5840 113350 6340
rect 113430 5840 113460 6340
rect 113540 5840 113570 6340
rect 113650 5840 113680 6340
rect 113920 5840 113950 6340
rect 114030 5840 114060 6340
rect 114140 5840 114170 6340
rect 114250 5840 114280 6340
rect 114360 5840 114390 6340
rect 114470 5840 114500 6340
rect 117040 5110 117070 6310
rect 117150 5110 117180 6310
rect 117260 5110 117290 6310
rect 117370 5110 117400 6310
rect 117480 5110 117510 6310
rect 117590 5110 117620 6310
rect 117700 5110 117730 6310
rect 117810 5110 117840 6310
rect 117920 5110 117950 6310
rect 118030 5110 118060 6310
rect 118140 5110 118170 6310
rect 118250 5110 118280 6310
rect 109320 3360 109350 3760
rect 109430 3360 109460 3760
rect 109540 3360 109570 3760
rect 109650 3360 109680 3760
rect 109760 3360 109790 3760
rect 109870 3360 109900 3760
rect 109980 3360 110010 3760
rect 110090 3360 110120 3760
rect 110200 3360 110230 3760
rect 110310 3360 110340 3760
rect 110420 3360 110450 3760
rect 110530 3360 110560 3760
rect 117040 3360 117070 3760
rect 117150 3360 117180 3760
rect 117260 3360 117290 3760
rect 117370 3360 117400 3760
rect 117480 3360 117510 3760
rect 117590 3360 117620 3760
rect 117700 3360 117730 3760
rect 117810 3360 117840 3760
rect 117920 3360 117950 3760
rect 118030 3360 118060 3760
rect 118140 3360 118170 3760
rect 118250 3360 118280 3760
<< ndiff >>
rect 113540 5100 113620 5130
rect 113540 4660 113560 5100
rect 113600 4660 113620 5100
rect 113540 4630 113620 4660
rect 113650 5100 113730 5130
rect 113650 4660 113670 5100
rect 113710 4660 113730 5100
rect 113650 4630 113730 4660
rect 113760 5100 113840 5130
rect 113760 4660 113780 5100
rect 113820 4660 113840 5100
rect 113760 4630 113840 4660
rect 113870 5100 113950 5130
rect 113870 4660 113890 5100
rect 113930 4660 113950 5100
rect 113870 4630 113950 4660
rect 113980 5100 114060 5130
rect 113980 4660 114000 5100
rect 114040 4660 114060 5100
rect 113980 4630 114060 4660
rect 112060 3780 112140 3810
rect 112060 3540 112080 3780
rect 112120 3540 112140 3780
rect 112060 3510 112140 3540
rect 112170 3780 112250 3810
rect 112170 3540 112190 3780
rect 112230 3540 112250 3780
rect 112170 3510 112250 3540
rect 112280 3780 112360 3810
rect 112280 3540 112300 3780
rect 112340 3540 112360 3780
rect 112280 3510 112360 3540
rect 112390 3780 112470 3810
rect 112390 3540 112410 3780
rect 112450 3540 112470 3780
rect 112390 3510 112470 3540
rect 112500 3780 112580 3810
rect 112500 3540 112520 3780
rect 112560 3540 112580 3780
rect 112500 3510 112580 3540
rect 112610 3780 112690 3810
rect 112610 3540 112630 3780
rect 112670 3540 112690 3780
rect 112610 3510 112690 3540
rect 112720 3780 112800 3810
rect 112720 3540 112740 3780
rect 112780 3540 112800 3780
rect 112720 3510 112800 3540
rect 112830 3780 112910 3810
rect 112830 3540 112850 3780
rect 112890 3540 112910 3780
rect 112830 3510 112910 3540
rect 112940 3780 113020 3810
rect 112940 3540 112960 3780
rect 113000 3540 113020 3780
rect 112940 3510 113020 3540
rect 113050 3780 113130 3810
rect 113050 3540 113070 3780
rect 113110 3540 113130 3780
rect 113050 3510 113130 3540
rect 113160 3780 113240 3810
rect 113160 3540 113180 3780
rect 113220 3540 113240 3780
rect 113160 3510 113240 3540
rect 113270 3780 113350 3810
rect 113270 3540 113290 3780
rect 113330 3540 113350 3780
rect 113270 3510 113350 3540
rect 113380 3780 113460 3810
rect 113380 3540 113400 3780
rect 113440 3540 113460 3780
rect 113380 3510 113460 3540
rect 114140 3780 114220 3810
rect 114140 3540 114160 3780
rect 114200 3540 114220 3780
rect 114140 3510 114220 3540
rect 114250 3780 114330 3810
rect 114250 3540 114270 3780
rect 114310 3540 114330 3780
rect 114250 3510 114330 3540
rect 114360 3780 114440 3810
rect 114360 3540 114380 3780
rect 114420 3540 114440 3780
rect 114360 3510 114440 3540
rect 114470 3780 114550 3810
rect 114470 3540 114490 3780
rect 114530 3540 114550 3780
rect 114470 3510 114550 3540
rect 114580 3780 114660 3810
rect 114580 3540 114600 3780
rect 114640 3540 114660 3780
rect 114580 3510 114660 3540
rect 114690 3780 114770 3810
rect 114690 3540 114710 3780
rect 114750 3540 114770 3780
rect 114690 3510 114770 3540
rect 114800 3780 114880 3810
rect 114800 3540 114820 3780
rect 114860 3540 114880 3780
rect 114800 3510 114880 3540
rect 114910 3780 114990 3810
rect 114910 3540 114930 3780
rect 114970 3540 114990 3780
rect 114910 3510 114990 3540
rect 115020 3780 115100 3810
rect 115020 3540 115040 3780
rect 115080 3540 115100 3780
rect 115020 3510 115100 3540
rect 115130 3780 115210 3810
rect 115130 3540 115150 3780
rect 115190 3540 115210 3780
rect 115130 3510 115210 3540
rect 115240 3780 115320 3810
rect 115240 3540 115260 3780
rect 115300 3540 115320 3780
rect 115240 3510 115320 3540
rect 115350 3780 115430 3810
rect 115350 3540 115370 3780
rect 115410 3540 115430 3780
rect 115350 3510 115430 3540
rect 115460 3780 115540 3810
rect 115460 3540 115480 3780
rect 115520 3540 115540 3780
rect 115460 3510 115540 3540
rect 109240 2850 109320 2880
rect 109240 2310 109260 2850
rect 109300 2310 109320 2850
rect 109240 2280 109320 2310
rect 109350 2850 109430 2880
rect 109350 2310 109370 2850
rect 109410 2310 109430 2850
rect 109350 2280 109430 2310
rect 109460 2850 109540 2880
rect 109460 2310 109480 2850
rect 109520 2310 109540 2850
rect 109460 2280 109540 2310
rect 109570 2850 109650 2880
rect 109570 2310 109590 2850
rect 109630 2310 109650 2850
rect 109570 2280 109650 2310
rect 109680 2850 109760 2880
rect 109680 2310 109700 2850
rect 109740 2310 109760 2850
rect 109680 2280 109760 2310
rect 109790 2850 109870 2880
rect 109790 2310 109810 2850
rect 109850 2310 109870 2850
rect 109790 2280 109870 2310
rect 109900 2850 109980 2880
rect 109900 2310 109920 2850
rect 109960 2310 109980 2850
rect 109900 2280 109980 2310
rect 110010 2850 110090 2880
rect 110010 2310 110030 2850
rect 110070 2310 110090 2850
rect 110010 2280 110090 2310
rect 110120 2850 110200 2880
rect 110120 2310 110140 2850
rect 110180 2310 110200 2850
rect 110120 2280 110200 2310
rect 110230 2850 110310 2880
rect 110230 2310 110250 2850
rect 110290 2310 110310 2850
rect 110230 2280 110310 2310
rect 110340 2850 110420 2880
rect 110340 2310 110360 2850
rect 110400 2310 110420 2850
rect 110340 2280 110420 2310
rect 110450 2850 110530 2880
rect 110450 2310 110470 2850
rect 110510 2310 110530 2850
rect 110450 2280 110530 2310
rect 110560 2850 110640 2880
rect 110560 2310 110580 2850
rect 110620 2310 110640 2850
rect 116960 2850 117040 2880
rect 110560 2280 110640 2310
rect 112060 2410 112140 2440
rect 112060 2170 112080 2410
rect 112120 2170 112140 2410
rect 112060 2140 112140 2170
rect 112170 2410 112250 2440
rect 112170 2170 112190 2410
rect 112230 2170 112250 2410
rect 112170 2140 112250 2170
rect 112280 2410 112360 2440
rect 112280 2170 112300 2410
rect 112340 2170 112360 2410
rect 112280 2140 112360 2170
rect 112390 2410 112470 2440
rect 112390 2170 112410 2410
rect 112450 2170 112470 2410
rect 112390 2140 112470 2170
rect 112500 2410 112580 2440
rect 112500 2170 112520 2410
rect 112560 2170 112580 2410
rect 112500 2140 112580 2170
rect 112610 2410 112690 2440
rect 112610 2170 112630 2410
rect 112670 2170 112690 2410
rect 112610 2140 112690 2170
rect 112720 2410 112800 2440
rect 112720 2170 112740 2410
rect 112780 2170 112800 2410
rect 112720 2140 112800 2170
rect 112830 2410 112910 2440
rect 112830 2170 112850 2410
rect 112890 2170 112910 2410
rect 112830 2140 112910 2170
rect 112940 2410 113020 2440
rect 112940 2170 112960 2410
rect 113000 2170 113020 2410
rect 112940 2140 113020 2170
rect 113050 2410 113130 2440
rect 113050 2170 113070 2410
rect 113110 2170 113130 2410
rect 113050 2140 113130 2170
rect 113160 2410 113240 2440
rect 113160 2170 113180 2410
rect 113220 2170 113240 2410
rect 113160 2140 113240 2170
rect 113270 2410 113350 2440
rect 113270 2170 113290 2410
rect 113330 2170 113350 2410
rect 113270 2140 113350 2170
rect 113380 2410 113460 2440
rect 113540 2410 113620 2440
rect 113380 2170 113400 2410
rect 113440 2170 113460 2410
rect 113540 2170 113560 2410
rect 113600 2170 113620 2410
rect 113380 2140 113460 2170
rect 113540 2140 113620 2170
rect 113650 2410 113730 2440
rect 113650 2170 113670 2410
rect 113710 2170 113730 2410
rect 113650 2140 113730 2170
rect 113760 2410 113840 2440
rect 113760 2170 113780 2410
rect 113820 2170 113840 2410
rect 113760 2140 113840 2170
rect 113870 2410 113950 2440
rect 113870 2170 113890 2410
rect 113930 2170 113950 2410
rect 113870 2140 113950 2170
rect 113980 2410 114060 2440
rect 114140 2410 114220 2440
rect 113980 2170 114000 2410
rect 114040 2170 114060 2410
rect 114140 2170 114160 2410
rect 114200 2170 114220 2410
rect 113980 2140 114060 2170
rect 114140 2140 114220 2170
rect 114250 2410 114330 2440
rect 114250 2170 114270 2410
rect 114310 2170 114330 2410
rect 114250 2140 114330 2170
rect 114360 2410 114440 2440
rect 114360 2170 114380 2410
rect 114420 2170 114440 2410
rect 114360 2140 114440 2170
rect 114470 2410 114550 2440
rect 114470 2170 114490 2410
rect 114530 2170 114550 2410
rect 114470 2140 114550 2170
rect 114580 2410 114660 2440
rect 114580 2170 114600 2410
rect 114640 2170 114660 2410
rect 114580 2140 114660 2170
rect 114690 2410 114770 2440
rect 114690 2170 114710 2410
rect 114750 2170 114770 2410
rect 114690 2140 114770 2170
rect 114800 2410 114880 2440
rect 114800 2170 114820 2410
rect 114860 2170 114880 2410
rect 114800 2140 114880 2170
rect 114910 2410 114990 2440
rect 114910 2170 114930 2410
rect 114970 2170 114990 2410
rect 114910 2140 114990 2170
rect 115020 2410 115100 2440
rect 115020 2170 115040 2410
rect 115080 2170 115100 2410
rect 115020 2140 115100 2170
rect 115130 2410 115210 2440
rect 115130 2170 115150 2410
rect 115190 2170 115210 2410
rect 115130 2140 115210 2170
rect 115240 2410 115320 2440
rect 115240 2170 115260 2410
rect 115300 2170 115320 2410
rect 115240 2140 115320 2170
rect 115350 2410 115430 2440
rect 115350 2170 115370 2410
rect 115410 2170 115430 2410
rect 115350 2140 115430 2170
rect 115460 2410 115540 2440
rect 115460 2170 115480 2410
rect 115520 2170 115540 2410
rect 116960 2310 116980 2850
rect 117020 2310 117040 2850
rect 116960 2280 117040 2310
rect 117070 2850 117150 2880
rect 117070 2310 117090 2850
rect 117130 2310 117150 2850
rect 117070 2280 117150 2310
rect 117180 2850 117260 2880
rect 117180 2310 117200 2850
rect 117240 2310 117260 2850
rect 117180 2280 117260 2310
rect 117290 2850 117370 2880
rect 117290 2310 117310 2850
rect 117350 2310 117370 2850
rect 117290 2280 117370 2310
rect 117400 2850 117480 2880
rect 117400 2310 117420 2850
rect 117460 2310 117480 2850
rect 117400 2280 117480 2310
rect 117510 2850 117590 2880
rect 117510 2310 117530 2850
rect 117570 2310 117590 2850
rect 117510 2280 117590 2310
rect 117620 2850 117700 2880
rect 117620 2310 117640 2850
rect 117680 2310 117700 2850
rect 117620 2280 117700 2310
rect 117730 2850 117810 2880
rect 117730 2310 117750 2850
rect 117790 2310 117810 2850
rect 117730 2280 117810 2310
rect 117840 2850 117920 2880
rect 117840 2310 117860 2850
rect 117900 2310 117920 2850
rect 117840 2280 117920 2310
rect 117950 2850 118030 2880
rect 117950 2310 117970 2850
rect 118010 2310 118030 2850
rect 117950 2280 118030 2310
rect 118060 2850 118140 2880
rect 118060 2310 118080 2850
rect 118120 2310 118140 2850
rect 118060 2280 118140 2310
rect 118170 2850 118250 2880
rect 118170 2310 118190 2850
rect 118230 2310 118250 2850
rect 118170 2280 118250 2310
rect 118280 2850 118360 2880
rect 118280 2310 118300 2850
rect 118340 2310 118360 2850
rect 118280 2280 118360 2310
rect 115460 2140 115540 2170
rect 112440 880 112520 910
rect 109300 650 109380 680
rect 109300 -690 109320 650
rect 109360 -690 109380 650
rect 109300 -720 109380 -690
rect 109500 650 109580 680
rect 109500 -690 109520 650
rect 109560 -690 109580 650
rect 109500 -720 109580 -690
rect 109700 650 109780 680
rect 109700 -690 109720 650
rect 109760 -690 109780 650
rect 109700 -720 109780 -690
rect 109900 650 109980 680
rect 109900 -690 109920 650
rect 109960 -690 109980 650
rect 109900 -720 109980 -690
rect 110100 650 110180 680
rect 110100 -690 110120 650
rect 110160 -690 110180 650
rect 110100 -720 110180 -690
rect 110300 650 110380 680
rect 110300 -690 110320 650
rect 110360 -690 110380 650
rect 110300 -720 110380 -690
rect 110500 650 110580 680
rect 110500 -690 110520 650
rect 110560 -690 110580 650
rect 112440 440 112460 880
rect 112500 440 112520 880
rect 112440 410 112520 440
rect 112550 880 112630 910
rect 112550 440 112570 880
rect 112610 440 112630 880
rect 112550 410 112630 440
rect 112660 880 112740 910
rect 112660 440 112680 880
rect 112720 440 112740 880
rect 112660 410 112740 440
rect 112770 880 112850 910
rect 112770 440 112790 880
rect 112830 440 112850 880
rect 112770 410 112850 440
rect 112880 880 112960 910
rect 112880 440 112900 880
rect 112940 440 112960 880
rect 112880 410 112960 440
rect 112990 880 113070 910
rect 112990 440 113010 880
rect 113050 440 113070 880
rect 112990 410 113070 440
rect 113100 880 113180 910
rect 113100 440 113120 880
rect 113160 440 113180 880
rect 113100 410 113180 440
rect 113210 880 113290 910
rect 113210 440 113230 880
rect 113270 440 113290 880
rect 113210 410 113290 440
rect 113320 880 113400 910
rect 113320 440 113340 880
rect 113380 440 113400 880
rect 113320 410 113400 440
rect 113430 880 113510 910
rect 113430 440 113450 880
rect 113490 440 113510 880
rect 113430 410 113510 440
rect 113540 880 113620 910
rect 113540 440 113560 880
rect 113600 440 113620 880
rect 113540 410 113620 440
rect 113650 880 113730 910
rect 113650 440 113670 880
rect 113710 440 113730 880
rect 113650 410 113730 440
rect 113760 880 113840 910
rect 113760 440 113780 880
rect 113820 440 113840 880
rect 113760 410 113840 440
rect 113870 880 113950 910
rect 113870 440 113890 880
rect 113930 440 113950 880
rect 113870 410 113950 440
rect 113980 880 114060 910
rect 113980 440 114000 880
rect 114040 440 114060 880
rect 113980 410 114060 440
rect 114090 880 114170 910
rect 114090 440 114110 880
rect 114150 440 114170 880
rect 114090 410 114170 440
rect 114200 880 114280 910
rect 114200 440 114220 880
rect 114260 440 114280 880
rect 114200 410 114280 440
rect 114310 880 114390 910
rect 114310 440 114330 880
rect 114370 440 114390 880
rect 114310 410 114390 440
rect 114420 880 114500 910
rect 114420 440 114440 880
rect 114480 440 114500 880
rect 114420 410 114500 440
rect 114530 880 114610 910
rect 114530 440 114550 880
rect 114590 440 114610 880
rect 114530 410 114610 440
rect 114640 880 114720 910
rect 114640 440 114660 880
rect 114700 440 114720 880
rect 114640 410 114720 440
rect 114750 880 114830 910
rect 114750 440 114770 880
rect 114810 440 114830 880
rect 114750 410 114830 440
rect 114860 880 114940 910
rect 114860 440 114880 880
rect 114920 440 114940 880
rect 114860 410 114940 440
rect 114970 880 115050 910
rect 114970 440 114990 880
rect 115030 440 115050 880
rect 114970 410 115050 440
rect 117020 650 117100 680
rect 110500 -720 110580 -690
rect 112860 -630 112940 -600
rect 112860 -870 112880 -630
rect 112920 -870 112940 -630
rect 112860 -900 112940 -870
rect 112970 -630 113050 -600
rect 112970 -870 112990 -630
rect 113030 -870 113050 -630
rect 112970 -900 113050 -870
rect 113080 -630 113160 -600
rect 113080 -870 113100 -630
rect 113140 -870 113160 -630
rect 113080 -900 113160 -870
rect 113190 -630 113270 -600
rect 113190 -870 113210 -630
rect 113250 -870 113270 -630
rect 113190 -900 113270 -870
rect 113300 -630 113380 -600
rect 113300 -870 113320 -630
rect 113360 -870 113380 -630
rect 113300 -900 113380 -870
rect 113410 -630 113490 -600
rect 113410 -870 113430 -630
rect 113470 -870 113490 -630
rect 113410 -900 113490 -870
rect 113520 -630 113600 -600
rect 113520 -870 113540 -630
rect 113580 -870 113600 -630
rect 113520 -900 113600 -870
rect 113740 -630 113820 -600
rect 113740 -870 113760 -630
rect 113800 -870 113820 -630
rect 113740 -900 113820 -870
rect 114420 -650 114500 -600
rect 114420 -850 114440 -650
rect 114480 -850 114500 -650
rect 117020 -690 117040 650
rect 117080 -690 117100 650
rect 117020 -720 117100 -690
rect 117220 650 117300 680
rect 117220 -690 117240 650
rect 117280 -690 117300 650
rect 117220 -720 117300 -690
rect 117420 650 117500 680
rect 117420 -690 117440 650
rect 117480 -690 117500 650
rect 117420 -720 117500 -690
rect 117620 650 117700 680
rect 117620 -690 117640 650
rect 117680 -690 117700 650
rect 117620 -720 117700 -690
rect 117820 650 117900 680
rect 117820 -690 117840 650
rect 117880 -690 117900 650
rect 117820 -720 117900 -690
rect 118020 650 118100 680
rect 118020 -690 118040 650
rect 118080 -690 118100 650
rect 118020 -720 118100 -690
rect 118220 650 118300 680
rect 118220 -690 118240 650
rect 118280 -690 118300 650
rect 118220 -720 118300 -690
rect 114420 -900 114500 -850
<< pdiff >>
rect 112170 9730 112250 9760
rect 112170 9090 112190 9730
rect 112230 9090 112250 9730
rect 112170 9060 112250 9090
rect 112290 9730 112370 9760
rect 112290 9090 112310 9730
rect 112350 9090 112370 9730
rect 112290 9060 112370 9090
rect 112410 9730 112490 9760
rect 112410 9090 112430 9730
rect 112470 9090 112490 9730
rect 112410 9060 112490 9090
rect 112530 9730 112610 9760
rect 112530 9090 112550 9730
rect 112590 9090 112610 9730
rect 114050 9730 114130 9760
rect 112530 9060 112610 9090
rect 113110 9390 113190 9420
rect 113110 9090 113130 9390
rect 113170 9090 113190 9390
rect 113110 9060 113190 9090
rect 113230 9390 113310 9420
rect 113230 9090 113250 9390
rect 113290 9090 113310 9390
rect 113230 9060 113310 9090
rect 113350 9390 113430 9420
rect 113350 9090 113370 9390
rect 113410 9090 113430 9390
rect 113350 9060 113430 9090
rect 113470 9390 113550 9420
rect 113470 9090 113490 9390
rect 113530 9090 113550 9390
rect 113470 9060 113550 9090
rect 114050 9090 114070 9730
rect 114110 9090 114130 9730
rect 114050 9060 114130 9090
rect 114170 9730 114250 9760
rect 114170 9090 114190 9730
rect 114230 9090 114250 9730
rect 114170 9060 114250 9090
rect 114290 9730 114370 9760
rect 114290 9090 114310 9730
rect 114350 9090 114370 9730
rect 114290 9060 114370 9090
rect 114410 9730 114490 9760
rect 114410 9090 114430 9730
rect 114470 9090 114490 9730
rect 114410 9060 114490 9090
rect 114990 9730 115070 9760
rect 114990 9090 115010 9730
rect 115050 9090 115070 9730
rect 114990 9060 115070 9090
rect 115110 9730 115190 9760
rect 115110 9090 115130 9730
rect 115170 9090 115190 9730
rect 115110 9060 115190 9090
rect 115230 9730 115310 9760
rect 115230 9090 115250 9730
rect 115290 9090 115310 9730
rect 115230 9060 115310 9090
rect 115350 9730 115430 9760
rect 115350 9090 115370 9730
rect 115410 9090 115430 9730
rect 115350 9060 115430 9090
rect 109180 7730 109260 7760
rect 109180 7090 109200 7730
rect 109240 7090 109260 7730
rect 109180 7060 109260 7090
rect 109300 7730 109380 7760
rect 109300 7090 109320 7730
rect 109360 7090 109380 7730
rect 109300 7060 109380 7090
rect 109420 7730 109500 7760
rect 109420 7090 109440 7730
rect 109480 7090 109500 7730
rect 109420 7060 109500 7090
rect 109540 7730 109620 7760
rect 109540 7090 109560 7730
rect 109600 7090 109620 7730
rect 109540 7060 109620 7090
rect 109660 7730 109740 7760
rect 109660 7090 109680 7730
rect 109720 7090 109740 7730
rect 109660 7060 109740 7090
rect 109780 7730 109860 7760
rect 109780 7090 109800 7730
rect 109840 7090 109860 7730
rect 109780 7060 109860 7090
rect 109900 7730 109980 7760
rect 109900 7090 109920 7730
rect 109960 7090 109980 7730
rect 109900 7060 109980 7090
rect 110020 7730 110100 7760
rect 110020 7090 110040 7730
rect 110080 7090 110100 7730
rect 110020 7060 110100 7090
rect 110140 7730 110220 7760
rect 110140 7090 110160 7730
rect 110200 7090 110220 7730
rect 110140 7060 110220 7090
rect 110260 7730 110340 7760
rect 110260 7090 110280 7730
rect 110320 7090 110340 7730
rect 110260 7060 110340 7090
rect 110380 7730 110460 7760
rect 110380 7090 110400 7730
rect 110440 7090 110460 7730
rect 110380 7060 110460 7090
rect 110500 7730 110580 7760
rect 110500 7090 110520 7730
rect 110560 7090 110580 7730
rect 110500 7060 110580 7090
rect 110620 7730 110700 7760
rect 110620 7090 110640 7730
rect 110680 7090 110700 7730
rect 110620 7060 110700 7090
rect 112010 7730 112090 7760
rect 112010 7090 112030 7730
rect 112070 7090 112090 7730
rect 112010 7060 112090 7090
rect 112130 7730 112210 7760
rect 112130 7090 112150 7730
rect 112190 7090 112210 7730
rect 112130 7060 112210 7090
rect 112250 7730 112330 7760
rect 112250 7090 112270 7730
rect 112310 7090 112330 7730
rect 112250 7060 112330 7090
rect 112370 7730 112450 7760
rect 112370 7090 112390 7730
rect 112430 7090 112450 7730
rect 112370 7060 112450 7090
rect 112490 7730 112570 7760
rect 112490 7090 112510 7730
rect 112550 7090 112570 7730
rect 112490 7060 112570 7090
rect 112610 7730 112690 7760
rect 112610 7090 112630 7730
rect 112670 7090 112690 7730
rect 112610 7060 112690 7090
rect 112730 7730 112810 7760
rect 112730 7090 112750 7730
rect 112790 7090 112810 7730
rect 112730 7060 112810 7090
rect 112850 7730 112930 7760
rect 112850 7090 112870 7730
rect 112910 7090 112930 7730
rect 112850 7060 112930 7090
rect 112970 7730 113050 7760
rect 112970 7090 112990 7730
rect 113030 7090 113050 7730
rect 112970 7060 113050 7090
rect 113090 7730 113170 7760
rect 113090 7090 113110 7730
rect 113150 7090 113170 7730
rect 113090 7060 113170 7090
rect 113210 7730 113290 7760
rect 113210 7090 113230 7730
rect 113270 7090 113290 7730
rect 113210 7060 113290 7090
rect 113330 7730 113410 7760
rect 113330 7090 113350 7730
rect 113390 7090 113410 7730
rect 113330 7060 113410 7090
rect 113450 7730 113530 7760
rect 113450 7090 113470 7730
rect 113510 7090 113530 7730
rect 113450 7060 113530 7090
rect 114070 7730 114150 7760
rect 114070 7090 114090 7730
rect 114130 7090 114150 7730
rect 114070 7060 114150 7090
rect 114190 7730 114270 7760
rect 114190 7090 114210 7730
rect 114250 7090 114270 7730
rect 114190 7060 114270 7090
rect 114310 7730 114390 7760
rect 114310 7090 114330 7730
rect 114370 7090 114390 7730
rect 114310 7060 114390 7090
rect 114430 7730 114510 7760
rect 114430 7090 114450 7730
rect 114490 7090 114510 7730
rect 114430 7060 114510 7090
rect 114550 7730 114630 7760
rect 114550 7090 114570 7730
rect 114610 7090 114630 7730
rect 114550 7060 114630 7090
rect 114670 7730 114750 7760
rect 114670 7090 114690 7730
rect 114730 7090 114750 7730
rect 114670 7060 114750 7090
rect 114790 7730 114870 7760
rect 114790 7090 114810 7730
rect 114850 7090 114870 7730
rect 114790 7060 114870 7090
rect 114910 7730 114990 7760
rect 114910 7090 114930 7730
rect 114970 7090 114990 7730
rect 114910 7060 114990 7090
rect 115030 7730 115110 7760
rect 115030 7090 115050 7730
rect 115090 7090 115110 7730
rect 115030 7060 115110 7090
rect 115150 7730 115230 7760
rect 115150 7090 115170 7730
rect 115210 7090 115230 7730
rect 115150 7060 115230 7090
rect 115270 7730 115350 7760
rect 115270 7090 115290 7730
rect 115330 7090 115350 7730
rect 115270 7060 115350 7090
rect 115390 7730 115470 7760
rect 115390 7090 115410 7730
rect 115450 7090 115470 7730
rect 115390 7060 115470 7090
rect 115510 7730 115590 7760
rect 115510 7090 115530 7730
rect 115570 7090 115590 7730
rect 115510 7060 115590 7090
rect 116900 7730 116980 7760
rect 116900 7090 116920 7730
rect 116960 7090 116980 7730
rect 116900 7060 116980 7090
rect 117020 7730 117100 7760
rect 117020 7090 117040 7730
rect 117080 7090 117100 7730
rect 117020 7060 117100 7090
rect 117140 7730 117220 7760
rect 117140 7090 117160 7730
rect 117200 7090 117220 7730
rect 117140 7060 117220 7090
rect 117260 7730 117340 7760
rect 117260 7090 117280 7730
rect 117320 7090 117340 7730
rect 117260 7060 117340 7090
rect 117380 7730 117460 7760
rect 117380 7090 117400 7730
rect 117440 7090 117460 7730
rect 117380 7060 117460 7090
rect 117500 7730 117580 7760
rect 117500 7090 117520 7730
rect 117560 7090 117580 7730
rect 117500 7060 117580 7090
rect 117620 7730 117700 7760
rect 117620 7090 117640 7730
rect 117680 7090 117700 7730
rect 117620 7060 117700 7090
rect 117740 7730 117820 7760
rect 117740 7090 117760 7730
rect 117800 7090 117820 7730
rect 117740 7060 117820 7090
rect 117860 7730 117940 7760
rect 117860 7090 117880 7730
rect 117920 7090 117940 7730
rect 117860 7060 117940 7090
rect 117980 7730 118060 7760
rect 117980 7090 118000 7730
rect 118040 7090 118060 7730
rect 117980 7060 118060 7090
rect 118100 7730 118180 7760
rect 118100 7090 118120 7730
rect 118160 7090 118180 7730
rect 118100 7060 118180 7090
rect 118220 7730 118300 7760
rect 118220 7090 118240 7730
rect 118280 7090 118300 7730
rect 118220 7060 118300 7090
rect 118340 7730 118420 7760
rect 118340 7090 118360 7730
rect 118400 7090 118420 7730
rect 118340 7060 118420 7090
rect 113020 6310 113100 6340
rect 109240 6280 109320 6310
rect 109240 5140 109260 6280
rect 109300 5140 109320 6280
rect 109240 5110 109320 5140
rect 109350 6280 109430 6310
rect 109350 5140 109370 6280
rect 109410 5140 109430 6280
rect 109350 5110 109430 5140
rect 109460 6280 109540 6310
rect 109460 5140 109480 6280
rect 109520 5140 109540 6280
rect 109460 5110 109540 5140
rect 109570 6280 109650 6310
rect 109570 5140 109590 6280
rect 109630 5140 109650 6280
rect 109570 5110 109650 5140
rect 109680 6280 109760 6310
rect 109680 5140 109700 6280
rect 109740 5140 109760 6280
rect 109680 5110 109760 5140
rect 109790 6280 109870 6310
rect 109790 5140 109810 6280
rect 109850 5140 109870 6280
rect 109790 5110 109870 5140
rect 109900 6280 109980 6310
rect 109900 5140 109920 6280
rect 109960 5140 109980 6280
rect 109900 5110 109980 5140
rect 110010 6280 110090 6310
rect 110010 5140 110030 6280
rect 110070 5140 110090 6280
rect 110010 5110 110090 5140
rect 110120 6280 110200 6310
rect 110120 5140 110140 6280
rect 110180 5140 110200 6280
rect 110120 5110 110200 5140
rect 110230 6280 110310 6310
rect 110230 5140 110250 6280
rect 110290 5140 110310 6280
rect 110230 5110 110310 5140
rect 110340 6280 110420 6310
rect 110340 5140 110360 6280
rect 110400 5140 110420 6280
rect 110340 5110 110420 5140
rect 110450 6280 110530 6310
rect 110450 5140 110470 6280
rect 110510 5140 110530 6280
rect 110450 5110 110530 5140
rect 110560 6280 110640 6310
rect 110560 5140 110580 6280
rect 110620 5140 110640 6280
rect 113020 6270 113040 6310
rect 113080 6270 113100 6310
rect 113020 6210 113100 6270
rect 113020 6170 113040 6210
rect 113080 6170 113100 6210
rect 113020 6110 113100 6170
rect 113020 6070 113040 6110
rect 113080 6070 113100 6110
rect 113020 6010 113100 6070
rect 113020 5970 113040 6010
rect 113080 5970 113100 6010
rect 113020 5910 113100 5970
rect 113020 5870 113040 5910
rect 113080 5870 113100 5910
rect 113020 5840 113100 5870
rect 113130 6310 113210 6340
rect 113130 6270 113150 6310
rect 113190 6270 113210 6310
rect 113130 6210 113210 6270
rect 113130 6170 113150 6210
rect 113190 6170 113210 6210
rect 113130 6110 113210 6170
rect 113130 6070 113150 6110
rect 113190 6070 113210 6110
rect 113130 6010 113210 6070
rect 113130 5970 113150 6010
rect 113190 5970 113210 6010
rect 113130 5910 113210 5970
rect 113130 5870 113150 5910
rect 113190 5870 113210 5910
rect 113130 5840 113210 5870
rect 113240 6310 113320 6340
rect 113240 6270 113260 6310
rect 113300 6270 113320 6310
rect 113240 6210 113320 6270
rect 113240 6170 113260 6210
rect 113300 6170 113320 6210
rect 113240 6110 113320 6170
rect 113240 6070 113260 6110
rect 113300 6070 113320 6110
rect 113240 6010 113320 6070
rect 113240 5970 113260 6010
rect 113300 5970 113320 6010
rect 113240 5910 113320 5970
rect 113240 5870 113260 5910
rect 113300 5870 113320 5910
rect 113240 5840 113320 5870
rect 113350 6310 113430 6340
rect 113350 6270 113370 6310
rect 113410 6270 113430 6310
rect 113350 6210 113430 6270
rect 113350 6170 113370 6210
rect 113410 6170 113430 6210
rect 113350 6110 113430 6170
rect 113350 6070 113370 6110
rect 113410 6070 113430 6110
rect 113350 6010 113430 6070
rect 113350 5970 113370 6010
rect 113410 5970 113430 6010
rect 113350 5910 113430 5970
rect 113350 5870 113370 5910
rect 113410 5870 113430 5910
rect 113350 5840 113430 5870
rect 113460 6310 113540 6340
rect 113460 6270 113480 6310
rect 113520 6270 113540 6310
rect 113460 6210 113540 6270
rect 113460 6170 113480 6210
rect 113520 6170 113540 6210
rect 113460 6110 113540 6170
rect 113460 6070 113480 6110
rect 113520 6070 113540 6110
rect 113460 6010 113540 6070
rect 113460 5970 113480 6010
rect 113520 5970 113540 6010
rect 113460 5910 113540 5970
rect 113460 5870 113480 5910
rect 113520 5870 113540 5910
rect 113460 5840 113540 5870
rect 113570 6310 113650 6340
rect 113570 6270 113590 6310
rect 113630 6270 113650 6310
rect 113570 6210 113650 6270
rect 113570 6170 113590 6210
rect 113630 6170 113650 6210
rect 113570 6110 113650 6170
rect 113570 6070 113590 6110
rect 113630 6070 113650 6110
rect 113570 6010 113650 6070
rect 113570 5970 113590 6010
rect 113630 5970 113650 6010
rect 113570 5910 113650 5970
rect 113570 5870 113590 5910
rect 113630 5870 113650 5910
rect 113570 5840 113650 5870
rect 113680 6310 113760 6340
rect 113840 6310 113920 6340
rect 113680 6270 113700 6310
rect 113740 6270 113760 6310
rect 113840 6270 113860 6310
rect 113900 6270 113920 6310
rect 113680 6210 113760 6270
rect 113840 6210 113920 6270
rect 113680 6170 113700 6210
rect 113740 6170 113760 6210
rect 113840 6170 113860 6210
rect 113900 6170 113920 6210
rect 113680 6110 113760 6170
rect 113840 6110 113920 6170
rect 113680 6070 113700 6110
rect 113740 6070 113760 6110
rect 113840 6070 113860 6110
rect 113900 6070 113920 6110
rect 113680 6010 113760 6070
rect 113840 6010 113920 6070
rect 113680 5970 113700 6010
rect 113740 5970 113760 6010
rect 113840 5970 113860 6010
rect 113900 5970 113920 6010
rect 113680 5910 113760 5970
rect 113840 5910 113920 5970
rect 113680 5870 113700 5910
rect 113740 5870 113760 5910
rect 113840 5870 113860 5910
rect 113900 5870 113920 5910
rect 113680 5840 113760 5870
rect 113840 5840 113920 5870
rect 113950 6310 114030 6340
rect 113950 6270 113970 6310
rect 114010 6270 114030 6310
rect 113950 6210 114030 6270
rect 113950 6170 113970 6210
rect 114010 6170 114030 6210
rect 113950 6110 114030 6170
rect 113950 6070 113970 6110
rect 114010 6070 114030 6110
rect 113950 6010 114030 6070
rect 113950 5970 113970 6010
rect 114010 5970 114030 6010
rect 113950 5910 114030 5970
rect 113950 5870 113970 5910
rect 114010 5870 114030 5910
rect 113950 5840 114030 5870
rect 114060 6310 114140 6340
rect 114060 6270 114080 6310
rect 114120 6270 114140 6310
rect 114060 6210 114140 6270
rect 114060 6170 114080 6210
rect 114120 6170 114140 6210
rect 114060 6110 114140 6170
rect 114060 6070 114080 6110
rect 114120 6070 114140 6110
rect 114060 6010 114140 6070
rect 114060 5970 114080 6010
rect 114120 5970 114140 6010
rect 114060 5910 114140 5970
rect 114060 5870 114080 5910
rect 114120 5870 114140 5910
rect 114060 5840 114140 5870
rect 114170 6310 114250 6340
rect 114170 6270 114190 6310
rect 114230 6270 114250 6310
rect 114170 6210 114250 6270
rect 114170 6170 114190 6210
rect 114230 6170 114250 6210
rect 114170 6110 114250 6170
rect 114170 6070 114190 6110
rect 114230 6070 114250 6110
rect 114170 6010 114250 6070
rect 114170 5970 114190 6010
rect 114230 5970 114250 6010
rect 114170 5910 114250 5970
rect 114170 5870 114190 5910
rect 114230 5870 114250 5910
rect 114170 5840 114250 5870
rect 114280 6310 114360 6340
rect 114280 6270 114300 6310
rect 114340 6270 114360 6310
rect 114280 6210 114360 6270
rect 114280 6170 114300 6210
rect 114340 6170 114360 6210
rect 114280 6110 114360 6170
rect 114280 6070 114300 6110
rect 114340 6070 114360 6110
rect 114280 6010 114360 6070
rect 114280 5970 114300 6010
rect 114340 5970 114360 6010
rect 114280 5910 114360 5970
rect 114280 5870 114300 5910
rect 114340 5870 114360 5910
rect 114280 5840 114360 5870
rect 114390 6310 114470 6340
rect 114390 6270 114410 6310
rect 114450 6270 114470 6310
rect 114390 6210 114470 6270
rect 114390 6170 114410 6210
rect 114450 6170 114470 6210
rect 114390 6110 114470 6170
rect 114390 6070 114410 6110
rect 114450 6070 114470 6110
rect 114390 6010 114470 6070
rect 114390 5970 114410 6010
rect 114450 5970 114470 6010
rect 114390 5910 114470 5970
rect 114390 5870 114410 5910
rect 114450 5870 114470 5910
rect 114390 5840 114470 5870
rect 114500 6310 114580 6340
rect 114500 6270 114520 6310
rect 114560 6270 114580 6310
rect 114500 6210 114580 6270
rect 114500 6170 114520 6210
rect 114560 6170 114580 6210
rect 114500 6110 114580 6170
rect 114500 6070 114520 6110
rect 114560 6070 114580 6110
rect 114500 6010 114580 6070
rect 114500 5970 114520 6010
rect 114560 5970 114580 6010
rect 114500 5910 114580 5970
rect 114500 5870 114520 5910
rect 114560 5870 114580 5910
rect 114500 5840 114580 5870
rect 116960 6280 117040 6310
rect 110560 5110 110640 5140
rect 116960 5140 116980 6280
rect 117020 5140 117040 6280
rect 116960 5110 117040 5140
rect 117070 6280 117150 6310
rect 117070 5140 117090 6280
rect 117130 5140 117150 6280
rect 117070 5110 117150 5140
rect 117180 6280 117260 6310
rect 117180 5140 117200 6280
rect 117240 5140 117260 6280
rect 117180 5110 117260 5140
rect 117290 6280 117370 6310
rect 117290 5140 117310 6280
rect 117350 5140 117370 6280
rect 117290 5110 117370 5140
rect 117400 6280 117480 6310
rect 117400 5140 117420 6280
rect 117460 5140 117480 6280
rect 117400 5110 117480 5140
rect 117510 6280 117590 6310
rect 117510 5140 117530 6280
rect 117570 5140 117590 6280
rect 117510 5110 117590 5140
rect 117620 6280 117700 6310
rect 117620 5140 117640 6280
rect 117680 5140 117700 6280
rect 117620 5110 117700 5140
rect 117730 6280 117810 6310
rect 117730 5140 117750 6280
rect 117790 5140 117810 6280
rect 117730 5110 117810 5140
rect 117840 6280 117920 6310
rect 117840 5140 117860 6280
rect 117900 5140 117920 6280
rect 117840 5110 117920 5140
rect 117950 6280 118030 6310
rect 117950 5140 117970 6280
rect 118010 5140 118030 6280
rect 117950 5110 118030 5140
rect 118060 6280 118140 6310
rect 118060 5140 118080 6280
rect 118120 5140 118140 6280
rect 118060 5110 118140 5140
rect 118170 6280 118250 6310
rect 118170 5140 118190 6280
rect 118230 5140 118250 6280
rect 118170 5110 118250 5140
rect 118280 6280 118360 6310
rect 118280 5140 118300 6280
rect 118340 5140 118360 6280
rect 118280 5110 118360 5140
rect 109240 3730 109320 3760
rect 109240 3390 109260 3730
rect 109300 3390 109320 3730
rect 109240 3360 109320 3390
rect 109350 3730 109430 3760
rect 109350 3390 109370 3730
rect 109410 3390 109430 3730
rect 109350 3360 109430 3390
rect 109460 3730 109540 3760
rect 109460 3390 109480 3730
rect 109520 3390 109540 3730
rect 109460 3360 109540 3390
rect 109570 3730 109650 3760
rect 109570 3390 109590 3730
rect 109630 3390 109650 3730
rect 109570 3360 109650 3390
rect 109680 3730 109760 3760
rect 109680 3390 109700 3730
rect 109740 3390 109760 3730
rect 109680 3360 109760 3390
rect 109790 3730 109870 3760
rect 109790 3390 109810 3730
rect 109850 3390 109870 3730
rect 109790 3360 109870 3390
rect 109900 3730 109980 3760
rect 109900 3390 109920 3730
rect 109960 3390 109980 3730
rect 109900 3360 109980 3390
rect 110010 3730 110090 3760
rect 110010 3390 110030 3730
rect 110070 3390 110090 3730
rect 110010 3360 110090 3390
rect 110120 3730 110200 3760
rect 110120 3390 110140 3730
rect 110180 3390 110200 3730
rect 110120 3360 110200 3390
rect 110230 3730 110310 3760
rect 110230 3390 110250 3730
rect 110290 3390 110310 3730
rect 110230 3360 110310 3390
rect 110340 3730 110420 3760
rect 110340 3390 110360 3730
rect 110400 3390 110420 3730
rect 110340 3360 110420 3390
rect 110450 3730 110530 3760
rect 110450 3390 110470 3730
rect 110510 3390 110530 3730
rect 110450 3360 110530 3390
rect 110560 3730 110640 3760
rect 110560 3390 110580 3730
rect 110620 3390 110640 3730
rect 116960 3730 117040 3760
rect 110560 3360 110640 3390
rect 116960 3390 116980 3730
rect 117020 3390 117040 3730
rect 116960 3360 117040 3390
rect 117070 3730 117150 3760
rect 117070 3390 117090 3730
rect 117130 3390 117150 3730
rect 117070 3360 117150 3390
rect 117180 3730 117260 3760
rect 117180 3390 117200 3730
rect 117240 3390 117260 3730
rect 117180 3360 117260 3390
rect 117290 3730 117370 3760
rect 117290 3390 117310 3730
rect 117350 3390 117370 3730
rect 117290 3360 117370 3390
rect 117400 3730 117480 3760
rect 117400 3390 117420 3730
rect 117460 3390 117480 3730
rect 117400 3360 117480 3390
rect 117510 3730 117590 3760
rect 117510 3390 117530 3730
rect 117570 3390 117590 3730
rect 117510 3360 117590 3390
rect 117620 3730 117700 3760
rect 117620 3390 117640 3730
rect 117680 3390 117700 3730
rect 117620 3360 117700 3390
rect 117730 3730 117810 3760
rect 117730 3390 117750 3730
rect 117790 3390 117810 3730
rect 117730 3360 117810 3390
rect 117840 3730 117920 3760
rect 117840 3390 117860 3730
rect 117900 3390 117920 3730
rect 117840 3360 117920 3390
rect 117950 3730 118030 3760
rect 117950 3390 117970 3730
rect 118010 3390 118030 3730
rect 117950 3360 118030 3390
rect 118060 3730 118140 3760
rect 118060 3390 118080 3730
rect 118120 3390 118140 3730
rect 118060 3360 118140 3390
rect 118170 3730 118250 3760
rect 118170 3390 118190 3730
rect 118230 3390 118250 3730
rect 118170 3360 118250 3390
rect 118280 3730 118360 3760
rect 118280 3390 118300 3730
rect 118340 3390 118360 3730
rect 118280 3360 118360 3390
<< ndiffc >>
rect 113560 4660 113600 5100
rect 113670 4660 113710 5100
rect 113780 4660 113820 5100
rect 113890 4660 113930 5100
rect 114000 4660 114040 5100
rect 112080 3540 112120 3780
rect 112190 3540 112230 3780
rect 112300 3540 112340 3780
rect 112410 3540 112450 3780
rect 112520 3540 112560 3780
rect 112630 3540 112670 3780
rect 112740 3540 112780 3780
rect 112850 3540 112890 3780
rect 112960 3540 113000 3780
rect 113070 3540 113110 3780
rect 113180 3540 113220 3780
rect 113290 3540 113330 3780
rect 113400 3540 113440 3780
rect 114160 3540 114200 3780
rect 114270 3540 114310 3780
rect 114380 3540 114420 3780
rect 114490 3540 114530 3780
rect 114600 3540 114640 3780
rect 114710 3540 114750 3780
rect 114820 3540 114860 3780
rect 114930 3540 114970 3780
rect 115040 3540 115080 3780
rect 115150 3540 115190 3780
rect 115260 3540 115300 3780
rect 115370 3540 115410 3780
rect 115480 3540 115520 3780
rect 109260 2310 109300 2850
rect 109370 2310 109410 2850
rect 109480 2310 109520 2850
rect 109590 2310 109630 2850
rect 109700 2310 109740 2850
rect 109810 2310 109850 2850
rect 109920 2310 109960 2850
rect 110030 2310 110070 2850
rect 110140 2310 110180 2850
rect 110250 2310 110290 2850
rect 110360 2310 110400 2850
rect 110470 2310 110510 2850
rect 110580 2310 110620 2850
rect 112080 2170 112120 2410
rect 112190 2170 112230 2410
rect 112300 2170 112340 2410
rect 112410 2170 112450 2410
rect 112520 2170 112560 2410
rect 112630 2170 112670 2410
rect 112740 2170 112780 2410
rect 112850 2170 112890 2410
rect 112960 2170 113000 2410
rect 113070 2170 113110 2410
rect 113180 2170 113220 2410
rect 113290 2170 113330 2410
rect 113400 2170 113440 2410
rect 113560 2170 113600 2410
rect 113670 2170 113710 2410
rect 113780 2170 113820 2410
rect 113890 2170 113930 2410
rect 114000 2170 114040 2410
rect 114160 2170 114200 2410
rect 114270 2170 114310 2410
rect 114380 2170 114420 2410
rect 114490 2170 114530 2410
rect 114600 2170 114640 2410
rect 114710 2170 114750 2410
rect 114820 2170 114860 2410
rect 114930 2170 114970 2410
rect 115040 2170 115080 2410
rect 115150 2170 115190 2410
rect 115260 2170 115300 2410
rect 115370 2170 115410 2410
rect 115480 2170 115520 2410
rect 116980 2310 117020 2850
rect 117090 2310 117130 2850
rect 117200 2310 117240 2850
rect 117310 2310 117350 2850
rect 117420 2310 117460 2850
rect 117530 2310 117570 2850
rect 117640 2310 117680 2850
rect 117750 2310 117790 2850
rect 117860 2310 117900 2850
rect 117970 2310 118010 2850
rect 118080 2310 118120 2850
rect 118190 2310 118230 2850
rect 118300 2310 118340 2850
rect 109320 -690 109360 650
rect 109520 -690 109560 650
rect 109720 -690 109760 650
rect 109920 -690 109960 650
rect 110120 -690 110160 650
rect 110320 -690 110360 650
rect 110520 -690 110560 650
rect 112460 440 112500 880
rect 112570 440 112610 880
rect 112680 440 112720 880
rect 112790 440 112830 880
rect 112900 440 112940 880
rect 113010 440 113050 880
rect 113120 440 113160 880
rect 113230 440 113270 880
rect 113340 440 113380 880
rect 113450 440 113490 880
rect 113560 440 113600 880
rect 113670 440 113710 880
rect 113780 440 113820 880
rect 113890 440 113930 880
rect 114000 440 114040 880
rect 114110 440 114150 880
rect 114220 440 114260 880
rect 114330 440 114370 880
rect 114440 440 114480 880
rect 114550 440 114590 880
rect 114660 440 114700 880
rect 114770 440 114810 880
rect 114880 440 114920 880
rect 114990 440 115030 880
rect 112880 -870 112920 -630
rect 112990 -870 113030 -630
rect 113100 -870 113140 -630
rect 113210 -870 113250 -630
rect 113320 -870 113360 -630
rect 113430 -870 113470 -630
rect 113540 -870 113580 -630
rect 113760 -870 113800 -630
rect 114440 -850 114480 -650
rect 117040 -690 117080 650
rect 117240 -690 117280 650
rect 117440 -690 117480 650
rect 117640 -690 117680 650
rect 117840 -690 117880 650
rect 118040 -690 118080 650
rect 118240 -690 118280 650
<< pdiffc >>
rect 112190 9090 112230 9730
rect 112310 9090 112350 9730
rect 112430 9090 112470 9730
rect 112550 9090 112590 9730
rect 113130 9090 113170 9390
rect 113250 9090 113290 9390
rect 113370 9090 113410 9390
rect 113490 9090 113530 9390
rect 114070 9090 114110 9730
rect 114190 9090 114230 9730
rect 114310 9090 114350 9730
rect 114430 9090 114470 9730
rect 115010 9090 115050 9730
rect 115130 9090 115170 9730
rect 115250 9090 115290 9730
rect 115370 9090 115410 9730
rect 109200 7090 109240 7730
rect 109320 7090 109360 7730
rect 109440 7090 109480 7730
rect 109560 7090 109600 7730
rect 109680 7090 109720 7730
rect 109800 7090 109840 7730
rect 109920 7090 109960 7730
rect 110040 7090 110080 7730
rect 110160 7090 110200 7730
rect 110280 7090 110320 7730
rect 110400 7090 110440 7730
rect 110520 7090 110560 7730
rect 110640 7090 110680 7730
rect 112030 7090 112070 7730
rect 112150 7090 112190 7730
rect 112270 7090 112310 7730
rect 112390 7090 112430 7730
rect 112510 7090 112550 7730
rect 112630 7090 112670 7730
rect 112750 7090 112790 7730
rect 112870 7090 112910 7730
rect 112990 7090 113030 7730
rect 113110 7090 113150 7730
rect 113230 7090 113270 7730
rect 113350 7090 113390 7730
rect 113470 7090 113510 7730
rect 114090 7090 114130 7730
rect 114210 7090 114250 7730
rect 114330 7090 114370 7730
rect 114450 7090 114490 7730
rect 114570 7090 114610 7730
rect 114690 7090 114730 7730
rect 114810 7090 114850 7730
rect 114930 7090 114970 7730
rect 115050 7090 115090 7730
rect 115170 7090 115210 7730
rect 115290 7090 115330 7730
rect 115410 7090 115450 7730
rect 115530 7090 115570 7730
rect 116920 7090 116960 7730
rect 117040 7090 117080 7730
rect 117160 7090 117200 7730
rect 117280 7090 117320 7730
rect 117400 7090 117440 7730
rect 117520 7090 117560 7730
rect 117640 7090 117680 7730
rect 117760 7090 117800 7730
rect 117880 7090 117920 7730
rect 118000 7090 118040 7730
rect 118120 7090 118160 7730
rect 118240 7090 118280 7730
rect 118360 7090 118400 7730
rect 109260 5140 109300 6280
rect 109370 5140 109410 6280
rect 109480 5140 109520 6280
rect 109590 5140 109630 6280
rect 109700 5140 109740 6280
rect 109810 5140 109850 6280
rect 109920 5140 109960 6280
rect 110030 5140 110070 6280
rect 110140 5140 110180 6280
rect 110250 5140 110290 6280
rect 110360 5140 110400 6280
rect 110470 5140 110510 6280
rect 110580 5140 110620 6280
rect 113040 6270 113080 6310
rect 113040 6170 113080 6210
rect 113040 6070 113080 6110
rect 113040 5970 113080 6010
rect 113040 5870 113080 5910
rect 113150 6270 113190 6310
rect 113150 6170 113190 6210
rect 113150 6070 113190 6110
rect 113150 5970 113190 6010
rect 113150 5870 113190 5910
rect 113260 6270 113300 6310
rect 113260 6170 113300 6210
rect 113260 6070 113300 6110
rect 113260 5970 113300 6010
rect 113260 5870 113300 5910
rect 113370 6270 113410 6310
rect 113370 6170 113410 6210
rect 113370 6070 113410 6110
rect 113370 5970 113410 6010
rect 113370 5870 113410 5910
rect 113480 6270 113520 6310
rect 113480 6170 113520 6210
rect 113480 6070 113520 6110
rect 113480 5970 113520 6010
rect 113480 5870 113520 5910
rect 113590 6270 113630 6310
rect 113590 6170 113630 6210
rect 113590 6070 113630 6110
rect 113590 5970 113630 6010
rect 113590 5870 113630 5910
rect 113700 6270 113740 6310
rect 113860 6270 113900 6310
rect 113700 6170 113740 6210
rect 113860 6170 113900 6210
rect 113700 6070 113740 6110
rect 113860 6070 113900 6110
rect 113700 5970 113740 6010
rect 113860 5970 113900 6010
rect 113700 5870 113740 5910
rect 113860 5870 113900 5910
rect 113970 6270 114010 6310
rect 113970 6170 114010 6210
rect 113970 6070 114010 6110
rect 113970 5970 114010 6010
rect 113970 5870 114010 5910
rect 114080 6270 114120 6310
rect 114080 6170 114120 6210
rect 114080 6070 114120 6110
rect 114080 5970 114120 6010
rect 114080 5870 114120 5910
rect 114190 6270 114230 6310
rect 114190 6170 114230 6210
rect 114190 6070 114230 6110
rect 114190 5970 114230 6010
rect 114190 5870 114230 5910
rect 114300 6270 114340 6310
rect 114300 6170 114340 6210
rect 114300 6070 114340 6110
rect 114300 5970 114340 6010
rect 114300 5870 114340 5910
rect 114410 6270 114450 6310
rect 114410 6170 114450 6210
rect 114410 6070 114450 6110
rect 114410 5970 114450 6010
rect 114410 5870 114450 5910
rect 114520 6270 114560 6310
rect 114520 6170 114560 6210
rect 114520 6070 114560 6110
rect 114520 5970 114560 6010
rect 114520 5870 114560 5910
rect 116980 5140 117020 6280
rect 117090 5140 117130 6280
rect 117200 5140 117240 6280
rect 117310 5140 117350 6280
rect 117420 5140 117460 6280
rect 117530 5140 117570 6280
rect 117640 5140 117680 6280
rect 117750 5140 117790 6280
rect 117860 5140 117900 6280
rect 117970 5140 118010 6280
rect 118080 5140 118120 6280
rect 118190 5140 118230 6280
rect 118300 5140 118340 6280
rect 109260 3390 109300 3730
rect 109370 3390 109410 3730
rect 109480 3390 109520 3730
rect 109590 3390 109630 3730
rect 109700 3390 109740 3730
rect 109810 3390 109850 3730
rect 109920 3390 109960 3730
rect 110030 3390 110070 3730
rect 110140 3390 110180 3730
rect 110250 3390 110290 3730
rect 110360 3390 110400 3730
rect 110470 3390 110510 3730
rect 110580 3390 110620 3730
rect 116980 3390 117020 3730
rect 117090 3390 117130 3730
rect 117200 3390 117240 3730
rect 117310 3390 117350 3730
rect 117420 3390 117460 3730
rect 117530 3390 117570 3730
rect 117640 3390 117680 3730
rect 117750 3390 117790 3730
rect 117860 3390 117900 3730
rect 117970 3390 118010 3730
rect 118080 3390 118120 3730
rect 118190 3390 118230 3730
rect 118300 3390 118340 3730
<< psubdiff >>
rect 113460 5100 113540 5130
rect 113460 4660 113480 5100
rect 113520 4660 113540 5100
rect 113460 4630 113540 4660
rect 114060 5100 114140 5130
rect 114060 4660 114080 5100
rect 114120 4660 114140 5100
rect 114060 4630 114140 4660
rect 111980 3780 112060 3810
rect 111980 3540 112000 3780
rect 112040 3540 112060 3780
rect 111980 3510 112060 3540
rect 113460 3780 113540 3810
rect 113460 3540 113480 3780
rect 113520 3540 113540 3780
rect 113460 3510 113540 3540
rect 114060 3780 114140 3810
rect 114060 3540 114080 3780
rect 114120 3540 114140 3780
rect 114060 3510 114140 3540
rect 115540 3780 115620 3810
rect 115540 3540 115560 3780
rect 115600 3540 115620 3780
rect 115540 3510 115620 3540
rect 109160 2850 109240 2880
rect 109160 2310 109180 2850
rect 109220 2310 109240 2850
rect 109160 2280 109240 2310
rect 110640 2850 110720 2880
rect 110640 2310 110660 2850
rect 110700 2310 110720 2850
rect 116880 2850 116960 2880
rect 110640 2280 110720 2310
rect 111980 2410 112060 2440
rect 111980 2170 112000 2410
rect 112040 2170 112060 2410
rect 111980 2140 112060 2170
rect 113460 2410 113540 2440
rect 113460 2170 113480 2410
rect 113520 2170 113540 2410
rect 113460 2140 113540 2170
rect 114060 2410 114140 2440
rect 114060 2170 114080 2410
rect 114120 2170 114140 2410
rect 114060 2140 114140 2170
rect 115540 2410 115620 2440
rect 115540 2170 115560 2410
rect 115600 2170 115620 2410
rect 116880 2310 116900 2850
rect 116940 2310 116960 2850
rect 116880 2280 116960 2310
rect 118360 2850 118440 2880
rect 118360 2310 118380 2850
rect 118420 2310 118440 2850
rect 118360 2280 118440 2310
rect 115540 2140 115620 2170
rect 112360 880 112440 910
rect 109220 650 109300 680
rect 109220 -690 109240 650
rect 109280 -690 109300 650
rect 109220 -720 109300 -690
rect 110580 650 110660 680
rect 110580 -690 110600 650
rect 110640 -690 110660 650
rect 112360 440 112380 880
rect 112420 440 112440 880
rect 112360 410 112440 440
rect 115050 880 115130 910
rect 115050 440 115070 880
rect 115110 440 115130 880
rect 115050 410 115130 440
rect 116940 650 117020 680
rect 110580 -720 110660 -690
rect 112780 -630 112860 -600
rect 112780 -870 112800 -630
rect 112840 -870 112860 -630
rect 112780 -900 112860 -870
rect 113600 -630 113680 -600
rect 113600 -870 113620 -630
rect 113660 -870 113680 -630
rect 113600 -900 113680 -870
rect 116940 -690 116960 650
rect 117000 -690 117020 650
rect 116940 -720 117020 -690
rect 118300 650 118380 680
rect 118300 -690 118320 650
rect 118360 -690 118380 650
rect 118300 -720 118380 -690
<< nsubdiff >>
rect 112090 9730 112170 9760
rect 112090 9090 112110 9730
rect 112150 9090 112170 9730
rect 112090 9060 112170 9090
rect 112610 9730 112690 9760
rect 112610 9090 112630 9730
rect 112670 9090 112690 9730
rect 113970 9730 114050 9760
rect 112610 9060 112690 9090
rect 113030 9390 113110 9420
rect 113030 9090 113050 9390
rect 113090 9090 113110 9390
rect 113030 9060 113110 9090
rect 113550 9390 113630 9420
rect 113550 9090 113570 9390
rect 113610 9090 113630 9390
rect 113550 9060 113630 9090
rect 113970 9090 113990 9730
rect 114030 9090 114050 9730
rect 113970 9060 114050 9090
rect 114490 9730 114570 9760
rect 114490 9090 114510 9730
rect 114550 9090 114570 9730
rect 114490 9060 114570 9090
rect 114910 9730 114990 9760
rect 114910 9090 114930 9730
rect 114970 9090 114990 9730
rect 114910 9060 114990 9090
rect 115430 9730 115510 9760
rect 115430 9090 115450 9730
rect 115490 9090 115510 9730
rect 115430 9060 115510 9090
rect 109100 7730 109180 7760
rect 109100 7090 109120 7730
rect 109160 7090 109180 7730
rect 109100 7060 109180 7090
rect 110700 7730 110780 7760
rect 110700 7090 110720 7730
rect 110760 7090 110780 7730
rect 110700 7060 110780 7090
rect 111930 7730 112010 7760
rect 111930 7090 111950 7730
rect 111990 7090 112010 7730
rect 111930 7060 112010 7090
rect 113530 7730 113610 7760
rect 113530 7090 113550 7730
rect 113590 7090 113610 7730
rect 113530 7060 113610 7090
rect 113990 7730 114070 7760
rect 113990 7090 114010 7730
rect 114050 7090 114070 7730
rect 113990 7060 114070 7090
rect 115590 7730 115670 7760
rect 115590 7090 115610 7730
rect 115650 7090 115670 7730
rect 115590 7060 115670 7090
rect 116820 7730 116900 7760
rect 116820 7090 116840 7730
rect 116880 7090 116900 7730
rect 116820 7060 116900 7090
rect 118420 7730 118500 7760
rect 118420 7090 118440 7730
rect 118480 7090 118500 7730
rect 118420 7060 118500 7090
rect 112940 6310 113020 6340
rect 109160 6280 109240 6310
rect 109160 5140 109180 6280
rect 109220 5140 109240 6280
rect 109160 5110 109240 5140
rect 110640 6280 110720 6310
rect 110640 5140 110660 6280
rect 110700 5140 110720 6280
rect 112940 6270 112960 6310
rect 113000 6270 113020 6310
rect 112940 6210 113020 6270
rect 112940 6170 112960 6210
rect 113000 6170 113020 6210
rect 112940 6110 113020 6170
rect 112940 6070 112960 6110
rect 113000 6070 113020 6110
rect 112940 6010 113020 6070
rect 112940 5970 112960 6010
rect 113000 5970 113020 6010
rect 112940 5910 113020 5970
rect 112940 5870 112960 5910
rect 113000 5870 113020 5910
rect 112940 5840 113020 5870
rect 113760 6310 113840 6340
rect 113760 6270 113780 6310
rect 113820 6270 113840 6310
rect 113760 6210 113840 6270
rect 113760 6170 113780 6210
rect 113820 6170 113840 6210
rect 113760 6110 113840 6170
rect 113760 6070 113780 6110
rect 113820 6070 113840 6110
rect 113760 6010 113840 6070
rect 113760 5970 113780 6010
rect 113820 5970 113840 6010
rect 113760 5910 113840 5970
rect 113760 5870 113780 5910
rect 113820 5870 113840 5910
rect 113760 5840 113840 5870
rect 114580 6310 114660 6340
rect 114580 6270 114600 6310
rect 114640 6270 114660 6310
rect 114580 6210 114660 6270
rect 114580 6170 114600 6210
rect 114640 6170 114660 6210
rect 114580 6110 114660 6170
rect 114580 6070 114600 6110
rect 114640 6070 114660 6110
rect 114580 6010 114660 6070
rect 114580 5970 114600 6010
rect 114640 5970 114660 6010
rect 114580 5910 114660 5970
rect 114580 5870 114600 5910
rect 114640 5870 114660 5910
rect 114580 5840 114660 5870
rect 116880 6280 116960 6310
rect 110640 5110 110720 5140
rect 116880 5140 116900 6280
rect 116940 5140 116960 6280
rect 116880 5110 116960 5140
rect 118360 6280 118440 6310
rect 118360 5140 118380 6280
rect 118420 5140 118440 6280
rect 118360 5110 118440 5140
rect 109160 3730 109240 3760
rect 109160 3390 109180 3730
rect 109220 3390 109240 3730
rect 109160 3360 109240 3390
rect 110640 3730 110720 3760
rect 110640 3390 110660 3730
rect 110700 3390 110720 3730
rect 116880 3730 116960 3760
rect 110640 3360 110720 3390
rect 116880 3390 116900 3730
rect 116940 3390 116960 3730
rect 116880 3360 116960 3390
rect 118360 3730 118440 3760
rect 118360 3390 118380 3730
rect 118420 3390 118440 3730
rect 118360 3360 118440 3390
<< psubdiffcont >>
rect 113480 4660 113520 5100
rect 114080 4660 114120 5100
rect 112000 3540 112040 3780
rect 113480 3540 113520 3780
rect 114080 3540 114120 3780
rect 115560 3540 115600 3780
rect 109180 2310 109220 2850
rect 110660 2310 110700 2850
rect 112000 2170 112040 2410
rect 113480 2170 113520 2410
rect 114080 2170 114120 2410
rect 115560 2170 115600 2410
rect 116900 2310 116940 2850
rect 118380 2310 118420 2850
rect 109240 -690 109280 650
rect 110600 -690 110640 650
rect 112380 440 112420 880
rect 115070 440 115110 880
rect 112800 -870 112840 -630
rect 113620 -870 113660 -630
rect 116960 -690 117000 650
rect 118320 -690 118360 650
<< nsubdiffcont >>
rect 112110 9090 112150 9730
rect 112630 9090 112670 9730
rect 113050 9090 113090 9390
rect 113570 9090 113610 9390
rect 113990 9090 114030 9730
rect 114510 9090 114550 9730
rect 114930 9090 114970 9730
rect 115450 9090 115490 9730
rect 109120 7090 109160 7730
rect 110720 7090 110760 7730
rect 111950 7090 111990 7730
rect 113550 7090 113590 7730
rect 114010 7090 114050 7730
rect 115610 7090 115650 7730
rect 116840 7090 116880 7730
rect 118440 7090 118480 7730
rect 109180 5140 109220 6280
rect 110660 5140 110700 6280
rect 112960 6270 113000 6310
rect 112960 6170 113000 6210
rect 112960 6070 113000 6110
rect 112960 5970 113000 6010
rect 112960 5870 113000 5910
rect 113780 6270 113820 6310
rect 113780 6170 113820 6210
rect 113780 6070 113820 6110
rect 113780 5970 113820 6010
rect 113780 5870 113820 5910
rect 114600 6270 114640 6310
rect 114600 6170 114640 6210
rect 114600 6070 114640 6110
rect 114600 5970 114640 6010
rect 114600 5870 114640 5910
rect 116900 5140 116940 6280
rect 118380 5140 118420 6280
rect 109180 3390 109220 3730
rect 110660 3390 110700 3730
rect 116900 3390 116940 3730
rect 118380 3390 118420 3730
<< poly >>
rect 112170 9850 112250 9870
rect 112170 9810 112190 9850
rect 112230 9820 112250 9850
rect 112530 9850 112610 9870
rect 112530 9820 112550 9850
rect 112230 9810 112290 9820
rect 112170 9790 112290 9810
rect 112490 9810 112550 9820
rect 112590 9810 112610 9850
rect 112490 9790 112610 9810
rect 114050 9850 114130 9870
rect 114050 9810 114070 9850
rect 114110 9820 114130 9850
rect 114410 9850 114490 9870
rect 114410 9820 114430 9850
rect 114110 9810 114170 9820
rect 114050 9790 114170 9810
rect 114370 9810 114430 9820
rect 114470 9810 114490 9850
rect 114370 9790 114490 9810
rect 114990 9850 115070 9870
rect 114990 9810 115010 9850
rect 115050 9820 115070 9850
rect 115350 9850 115430 9870
rect 115350 9820 115370 9850
rect 115050 9810 115110 9820
rect 114990 9790 115110 9810
rect 115310 9810 115370 9820
rect 115410 9810 115430 9850
rect 115310 9790 115430 9810
rect 112250 9760 112290 9790
rect 112370 9760 112410 9790
rect 112490 9760 112530 9790
rect 114130 9760 114170 9790
rect 114250 9760 114290 9790
rect 114370 9760 114410 9790
rect 115070 9760 115110 9790
rect 115190 9760 115230 9790
rect 115310 9760 115350 9790
rect 113110 9510 113190 9530
rect 113110 9470 113130 9510
rect 113170 9480 113190 9510
rect 113470 9510 113550 9530
rect 113470 9480 113490 9510
rect 113170 9470 113230 9480
rect 113110 9450 113230 9470
rect 113430 9470 113490 9480
rect 113530 9470 113550 9510
rect 113430 9450 113550 9470
rect 113190 9420 113230 9450
rect 113310 9420 113350 9450
rect 113430 9420 113470 9450
rect 112250 9030 112290 9060
rect 112370 8970 112410 9060
rect 112490 9030 112530 9060
rect 113190 9030 113230 9060
rect 113310 8970 113350 9060
rect 113430 9030 113470 9060
rect 114130 9030 114170 9060
rect 112300 8950 112410 8970
rect 112300 8910 112320 8950
rect 112360 8910 112410 8950
rect 112300 8890 112410 8910
rect 113260 8950 113350 8970
rect 113260 8910 113270 8950
rect 113310 8940 113350 8950
rect 114250 8970 114290 9060
rect 114370 9030 114410 9060
rect 115070 9030 115110 9060
rect 114250 8950 114340 8970
rect 115190 8950 115230 9060
rect 115310 9030 115350 9060
rect 114250 8940 114290 8950
rect 113310 8910 113320 8940
rect 113260 8890 113320 8910
rect 114280 8910 114290 8940
rect 114330 8910 114340 8950
rect 114280 8890 114340 8910
rect 115152 8930 115230 8950
rect 115152 8890 115162 8930
rect 115202 8920 115230 8930
rect 115202 8890 115212 8920
rect 115152 8870 115212 8890
rect 112020 7850 112080 7870
rect 112020 7810 112030 7850
rect 112070 7820 112080 7850
rect 113460 7850 113520 7870
rect 113460 7820 113470 7850
rect 112070 7810 112130 7820
rect 112020 7790 112130 7810
rect 113410 7810 113470 7820
rect 113510 7810 113520 7850
rect 113410 7790 113520 7810
rect 114080 7850 114140 7870
rect 114080 7810 114090 7850
rect 114130 7820 114140 7850
rect 115520 7850 115580 7870
rect 115520 7820 115530 7850
rect 114130 7810 114190 7820
rect 114080 7790 114190 7810
rect 115470 7810 115530 7820
rect 115570 7810 115580 7850
rect 115470 7790 115580 7810
rect 116900 7850 116980 7870
rect 116900 7810 116920 7850
rect 116960 7820 116980 7850
rect 118340 7850 118420 7870
rect 118340 7820 118360 7850
rect 116960 7810 117020 7820
rect 116900 7790 117020 7810
rect 118300 7810 118360 7820
rect 118400 7810 118420 7850
rect 118300 7790 118420 7810
rect 109260 7760 109300 7790
rect 109380 7760 109420 7790
rect 109500 7760 109540 7790
rect 109620 7760 109660 7790
rect 109740 7760 109780 7790
rect 109860 7760 109900 7790
rect 109980 7760 110020 7790
rect 110100 7760 110140 7790
rect 110220 7760 110260 7790
rect 110340 7760 110380 7790
rect 110460 7760 110500 7790
rect 110580 7760 110620 7790
rect 112090 7760 112130 7790
rect 112210 7760 112250 7790
rect 112330 7760 112370 7790
rect 112450 7760 112490 7790
rect 112570 7760 112610 7790
rect 112690 7760 112730 7790
rect 112810 7760 112850 7790
rect 112930 7760 112970 7790
rect 113050 7760 113090 7790
rect 113170 7760 113210 7790
rect 113290 7760 113330 7790
rect 113410 7760 113450 7790
rect 114150 7760 114190 7790
rect 114270 7760 114310 7790
rect 114390 7760 114430 7790
rect 114510 7760 114550 7790
rect 114630 7760 114670 7790
rect 114750 7760 114790 7790
rect 114870 7760 114910 7790
rect 114990 7760 115030 7790
rect 115110 7760 115150 7790
rect 115230 7760 115270 7790
rect 115350 7760 115390 7790
rect 115470 7760 115510 7790
rect 116980 7760 117020 7790
rect 117100 7760 117140 7790
rect 117220 7760 117260 7790
rect 117340 7760 117380 7790
rect 117460 7760 117500 7790
rect 117580 7760 117620 7790
rect 117700 7760 117740 7790
rect 117820 7760 117860 7790
rect 117940 7760 117980 7790
rect 118060 7760 118100 7790
rect 118180 7760 118220 7790
rect 118300 7760 118340 7790
rect 109260 7030 109300 7060
rect 109380 6950 109420 7060
rect 109500 6950 109540 7060
rect 109620 6950 109660 7060
rect 109740 6950 109780 7060
rect 109860 6950 109900 7060
rect 109980 6950 110020 7060
rect 110100 6950 110140 7060
rect 110220 6950 110260 7060
rect 110340 6950 110380 7060
rect 110460 6950 110500 7060
rect 110580 7030 110620 7060
rect 112090 7030 112130 7060
rect 112210 6950 112250 7060
rect 112330 6950 112370 7060
rect 112450 6950 112490 7060
rect 112570 6950 112610 7060
rect 112690 6950 112730 7060
rect 112810 6950 112850 7060
rect 112930 6950 112970 7060
rect 113050 6950 113090 7060
rect 113170 6950 113210 7060
rect 113290 6950 113330 7060
rect 113410 7030 113450 7060
rect 114150 7030 114190 7060
rect 114270 6950 114310 7060
rect 114390 6950 114430 7060
rect 114510 6950 114550 7060
rect 114630 6950 114670 7060
rect 114750 6950 114790 7060
rect 114870 6950 114910 7060
rect 114990 6950 115030 7060
rect 115110 6950 115150 7060
rect 115230 6950 115270 7060
rect 115350 6950 115390 7060
rect 115470 7030 115510 7060
rect 116980 7030 117020 7060
rect 116910 7010 117020 7030
rect 116910 6970 116920 7010
rect 116960 7000 117020 7010
rect 116960 6970 116970 7000
rect 116910 6950 116970 6970
rect 117100 6950 117140 7060
rect 117220 6950 117260 7060
rect 117340 6950 117380 7060
rect 117460 6950 117500 7060
rect 117580 6950 117620 7060
rect 117700 6950 117740 7060
rect 117820 6950 117860 7060
rect 117940 6950 117980 7060
rect 118060 6950 118100 7060
rect 118180 6950 118220 7060
rect 118300 7030 118340 7060
rect 118300 7010 118410 7030
rect 118300 7000 118360 7010
rect 118350 6970 118360 7000
rect 118400 6970 118410 7010
rect 118350 6950 118410 6970
rect 109370 6930 109430 6950
rect 109370 6890 109380 6930
rect 109420 6890 109430 6930
rect 109370 6870 109430 6890
rect 109490 6930 109550 6950
rect 109490 6890 109500 6930
rect 109540 6890 109550 6930
rect 109490 6870 109550 6890
rect 109610 6930 109670 6950
rect 109610 6890 109620 6930
rect 109660 6890 109670 6930
rect 109610 6870 109670 6890
rect 109730 6930 109790 6950
rect 109730 6890 109740 6930
rect 109780 6890 109790 6930
rect 109730 6870 109790 6890
rect 109850 6930 109910 6950
rect 109850 6890 109860 6930
rect 109900 6890 109910 6930
rect 109850 6870 109910 6890
rect 109970 6930 110030 6950
rect 109970 6890 109980 6930
rect 110020 6890 110030 6930
rect 109970 6870 110030 6890
rect 110090 6930 110150 6950
rect 110090 6890 110100 6930
rect 110140 6890 110150 6930
rect 110090 6870 110150 6890
rect 110210 6930 110270 6950
rect 110210 6890 110220 6930
rect 110260 6890 110270 6930
rect 110210 6870 110270 6890
rect 110330 6930 110390 6950
rect 110330 6890 110340 6930
rect 110380 6890 110390 6930
rect 110330 6870 110390 6890
rect 110450 6930 110510 6950
rect 110450 6890 110460 6930
rect 110500 6890 110510 6930
rect 110450 6870 110510 6890
rect 112200 6930 112260 6950
rect 112200 6890 112210 6930
rect 112250 6890 112260 6930
rect 112200 6870 112260 6890
rect 112320 6930 112380 6950
rect 112320 6890 112330 6930
rect 112370 6890 112380 6930
rect 112320 6870 112380 6890
rect 112440 6930 112500 6950
rect 112440 6890 112450 6930
rect 112490 6890 112500 6930
rect 112440 6870 112500 6890
rect 112560 6930 112620 6950
rect 112560 6890 112570 6930
rect 112610 6890 112620 6930
rect 112560 6870 112620 6890
rect 112680 6930 112740 6950
rect 112680 6890 112690 6930
rect 112730 6890 112740 6930
rect 112680 6870 112740 6890
rect 112800 6930 112860 6950
rect 112800 6890 112810 6930
rect 112850 6890 112860 6930
rect 112800 6870 112860 6890
rect 112920 6930 112980 6950
rect 112920 6890 112930 6930
rect 112970 6890 112980 6930
rect 112920 6870 112980 6890
rect 113040 6930 113100 6950
rect 113040 6890 113050 6930
rect 113090 6890 113100 6930
rect 113040 6870 113100 6890
rect 113160 6930 113220 6950
rect 113160 6890 113170 6930
rect 113210 6890 113220 6930
rect 113160 6870 113220 6890
rect 113280 6930 113340 6950
rect 113280 6890 113290 6930
rect 113330 6890 113340 6930
rect 113280 6870 113340 6890
rect 114260 6930 114320 6950
rect 114260 6890 114270 6930
rect 114310 6890 114320 6930
rect 114260 6870 114320 6890
rect 114380 6930 114440 6950
rect 114380 6890 114390 6930
rect 114430 6890 114440 6930
rect 114380 6870 114440 6890
rect 114500 6930 114560 6950
rect 114500 6890 114510 6930
rect 114550 6890 114560 6930
rect 114500 6870 114560 6890
rect 114620 6930 114680 6950
rect 114620 6890 114630 6930
rect 114670 6890 114680 6930
rect 114620 6870 114680 6890
rect 114740 6930 114800 6950
rect 114740 6890 114750 6930
rect 114790 6890 114800 6930
rect 114740 6870 114800 6890
rect 114860 6930 114920 6950
rect 114860 6890 114870 6930
rect 114910 6890 114920 6930
rect 114860 6870 114920 6890
rect 114980 6930 115040 6950
rect 114980 6890 114990 6930
rect 115030 6890 115040 6930
rect 114980 6870 115040 6890
rect 115100 6930 115160 6950
rect 115100 6890 115110 6930
rect 115150 6890 115160 6930
rect 115100 6870 115160 6890
rect 115220 6930 115280 6950
rect 115220 6890 115230 6930
rect 115270 6890 115280 6930
rect 115220 6870 115280 6890
rect 115340 6930 115400 6950
rect 115340 6890 115350 6930
rect 115390 6890 115400 6930
rect 115340 6870 115400 6890
rect 117090 6930 117150 6950
rect 117090 6890 117100 6930
rect 117140 6890 117150 6930
rect 117090 6870 117150 6890
rect 117210 6930 117270 6950
rect 117210 6890 117220 6930
rect 117260 6890 117270 6930
rect 117210 6870 117270 6890
rect 117330 6930 117390 6950
rect 117330 6890 117340 6930
rect 117380 6890 117390 6930
rect 117330 6870 117390 6890
rect 117450 6930 117510 6950
rect 117450 6890 117460 6930
rect 117500 6890 117510 6930
rect 117450 6870 117510 6890
rect 117570 6930 117630 6950
rect 117570 6890 117580 6930
rect 117620 6890 117630 6930
rect 117570 6870 117630 6890
rect 117690 6930 117750 6950
rect 117690 6890 117700 6930
rect 117740 6890 117750 6930
rect 117690 6870 117750 6890
rect 117810 6930 117870 6950
rect 117810 6890 117820 6930
rect 117860 6890 117870 6930
rect 117810 6870 117870 6890
rect 117930 6930 117990 6950
rect 117930 6890 117940 6930
rect 117980 6890 117990 6930
rect 117930 6870 117990 6890
rect 118050 6930 118110 6950
rect 118050 6890 118060 6930
rect 118100 6890 118110 6930
rect 118050 6870 118110 6890
rect 118170 6930 118230 6950
rect 118170 6890 118180 6930
rect 118220 6890 118230 6930
rect 118170 6870 118230 6890
rect 113020 6540 113100 6560
rect 113020 6500 113040 6540
rect 113080 6510 113100 6540
rect 113680 6540 113760 6560
rect 113680 6510 113700 6540
rect 113080 6500 113130 6510
rect 113020 6480 113130 6500
rect 109250 6400 109310 6420
rect 109250 6360 109260 6400
rect 109300 6370 109310 6400
rect 110570 6400 110630 6420
rect 110570 6370 110580 6400
rect 109300 6360 109350 6370
rect 109250 6340 109350 6360
rect 110530 6360 110580 6370
rect 110620 6360 110630 6400
rect 110530 6340 110630 6360
rect 113100 6340 113130 6480
rect 113650 6500 113700 6510
rect 113740 6500 113760 6540
rect 113650 6480 113760 6500
rect 113840 6540 113920 6560
rect 113840 6500 113860 6540
rect 113900 6510 113920 6540
rect 114500 6540 114580 6560
rect 114500 6510 114520 6540
rect 113900 6500 113950 6510
rect 113840 6480 113950 6500
rect 113210 6340 113240 6370
rect 113320 6340 113350 6370
rect 113430 6340 113460 6370
rect 113540 6340 113570 6370
rect 113650 6340 113680 6480
rect 113920 6340 113950 6480
rect 114470 6500 114520 6510
rect 114560 6500 114580 6540
rect 114470 6480 114580 6500
rect 114030 6340 114060 6370
rect 114140 6340 114170 6370
rect 114250 6340 114280 6370
rect 114360 6340 114390 6370
rect 114470 6340 114500 6480
rect 116970 6400 117030 6420
rect 116970 6360 116980 6400
rect 117020 6370 117030 6400
rect 118290 6400 118350 6420
rect 118290 6370 118300 6400
rect 117020 6360 117070 6370
rect 116970 6340 117070 6360
rect 118250 6360 118300 6370
rect 118340 6360 118350 6400
rect 118250 6340 118350 6360
rect 109320 6310 109350 6340
rect 109430 6310 109460 6340
rect 109540 6310 109570 6340
rect 109650 6310 109680 6340
rect 109760 6310 109790 6340
rect 109870 6310 109900 6340
rect 109980 6310 110010 6340
rect 110090 6310 110120 6340
rect 110200 6310 110230 6340
rect 110310 6310 110340 6340
rect 110420 6310 110450 6340
rect 110530 6310 110560 6340
rect 117040 6310 117070 6340
rect 117150 6310 117180 6340
rect 117260 6310 117290 6340
rect 117370 6310 117400 6340
rect 117480 6310 117510 6340
rect 117590 6310 117620 6340
rect 117700 6310 117730 6340
rect 117810 6310 117840 6340
rect 117920 6310 117950 6340
rect 118030 6310 118060 6340
rect 118140 6310 118170 6340
rect 118250 6310 118280 6340
rect 113100 5810 113130 5840
rect 113210 5810 113240 5840
rect 113320 5820 113350 5840
rect 113430 5820 113460 5840
rect 113210 5790 113274 5810
rect 113320 5790 113460 5820
rect 113540 5810 113570 5840
rect 113650 5810 113680 5840
rect 113920 5810 113950 5840
rect 114030 5810 114060 5840
rect 114140 5820 114170 5840
rect 114250 5820 114280 5840
rect 113506 5790 113570 5810
rect 114030 5790 114094 5810
rect 114140 5790 114280 5820
rect 114360 5810 114390 5840
rect 114470 5810 114500 5840
rect 114326 5790 114390 5810
rect 113214 5750 113224 5790
rect 113264 5750 113274 5790
rect 113214 5730 113274 5750
rect 113350 5750 113370 5790
rect 113410 5750 113430 5790
rect 113350 5730 113430 5750
rect 113506 5750 113516 5790
rect 113556 5750 113566 5790
rect 113506 5730 113566 5750
rect 114034 5750 114044 5790
rect 114084 5750 114094 5790
rect 114034 5730 114094 5750
rect 114170 5750 114190 5790
rect 114230 5750 114250 5790
rect 114170 5730 114250 5750
rect 114326 5750 114336 5790
rect 114376 5750 114386 5790
rect 114326 5730 114386 5750
rect 113700 5220 113780 5240
rect 113700 5180 113720 5220
rect 113760 5180 113780 5220
rect 113700 5160 113870 5180
rect 113620 5130 113650 5160
rect 113730 5150 113870 5160
rect 113730 5130 113760 5150
rect 113840 5130 113870 5150
rect 113950 5130 113980 5160
rect 109320 5080 109350 5110
rect 109430 5090 109460 5110
rect 109540 5090 109570 5110
rect 109650 5090 109680 5110
rect 109760 5090 109790 5110
rect 109870 5090 109900 5110
rect 109980 5090 110010 5110
rect 110090 5090 110120 5110
rect 110200 5090 110230 5110
rect 110310 5090 110340 5110
rect 110420 5090 110450 5110
rect 109430 5060 110450 5090
rect 110530 5080 110560 5110
rect 109910 5020 109920 5060
rect 109960 5020 109970 5060
rect 109910 4950 109970 5020
rect 109900 4930 109980 4950
rect 109900 4890 109920 4930
rect 109960 4890 109980 4930
rect 109900 4850 109980 4890
rect 109900 4810 109920 4850
rect 109960 4810 109980 4850
rect 109900 4770 109980 4810
rect 109900 4730 109920 4770
rect 109960 4730 109980 4770
rect 109900 4710 109980 4730
rect 117040 5080 117070 5110
rect 117150 5090 117180 5110
rect 117260 5090 117290 5110
rect 117370 5090 117400 5110
rect 117480 5090 117510 5110
rect 117590 5090 117620 5110
rect 117700 5090 117730 5110
rect 117810 5090 117840 5110
rect 117920 5090 117950 5110
rect 118030 5090 118060 5110
rect 118140 5090 118170 5110
rect 117150 5060 118170 5090
rect 118250 5080 118280 5110
rect 117630 5020 117640 5060
rect 117680 5020 117690 5060
rect 117630 4950 117690 5020
rect 117620 4930 117700 4950
rect 117620 4890 117640 4930
rect 117680 4890 117700 4930
rect 117620 4850 117700 4890
rect 117620 4810 117640 4850
rect 117680 4810 117700 4850
rect 117620 4770 117700 4810
rect 117620 4730 117640 4770
rect 117680 4730 117700 4770
rect 117620 4710 117700 4730
rect 113620 4600 113650 4630
rect 113730 4600 113760 4630
rect 113840 4600 113870 4630
rect 113950 4600 113980 4630
rect 113540 4580 113650 4600
rect 113540 4540 113560 4580
rect 113600 4570 113650 4580
rect 113950 4580 114060 4600
rect 113950 4570 114000 4580
rect 113600 4540 113620 4570
rect 113540 4520 113620 4540
rect 113980 4540 114000 4570
rect 114040 4540 114060 4580
rect 113980 4520 114060 4540
rect 112232 3900 112298 3920
rect 109250 3850 109310 3870
rect 109250 3810 109260 3850
rect 109300 3820 109310 3850
rect 110570 3850 110630 3870
rect 110570 3820 110580 3850
rect 109300 3810 109350 3820
rect 109250 3790 109350 3810
rect 110530 3810 110580 3820
rect 110620 3810 110630 3850
rect 112232 3860 112245 3900
rect 112285 3860 112298 3900
rect 112232 3840 112298 3860
rect 112342 3900 112408 3920
rect 112342 3860 112355 3900
rect 112395 3860 112408 3900
rect 112342 3840 112408 3860
rect 112452 3900 112518 3920
rect 112452 3860 112465 3900
rect 112505 3860 112518 3900
rect 112452 3840 112518 3860
rect 112562 3900 112628 3920
rect 112562 3860 112575 3900
rect 112615 3860 112628 3900
rect 112562 3840 112628 3860
rect 112672 3900 112738 3920
rect 112672 3860 112685 3900
rect 112725 3860 112738 3900
rect 112672 3840 112738 3860
rect 112782 3900 112848 3920
rect 112782 3860 112795 3900
rect 112835 3860 112848 3900
rect 112782 3840 112848 3860
rect 112892 3900 112958 3920
rect 112892 3860 112905 3900
rect 112945 3860 112958 3900
rect 112892 3840 112958 3860
rect 113002 3900 113068 3920
rect 113002 3860 113015 3900
rect 113055 3860 113068 3900
rect 113002 3840 113068 3860
rect 113112 3900 113178 3920
rect 113112 3860 113125 3900
rect 113165 3860 113178 3900
rect 113112 3840 113178 3860
rect 113222 3900 113288 3920
rect 113222 3860 113235 3900
rect 113275 3860 113288 3900
rect 113222 3840 113288 3860
rect 114312 3900 114378 3920
rect 114312 3860 114325 3900
rect 114365 3860 114378 3900
rect 114312 3840 114378 3860
rect 114422 3900 114488 3920
rect 114422 3860 114435 3900
rect 114475 3860 114488 3900
rect 114422 3840 114488 3860
rect 114532 3900 114598 3920
rect 114532 3860 114545 3900
rect 114585 3860 114598 3900
rect 114532 3840 114598 3860
rect 114642 3900 114708 3920
rect 114642 3860 114655 3900
rect 114695 3860 114708 3900
rect 114642 3840 114708 3860
rect 114752 3900 114818 3920
rect 114752 3860 114765 3900
rect 114805 3860 114818 3900
rect 114752 3840 114818 3860
rect 114862 3900 114928 3920
rect 114862 3860 114875 3900
rect 114915 3860 114928 3900
rect 114862 3840 114928 3860
rect 114972 3900 115038 3920
rect 114972 3860 114985 3900
rect 115025 3860 115038 3900
rect 114972 3840 115038 3860
rect 115082 3900 115148 3920
rect 115082 3860 115095 3900
rect 115135 3860 115148 3900
rect 115082 3840 115148 3860
rect 115192 3900 115258 3920
rect 115192 3860 115205 3900
rect 115245 3860 115258 3900
rect 115192 3840 115258 3860
rect 115302 3900 115368 3920
rect 115302 3860 115315 3900
rect 115355 3860 115368 3900
rect 115302 3840 115368 3860
rect 116970 3850 117030 3870
rect 112140 3810 112170 3840
rect 112250 3810 112280 3840
rect 112360 3810 112390 3840
rect 112470 3810 112500 3840
rect 112580 3810 112610 3840
rect 112690 3810 112720 3840
rect 112800 3810 112830 3840
rect 112910 3810 112940 3840
rect 113020 3810 113050 3840
rect 113130 3810 113160 3840
rect 113240 3810 113270 3840
rect 113350 3810 113380 3840
rect 114220 3810 114250 3840
rect 114330 3810 114360 3840
rect 114440 3810 114470 3840
rect 114550 3810 114580 3840
rect 114660 3810 114690 3840
rect 114770 3810 114800 3840
rect 114880 3810 114910 3840
rect 114990 3810 115020 3840
rect 115100 3810 115130 3840
rect 115210 3810 115240 3840
rect 115320 3810 115350 3840
rect 115430 3810 115460 3840
rect 116970 3810 116980 3850
rect 117020 3820 117030 3850
rect 118290 3850 118350 3870
rect 118290 3820 118300 3850
rect 117020 3810 117070 3820
rect 110530 3790 110630 3810
rect 109320 3760 109350 3790
rect 109430 3760 109460 3790
rect 109540 3760 109570 3790
rect 109650 3760 109680 3790
rect 109760 3760 109790 3790
rect 109870 3760 109900 3790
rect 109980 3760 110010 3790
rect 110090 3760 110120 3790
rect 110200 3760 110230 3790
rect 110310 3760 110340 3790
rect 110420 3760 110450 3790
rect 110530 3760 110560 3790
rect 116970 3790 117070 3810
rect 118250 3810 118300 3820
rect 118340 3810 118350 3850
rect 118250 3790 118350 3810
rect 117040 3760 117070 3790
rect 117150 3760 117180 3790
rect 117260 3760 117290 3790
rect 117370 3760 117400 3790
rect 117480 3760 117510 3790
rect 117590 3760 117620 3790
rect 117700 3760 117730 3790
rect 117810 3760 117840 3790
rect 117920 3760 117950 3790
rect 118030 3760 118060 3790
rect 118140 3760 118170 3790
rect 118250 3760 118280 3790
rect 112140 3480 112170 3510
rect 112250 3480 112280 3510
rect 112360 3480 112390 3510
rect 112470 3480 112500 3510
rect 112580 3480 112610 3510
rect 112690 3480 112720 3510
rect 112800 3480 112830 3510
rect 112910 3480 112940 3510
rect 113020 3480 113050 3510
rect 113130 3480 113160 3510
rect 113240 3480 113270 3510
rect 113350 3480 113380 3510
rect 114220 3480 114250 3510
rect 114330 3480 114360 3510
rect 114440 3480 114470 3510
rect 114550 3480 114580 3510
rect 114660 3480 114690 3510
rect 114770 3480 114800 3510
rect 114880 3480 114910 3510
rect 114990 3480 115020 3510
rect 115100 3480 115130 3510
rect 115210 3480 115240 3510
rect 115320 3480 115350 3510
rect 115430 3480 115460 3510
rect 112070 3460 112170 3480
rect 112070 3420 112080 3460
rect 112120 3450 112170 3460
rect 113350 3460 113450 3480
rect 113350 3450 113400 3460
rect 112120 3420 112130 3450
rect 112070 3400 112130 3420
rect 113390 3420 113400 3450
rect 113440 3420 113450 3460
rect 113390 3400 113450 3420
rect 114150 3460 114250 3480
rect 114150 3420 114160 3460
rect 114200 3450 114250 3460
rect 115430 3460 115530 3480
rect 115430 3450 115480 3460
rect 114200 3420 114210 3450
rect 114150 3400 114210 3420
rect 115470 3420 115480 3450
rect 115520 3420 115530 3460
rect 115470 3400 115530 3420
rect 109320 3330 109350 3360
rect 109430 3340 109460 3360
rect 109540 3340 109570 3360
rect 109650 3340 109680 3360
rect 109760 3340 109790 3360
rect 109870 3340 109900 3360
rect 109980 3340 110010 3360
rect 110090 3340 110120 3360
rect 110200 3340 110230 3360
rect 110310 3340 110340 3360
rect 110420 3340 110450 3360
rect 109430 3310 110450 3340
rect 110530 3330 110560 3360
rect 117040 3330 117070 3360
rect 117150 3340 117180 3360
rect 117260 3340 117290 3360
rect 117370 3340 117400 3360
rect 117480 3340 117510 3360
rect 117590 3340 117620 3360
rect 117700 3340 117730 3360
rect 117810 3340 117840 3360
rect 117920 3340 117950 3360
rect 118030 3340 118060 3360
rect 118140 3340 118170 3360
rect 117150 3310 118170 3340
rect 118250 3330 118280 3360
rect 110240 3270 110250 3310
rect 110290 3270 110300 3310
rect 110240 3250 110300 3270
rect 117300 3270 117310 3310
rect 117350 3270 117360 3310
rect 117300 3250 117360 3270
rect 110250 3200 110290 3250
rect 117310 3200 117350 3250
rect 110230 3180 110310 3200
rect 110230 3140 110250 3180
rect 110290 3140 110310 3180
rect 110230 3100 110310 3140
rect 110230 3060 110250 3100
rect 110290 3060 110310 3100
rect 110230 3040 110310 3060
rect 117290 3180 117370 3200
rect 117290 3140 117310 3180
rect 117350 3140 117370 3180
rect 117290 3100 117370 3140
rect 117290 3060 117310 3100
rect 117350 3060 117370 3100
rect 117290 3040 117370 3060
rect 110250 2990 110290 3040
rect 117310 2990 117350 3040
rect 110240 2970 110300 2990
rect 110240 2930 110250 2970
rect 110290 2930 110300 2970
rect 117300 2970 117360 2990
rect 117300 2930 117310 2970
rect 117350 2930 117360 2970
rect 109320 2880 109350 2910
rect 109430 2900 110450 2930
rect 109430 2880 109460 2900
rect 109540 2880 109570 2900
rect 109650 2880 109680 2900
rect 109760 2880 109790 2900
rect 109870 2880 109900 2900
rect 109980 2880 110010 2900
rect 110090 2880 110120 2900
rect 110200 2880 110230 2900
rect 110310 2880 110340 2900
rect 110420 2880 110450 2900
rect 110530 2880 110560 2910
rect 117040 2880 117070 2910
rect 117150 2900 118170 2930
rect 117150 2880 117180 2900
rect 117260 2880 117290 2900
rect 117370 2880 117400 2900
rect 117480 2880 117510 2900
rect 117590 2880 117620 2900
rect 117700 2880 117730 2900
rect 117810 2880 117840 2900
rect 117920 2880 117950 2900
rect 118030 2880 118060 2900
rect 118140 2880 118170 2900
rect 118250 2880 118280 2910
rect 113380 2600 113440 2620
rect 112080 2580 112140 2600
rect 112080 2540 112090 2580
rect 112130 2550 112140 2580
rect 113380 2570 113390 2600
rect 113240 2560 113390 2570
rect 113430 2560 113440 2600
rect 112130 2540 112280 2550
rect 112080 2520 112280 2540
rect 112250 2490 112280 2520
rect 113240 2540 113440 2560
rect 113680 2600 113740 2620
rect 113680 2560 113690 2600
rect 113730 2570 113740 2600
rect 113860 2600 113920 2620
rect 113860 2570 113870 2600
rect 113730 2560 113760 2570
rect 113680 2540 113760 2560
rect 113240 2490 113270 2540
rect 112140 2440 112170 2470
rect 112250 2460 113270 2490
rect 112250 2440 112280 2460
rect 112360 2440 112390 2460
rect 112470 2440 112500 2460
rect 112580 2440 112610 2460
rect 112690 2440 112720 2460
rect 112800 2440 112830 2460
rect 112910 2440 112940 2460
rect 113020 2440 113050 2460
rect 113130 2440 113160 2460
rect 113240 2440 113270 2460
rect 113350 2440 113380 2470
rect 113620 2440 113650 2470
rect 113730 2440 113760 2540
rect 113840 2560 113870 2570
rect 113910 2560 113920 2600
rect 113840 2540 113920 2560
rect 114160 2600 114220 2620
rect 114160 2560 114170 2600
rect 114210 2570 114220 2600
rect 115460 2580 115520 2600
rect 114210 2560 114360 2570
rect 114160 2540 114360 2560
rect 115460 2550 115470 2580
rect 113840 2440 113870 2540
rect 114330 2490 114360 2540
rect 115320 2540 115470 2550
rect 115510 2540 115520 2580
rect 115320 2520 115520 2540
rect 115320 2490 115350 2520
rect 113950 2440 113980 2470
rect 114220 2440 114250 2470
rect 114330 2460 115350 2490
rect 114330 2440 114360 2460
rect 114440 2440 114470 2460
rect 114550 2440 114580 2460
rect 114660 2440 114690 2460
rect 114770 2440 114800 2460
rect 114880 2440 114910 2460
rect 114990 2440 115020 2460
rect 115100 2440 115130 2460
rect 115210 2440 115240 2460
rect 115320 2440 115350 2460
rect 115430 2440 115460 2470
rect 109320 2250 109350 2280
rect 109430 2250 109460 2280
rect 109540 2250 109570 2280
rect 109650 2250 109680 2280
rect 109760 2250 109790 2280
rect 109870 2250 109900 2280
rect 109980 2250 110010 2280
rect 110090 2250 110120 2280
rect 110200 2250 110230 2280
rect 110310 2250 110340 2280
rect 110420 2250 110450 2280
rect 110530 2250 110560 2280
rect 109250 2230 109350 2250
rect 109250 2190 109260 2230
rect 109300 2220 109350 2230
rect 110530 2230 110630 2250
rect 110530 2220 110580 2230
rect 109300 2190 109310 2220
rect 109250 2160 109310 2190
rect 110570 2190 110580 2220
rect 110620 2190 110630 2230
rect 110570 2160 110630 2190
rect 117040 2250 117070 2280
rect 117150 2250 117180 2280
rect 117260 2250 117290 2280
rect 117370 2250 117400 2280
rect 117480 2250 117510 2280
rect 117590 2250 117620 2280
rect 117700 2250 117730 2280
rect 117810 2250 117840 2280
rect 117920 2250 117950 2280
rect 118030 2250 118060 2280
rect 118140 2250 118170 2280
rect 118250 2250 118280 2280
rect 116970 2230 117070 2250
rect 116970 2190 116980 2230
rect 117020 2220 117070 2230
rect 118250 2230 118350 2250
rect 118250 2220 118300 2230
rect 117020 2190 117030 2220
rect 116970 2160 117030 2190
rect 118290 2190 118300 2220
rect 118340 2190 118350 2230
rect 118290 2170 118350 2190
rect 112140 2110 112170 2140
rect 112250 2110 112280 2140
rect 112360 2110 112390 2140
rect 112470 2110 112500 2140
rect 112580 2110 112610 2140
rect 112690 2110 112720 2140
rect 112800 2110 112830 2140
rect 112910 2110 112940 2140
rect 113020 2110 113050 2140
rect 113130 2110 113160 2140
rect 113240 2110 113270 2140
rect 113350 2110 113380 2140
rect 113620 2110 113650 2140
rect 113730 2110 113760 2140
rect 113840 2110 113870 2140
rect 113950 2110 113980 2140
rect 114220 2110 114250 2140
rect 114330 2110 114360 2140
rect 114440 2110 114470 2140
rect 114550 2110 114580 2140
rect 114660 2110 114690 2140
rect 114770 2110 114800 2140
rect 114880 2110 114910 2140
rect 114990 2110 115020 2140
rect 115100 2110 115130 2140
rect 115210 2110 115240 2140
rect 115320 2110 115350 2140
rect 115430 2110 115460 2140
rect 112070 2090 112170 2110
rect 112070 2050 112080 2090
rect 112120 2080 112170 2090
rect 113350 2090 113650 2110
rect 113350 2080 113480 2090
rect 112120 2050 112130 2080
rect 112070 2030 112130 2050
rect 113470 2050 113480 2080
rect 113520 2080 113650 2090
rect 113950 2090 114250 2110
rect 113950 2080 114080 2090
rect 113520 2050 113530 2080
rect 113470 2030 113530 2050
rect 114070 2050 114080 2080
rect 114120 2080 114250 2090
rect 115430 2090 115530 2110
rect 115430 2080 115480 2090
rect 114120 2050 114130 2080
rect 114070 2030 114130 2050
rect 115470 2050 115480 2080
rect 115520 2050 115530 2090
rect 115470 2030 115530 2050
rect 113650 1000 113730 1020
rect 113650 960 113670 1000
rect 113710 960 113730 1000
rect 113870 1000 113950 1020
rect 113870 960 113890 1000
rect 113930 960 113950 1000
rect 112520 910 112550 940
rect 112630 930 114750 960
rect 112630 910 112660 930
rect 112740 910 112770 930
rect 112850 910 112880 930
rect 112960 910 112990 930
rect 113070 910 113100 930
rect 113180 910 113210 930
rect 113290 910 113320 930
rect 113400 910 113430 930
rect 113510 910 113540 930
rect 113620 910 113650 930
rect 113730 910 113760 930
rect 113840 910 113870 930
rect 113950 910 113980 930
rect 114060 910 114090 930
rect 114170 910 114200 930
rect 114280 910 114310 930
rect 114390 910 114420 930
rect 114500 910 114530 930
rect 114610 910 114640 930
rect 114720 910 114750 930
rect 114830 910 114860 940
rect 114940 910 114970 940
rect 109600 760 109680 780
rect 109600 730 109620 760
rect 109580 720 109620 730
rect 109660 730 109680 760
rect 109800 760 109880 780
rect 109800 730 109820 760
rect 109660 720 109820 730
rect 109860 730 109880 760
rect 110000 760 110080 780
rect 110000 730 110020 760
rect 109860 720 110020 730
rect 110060 730 110080 760
rect 110200 760 110280 780
rect 110200 730 110220 760
rect 110060 720 110220 730
rect 110260 730 110280 760
rect 110260 720 110300 730
rect 109380 680 109500 710
rect 109580 700 110300 720
rect 109580 680 109700 700
rect 109780 680 109900 700
rect 109980 680 110100 700
rect 110180 680 110300 700
rect 110380 680 110500 710
rect 117320 760 117400 780
rect 117320 720 117340 760
rect 117380 720 117400 760
rect 117320 710 117400 720
rect 117520 760 117600 780
rect 117520 720 117540 760
rect 117580 720 117600 760
rect 117520 710 117600 720
rect 117720 760 117800 780
rect 117720 720 117740 760
rect 117780 720 117800 760
rect 117720 710 117800 720
rect 117920 760 118000 780
rect 117920 720 117940 760
rect 117980 720 118000 760
rect 117920 710 118000 720
rect 117100 680 117220 710
rect 117300 680 117420 710
rect 117500 680 117620 710
rect 117700 680 117820 710
rect 117900 680 118020 710
rect 118100 680 118220 710
rect 112520 380 112550 410
rect 112630 380 112660 410
rect 112740 380 112770 410
rect 112850 380 112880 410
rect 112960 380 112990 410
rect 113070 380 113100 410
rect 113180 380 113210 410
rect 113290 380 113320 410
rect 113400 380 113430 410
rect 113510 380 113540 410
rect 113620 380 113650 410
rect 113730 380 113760 410
rect 113840 380 113870 410
rect 113950 380 113980 410
rect 114060 380 114090 410
rect 114170 380 114200 410
rect 114280 380 114310 410
rect 114390 380 114420 410
rect 114500 380 114530 410
rect 114610 380 114640 410
rect 114720 380 114750 410
rect 112440 360 112550 380
rect 112440 320 112460 360
rect 112500 350 112550 360
rect 112500 320 112520 350
rect 112440 300 112520 320
rect 114830 0 114860 410
rect 114940 380 114970 410
rect 114940 360 115050 380
rect 114940 350 114990 360
rect 114970 320 114990 350
rect 115030 320 115050 360
rect 114970 300 115050 320
rect 114830 -20 114910 0
rect 114830 -60 114850 -20
rect 114890 -60 114910 -20
rect 114830 -80 114910 -60
rect 113190 -510 113270 -490
rect 113190 -550 113210 -510
rect 113250 -550 113270 -510
rect 114080 -510 114160 -490
rect 114080 -550 114100 -510
rect 114140 -550 114160 -510
rect 112940 -600 112970 -570
rect 113050 -580 113410 -550
rect 114080 -570 114160 -550
rect 113050 -600 113080 -580
rect 113160 -600 113190 -580
rect 113270 -600 113300 -580
rect 113380 -600 113410 -580
rect 113490 -600 113520 -570
rect 113820 -600 114420 -570
rect 109380 -750 109500 -720
rect 109580 -750 109700 -720
rect 109780 -750 109900 -720
rect 109980 -750 110100 -720
rect 110180 -750 110300 -720
rect 110380 -750 110500 -720
rect 109310 -770 109500 -750
rect 109310 -810 109320 -770
rect 109360 -780 109500 -770
rect 110380 -770 110570 -750
rect 110380 -780 110520 -770
rect 109360 -810 109370 -780
rect 109310 -830 109370 -810
rect 110510 -810 110520 -780
rect 110560 -810 110570 -770
rect 110510 -830 110570 -810
rect 117100 -750 117220 -720
rect 117300 -750 117420 -720
rect 117500 -750 117620 -720
rect 117700 -750 117820 -720
rect 117900 -750 118020 -720
rect 118100 -750 118220 -720
rect 117030 -770 117220 -750
rect 117030 -810 117040 -770
rect 117080 -780 117220 -770
rect 118100 -770 118290 -750
rect 118100 -780 118240 -770
rect 117080 -810 117090 -780
rect 117030 -830 117090 -810
rect 118230 -810 118240 -780
rect 118280 -810 118290 -770
rect 118230 -830 118290 -810
rect 112940 -930 112970 -900
rect 113050 -930 113080 -900
rect 113160 -930 113190 -900
rect 113270 -930 113300 -900
rect 113380 -930 113410 -900
rect 113490 -930 113520 -900
rect 113820 -930 114420 -900
rect 112870 -950 112970 -930
rect 112870 -990 112880 -950
rect 112920 -960 112970 -950
rect 113490 -950 113590 -930
rect 113490 -960 113540 -950
rect 112920 -990 112930 -960
rect 112870 -1010 112930 -990
rect 113530 -990 113540 -960
rect 113580 -990 113590 -950
rect 113530 -1010 113590 -990
rect 114080 -950 114160 -930
rect 114080 -990 114100 -950
rect 114140 -990 114160 -950
rect 114080 -1010 114160 -990
<< polycont >>
rect 112190 9810 112230 9850
rect 112550 9810 112590 9850
rect 114070 9810 114110 9850
rect 114430 9810 114470 9850
rect 115010 9810 115050 9850
rect 115370 9810 115410 9850
rect 113130 9470 113170 9510
rect 113490 9470 113530 9510
rect 112320 8910 112360 8950
rect 113270 8910 113310 8950
rect 114290 8910 114330 8950
rect 115162 8890 115202 8930
rect 112030 7810 112070 7850
rect 113470 7810 113510 7850
rect 114090 7810 114130 7850
rect 115530 7810 115570 7850
rect 116920 7810 116960 7850
rect 118360 7810 118400 7850
rect 116920 6970 116960 7010
rect 118360 6970 118400 7010
rect 109380 6890 109420 6930
rect 109500 6890 109540 6930
rect 109620 6890 109660 6930
rect 109740 6890 109780 6930
rect 109860 6890 109900 6930
rect 109980 6890 110020 6930
rect 110100 6890 110140 6930
rect 110220 6890 110260 6930
rect 110340 6890 110380 6930
rect 110460 6890 110500 6930
rect 112210 6890 112250 6930
rect 112330 6890 112370 6930
rect 112450 6890 112490 6930
rect 112570 6890 112610 6930
rect 112690 6890 112730 6930
rect 112810 6890 112850 6930
rect 112930 6890 112970 6930
rect 113050 6890 113090 6930
rect 113170 6890 113210 6930
rect 113290 6890 113330 6930
rect 114270 6890 114310 6930
rect 114390 6890 114430 6930
rect 114510 6890 114550 6930
rect 114630 6890 114670 6930
rect 114750 6890 114790 6930
rect 114870 6890 114910 6930
rect 114990 6890 115030 6930
rect 115110 6890 115150 6930
rect 115230 6890 115270 6930
rect 115350 6890 115390 6930
rect 117100 6890 117140 6930
rect 117220 6890 117260 6930
rect 117340 6890 117380 6930
rect 117460 6890 117500 6930
rect 117580 6890 117620 6930
rect 117700 6890 117740 6930
rect 117820 6890 117860 6930
rect 117940 6890 117980 6930
rect 118060 6890 118100 6930
rect 118180 6890 118220 6930
rect 113040 6500 113080 6540
rect 109260 6360 109300 6400
rect 110580 6360 110620 6400
rect 113700 6500 113740 6540
rect 113860 6500 113900 6540
rect 114520 6500 114560 6540
rect 116980 6360 117020 6400
rect 118300 6360 118340 6400
rect 113224 5750 113264 5790
rect 113370 5750 113410 5790
rect 113516 5750 113556 5790
rect 114044 5750 114084 5790
rect 114190 5750 114230 5790
rect 114336 5750 114376 5790
rect 113720 5180 113760 5220
rect 109920 5020 109960 5060
rect 109920 4890 109960 4930
rect 109920 4810 109960 4850
rect 109920 4730 109960 4770
rect 117640 5020 117680 5060
rect 117640 4890 117680 4930
rect 117640 4810 117680 4850
rect 117640 4730 117680 4770
rect 113560 4540 113600 4580
rect 114000 4540 114040 4580
rect 109260 3810 109300 3850
rect 110580 3810 110620 3850
rect 112245 3860 112285 3900
rect 112355 3860 112395 3900
rect 112465 3860 112505 3900
rect 112575 3860 112615 3900
rect 112685 3860 112725 3900
rect 112795 3860 112835 3900
rect 112905 3860 112945 3900
rect 113015 3860 113055 3900
rect 113125 3860 113165 3900
rect 113235 3860 113275 3900
rect 114325 3860 114365 3900
rect 114435 3860 114475 3900
rect 114545 3860 114585 3900
rect 114655 3860 114695 3900
rect 114765 3860 114805 3900
rect 114875 3860 114915 3900
rect 114985 3860 115025 3900
rect 115095 3860 115135 3900
rect 115205 3860 115245 3900
rect 115315 3860 115355 3900
rect 116980 3810 117020 3850
rect 118300 3810 118340 3850
rect 112080 3420 112120 3460
rect 113400 3420 113440 3460
rect 114160 3420 114200 3460
rect 115480 3420 115520 3460
rect 110250 3270 110290 3310
rect 117310 3270 117350 3310
rect 110250 3140 110290 3180
rect 110250 3060 110290 3100
rect 117310 3140 117350 3180
rect 117310 3060 117350 3100
rect 110250 2930 110290 2970
rect 117310 2930 117350 2970
rect 112090 2540 112130 2580
rect 113390 2560 113430 2600
rect 113690 2560 113730 2600
rect 113870 2560 113910 2600
rect 114170 2560 114210 2600
rect 115470 2540 115510 2580
rect 109260 2190 109300 2230
rect 110580 2190 110620 2230
rect 116980 2190 117020 2230
rect 118300 2190 118340 2230
rect 112080 2050 112120 2090
rect 113480 2050 113520 2090
rect 114080 2050 114120 2090
rect 115480 2050 115520 2090
rect 113670 960 113710 1000
rect 113890 960 113930 1000
rect 109620 720 109660 760
rect 109820 720 109860 760
rect 110020 720 110060 760
rect 110220 720 110260 760
rect 117340 720 117380 760
rect 117540 720 117580 760
rect 117740 720 117780 760
rect 117940 720 117980 760
rect 112460 320 112500 360
rect 114990 320 115030 360
rect 114850 -60 114890 -20
rect 113210 -550 113250 -510
rect 114100 -550 114140 -510
rect 109320 -810 109360 -770
rect 110520 -810 110560 -770
rect 117040 -810 117080 -770
rect 118240 -810 118280 -770
rect 112880 -990 112920 -950
rect 113540 -990 113580 -950
rect 114100 -990 114140 -950
<< xpolycontact >>
rect 108408 5880 108690 6320
rect 108408 5190 108690 5630
rect 118910 5880 119192 6320
rect 118910 5190 119192 5630
rect 108510 3088 108580 3528
rect 108510 2330 108580 2770
rect 108630 3088 108700 3528
rect 108630 2330 108700 2770
rect 108750 3088 108820 3528
rect 108750 2330 108820 2770
rect 108870 3088 108940 3528
rect 118660 3088 118730 3528
rect 108870 2330 108940 2770
rect 118660 2330 118730 2770
rect 118780 3088 118850 3528
rect 118780 2330 118850 2770
rect 118900 3088 118970 3528
rect 118900 2330 118970 2770
rect 119020 3088 119090 3528
rect 119020 2330 119090 2770
rect 108650 140 108720 580
rect 108650 -794 108720 -354
rect 108770 140 108840 580
rect 108770 -794 108840 -354
rect 118760 140 118830 580
rect 118760 -794 118830 -354
rect 118880 140 118950 580
rect 118880 -794 118950 -354
<< ppolyres >>
rect 108408 5630 108690 5880
rect 118910 5630 119192 5880
<< xpolyres >>
rect 108510 2770 108580 3088
rect 108630 2770 108700 3088
rect 108750 2770 108820 3088
rect 108870 2770 108940 3088
rect 118660 2770 118730 3088
rect 118780 2770 118850 3088
rect 118900 2770 118970 3088
rect 119020 2770 119090 3088
rect 108650 -354 108720 140
rect 108770 -354 108840 140
rect 118760 -354 118830 140
rect 118880 -354 118950 140
<< locali >>
rect 112170 9850 112250 9870
rect 112170 9810 112190 9850
rect 112230 9810 112250 9850
rect 112170 9790 112250 9810
rect 112530 9850 112610 9870
rect 112530 9810 112550 9850
rect 112590 9810 112610 9850
rect 112530 9790 112610 9810
rect 114050 9850 114130 9870
rect 114050 9810 114070 9850
rect 114110 9810 114130 9850
rect 114050 9790 114130 9810
rect 114410 9850 114490 9870
rect 114410 9810 114430 9850
rect 114470 9810 114490 9850
rect 114410 9790 114490 9810
rect 114990 9850 115070 9870
rect 114990 9810 115010 9850
rect 115050 9810 115070 9850
rect 114990 9790 115070 9810
rect 115350 9850 115430 9870
rect 115350 9810 115370 9850
rect 115410 9810 115430 9850
rect 115350 9790 115430 9810
rect 112100 9730 112240 9750
rect 112100 9090 112110 9730
rect 112150 9090 112190 9730
rect 112230 9090 112240 9730
rect 112100 9070 112240 9090
rect 112300 9730 112360 9750
rect 112300 9090 112310 9730
rect 112350 9090 112360 9730
rect 112300 9070 112360 9090
rect 112420 9730 112480 9750
rect 112420 9090 112430 9730
rect 112470 9090 112480 9730
rect 112420 9070 112480 9090
rect 112540 9730 112680 9750
rect 112540 9090 112550 9730
rect 112590 9090 112630 9730
rect 112670 9090 112680 9730
rect 113980 9730 114120 9750
rect 113110 9510 113190 9530
rect 113110 9470 113130 9510
rect 113170 9470 113190 9510
rect 113110 9450 113190 9470
rect 113470 9510 113550 9530
rect 113470 9470 113490 9510
rect 113530 9470 113550 9510
rect 113470 9450 113550 9470
rect 112540 9070 112680 9090
rect 113040 9390 113180 9410
rect 113040 9090 113050 9390
rect 113090 9090 113130 9390
rect 113170 9090 113180 9390
rect 113040 9070 113180 9090
rect 113240 9390 113300 9410
rect 113240 9090 113250 9390
rect 113290 9090 113300 9390
rect 113240 9070 113300 9090
rect 113360 9390 113420 9410
rect 113360 9090 113370 9390
rect 113410 9090 113420 9390
rect 113360 9070 113420 9090
rect 113480 9390 113620 9410
rect 113480 9090 113490 9390
rect 113530 9090 113570 9390
rect 113610 9090 113620 9390
rect 113480 9070 113620 9090
rect 113980 9090 113990 9730
rect 114030 9090 114070 9730
rect 114110 9090 114120 9730
rect 113980 9070 114120 9090
rect 114180 9730 114240 9750
rect 114180 9090 114190 9730
rect 114230 9090 114240 9730
rect 114180 9070 114240 9090
rect 114300 9730 114360 9750
rect 114300 9090 114310 9730
rect 114350 9090 114360 9730
rect 114300 9070 114360 9090
rect 114420 9730 114560 9750
rect 114420 9090 114430 9730
rect 114470 9090 114510 9730
rect 114550 9090 114560 9730
rect 114420 9070 114560 9090
rect 114920 9730 115060 9750
rect 114920 9090 114930 9730
rect 114970 9090 115010 9730
rect 115050 9090 115060 9730
rect 114920 9070 115060 9090
rect 115120 9730 115180 9750
rect 115120 9090 115130 9730
rect 115170 9090 115180 9730
rect 115120 9070 115180 9090
rect 115240 9730 115300 9750
rect 115240 9090 115250 9730
rect 115290 9090 115300 9730
rect 115240 9070 115300 9090
rect 115360 9730 115500 9750
rect 115360 9090 115370 9730
rect 115410 9090 115450 9730
rect 115490 9090 115500 9730
rect 115360 9070 115500 9090
rect 112300 8950 112380 8970
rect 112300 8910 112320 8950
rect 112360 8910 112380 8950
rect 112300 8890 112380 8910
rect 113260 8950 113320 8970
rect 113260 8910 113270 8950
rect 113310 8910 113320 8950
rect 113260 8890 113320 8910
rect 114280 8950 114340 8970
rect 114280 8910 114290 8950
rect 114330 8910 114340 8950
rect 114280 8890 114340 8910
rect 115152 8930 115212 8950
rect 115152 8890 115162 8930
rect 115202 8890 115212 8930
rect 115152 8870 115212 8890
rect 112020 7850 112080 7870
rect 112020 7810 112030 7850
rect 112070 7810 112080 7850
rect 112020 7790 112080 7810
rect 113460 7850 113520 7870
rect 113460 7810 113470 7850
rect 113510 7810 113520 7850
rect 113460 7790 113520 7810
rect 114080 7850 114140 7870
rect 114080 7810 114090 7850
rect 114130 7810 114140 7850
rect 114080 7790 114140 7810
rect 115520 7850 115580 7870
rect 115520 7810 115530 7850
rect 115570 7810 115580 7850
rect 115520 7790 115580 7810
rect 116900 7850 116980 7870
rect 116900 7810 116920 7850
rect 116960 7810 116980 7850
rect 116900 7790 116980 7810
rect 118340 7850 118420 7870
rect 118340 7810 118360 7850
rect 118400 7810 118420 7850
rect 118340 7790 118420 7810
rect 109110 7730 109250 7750
rect 109110 7090 109120 7730
rect 109160 7090 109200 7730
rect 109240 7090 109250 7730
rect 109110 7070 109250 7090
rect 109310 7730 109370 7750
rect 109310 7090 109320 7730
rect 109360 7090 109370 7730
rect 109310 7070 109370 7090
rect 109430 7730 109490 7750
rect 109430 7090 109440 7730
rect 109480 7090 109490 7730
rect 109430 7070 109490 7090
rect 109550 7730 109610 7750
rect 109550 7090 109560 7730
rect 109600 7090 109610 7730
rect 109550 7070 109610 7090
rect 109670 7730 109730 7750
rect 109670 7090 109680 7730
rect 109720 7090 109730 7730
rect 109670 7070 109730 7090
rect 109790 7730 109850 7750
rect 109790 7090 109800 7730
rect 109840 7090 109850 7730
rect 109790 7070 109850 7090
rect 109910 7730 109970 7750
rect 109910 7090 109920 7730
rect 109960 7090 109970 7730
rect 109910 7070 109970 7090
rect 110030 7730 110090 7750
rect 110030 7090 110040 7730
rect 110080 7090 110090 7730
rect 110030 7070 110090 7090
rect 110150 7730 110210 7750
rect 110150 7090 110160 7730
rect 110200 7090 110210 7730
rect 110150 7070 110210 7090
rect 110270 7730 110330 7750
rect 110270 7090 110280 7730
rect 110320 7090 110330 7730
rect 110270 7070 110330 7090
rect 110390 7730 110450 7750
rect 110390 7090 110400 7730
rect 110440 7090 110450 7730
rect 110390 7070 110450 7090
rect 110510 7730 110570 7750
rect 110510 7090 110520 7730
rect 110560 7090 110570 7730
rect 110510 7070 110570 7090
rect 110630 7730 110770 7750
rect 110630 7090 110640 7730
rect 110680 7090 110720 7730
rect 110760 7090 110770 7730
rect 110630 7070 110770 7090
rect 111940 7730 112080 7750
rect 111940 7090 111950 7730
rect 111990 7090 112030 7730
rect 112070 7090 112080 7730
rect 111940 7070 112080 7090
rect 112140 7730 112200 7750
rect 112140 7090 112150 7730
rect 112190 7090 112200 7730
rect 112140 7070 112200 7090
rect 112260 7730 112320 7750
rect 112260 7090 112270 7730
rect 112310 7090 112320 7730
rect 112260 7070 112320 7090
rect 112380 7730 112440 7750
rect 112380 7090 112390 7730
rect 112430 7090 112440 7730
rect 112380 7070 112440 7090
rect 112500 7730 112560 7750
rect 112500 7090 112510 7730
rect 112550 7090 112560 7730
rect 112500 7070 112560 7090
rect 112620 7730 112680 7750
rect 112620 7090 112630 7730
rect 112670 7090 112680 7730
rect 112620 7070 112680 7090
rect 112740 7730 112800 7750
rect 112740 7090 112750 7730
rect 112790 7090 112800 7730
rect 112740 7070 112800 7090
rect 112860 7730 112920 7750
rect 112860 7090 112870 7730
rect 112910 7090 112920 7730
rect 112860 7070 112920 7090
rect 112980 7730 113040 7750
rect 112980 7090 112990 7730
rect 113030 7090 113040 7730
rect 112980 7070 113040 7090
rect 113100 7730 113160 7750
rect 113100 7090 113110 7730
rect 113150 7090 113160 7730
rect 113100 7070 113160 7090
rect 113220 7730 113280 7750
rect 113220 7090 113230 7730
rect 113270 7090 113280 7730
rect 113220 7070 113280 7090
rect 113340 7730 113400 7750
rect 113340 7090 113350 7730
rect 113390 7090 113400 7730
rect 113340 7070 113400 7090
rect 113460 7730 113600 7750
rect 113460 7090 113470 7730
rect 113510 7090 113550 7730
rect 113590 7090 113600 7730
rect 113460 7070 113600 7090
rect 114000 7730 114140 7750
rect 114000 7090 114010 7730
rect 114050 7090 114090 7730
rect 114130 7090 114140 7730
rect 114000 7070 114140 7090
rect 114200 7730 114260 7750
rect 114200 7090 114210 7730
rect 114250 7090 114260 7730
rect 114200 7070 114260 7090
rect 114320 7730 114380 7750
rect 114320 7090 114330 7730
rect 114370 7090 114380 7730
rect 114320 7070 114380 7090
rect 114440 7730 114500 7750
rect 114440 7090 114450 7730
rect 114490 7090 114500 7730
rect 114440 7070 114500 7090
rect 114560 7730 114620 7750
rect 114560 7090 114570 7730
rect 114610 7090 114620 7730
rect 114560 7070 114620 7090
rect 114680 7730 114740 7750
rect 114680 7090 114690 7730
rect 114730 7090 114740 7730
rect 114680 7070 114740 7090
rect 114800 7730 114860 7750
rect 114800 7090 114810 7730
rect 114850 7090 114860 7730
rect 114800 7070 114860 7090
rect 114920 7730 114980 7750
rect 114920 7090 114930 7730
rect 114970 7090 114980 7730
rect 114920 7070 114980 7090
rect 115040 7730 115100 7750
rect 115040 7090 115050 7730
rect 115090 7090 115100 7730
rect 115040 7070 115100 7090
rect 115160 7730 115220 7750
rect 115160 7090 115170 7730
rect 115210 7090 115220 7730
rect 115160 7070 115220 7090
rect 115280 7730 115340 7750
rect 115280 7090 115290 7730
rect 115330 7090 115340 7730
rect 115280 7070 115340 7090
rect 115400 7730 115460 7750
rect 115400 7090 115410 7730
rect 115450 7090 115460 7730
rect 115400 7070 115460 7090
rect 115520 7730 115660 7750
rect 115520 7090 115530 7730
rect 115570 7090 115610 7730
rect 115650 7090 115660 7730
rect 115520 7070 115660 7090
rect 116830 7730 116970 7750
rect 116830 7090 116840 7730
rect 116880 7090 116920 7730
rect 116960 7090 116970 7730
rect 116830 7070 116970 7090
rect 117030 7730 117090 7750
rect 117030 7090 117040 7730
rect 117080 7090 117090 7730
rect 117030 7070 117090 7090
rect 117150 7730 117210 7750
rect 117150 7090 117160 7730
rect 117200 7090 117210 7730
rect 117150 7070 117210 7090
rect 117270 7730 117330 7750
rect 117270 7090 117280 7730
rect 117320 7090 117330 7730
rect 117270 7070 117330 7090
rect 117390 7730 117450 7750
rect 117390 7090 117400 7730
rect 117440 7090 117450 7730
rect 117390 7070 117450 7090
rect 117510 7730 117570 7750
rect 117510 7090 117520 7730
rect 117560 7090 117570 7730
rect 117510 7070 117570 7090
rect 117630 7730 117690 7750
rect 117630 7090 117640 7730
rect 117680 7090 117690 7730
rect 117630 7070 117690 7090
rect 117750 7730 117810 7750
rect 117750 7090 117760 7730
rect 117800 7090 117810 7730
rect 117750 7070 117810 7090
rect 117870 7730 117930 7750
rect 117870 7090 117880 7730
rect 117920 7090 117930 7730
rect 117870 7070 117930 7090
rect 117990 7730 118050 7750
rect 117990 7090 118000 7730
rect 118040 7090 118050 7730
rect 117990 7070 118050 7090
rect 118110 7730 118170 7750
rect 118110 7090 118120 7730
rect 118160 7090 118170 7730
rect 118110 7070 118170 7090
rect 118230 7730 118290 7750
rect 118230 7090 118240 7730
rect 118280 7090 118290 7730
rect 118230 7070 118290 7090
rect 118350 7730 118490 7750
rect 118350 7090 118360 7730
rect 118400 7090 118440 7730
rect 118480 7090 118490 7730
rect 118350 7070 118490 7090
rect 116910 7010 116970 7030
rect 116910 6970 116920 7010
rect 116960 6970 116970 7010
rect 116910 6950 116970 6970
rect 118350 7010 118410 7030
rect 118350 6970 118360 7010
rect 118400 6970 118410 7010
rect 118350 6950 118410 6970
rect 109370 6930 109430 6950
rect 109370 6890 109380 6930
rect 109420 6890 109430 6930
rect 109370 6870 109430 6890
rect 109490 6930 109550 6950
rect 109490 6890 109500 6930
rect 109540 6890 109550 6930
rect 109490 6870 109550 6890
rect 109610 6930 109670 6950
rect 109610 6890 109620 6930
rect 109660 6890 109670 6930
rect 109610 6870 109670 6890
rect 109730 6930 109790 6950
rect 109730 6890 109740 6930
rect 109780 6890 109790 6930
rect 109730 6870 109790 6890
rect 109850 6930 109910 6950
rect 109850 6890 109860 6930
rect 109900 6890 109910 6930
rect 109850 6870 109910 6890
rect 109970 6930 110030 6950
rect 109970 6890 109980 6930
rect 110020 6890 110030 6930
rect 109970 6870 110030 6890
rect 110090 6930 110150 6950
rect 110090 6890 110100 6930
rect 110140 6890 110150 6930
rect 110090 6870 110150 6890
rect 110210 6930 110270 6950
rect 110210 6890 110220 6930
rect 110260 6890 110270 6930
rect 110210 6870 110270 6890
rect 110330 6930 110390 6950
rect 110330 6890 110340 6930
rect 110380 6890 110390 6930
rect 110330 6870 110390 6890
rect 110450 6930 110510 6950
rect 110450 6890 110460 6930
rect 110500 6890 110510 6930
rect 110450 6870 110510 6890
rect 112200 6930 112260 6950
rect 112200 6890 112210 6930
rect 112250 6890 112260 6930
rect 112200 6870 112260 6890
rect 112320 6930 112380 6950
rect 112320 6890 112330 6930
rect 112370 6890 112380 6930
rect 112320 6870 112380 6890
rect 112440 6930 112500 6950
rect 112440 6890 112450 6930
rect 112490 6890 112500 6930
rect 112440 6870 112500 6890
rect 112560 6930 112620 6950
rect 112560 6890 112570 6930
rect 112610 6890 112620 6930
rect 112560 6870 112620 6890
rect 112680 6930 112740 6950
rect 112680 6890 112690 6930
rect 112730 6890 112740 6930
rect 112680 6870 112740 6890
rect 112800 6930 112860 6950
rect 112800 6890 112810 6930
rect 112850 6890 112860 6930
rect 112800 6870 112860 6890
rect 112920 6930 112980 6950
rect 112920 6890 112930 6930
rect 112970 6890 112980 6930
rect 112920 6870 112980 6890
rect 113040 6930 113100 6950
rect 113040 6890 113050 6930
rect 113090 6890 113100 6930
rect 113040 6870 113100 6890
rect 113160 6930 113220 6950
rect 113160 6890 113170 6930
rect 113210 6890 113220 6930
rect 113160 6870 113220 6890
rect 113280 6930 113340 6950
rect 113280 6890 113290 6930
rect 113330 6890 113340 6930
rect 113280 6870 113340 6890
rect 114260 6930 114320 6950
rect 114260 6890 114270 6930
rect 114310 6890 114320 6930
rect 114260 6870 114320 6890
rect 114380 6930 114440 6950
rect 114380 6890 114390 6930
rect 114430 6890 114440 6930
rect 114380 6870 114440 6890
rect 114500 6930 114560 6950
rect 114500 6890 114510 6930
rect 114550 6890 114560 6930
rect 114500 6870 114560 6890
rect 114620 6930 114680 6950
rect 114620 6890 114630 6930
rect 114670 6890 114680 6930
rect 114620 6870 114680 6890
rect 114740 6930 114800 6950
rect 114740 6890 114750 6930
rect 114790 6890 114800 6930
rect 114740 6870 114800 6890
rect 114860 6930 114920 6950
rect 114860 6890 114870 6930
rect 114910 6890 114920 6930
rect 114860 6870 114920 6890
rect 114980 6930 115040 6950
rect 114980 6890 114990 6930
rect 115030 6890 115040 6930
rect 114980 6870 115040 6890
rect 115100 6930 115160 6950
rect 115100 6890 115110 6930
rect 115150 6890 115160 6930
rect 115100 6870 115160 6890
rect 115220 6930 115280 6950
rect 115220 6890 115230 6930
rect 115270 6890 115280 6930
rect 115220 6870 115280 6890
rect 115340 6930 115400 6950
rect 115340 6890 115350 6930
rect 115390 6890 115400 6930
rect 115340 6870 115400 6890
rect 117090 6930 117150 6950
rect 117090 6890 117100 6930
rect 117140 6890 117150 6930
rect 117090 6870 117150 6890
rect 117210 6930 117270 6950
rect 117210 6890 117220 6930
rect 117260 6890 117270 6930
rect 117210 6870 117270 6890
rect 117330 6930 117390 6950
rect 117330 6890 117340 6930
rect 117380 6890 117390 6930
rect 117330 6870 117390 6890
rect 117450 6930 117510 6950
rect 117450 6890 117460 6930
rect 117500 6890 117510 6930
rect 117450 6870 117510 6890
rect 117570 6930 117630 6950
rect 117570 6890 117580 6930
rect 117620 6890 117630 6930
rect 117570 6870 117630 6890
rect 117690 6930 117750 6950
rect 117690 6890 117700 6930
rect 117740 6890 117750 6930
rect 117690 6870 117750 6890
rect 117810 6930 117870 6950
rect 117810 6890 117820 6930
rect 117860 6890 117870 6930
rect 117810 6870 117870 6890
rect 117930 6930 117990 6950
rect 117930 6890 117940 6930
rect 117980 6890 117990 6930
rect 117930 6870 117990 6890
rect 118050 6930 118110 6950
rect 118050 6890 118060 6930
rect 118100 6890 118110 6930
rect 118050 6870 118110 6890
rect 118170 6930 118230 6950
rect 118170 6890 118180 6930
rect 118220 6890 118230 6930
rect 118170 6870 118230 6890
rect 113020 6540 113100 6560
rect 113020 6500 113040 6540
rect 113080 6500 113100 6540
rect 113020 6480 113100 6500
rect 113360 6540 113420 6560
rect 113360 6500 113370 6540
rect 113410 6500 113420 6540
rect 113360 6480 113420 6500
rect 113680 6540 113760 6560
rect 113680 6500 113700 6540
rect 113740 6500 113760 6540
rect 113680 6480 113760 6500
rect 113840 6540 113920 6560
rect 113840 6500 113860 6540
rect 113900 6500 113920 6540
rect 113840 6480 113920 6500
rect 114180 6540 114240 6560
rect 114180 6500 114190 6540
rect 114230 6500 114240 6540
rect 114180 6480 114240 6500
rect 114500 6540 114580 6560
rect 114500 6500 114520 6540
rect 114560 6500 114580 6540
rect 114500 6480 114580 6500
rect 109250 6400 109310 6420
rect 108408 6380 108690 6400
rect 108408 6340 108420 6380
rect 108460 6340 108530 6380
rect 108570 6340 108640 6380
rect 108680 6340 108690 6380
rect 109250 6360 109260 6400
rect 109300 6360 109310 6400
rect 109250 6340 109310 6360
rect 110570 6400 110630 6420
rect 110570 6360 110580 6400
rect 110620 6360 110630 6400
rect 110570 6340 110630 6360
rect 108408 6320 108690 6340
rect 113040 6330 113080 6480
rect 113240 6430 113320 6450
rect 113240 6390 113260 6430
rect 113300 6390 113320 6430
rect 113240 6370 113320 6390
rect 113260 6330 113300 6370
rect 113370 6330 113410 6480
rect 113460 6430 113540 6450
rect 113460 6390 113480 6430
rect 113520 6390 113540 6430
rect 113460 6370 113540 6390
rect 113480 6330 113520 6370
rect 113700 6330 113740 6480
rect 113860 6330 113900 6480
rect 114060 6430 114140 6450
rect 114060 6390 114080 6430
rect 114120 6390 114140 6430
rect 114060 6370 114140 6390
rect 114080 6330 114120 6370
rect 114190 6330 114230 6480
rect 114280 6430 114360 6450
rect 114280 6390 114300 6430
rect 114340 6390 114360 6430
rect 114280 6370 114360 6390
rect 114300 6330 114340 6370
rect 114520 6330 114560 6480
rect 116970 6400 117030 6420
rect 116970 6360 116980 6400
rect 117020 6360 117030 6400
rect 116970 6340 117030 6360
rect 118290 6400 118350 6420
rect 118290 6360 118300 6400
rect 118340 6360 118350 6400
rect 118290 6340 118350 6360
rect 118910 6380 119192 6400
rect 118910 6340 118920 6380
rect 118960 6340 119030 6380
rect 119070 6340 119140 6380
rect 119180 6340 119192 6380
rect 112950 6310 113090 6330
rect 109170 6280 109310 6300
rect 108408 5170 108690 5190
rect 108408 5130 108420 5170
rect 108460 5130 108530 5170
rect 108570 5130 108640 5170
rect 108680 5130 108690 5170
rect 108408 5110 108690 5130
rect 109170 5140 109180 6280
rect 109220 5140 109260 6280
rect 109300 5140 109310 6280
rect 109170 5120 109310 5140
rect 109360 6280 109420 6300
rect 109360 5140 109370 6280
rect 109410 5140 109420 6280
rect 109360 5120 109420 5140
rect 109470 6280 109530 6300
rect 109470 5140 109480 6280
rect 109520 5140 109530 6280
rect 109470 5120 109530 5140
rect 109580 6280 109640 6300
rect 109580 5140 109590 6280
rect 109630 5140 109640 6280
rect 109580 5120 109640 5140
rect 109690 6280 109750 6300
rect 109690 5140 109700 6280
rect 109740 5140 109750 6280
rect 109690 5120 109750 5140
rect 109800 6280 109860 6300
rect 109800 5140 109810 6280
rect 109850 5140 109860 6280
rect 109800 5120 109860 5140
rect 109910 6280 109970 6300
rect 109910 5140 109920 6280
rect 109960 5140 109970 6280
rect 109910 5120 109970 5140
rect 110020 6280 110080 6300
rect 110020 5140 110030 6280
rect 110070 5140 110080 6280
rect 110020 5120 110080 5140
rect 110130 6280 110190 6300
rect 110130 5140 110140 6280
rect 110180 5140 110190 6280
rect 110130 5120 110190 5140
rect 110240 6280 110300 6300
rect 110240 5140 110250 6280
rect 110290 5140 110300 6280
rect 110240 5120 110300 5140
rect 110350 6280 110410 6300
rect 110350 5140 110360 6280
rect 110400 5140 110410 6280
rect 110350 5120 110410 5140
rect 110460 6280 110520 6300
rect 110460 5140 110470 6280
rect 110510 5140 110520 6280
rect 110460 5120 110520 5140
rect 110570 6280 110710 6300
rect 110570 5140 110580 6280
rect 110620 5140 110660 6280
rect 110700 5140 110710 6280
rect 112950 6270 112960 6310
rect 113000 6270 113040 6310
rect 113080 6270 113090 6310
rect 112950 6210 113090 6270
rect 112950 6170 112960 6210
rect 113000 6170 113040 6210
rect 113080 6170 113090 6210
rect 112950 6110 113090 6170
rect 112950 6070 112960 6110
rect 113000 6070 113040 6110
rect 113080 6070 113090 6110
rect 112950 6010 113090 6070
rect 112950 5970 112960 6010
rect 113000 5970 113040 6010
rect 113080 5970 113090 6010
rect 112950 5910 113090 5970
rect 112950 5870 112960 5910
rect 113000 5870 113040 5910
rect 113080 5870 113090 5910
rect 112950 5850 113090 5870
rect 113140 6310 113200 6330
rect 113140 6270 113150 6310
rect 113190 6270 113200 6310
rect 113140 6210 113200 6270
rect 113140 6170 113150 6210
rect 113190 6170 113200 6210
rect 113140 6110 113200 6170
rect 113140 6070 113150 6110
rect 113190 6070 113200 6110
rect 113140 6010 113200 6070
rect 113140 5970 113150 6010
rect 113190 5970 113200 6010
rect 113140 5910 113200 5970
rect 113140 5870 113150 5910
rect 113190 5870 113200 5910
rect 113140 5850 113200 5870
rect 113250 6310 113310 6330
rect 113250 6270 113260 6310
rect 113300 6270 113310 6310
rect 113250 6210 113310 6270
rect 113250 6170 113260 6210
rect 113300 6170 113310 6210
rect 113250 6110 113310 6170
rect 113250 6070 113260 6110
rect 113300 6070 113310 6110
rect 113250 6010 113310 6070
rect 113250 5970 113260 6010
rect 113300 5970 113310 6010
rect 113250 5910 113310 5970
rect 113250 5870 113260 5910
rect 113300 5870 113310 5910
rect 113250 5850 113310 5870
rect 113360 6310 113420 6330
rect 113360 6270 113370 6310
rect 113410 6270 113420 6310
rect 113360 6210 113420 6270
rect 113360 6170 113370 6210
rect 113410 6170 113420 6210
rect 113360 6110 113420 6170
rect 113360 6070 113370 6110
rect 113410 6070 113420 6110
rect 113360 6010 113420 6070
rect 113360 5970 113370 6010
rect 113410 5970 113420 6010
rect 113360 5910 113420 5970
rect 113360 5870 113370 5910
rect 113410 5870 113420 5910
rect 113360 5850 113420 5870
rect 113470 6310 113530 6330
rect 113470 6270 113480 6310
rect 113520 6270 113530 6310
rect 113470 6210 113530 6270
rect 113470 6170 113480 6210
rect 113520 6170 113530 6210
rect 113470 6110 113530 6170
rect 113470 6070 113480 6110
rect 113520 6070 113530 6110
rect 113470 6010 113530 6070
rect 113470 5970 113480 6010
rect 113520 5970 113530 6010
rect 113470 5910 113530 5970
rect 113470 5870 113480 5910
rect 113520 5870 113530 5910
rect 113470 5850 113530 5870
rect 113580 6310 113640 6330
rect 113580 6270 113590 6310
rect 113630 6270 113640 6310
rect 113580 6210 113640 6270
rect 113580 6170 113590 6210
rect 113630 6170 113640 6210
rect 113580 6110 113640 6170
rect 113580 6070 113590 6110
rect 113630 6070 113640 6110
rect 113580 6010 113640 6070
rect 113580 5970 113590 6010
rect 113630 5970 113640 6010
rect 113580 5910 113640 5970
rect 113580 5870 113590 5910
rect 113630 5870 113640 5910
rect 113580 5850 113640 5870
rect 113690 6310 113910 6330
rect 113690 6270 113700 6310
rect 113740 6270 113780 6310
rect 113820 6270 113860 6310
rect 113900 6270 113910 6310
rect 113690 6210 113910 6270
rect 113690 6170 113700 6210
rect 113740 6170 113780 6210
rect 113820 6170 113860 6210
rect 113900 6170 113910 6210
rect 113690 6110 113910 6170
rect 113690 6070 113700 6110
rect 113740 6070 113780 6110
rect 113820 6070 113860 6110
rect 113900 6070 113910 6110
rect 113690 6010 113910 6070
rect 113690 5970 113700 6010
rect 113740 5970 113780 6010
rect 113820 5970 113860 6010
rect 113900 5970 113910 6010
rect 113690 5910 113910 5970
rect 113690 5870 113700 5910
rect 113740 5870 113780 5910
rect 113820 5870 113860 5910
rect 113900 5870 113910 5910
rect 113690 5850 113910 5870
rect 113960 6310 114020 6330
rect 113960 6270 113970 6310
rect 114010 6270 114020 6310
rect 113960 6210 114020 6270
rect 113960 6170 113970 6210
rect 114010 6170 114020 6210
rect 113960 6110 114020 6170
rect 113960 6070 113970 6110
rect 114010 6070 114020 6110
rect 113960 6010 114020 6070
rect 113960 5970 113970 6010
rect 114010 5970 114020 6010
rect 113960 5910 114020 5970
rect 113960 5870 113970 5910
rect 114010 5870 114020 5910
rect 113960 5850 114020 5870
rect 114070 6310 114130 6330
rect 114070 6270 114080 6310
rect 114120 6270 114130 6310
rect 114070 6210 114130 6270
rect 114070 6170 114080 6210
rect 114120 6170 114130 6210
rect 114070 6110 114130 6170
rect 114070 6070 114080 6110
rect 114120 6070 114130 6110
rect 114070 6010 114130 6070
rect 114070 5970 114080 6010
rect 114120 5970 114130 6010
rect 114070 5910 114130 5970
rect 114070 5870 114080 5910
rect 114120 5870 114130 5910
rect 114070 5850 114130 5870
rect 114180 6310 114240 6330
rect 114180 6270 114190 6310
rect 114230 6270 114240 6310
rect 114180 6210 114240 6270
rect 114180 6170 114190 6210
rect 114230 6170 114240 6210
rect 114180 6110 114240 6170
rect 114180 6070 114190 6110
rect 114230 6070 114240 6110
rect 114180 6010 114240 6070
rect 114180 5970 114190 6010
rect 114230 5970 114240 6010
rect 114180 5910 114240 5970
rect 114180 5870 114190 5910
rect 114230 5870 114240 5910
rect 114180 5850 114240 5870
rect 114290 6310 114350 6330
rect 114290 6270 114300 6310
rect 114340 6270 114350 6310
rect 114290 6210 114350 6270
rect 114290 6170 114300 6210
rect 114340 6170 114350 6210
rect 114290 6110 114350 6170
rect 114290 6070 114300 6110
rect 114340 6070 114350 6110
rect 114290 6010 114350 6070
rect 114290 5970 114300 6010
rect 114340 5970 114350 6010
rect 114290 5910 114350 5970
rect 114290 5870 114300 5910
rect 114340 5870 114350 5910
rect 114290 5850 114350 5870
rect 114400 6310 114460 6330
rect 114400 6270 114410 6310
rect 114450 6270 114460 6310
rect 114400 6210 114460 6270
rect 114400 6170 114410 6210
rect 114450 6170 114460 6210
rect 114400 6110 114460 6170
rect 114400 6070 114410 6110
rect 114450 6070 114460 6110
rect 114400 6010 114460 6070
rect 114400 5970 114410 6010
rect 114450 5970 114460 6010
rect 114400 5910 114460 5970
rect 114400 5870 114410 5910
rect 114450 5870 114460 5910
rect 114400 5850 114460 5870
rect 114510 6310 114650 6330
rect 114510 6270 114520 6310
rect 114560 6270 114600 6310
rect 114640 6270 114650 6310
rect 118910 6320 119192 6340
rect 114510 6210 114650 6270
rect 114510 6170 114520 6210
rect 114560 6170 114600 6210
rect 114640 6170 114650 6210
rect 114510 6110 114650 6170
rect 114510 6070 114520 6110
rect 114560 6070 114600 6110
rect 114640 6070 114650 6110
rect 114510 6010 114650 6070
rect 114510 5970 114520 6010
rect 114560 5970 114600 6010
rect 114640 5970 114650 6010
rect 114510 5910 114650 5970
rect 114510 5870 114520 5910
rect 114560 5870 114600 5910
rect 114640 5870 114650 5910
rect 114510 5850 114650 5870
rect 116890 6280 117030 6300
rect 113140 5830 113180 5850
rect 113120 5810 113180 5830
rect 113600 5830 113640 5850
rect 113960 5830 114000 5850
rect 113600 5810 113660 5830
rect 113120 5770 113130 5810
rect 113170 5770 113180 5810
rect 113120 5750 113180 5770
rect 113214 5790 113274 5810
rect 113214 5750 113224 5790
rect 113264 5750 113274 5790
rect 113214 5730 113274 5750
rect 113350 5790 113430 5810
rect 113350 5750 113370 5790
rect 113410 5750 113430 5790
rect 113350 5730 113430 5750
rect 113506 5790 113566 5810
rect 113506 5750 113516 5790
rect 113556 5750 113566 5790
rect 113600 5770 113610 5810
rect 113650 5770 113660 5810
rect 113600 5750 113660 5770
rect 113940 5810 114000 5830
rect 114420 5830 114460 5850
rect 114420 5810 114480 5830
rect 113940 5770 113950 5810
rect 113990 5770 114000 5810
rect 113940 5750 114000 5770
rect 114034 5790 114094 5810
rect 114034 5750 114044 5790
rect 114084 5750 114094 5790
rect 113506 5730 113566 5750
rect 114034 5730 114094 5750
rect 114170 5790 114250 5810
rect 114170 5750 114190 5790
rect 114230 5750 114250 5790
rect 114170 5730 114250 5750
rect 114326 5790 114386 5810
rect 114326 5750 114336 5790
rect 114376 5750 114386 5790
rect 114420 5770 114430 5810
rect 114470 5770 114480 5810
rect 114420 5750 114480 5770
rect 114326 5730 114386 5750
rect 113200 5650 113280 5670
rect 113200 5610 113220 5650
rect 113260 5610 113280 5650
rect 113200 5590 113280 5610
rect 114320 5650 114400 5670
rect 114320 5610 114340 5650
rect 114380 5610 114400 5650
rect 114320 5590 114400 5610
rect 113700 5220 113780 5240
rect 113700 5180 113720 5220
rect 113760 5180 113780 5220
rect 113700 5160 113780 5180
rect 113870 5220 113950 5240
rect 113870 5180 113890 5220
rect 113930 5180 113950 5220
rect 113870 5160 113950 5180
rect 110570 5120 110710 5140
rect 116890 5140 116900 6280
rect 116940 5140 116980 6280
rect 117020 5140 117030 6280
rect 116890 5120 117030 5140
rect 117080 6280 117140 6300
rect 117080 5140 117090 6280
rect 117130 5140 117140 6280
rect 117080 5120 117140 5140
rect 117190 6280 117250 6300
rect 117190 5140 117200 6280
rect 117240 5140 117250 6280
rect 117190 5120 117250 5140
rect 117300 6280 117360 6300
rect 117300 5140 117310 6280
rect 117350 5140 117360 6280
rect 117300 5120 117360 5140
rect 117410 6280 117470 6300
rect 117410 5140 117420 6280
rect 117460 5140 117470 6280
rect 117410 5120 117470 5140
rect 117520 6280 117580 6300
rect 117520 5140 117530 6280
rect 117570 5140 117580 6280
rect 117520 5120 117580 5140
rect 117630 6280 117690 6300
rect 117630 5140 117640 6280
rect 117680 5140 117690 6280
rect 117630 5120 117690 5140
rect 117740 6280 117800 6300
rect 117740 5140 117750 6280
rect 117790 5140 117800 6280
rect 117740 5120 117800 5140
rect 117850 6280 117910 6300
rect 117850 5140 117860 6280
rect 117900 5140 117910 6280
rect 117850 5120 117910 5140
rect 117960 6280 118020 6300
rect 117960 5140 117970 6280
rect 118010 5140 118020 6280
rect 117960 5120 118020 5140
rect 118070 6280 118130 6300
rect 118070 5140 118080 6280
rect 118120 5140 118130 6280
rect 118070 5120 118130 5140
rect 118180 6280 118240 6300
rect 118180 5140 118190 6280
rect 118230 5140 118240 6280
rect 118180 5120 118240 5140
rect 118290 6280 118430 6300
rect 118290 5140 118300 6280
rect 118340 5140 118380 6280
rect 118420 5140 118430 6280
rect 118290 5120 118430 5140
rect 118910 5170 119192 5190
rect 118910 5130 118920 5170
rect 118960 5130 119030 5170
rect 119070 5130 119140 5170
rect 119180 5130 119192 5170
rect 113470 5100 113610 5120
rect 109910 5060 109970 5080
rect 109910 5020 109920 5060
rect 109960 5020 109970 5060
rect 109910 5000 109970 5020
rect 109900 4930 109980 4950
rect 109900 4890 109920 4930
rect 109960 4890 109980 4930
rect 109900 4850 109980 4890
rect 109900 4810 109920 4850
rect 109960 4810 109980 4850
rect 109900 4770 109980 4810
rect 109900 4730 109920 4770
rect 109960 4730 109980 4770
rect 109900 4710 109980 4730
rect 113470 4660 113480 5100
rect 113520 4660 113560 5100
rect 113600 4660 113610 5100
rect 113470 4640 113610 4660
rect 113660 5100 113720 5120
rect 113660 4660 113670 5100
rect 113710 4660 113720 5100
rect 113660 4640 113720 4660
rect 113770 5100 113830 5120
rect 113770 4660 113780 5100
rect 113820 4660 113830 5100
rect 113770 4640 113830 4660
rect 113880 5100 113940 5120
rect 113880 4660 113890 5100
rect 113930 4660 113940 5100
rect 113880 4640 113940 4660
rect 113990 5100 114130 5120
rect 118910 5110 119192 5130
rect 113990 4660 114000 5100
rect 114040 4660 114080 5100
rect 114120 4660 114130 5100
rect 117630 5060 117690 5080
rect 117630 5020 117640 5060
rect 117680 5020 117690 5060
rect 117630 5000 117690 5020
rect 117620 4930 117700 4950
rect 117620 4890 117640 4930
rect 117680 4890 117700 4930
rect 117620 4850 117700 4890
rect 117620 4810 117640 4850
rect 117680 4810 117700 4850
rect 117620 4770 117700 4810
rect 117620 4730 117640 4770
rect 117680 4730 117700 4770
rect 117620 4710 117700 4730
rect 113990 4640 114130 4660
rect 113540 4580 113620 4600
rect 113540 4540 113560 4580
rect 113600 4540 113620 4580
rect 113540 4520 113620 4540
rect 113980 4580 114060 4600
rect 113980 4540 114000 4580
rect 114040 4540 114060 4580
rect 113980 4520 114060 4540
rect 112232 3900 112298 3920
rect 109250 3850 109310 3870
rect 109250 3810 109260 3850
rect 109300 3810 109310 3850
rect 109250 3790 109310 3810
rect 110570 3850 110630 3870
rect 110570 3810 110580 3850
rect 110620 3810 110630 3850
rect 112232 3860 112245 3900
rect 112285 3860 112298 3900
rect 112232 3840 112298 3860
rect 112342 3900 112408 3920
rect 112342 3860 112355 3900
rect 112395 3860 112408 3900
rect 112342 3840 112408 3860
rect 112452 3900 112518 3920
rect 112452 3860 112465 3900
rect 112505 3860 112518 3900
rect 112452 3840 112518 3860
rect 112562 3900 112628 3920
rect 112562 3860 112575 3900
rect 112615 3860 112628 3900
rect 112562 3840 112628 3860
rect 112672 3900 112738 3920
rect 112672 3860 112685 3900
rect 112725 3860 112738 3900
rect 112672 3840 112738 3860
rect 112782 3900 112848 3920
rect 112782 3860 112795 3900
rect 112835 3860 112848 3900
rect 112782 3840 112848 3860
rect 112892 3900 112958 3920
rect 112892 3860 112905 3900
rect 112945 3860 112958 3900
rect 112892 3840 112958 3860
rect 113002 3900 113068 3920
rect 113002 3860 113015 3900
rect 113055 3860 113068 3900
rect 113002 3840 113068 3860
rect 113112 3900 113178 3920
rect 113112 3860 113125 3900
rect 113165 3860 113178 3900
rect 113112 3840 113178 3860
rect 113222 3900 113288 3920
rect 113222 3860 113235 3900
rect 113275 3860 113288 3900
rect 113222 3840 113288 3860
rect 114312 3900 114378 3920
rect 114312 3860 114325 3900
rect 114365 3860 114378 3900
rect 114312 3840 114378 3860
rect 114422 3900 114488 3920
rect 114422 3860 114435 3900
rect 114475 3860 114488 3900
rect 114422 3840 114488 3860
rect 114532 3900 114598 3920
rect 114532 3860 114545 3900
rect 114585 3860 114598 3900
rect 114532 3840 114598 3860
rect 114642 3900 114708 3920
rect 114642 3860 114655 3900
rect 114695 3860 114708 3900
rect 114642 3840 114708 3860
rect 114752 3900 114818 3920
rect 114752 3860 114765 3900
rect 114805 3860 114818 3900
rect 114752 3840 114818 3860
rect 114862 3900 114928 3920
rect 114862 3860 114875 3900
rect 114915 3860 114928 3900
rect 114862 3840 114928 3860
rect 114972 3900 115038 3920
rect 114972 3860 114985 3900
rect 115025 3860 115038 3900
rect 114972 3840 115038 3860
rect 115082 3900 115148 3920
rect 115082 3860 115095 3900
rect 115135 3860 115148 3900
rect 115082 3840 115148 3860
rect 115192 3900 115258 3920
rect 115192 3860 115205 3900
rect 115245 3860 115258 3900
rect 115192 3840 115258 3860
rect 115302 3900 115368 3920
rect 115302 3860 115315 3900
rect 115355 3860 115368 3900
rect 115302 3840 115368 3860
rect 116970 3850 117030 3870
rect 110570 3790 110630 3810
rect 116970 3810 116980 3850
rect 117020 3810 117030 3850
rect 111990 3780 112130 3800
rect 109170 3730 109310 3750
rect 108510 3562 108940 3602
rect 108510 3528 108580 3562
rect 108870 3528 108940 3562
rect 108700 3428 108750 3528
rect 109170 3390 109180 3730
rect 109220 3390 109260 3730
rect 109300 3390 109310 3730
rect 109170 3370 109310 3390
rect 109360 3730 109420 3750
rect 109360 3390 109370 3730
rect 109410 3390 109420 3730
rect 109360 3370 109420 3390
rect 109470 3730 109530 3750
rect 109470 3390 109480 3730
rect 109520 3390 109530 3730
rect 109470 3370 109530 3390
rect 109580 3730 109640 3750
rect 109580 3390 109590 3730
rect 109630 3390 109640 3730
rect 109580 3370 109640 3390
rect 109690 3730 109750 3750
rect 109690 3390 109700 3730
rect 109740 3390 109750 3730
rect 109690 3370 109750 3390
rect 109800 3730 109860 3750
rect 109800 3390 109810 3730
rect 109850 3390 109860 3730
rect 109800 3370 109860 3390
rect 109910 3730 109970 3750
rect 109910 3390 109920 3730
rect 109960 3390 109970 3730
rect 109910 3370 109970 3390
rect 110020 3730 110080 3750
rect 110020 3390 110030 3730
rect 110070 3390 110080 3730
rect 110020 3370 110080 3390
rect 110130 3730 110190 3750
rect 110130 3390 110140 3730
rect 110180 3390 110190 3730
rect 110130 3370 110190 3390
rect 110240 3730 110300 3750
rect 110240 3390 110250 3730
rect 110290 3390 110300 3730
rect 110240 3370 110300 3390
rect 110350 3730 110410 3750
rect 110350 3390 110360 3730
rect 110400 3390 110410 3730
rect 110350 3370 110410 3390
rect 110460 3730 110520 3750
rect 110460 3390 110470 3730
rect 110510 3390 110520 3730
rect 110460 3370 110520 3390
rect 110570 3730 110710 3750
rect 110570 3390 110580 3730
rect 110620 3390 110660 3730
rect 110700 3390 110710 3730
rect 111990 3540 112000 3780
rect 112040 3540 112080 3780
rect 112120 3540 112130 3780
rect 111990 3520 112130 3540
rect 112180 3780 112240 3800
rect 112180 3540 112190 3780
rect 112230 3540 112240 3780
rect 112180 3520 112240 3540
rect 112290 3780 112350 3800
rect 112290 3540 112300 3780
rect 112340 3540 112350 3780
rect 112290 3520 112350 3540
rect 112400 3780 112460 3800
rect 112400 3540 112410 3780
rect 112450 3540 112460 3780
rect 112400 3520 112460 3540
rect 112510 3780 112570 3800
rect 112510 3540 112520 3780
rect 112560 3540 112570 3780
rect 112510 3520 112570 3540
rect 112620 3780 112680 3800
rect 112620 3540 112630 3780
rect 112670 3540 112680 3780
rect 112620 3520 112680 3540
rect 112730 3780 112790 3800
rect 112730 3540 112740 3780
rect 112780 3540 112790 3780
rect 112730 3520 112790 3540
rect 112840 3780 112900 3800
rect 112840 3540 112850 3780
rect 112890 3540 112900 3780
rect 112840 3520 112900 3540
rect 112950 3780 113010 3800
rect 112950 3540 112960 3780
rect 113000 3540 113010 3780
rect 112950 3520 113010 3540
rect 113060 3780 113120 3800
rect 113060 3540 113070 3780
rect 113110 3540 113120 3780
rect 113060 3520 113120 3540
rect 113170 3780 113230 3800
rect 113170 3540 113180 3780
rect 113220 3540 113230 3780
rect 113170 3520 113230 3540
rect 113280 3780 113340 3800
rect 113280 3540 113290 3780
rect 113330 3540 113340 3780
rect 113280 3520 113340 3540
rect 113390 3780 113530 3800
rect 113390 3540 113400 3780
rect 113440 3540 113480 3780
rect 113520 3540 113530 3780
rect 113390 3520 113530 3540
rect 114070 3780 114210 3800
rect 114070 3540 114080 3780
rect 114120 3540 114160 3780
rect 114200 3540 114210 3780
rect 114070 3520 114210 3540
rect 114260 3780 114320 3800
rect 114260 3540 114270 3780
rect 114310 3540 114320 3780
rect 114260 3520 114320 3540
rect 114370 3780 114430 3800
rect 114370 3540 114380 3780
rect 114420 3540 114430 3780
rect 114370 3520 114430 3540
rect 114480 3780 114540 3800
rect 114480 3540 114490 3780
rect 114530 3540 114540 3780
rect 114480 3520 114540 3540
rect 114590 3780 114650 3800
rect 114590 3540 114600 3780
rect 114640 3540 114650 3780
rect 114590 3520 114650 3540
rect 114700 3780 114760 3800
rect 114700 3540 114710 3780
rect 114750 3540 114760 3780
rect 114700 3520 114760 3540
rect 114810 3780 114870 3800
rect 114810 3540 114820 3780
rect 114860 3540 114870 3780
rect 114810 3520 114870 3540
rect 114920 3780 114980 3800
rect 114920 3540 114930 3780
rect 114970 3540 114980 3780
rect 114920 3520 114980 3540
rect 115030 3780 115090 3800
rect 115030 3540 115040 3780
rect 115080 3540 115090 3780
rect 115030 3520 115090 3540
rect 115140 3780 115200 3800
rect 115140 3540 115150 3780
rect 115190 3540 115200 3780
rect 115140 3520 115200 3540
rect 115250 3780 115310 3800
rect 115250 3540 115260 3780
rect 115300 3540 115310 3780
rect 115250 3520 115310 3540
rect 115360 3780 115420 3800
rect 115360 3540 115370 3780
rect 115410 3540 115420 3780
rect 115360 3520 115420 3540
rect 115470 3780 115610 3800
rect 116970 3790 117030 3810
rect 118290 3850 118350 3870
rect 118290 3810 118300 3850
rect 118340 3810 118350 3850
rect 118290 3790 118350 3810
rect 115470 3540 115480 3780
rect 115520 3540 115560 3780
rect 115600 3540 115610 3780
rect 115470 3520 115610 3540
rect 116890 3730 117030 3750
rect 112070 3460 112130 3520
rect 112070 3420 112080 3460
rect 112120 3420 112130 3460
rect 112070 3400 112130 3420
rect 113390 3460 113450 3480
rect 113390 3420 113400 3460
rect 113440 3420 113450 3460
rect 113390 3400 113450 3420
rect 114150 3460 114210 3480
rect 114150 3420 114160 3460
rect 114200 3420 114210 3460
rect 114150 3400 114210 3420
rect 115470 3460 115530 3520
rect 115470 3420 115480 3460
rect 115520 3420 115530 3460
rect 115470 3400 115530 3420
rect 110570 3370 110710 3390
rect 116890 3390 116900 3730
rect 116940 3390 116980 3730
rect 117020 3390 117030 3730
rect 116890 3370 117030 3390
rect 117080 3730 117140 3750
rect 117080 3390 117090 3730
rect 117130 3390 117140 3730
rect 117080 3370 117140 3390
rect 117190 3730 117250 3750
rect 117190 3390 117200 3730
rect 117240 3390 117250 3730
rect 117190 3370 117250 3390
rect 117300 3730 117360 3750
rect 117300 3390 117310 3730
rect 117350 3390 117360 3730
rect 117300 3370 117360 3390
rect 117410 3730 117470 3750
rect 117410 3390 117420 3730
rect 117460 3390 117470 3730
rect 117410 3370 117470 3390
rect 117520 3730 117580 3750
rect 117520 3390 117530 3730
rect 117570 3390 117580 3730
rect 117520 3370 117580 3390
rect 117630 3730 117690 3750
rect 117630 3390 117640 3730
rect 117680 3390 117690 3730
rect 117630 3370 117690 3390
rect 117740 3730 117800 3750
rect 117740 3390 117750 3730
rect 117790 3390 117800 3730
rect 117740 3370 117800 3390
rect 117850 3730 117910 3750
rect 117850 3390 117860 3730
rect 117900 3390 117910 3730
rect 117850 3370 117910 3390
rect 117960 3730 118020 3750
rect 117960 3390 117970 3730
rect 118010 3390 118020 3730
rect 117960 3370 118020 3390
rect 118070 3730 118130 3750
rect 118070 3390 118080 3730
rect 118120 3390 118130 3730
rect 118070 3370 118130 3390
rect 118180 3730 118240 3750
rect 118180 3390 118190 3730
rect 118230 3390 118240 3730
rect 118180 3370 118240 3390
rect 118290 3730 118430 3750
rect 118290 3390 118300 3730
rect 118340 3390 118380 3730
rect 118420 3390 118430 3730
rect 118290 3370 118430 3390
rect 118660 3562 119090 3602
rect 118660 3528 118730 3562
rect 119020 3528 119090 3562
rect 109460 3310 109540 3330
rect 109460 3270 109480 3310
rect 109520 3270 109540 3310
rect 109460 3250 109540 3270
rect 109680 3310 109760 3330
rect 109680 3270 109700 3310
rect 109740 3270 109760 3310
rect 109680 3250 109760 3270
rect 109900 3310 109980 3330
rect 109900 3270 109920 3310
rect 109960 3270 109980 3310
rect 109900 3250 109980 3270
rect 110120 3310 110200 3330
rect 110120 3270 110140 3310
rect 110180 3270 110200 3310
rect 110120 3250 110200 3270
rect 110240 3310 110300 3330
rect 110240 3270 110250 3310
rect 110290 3270 110300 3310
rect 110240 3250 110300 3270
rect 110340 3310 110420 3330
rect 110340 3270 110360 3310
rect 110400 3270 110420 3310
rect 110340 3250 110420 3270
rect 117180 3310 117260 3330
rect 117180 3270 117200 3310
rect 117240 3270 117260 3310
rect 117180 3250 117260 3270
rect 117300 3310 117360 3330
rect 117300 3270 117310 3310
rect 117350 3270 117360 3310
rect 117300 3250 117360 3270
rect 117400 3310 117480 3330
rect 117400 3270 117420 3310
rect 117460 3270 117480 3310
rect 117400 3250 117480 3270
rect 117620 3310 117700 3330
rect 117620 3270 117640 3310
rect 117680 3270 117700 3310
rect 117620 3250 117700 3270
rect 117840 3310 117920 3330
rect 117840 3270 117860 3310
rect 117900 3270 117920 3310
rect 117840 3250 117920 3270
rect 118060 3310 118140 3330
rect 118060 3270 118080 3310
rect 118120 3270 118140 3310
rect 118060 3250 118140 3270
rect 110230 3180 110310 3200
rect 110230 3140 110250 3180
rect 110290 3140 110310 3180
rect 110230 3100 110310 3140
rect 110230 3060 110250 3100
rect 110290 3060 110310 3100
rect 110230 3040 110310 3060
rect 117290 3180 117370 3200
rect 117290 3140 117310 3180
rect 117350 3140 117370 3180
rect 117290 3100 117370 3140
rect 117290 3060 117310 3100
rect 117350 3060 117370 3100
rect 118850 3428 118900 3528
rect 117290 3040 117370 3060
rect 110240 2970 110300 2990
rect 110240 2930 110250 2970
rect 110290 2930 110300 2970
rect 110240 2910 110300 2930
rect 117300 2970 117360 2990
rect 117300 2930 117310 2970
rect 117350 2930 117360 2970
rect 117300 2910 117360 2930
rect 109170 2850 109310 2870
rect 108510 2310 108580 2330
rect 108510 2260 108520 2310
rect 108570 2260 108580 2310
rect 108510 2240 108580 2260
rect 108630 2310 108700 2330
rect 108630 2260 108640 2310
rect 108690 2260 108700 2310
rect 108630 2240 108700 2260
rect 108750 2310 108820 2330
rect 108750 2260 108760 2310
rect 108810 2260 108820 2310
rect 108750 2240 108820 2260
rect 108870 2310 108940 2330
rect 108870 2260 108880 2310
rect 108930 2260 108940 2310
rect 109170 2310 109180 2850
rect 109220 2310 109260 2850
rect 109300 2310 109310 2850
rect 109170 2290 109310 2310
rect 109360 2850 109420 2870
rect 109360 2310 109370 2850
rect 109410 2310 109420 2850
rect 109360 2290 109420 2310
rect 109470 2850 109530 2870
rect 109470 2310 109480 2850
rect 109520 2310 109530 2850
rect 109470 2290 109530 2310
rect 109580 2850 109640 2870
rect 109580 2310 109590 2850
rect 109630 2310 109640 2850
rect 109580 2290 109640 2310
rect 109690 2850 109750 2870
rect 109690 2310 109700 2850
rect 109740 2310 109750 2850
rect 109690 2290 109750 2310
rect 109800 2850 109860 2870
rect 109800 2310 109810 2850
rect 109850 2310 109860 2850
rect 109800 2290 109860 2310
rect 109910 2850 109970 2870
rect 109910 2310 109920 2850
rect 109960 2310 109970 2850
rect 109910 2290 109970 2310
rect 110020 2850 110080 2870
rect 110020 2310 110030 2850
rect 110070 2310 110080 2850
rect 110020 2290 110080 2310
rect 110130 2850 110190 2870
rect 110130 2310 110140 2850
rect 110180 2310 110190 2850
rect 110130 2290 110190 2310
rect 110240 2850 110300 2870
rect 110240 2310 110250 2850
rect 110290 2310 110300 2850
rect 110240 2290 110300 2310
rect 110350 2850 110410 2870
rect 110350 2310 110360 2850
rect 110400 2310 110410 2850
rect 110350 2290 110410 2310
rect 110460 2850 110520 2870
rect 110460 2310 110470 2850
rect 110510 2310 110520 2850
rect 110460 2290 110520 2310
rect 110570 2850 110710 2870
rect 110570 2310 110580 2850
rect 110620 2310 110660 2850
rect 110700 2310 110710 2850
rect 116890 2850 117030 2870
rect 113380 2600 113440 2620
rect 112080 2580 112140 2600
rect 112080 2540 112090 2580
rect 112130 2540 112140 2580
rect 113380 2560 113390 2600
rect 113430 2560 113440 2600
rect 113380 2540 113440 2560
rect 113680 2600 113740 2620
rect 113680 2560 113690 2600
rect 113730 2560 113740 2600
rect 113680 2540 113740 2560
rect 113860 2600 113920 2620
rect 113860 2560 113870 2600
rect 113910 2560 113920 2600
rect 113860 2540 113920 2560
rect 114160 2600 114220 2620
rect 114160 2560 114170 2600
rect 114210 2560 114220 2600
rect 114160 2540 114220 2560
rect 115460 2580 115520 2600
rect 115460 2540 115470 2580
rect 115510 2540 115520 2580
rect 112080 2520 112140 2540
rect 115460 2520 115520 2540
rect 110570 2290 110710 2310
rect 111990 2410 112130 2430
rect 108870 2240 108940 2260
rect 109250 2230 109310 2250
rect 109250 2190 109260 2230
rect 109300 2190 109310 2230
rect 109250 2160 109310 2190
rect 110570 2230 110630 2250
rect 110570 2190 110580 2230
rect 110620 2190 110630 2230
rect 110570 2160 110630 2190
rect 111990 2170 112000 2410
rect 112040 2170 112080 2410
rect 112120 2170 112130 2410
rect 111990 2150 112130 2170
rect 112180 2410 112240 2430
rect 112180 2170 112190 2410
rect 112230 2170 112240 2410
rect 112180 2150 112240 2170
rect 112290 2410 112350 2430
rect 112290 2170 112300 2410
rect 112340 2170 112350 2410
rect 112290 2150 112350 2170
rect 112400 2410 112460 2430
rect 112400 2170 112410 2410
rect 112450 2170 112460 2410
rect 112400 2150 112460 2170
rect 112510 2410 112570 2430
rect 112510 2170 112520 2410
rect 112560 2170 112570 2410
rect 112510 2150 112570 2170
rect 112620 2410 112680 2430
rect 112620 2170 112630 2410
rect 112670 2170 112680 2410
rect 112620 2150 112680 2170
rect 112730 2410 112790 2430
rect 112730 2170 112740 2410
rect 112780 2170 112790 2410
rect 112730 2150 112790 2170
rect 112840 2410 112900 2430
rect 112840 2170 112850 2410
rect 112890 2170 112900 2410
rect 112840 2150 112900 2170
rect 112950 2410 113010 2430
rect 112950 2170 112960 2410
rect 113000 2170 113010 2410
rect 112950 2150 113010 2170
rect 113060 2410 113120 2430
rect 113060 2170 113070 2410
rect 113110 2170 113120 2410
rect 113060 2150 113120 2170
rect 113170 2410 113230 2430
rect 113170 2170 113180 2410
rect 113220 2170 113230 2410
rect 113170 2150 113230 2170
rect 113280 2410 113340 2430
rect 113280 2170 113290 2410
rect 113330 2170 113340 2410
rect 113280 2150 113340 2170
rect 113390 2410 113610 2430
rect 113390 2170 113400 2410
rect 113440 2170 113480 2410
rect 113520 2170 113560 2410
rect 113600 2170 113610 2410
rect 113390 2150 113610 2170
rect 113660 2410 113720 2430
rect 113660 2170 113670 2410
rect 113710 2170 113720 2410
rect 113660 2150 113720 2170
rect 113770 2410 113830 2430
rect 113770 2170 113780 2410
rect 113820 2170 113830 2410
rect 113770 2150 113830 2170
rect 113880 2410 113940 2430
rect 113880 2170 113890 2410
rect 113930 2170 113940 2410
rect 113880 2150 113940 2170
rect 113990 2410 114210 2430
rect 113990 2170 114000 2410
rect 114040 2170 114080 2410
rect 114120 2170 114160 2410
rect 114200 2170 114210 2410
rect 113990 2150 114210 2170
rect 114260 2410 114320 2430
rect 114260 2170 114270 2410
rect 114310 2170 114320 2410
rect 114260 2150 114320 2170
rect 114370 2410 114430 2430
rect 114370 2170 114380 2410
rect 114420 2170 114430 2410
rect 114370 2150 114430 2170
rect 114480 2410 114540 2430
rect 114480 2170 114490 2410
rect 114530 2170 114540 2410
rect 114480 2150 114540 2170
rect 114590 2410 114650 2430
rect 114590 2170 114600 2410
rect 114640 2170 114650 2410
rect 114590 2150 114650 2170
rect 114700 2410 114760 2430
rect 114700 2170 114710 2410
rect 114750 2170 114760 2410
rect 114700 2150 114760 2170
rect 114810 2410 114870 2430
rect 114810 2170 114820 2410
rect 114860 2170 114870 2410
rect 114810 2150 114870 2170
rect 114920 2410 114980 2430
rect 114920 2170 114930 2410
rect 114970 2170 114980 2410
rect 114920 2150 114980 2170
rect 115030 2410 115090 2430
rect 115030 2170 115040 2410
rect 115080 2170 115090 2410
rect 115030 2150 115090 2170
rect 115140 2410 115200 2430
rect 115140 2170 115150 2410
rect 115190 2170 115200 2410
rect 115140 2150 115200 2170
rect 115250 2410 115310 2430
rect 115250 2170 115260 2410
rect 115300 2170 115310 2410
rect 115250 2150 115310 2170
rect 115360 2410 115420 2430
rect 115360 2170 115370 2410
rect 115410 2170 115420 2410
rect 115360 2150 115420 2170
rect 115470 2410 115610 2430
rect 115470 2170 115480 2410
rect 115520 2170 115560 2410
rect 115600 2170 115610 2410
rect 116890 2310 116900 2850
rect 116940 2310 116980 2850
rect 117020 2310 117030 2850
rect 116890 2290 117030 2310
rect 117080 2850 117140 2870
rect 117080 2310 117090 2850
rect 117130 2310 117140 2850
rect 117080 2290 117140 2310
rect 117190 2850 117250 2870
rect 117190 2310 117200 2850
rect 117240 2310 117250 2850
rect 117190 2290 117250 2310
rect 117300 2850 117360 2870
rect 117300 2310 117310 2850
rect 117350 2310 117360 2850
rect 117300 2290 117360 2310
rect 117410 2850 117470 2870
rect 117410 2310 117420 2850
rect 117460 2310 117470 2850
rect 117410 2290 117470 2310
rect 117520 2850 117580 2870
rect 117520 2310 117530 2850
rect 117570 2310 117580 2850
rect 117520 2290 117580 2310
rect 117630 2850 117690 2870
rect 117630 2310 117640 2850
rect 117680 2310 117690 2850
rect 117630 2290 117690 2310
rect 117740 2850 117800 2870
rect 117740 2310 117750 2850
rect 117790 2310 117800 2850
rect 117740 2290 117800 2310
rect 117850 2850 117910 2870
rect 117850 2310 117860 2850
rect 117900 2310 117910 2850
rect 117850 2290 117910 2310
rect 117960 2850 118020 2870
rect 117960 2310 117970 2850
rect 118010 2310 118020 2850
rect 117960 2290 118020 2310
rect 118070 2850 118130 2870
rect 118070 2310 118080 2850
rect 118120 2310 118130 2850
rect 118070 2290 118130 2310
rect 118180 2850 118240 2870
rect 118180 2310 118190 2850
rect 118230 2310 118240 2850
rect 118180 2290 118240 2310
rect 118290 2850 118430 2870
rect 118290 2310 118300 2850
rect 118340 2310 118380 2850
rect 118420 2310 118430 2850
rect 118290 2290 118430 2310
rect 118660 2310 118730 2330
rect 118660 2260 118670 2310
rect 118720 2260 118730 2310
rect 115470 2150 115610 2170
rect 116970 2230 117030 2250
rect 116970 2190 116980 2230
rect 117020 2190 117030 2230
rect 116970 2160 117030 2190
rect 118290 2230 118350 2250
rect 118660 2240 118730 2260
rect 118780 2310 118850 2330
rect 118780 2260 118790 2310
rect 118840 2260 118850 2310
rect 118780 2240 118850 2260
rect 118900 2310 118970 2330
rect 118900 2260 118910 2310
rect 118960 2260 118970 2310
rect 118900 2240 118970 2260
rect 119020 2310 119090 2330
rect 119020 2260 119030 2310
rect 119080 2260 119090 2310
rect 119020 2240 119090 2260
rect 118290 2190 118300 2230
rect 118340 2190 118350 2230
rect 118290 2170 118350 2190
rect 112080 2110 112130 2150
rect 112070 2090 112130 2110
rect 112070 2050 112080 2090
rect 112120 2050 112130 2090
rect 112070 2030 112130 2050
rect 113470 2090 113530 2110
rect 113470 2050 113480 2090
rect 113520 2050 113530 2090
rect 113470 2030 113530 2050
rect 114070 2090 114130 2110
rect 114070 2050 114080 2090
rect 114120 2050 114130 2090
rect 114070 2030 114130 2050
rect 115470 2090 115530 2150
rect 115470 2050 115480 2090
rect 115520 2050 115530 2090
rect 115470 2030 115530 2050
rect 113650 1000 113730 1020
rect 113650 960 113670 1000
rect 113710 960 113730 1000
rect 113650 940 113730 960
rect 113870 1000 113950 1020
rect 113870 960 113890 1000
rect 113930 960 113950 1000
rect 113870 940 113950 960
rect 112370 880 112510 900
rect 109600 760 109680 780
rect 109600 720 109620 760
rect 109660 720 109680 760
rect 109600 700 109680 720
rect 109800 760 109880 780
rect 109800 720 109820 760
rect 109860 720 109880 760
rect 109800 700 109880 720
rect 110000 760 110080 780
rect 110000 720 110020 760
rect 110060 720 110080 760
rect 110000 700 110080 720
rect 110200 760 110280 780
rect 110200 720 110220 760
rect 110260 720 110280 760
rect 110200 700 110280 720
rect 108650 650 108720 670
rect 108650 600 108660 650
rect 108710 600 108720 650
rect 108650 580 108720 600
rect 108770 650 108840 670
rect 108770 600 108780 650
rect 108830 600 108840 650
rect 108770 580 108840 600
rect 109230 650 109370 670
rect 108720 -794 108770 -694
rect 109230 -690 109240 650
rect 109280 -690 109320 650
rect 109360 -690 109370 650
rect 109230 -710 109370 -690
rect 109510 650 109570 670
rect 109510 -690 109520 650
rect 109560 -690 109570 650
rect 109510 -710 109570 -690
rect 109710 650 109770 670
rect 109710 -690 109720 650
rect 109760 -690 109770 650
rect 109710 -710 109770 -690
rect 109910 650 109970 670
rect 109910 -690 109920 650
rect 109960 -690 109970 650
rect 109910 -710 109970 -690
rect 110110 650 110170 670
rect 110110 -690 110120 650
rect 110160 -690 110170 650
rect 110110 -710 110170 -690
rect 110310 650 110370 670
rect 110310 -690 110320 650
rect 110360 -690 110370 650
rect 110310 -710 110370 -690
rect 110510 650 110650 670
rect 110510 -690 110520 650
rect 110560 -690 110600 650
rect 110640 -690 110650 650
rect 112370 440 112380 880
rect 112420 440 112460 880
rect 112500 440 112510 880
rect 112370 420 112510 440
rect 112560 880 112620 900
rect 112560 440 112570 880
rect 112610 440 112620 880
rect 112560 420 112620 440
rect 112670 880 112730 900
rect 112670 440 112680 880
rect 112720 440 112730 880
rect 112670 420 112730 440
rect 112780 880 112840 900
rect 112780 440 112790 880
rect 112830 440 112840 880
rect 112780 420 112840 440
rect 112890 880 112950 900
rect 112890 440 112900 880
rect 112940 440 112950 880
rect 112890 420 112950 440
rect 113000 880 113060 900
rect 113000 440 113010 880
rect 113050 440 113060 880
rect 113000 420 113060 440
rect 113110 880 113170 900
rect 113110 440 113120 880
rect 113160 440 113170 880
rect 113110 420 113170 440
rect 113220 880 113280 900
rect 113220 440 113230 880
rect 113270 440 113280 880
rect 113220 420 113280 440
rect 113330 880 113390 900
rect 113330 440 113340 880
rect 113380 440 113390 880
rect 113330 420 113390 440
rect 113440 880 113500 900
rect 113440 440 113450 880
rect 113490 440 113500 880
rect 113440 420 113500 440
rect 113550 880 113610 900
rect 113550 440 113560 880
rect 113600 440 113610 880
rect 113550 420 113610 440
rect 113660 880 113720 900
rect 113660 440 113670 880
rect 113710 440 113720 880
rect 113660 420 113720 440
rect 113770 880 113830 900
rect 113770 440 113780 880
rect 113820 440 113830 880
rect 113770 420 113830 440
rect 113880 880 113940 900
rect 113880 440 113890 880
rect 113930 440 113940 880
rect 113880 420 113940 440
rect 113990 880 114050 900
rect 113990 440 114000 880
rect 114040 440 114050 880
rect 113990 420 114050 440
rect 114100 880 114160 900
rect 114100 440 114110 880
rect 114150 440 114160 880
rect 114100 420 114160 440
rect 114210 880 114270 900
rect 114210 440 114220 880
rect 114260 440 114270 880
rect 114210 420 114270 440
rect 114320 880 114380 900
rect 114320 440 114330 880
rect 114370 440 114380 880
rect 114320 420 114380 440
rect 114430 880 114490 900
rect 114430 440 114440 880
rect 114480 440 114490 880
rect 114430 420 114490 440
rect 114540 880 114600 900
rect 114540 440 114550 880
rect 114590 440 114600 880
rect 114540 420 114600 440
rect 114650 880 114710 900
rect 114650 440 114660 880
rect 114700 440 114710 880
rect 114650 420 114710 440
rect 114760 880 114820 900
rect 114760 440 114770 880
rect 114810 440 114820 880
rect 114760 420 114820 440
rect 114870 880 114930 900
rect 114870 440 114880 880
rect 114920 440 114930 880
rect 114870 420 114930 440
rect 114980 880 115120 900
rect 114980 440 114990 880
rect 115030 440 115070 880
rect 115110 440 115120 880
rect 117320 760 117400 780
rect 117320 720 117340 760
rect 117380 720 117400 760
rect 117320 700 117400 720
rect 117520 760 117600 780
rect 117520 720 117540 760
rect 117580 720 117600 760
rect 117520 700 117600 720
rect 117720 760 117800 780
rect 117720 720 117740 760
rect 117780 720 117800 760
rect 117720 700 117800 720
rect 117920 760 118000 780
rect 117920 720 117940 760
rect 117980 720 118000 760
rect 117920 700 118000 720
rect 114980 420 115120 440
rect 116950 650 117090 670
rect 112440 360 112520 380
rect 112440 320 112460 360
rect 112500 320 112520 360
rect 112440 300 112520 320
rect 114970 360 115050 380
rect 114970 320 114990 360
rect 115030 320 115050 360
rect 114970 300 115050 320
rect 114830 -20 114910 0
rect 114830 -60 114850 -20
rect 114890 -60 114910 -20
rect 114830 -80 114910 -60
rect 113190 -510 113270 -490
rect 113190 -550 113210 -510
rect 113250 -550 113270 -510
rect 113190 -570 113270 -550
rect 114080 -510 114160 -490
rect 114080 -550 114100 -510
rect 114140 -550 114160 -510
rect 114080 -570 114160 -550
rect 110510 -710 110650 -690
rect 112790 -630 112930 -610
rect 109310 -770 109370 -750
rect 109310 -810 109320 -770
rect 109360 -810 109370 -770
rect 109310 -830 109370 -810
rect 110510 -770 110570 -750
rect 110510 -810 110520 -770
rect 110560 -810 110570 -770
rect 110510 -830 110570 -810
rect 112790 -870 112800 -630
rect 112840 -870 112880 -630
rect 112920 -870 112930 -630
rect 112790 -890 112930 -870
rect 112980 -630 113040 -610
rect 112980 -870 112990 -630
rect 113030 -870 113040 -630
rect 112980 -890 113040 -870
rect 113090 -630 113150 -610
rect 113090 -870 113100 -630
rect 113140 -870 113150 -630
rect 113090 -890 113150 -870
rect 113200 -630 113260 -610
rect 113200 -870 113210 -630
rect 113250 -870 113260 -630
rect 113200 -890 113260 -870
rect 113310 -630 113370 -610
rect 113310 -870 113320 -630
rect 113360 -870 113370 -630
rect 113310 -890 113370 -870
rect 113420 -630 113480 -610
rect 113420 -870 113430 -630
rect 113470 -870 113480 -630
rect 113420 -890 113480 -870
rect 113530 -630 113670 -610
rect 113530 -870 113540 -630
rect 113580 -870 113620 -630
rect 113660 -870 113670 -630
rect 113530 -890 113670 -870
rect 113750 -630 113810 -610
rect 113750 -870 113760 -630
rect 113800 -870 113810 -630
rect 114430 -650 114490 -630
rect 114430 -850 114440 -650
rect 114480 -850 114490 -650
rect 116950 -690 116960 650
rect 117000 -690 117040 650
rect 117080 -690 117090 650
rect 116950 -710 117090 -690
rect 117230 650 117290 670
rect 117230 -690 117240 650
rect 117280 -690 117290 650
rect 117230 -710 117290 -690
rect 117430 650 117490 670
rect 117430 -690 117440 650
rect 117480 -690 117490 650
rect 117430 -710 117490 -690
rect 117630 650 117690 670
rect 117630 -690 117640 650
rect 117680 -690 117690 650
rect 117630 -710 117690 -690
rect 117830 650 117890 670
rect 117830 -690 117840 650
rect 117880 -690 117890 650
rect 117830 -710 117890 -690
rect 118030 650 118090 670
rect 118030 -690 118040 650
rect 118080 -690 118090 650
rect 118030 -710 118090 -690
rect 118230 650 118370 670
rect 118230 -690 118240 650
rect 118280 -690 118320 650
rect 118360 -690 118370 650
rect 118760 650 118830 670
rect 118760 600 118770 650
rect 118820 600 118830 650
rect 118760 580 118830 600
rect 118880 650 118950 670
rect 118880 600 118890 650
rect 118940 600 118950 650
rect 118880 580 118950 600
rect 118230 -710 118370 -690
rect 117030 -770 117090 -750
rect 117030 -810 117040 -770
rect 117080 -810 117090 -770
rect 117030 -830 117090 -810
rect 118230 -770 118290 -750
rect 118230 -810 118240 -770
rect 118280 -810 118290 -770
rect 118830 -794 118880 -694
rect 118230 -830 118290 -810
rect 114430 -870 114490 -850
rect 113750 -890 113810 -870
rect 112870 -950 112930 -930
rect 112870 -990 112880 -950
rect 112920 -990 112930 -950
rect 112870 -1010 112930 -990
rect 113530 -950 113590 -930
rect 113530 -990 113540 -950
rect 113580 -990 113590 -950
rect 113530 -1010 113590 -990
rect 114080 -950 114160 -930
rect 114080 -990 114100 -950
rect 114140 -990 114160 -950
rect 114080 -1010 114160 -990
<< viali >>
rect 112190 9810 112230 9850
rect 112550 9810 112590 9850
rect 114070 9810 114110 9850
rect 114430 9810 114470 9850
rect 115010 9810 115050 9850
rect 115370 9810 115410 9850
rect 112190 9090 112230 9730
rect 112310 9090 112350 9730
rect 112430 9090 112470 9730
rect 112550 9090 112590 9730
rect 113130 9470 113170 9510
rect 113490 9470 113530 9510
rect 113130 9090 113170 9390
rect 113250 9090 113290 9390
rect 113370 9090 113410 9390
rect 113490 9090 113530 9390
rect 114070 9090 114110 9730
rect 114190 9090 114230 9730
rect 114310 9090 114350 9730
rect 114430 9090 114470 9730
rect 115010 9090 115050 9730
rect 115130 9090 115170 9730
rect 115250 9090 115290 9730
rect 115370 9090 115410 9730
rect 112320 8910 112360 8950
rect 113270 8910 113310 8950
rect 114290 8910 114330 8950
rect 115162 8890 115202 8930
rect 112030 7810 112070 7850
rect 113470 7810 113510 7850
rect 114090 7810 114130 7850
rect 115530 7810 115570 7850
rect 116920 7810 116960 7850
rect 118360 7810 118400 7850
rect 109200 7090 109240 7730
rect 109320 7090 109360 7730
rect 109440 7090 109480 7730
rect 109560 7090 109600 7730
rect 109680 7090 109720 7730
rect 109800 7090 109840 7730
rect 109920 7090 109960 7730
rect 110040 7090 110080 7730
rect 110160 7090 110200 7730
rect 110280 7090 110320 7730
rect 110400 7090 110440 7730
rect 110520 7090 110560 7730
rect 110640 7090 110680 7730
rect 112030 7090 112070 7730
rect 112150 7090 112190 7730
rect 112270 7090 112310 7730
rect 112390 7090 112430 7730
rect 112510 7090 112550 7730
rect 112630 7090 112670 7730
rect 112750 7090 112790 7730
rect 112870 7090 112910 7730
rect 112990 7090 113030 7730
rect 113110 7090 113150 7730
rect 113230 7090 113270 7730
rect 113350 7090 113390 7730
rect 113470 7090 113510 7730
rect 114090 7090 114130 7730
rect 114210 7090 114250 7730
rect 114330 7090 114370 7730
rect 114450 7090 114490 7730
rect 114570 7090 114610 7730
rect 114690 7090 114730 7730
rect 114810 7090 114850 7730
rect 114930 7090 114970 7730
rect 115050 7090 115090 7730
rect 115170 7090 115210 7730
rect 115290 7090 115330 7730
rect 115410 7090 115450 7730
rect 115530 7090 115570 7730
rect 116920 7090 116960 7730
rect 117040 7090 117080 7730
rect 117160 7090 117200 7730
rect 117280 7090 117320 7730
rect 117400 7090 117440 7730
rect 117520 7090 117560 7730
rect 117640 7090 117680 7730
rect 117760 7090 117800 7730
rect 117880 7090 117920 7730
rect 118000 7090 118040 7730
rect 118120 7090 118160 7730
rect 118240 7090 118280 7730
rect 118360 7090 118400 7730
rect 116920 6970 116960 7010
rect 118360 6970 118400 7010
rect 109380 6890 109420 6930
rect 109500 6890 109540 6930
rect 109620 6890 109660 6930
rect 109740 6890 109780 6930
rect 109860 6890 109900 6930
rect 109980 6890 110020 6930
rect 110100 6890 110140 6930
rect 110220 6890 110260 6930
rect 110340 6890 110380 6930
rect 110460 6890 110500 6930
rect 112210 6890 112250 6930
rect 112330 6890 112370 6930
rect 112450 6890 112490 6930
rect 112570 6890 112610 6930
rect 112690 6890 112730 6930
rect 112810 6890 112850 6930
rect 112930 6890 112970 6930
rect 113050 6890 113090 6930
rect 113170 6890 113210 6930
rect 113290 6890 113330 6930
rect 114270 6890 114310 6930
rect 114390 6890 114430 6930
rect 114510 6890 114550 6930
rect 114630 6890 114670 6930
rect 114750 6890 114790 6930
rect 114870 6890 114910 6930
rect 114990 6890 115030 6930
rect 115110 6890 115150 6930
rect 115230 6890 115270 6930
rect 115350 6890 115390 6930
rect 117100 6890 117140 6930
rect 117220 6890 117260 6930
rect 117340 6890 117380 6930
rect 117460 6890 117500 6930
rect 117580 6890 117620 6930
rect 117700 6890 117740 6930
rect 117820 6890 117860 6930
rect 117940 6890 117980 6930
rect 118060 6890 118100 6930
rect 118180 6890 118220 6930
rect 113040 6500 113080 6540
rect 113370 6500 113410 6540
rect 113700 6500 113740 6540
rect 113860 6500 113900 6540
rect 114190 6500 114230 6540
rect 114520 6500 114560 6540
rect 108420 6340 108460 6380
rect 108530 6340 108570 6380
rect 108640 6340 108680 6380
rect 109260 6360 109300 6400
rect 110580 6360 110620 6400
rect 113260 6390 113300 6430
rect 113480 6390 113520 6430
rect 114080 6390 114120 6430
rect 114300 6390 114340 6430
rect 116980 6360 117020 6400
rect 118300 6360 118340 6400
rect 118920 6340 118960 6380
rect 119030 6340 119070 6380
rect 119140 6340 119180 6380
rect 108420 5130 108460 5170
rect 108530 5130 108570 5170
rect 108640 5130 108680 5170
rect 109260 5140 109300 6280
rect 109370 5140 109410 6280
rect 109480 5140 109520 6280
rect 109590 5140 109630 6280
rect 109700 5140 109740 6280
rect 109810 5140 109850 6280
rect 109920 5140 109960 6280
rect 110030 5140 110070 6280
rect 110140 5140 110180 6280
rect 110250 5140 110290 6280
rect 110360 5140 110400 6280
rect 110470 5140 110510 6280
rect 110580 5140 110620 6280
rect 113130 5770 113170 5810
rect 113224 5750 113264 5790
rect 113370 5750 113410 5790
rect 113516 5750 113556 5790
rect 113610 5770 113650 5810
rect 113950 5770 113990 5810
rect 114044 5750 114084 5790
rect 114190 5750 114230 5790
rect 114336 5750 114376 5790
rect 114430 5770 114470 5810
rect 113220 5610 113260 5650
rect 114340 5610 114380 5650
rect 113720 5180 113760 5220
rect 113890 5180 113930 5220
rect 116980 5140 117020 6280
rect 117090 5140 117130 6280
rect 117200 5140 117240 6280
rect 117310 5140 117350 6280
rect 117420 5140 117460 6280
rect 117530 5140 117570 6280
rect 117640 5140 117680 6280
rect 117750 5140 117790 6280
rect 117860 5140 117900 6280
rect 117970 5140 118010 6280
rect 118080 5140 118120 6280
rect 118190 5140 118230 6280
rect 118300 5140 118340 6280
rect 118920 5130 118960 5170
rect 119030 5130 119070 5170
rect 119140 5130 119180 5170
rect 109920 4890 109960 4930
rect 109920 4810 109960 4850
rect 109920 4730 109960 4770
rect 113560 4660 113600 5100
rect 113670 4660 113710 5100
rect 113780 4660 113820 5100
rect 113890 4660 113930 5100
rect 114000 4660 114040 5100
rect 117640 4890 117680 4930
rect 117640 4810 117680 4850
rect 117640 4730 117680 4770
rect 113560 4540 113600 4580
rect 114000 4540 114040 4580
rect 109260 3810 109300 3850
rect 110580 3810 110620 3850
rect 112245 3860 112285 3900
rect 112355 3860 112395 3900
rect 112465 3860 112505 3900
rect 112575 3860 112615 3900
rect 112685 3860 112725 3900
rect 112795 3860 112835 3900
rect 112905 3860 112945 3900
rect 113015 3860 113055 3900
rect 113125 3860 113165 3900
rect 113235 3860 113275 3900
rect 114325 3860 114365 3900
rect 114435 3860 114475 3900
rect 114545 3860 114585 3900
rect 114655 3860 114695 3900
rect 114765 3860 114805 3900
rect 114875 3860 114915 3900
rect 114985 3860 115025 3900
rect 115095 3860 115135 3900
rect 115205 3860 115245 3900
rect 115315 3860 115355 3900
rect 116980 3810 117020 3850
rect 109260 3390 109300 3730
rect 109370 3390 109410 3730
rect 109480 3390 109520 3730
rect 109590 3390 109630 3730
rect 109700 3390 109740 3730
rect 109810 3390 109850 3730
rect 109920 3390 109960 3730
rect 110030 3390 110070 3730
rect 110140 3390 110180 3730
rect 110250 3390 110290 3730
rect 110360 3390 110400 3730
rect 110470 3390 110510 3730
rect 110580 3390 110620 3730
rect 112080 3540 112120 3780
rect 112190 3540 112230 3780
rect 112300 3540 112340 3780
rect 112410 3540 112450 3780
rect 112520 3540 112560 3780
rect 112630 3540 112670 3780
rect 112740 3540 112780 3780
rect 112850 3540 112890 3780
rect 112960 3540 113000 3780
rect 113070 3540 113110 3780
rect 113180 3540 113220 3780
rect 113290 3540 113330 3780
rect 113400 3540 113440 3780
rect 114160 3540 114200 3780
rect 114270 3540 114310 3780
rect 114380 3540 114420 3780
rect 114490 3540 114530 3780
rect 114600 3540 114640 3780
rect 114710 3540 114750 3780
rect 114820 3540 114860 3780
rect 114930 3540 114970 3780
rect 115040 3540 115080 3780
rect 115150 3540 115190 3780
rect 115260 3540 115300 3780
rect 115370 3540 115410 3780
rect 118300 3810 118340 3850
rect 115480 3540 115520 3780
rect 112080 3420 112120 3460
rect 113400 3420 113440 3460
rect 114160 3420 114200 3460
rect 115480 3420 115520 3460
rect 116980 3390 117020 3730
rect 117090 3390 117130 3730
rect 117200 3390 117240 3730
rect 117310 3390 117350 3730
rect 117420 3390 117460 3730
rect 117530 3390 117570 3730
rect 117640 3390 117680 3730
rect 117750 3390 117790 3730
rect 117860 3390 117900 3730
rect 117970 3390 118010 3730
rect 118080 3390 118120 3730
rect 118190 3390 118230 3730
rect 118300 3390 118340 3730
rect 109480 3270 109520 3310
rect 109700 3270 109740 3310
rect 109920 3270 109960 3310
rect 110140 3270 110180 3310
rect 110360 3270 110400 3310
rect 117200 3270 117240 3310
rect 117420 3270 117460 3310
rect 117640 3270 117680 3310
rect 117860 3270 117900 3310
rect 118080 3270 118120 3310
rect 110250 3140 110290 3180
rect 110250 3060 110290 3100
rect 117310 3140 117350 3180
rect 117310 3060 117350 3100
rect 108520 2260 108570 2310
rect 108640 2260 108690 2310
rect 108760 2260 108810 2310
rect 108880 2260 108930 2310
rect 109260 2310 109300 2850
rect 109370 2310 109410 2850
rect 109480 2310 109520 2850
rect 109590 2310 109630 2850
rect 109700 2310 109740 2850
rect 109810 2310 109850 2850
rect 109920 2310 109960 2850
rect 110030 2310 110070 2850
rect 110140 2310 110180 2850
rect 110250 2310 110290 2850
rect 110360 2310 110400 2850
rect 110470 2310 110510 2850
rect 110580 2310 110620 2850
rect 112090 2540 112130 2580
rect 113390 2560 113430 2600
rect 113690 2560 113730 2600
rect 113870 2560 113910 2600
rect 114170 2560 114210 2600
rect 115470 2540 115510 2580
rect 109260 2190 109300 2230
rect 110580 2190 110620 2230
rect 112080 2170 112120 2410
rect 112190 2170 112230 2410
rect 112300 2170 112340 2410
rect 112410 2170 112450 2410
rect 112520 2170 112560 2410
rect 112630 2170 112670 2410
rect 112740 2170 112780 2410
rect 112850 2170 112890 2410
rect 112960 2170 113000 2410
rect 113070 2170 113110 2410
rect 113180 2170 113220 2410
rect 113290 2170 113330 2410
rect 113400 2170 113440 2410
rect 113560 2170 113600 2410
rect 113670 2170 113710 2410
rect 113780 2170 113820 2410
rect 113890 2170 113930 2410
rect 114000 2170 114040 2410
rect 114160 2170 114200 2410
rect 114270 2170 114310 2410
rect 114380 2170 114420 2410
rect 114490 2170 114530 2410
rect 114600 2170 114640 2410
rect 114710 2170 114750 2410
rect 114820 2170 114860 2410
rect 114930 2170 114970 2410
rect 115040 2170 115080 2410
rect 115150 2170 115190 2410
rect 115260 2170 115300 2410
rect 115370 2170 115410 2410
rect 115480 2170 115520 2410
rect 116980 2310 117020 2850
rect 117090 2310 117130 2850
rect 117200 2310 117240 2850
rect 117310 2310 117350 2850
rect 117420 2310 117460 2850
rect 117530 2310 117570 2850
rect 117640 2310 117680 2850
rect 117750 2310 117790 2850
rect 117860 2310 117900 2850
rect 117970 2310 118010 2850
rect 118080 2310 118120 2850
rect 118190 2310 118230 2850
rect 118300 2310 118340 2850
rect 118670 2260 118720 2310
rect 116980 2190 117020 2230
rect 118790 2260 118840 2310
rect 118910 2260 118960 2310
rect 119030 2260 119080 2310
rect 118300 2190 118340 2230
rect 112080 2050 112120 2090
rect 113480 2050 113520 2090
rect 114080 2050 114120 2090
rect 115480 2050 115520 2090
rect 113670 960 113710 1000
rect 113890 960 113930 1000
rect 109620 720 109660 760
rect 109820 720 109860 760
rect 110020 720 110060 760
rect 110220 720 110260 760
rect 108660 600 108710 650
rect 108780 600 108830 650
rect 109320 -690 109360 650
rect 109520 -690 109560 650
rect 109720 -690 109760 650
rect 109920 -690 109960 650
rect 110120 -690 110160 650
rect 110320 -690 110360 650
rect 110520 -690 110560 650
rect 112460 440 112500 880
rect 112570 440 112610 880
rect 112680 440 112720 880
rect 112790 440 112830 880
rect 112900 440 112940 880
rect 113010 440 113050 880
rect 113120 440 113160 880
rect 113230 440 113270 880
rect 113340 440 113380 880
rect 113450 440 113490 880
rect 113560 440 113600 880
rect 113670 440 113710 880
rect 113780 440 113820 880
rect 113890 440 113930 880
rect 114000 440 114040 880
rect 114110 440 114150 880
rect 114220 440 114260 880
rect 114330 440 114370 880
rect 114440 440 114480 880
rect 114550 440 114590 880
rect 114660 440 114700 880
rect 114770 440 114810 880
rect 114880 440 114920 880
rect 114990 440 115030 880
rect 117340 720 117380 760
rect 117540 720 117580 760
rect 117740 720 117780 760
rect 117940 720 117980 760
rect 112460 320 112500 360
rect 114990 320 115030 360
rect 114850 -60 114890 -20
rect 113210 -550 113250 -510
rect 114100 -550 114140 -510
rect 109320 -810 109360 -770
rect 110520 -810 110560 -770
rect 112880 -870 112920 -630
rect 112990 -870 113030 -630
rect 113100 -870 113140 -630
rect 113210 -870 113250 -630
rect 113320 -870 113360 -630
rect 113430 -870 113470 -630
rect 113540 -870 113580 -630
rect 113760 -870 113800 -630
rect 114440 -850 114480 -650
rect 117040 -690 117080 650
rect 117240 -690 117280 650
rect 117440 -690 117480 650
rect 117640 -690 117680 650
rect 117840 -690 117880 650
rect 118040 -690 118080 650
rect 118240 -690 118280 650
rect 118770 600 118820 650
rect 118890 600 118940 650
rect 117040 -810 117080 -770
rect 118240 -810 118280 -770
rect 112880 -990 112920 -950
rect 113540 -990 113580 -950
rect 114100 -990 114140 -950
<< metal1 >>
rect 104580 8640 104820 12220
rect 104580 8580 104590 8640
rect 104650 8580 104670 8640
rect 104730 8580 104750 8640
rect 104810 8580 104820 8640
rect 104580 8560 104820 8580
rect 104580 8500 104590 8560
rect 104650 8500 104670 8560
rect 104730 8500 104750 8560
rect 104810 8500 104820 8560
rect 104580 8480 104820 8500
rect 104580 8420 104590 8480
rect 104650 8420 104670 8480
rect 104730 8420 104750 8480
rect 104810 8420 104820 8480
rect 104580 8410 104820 8420
rect 105280 8640 105520 12220
rect 105280 8580 105290 8640
rect 105350 8580 105370 8640
rect 105430 8580 105450 8640
rect 105510 8580 105520 8640
rect 105280 8560 105520 8580
rect 105280 8500 105290 8560
rect 105350 8500 105370 8560
rect 105430 8500 105450 8560
rect 105510 8500 105520 8560
rect 105280 8480 105520 8500
rect 105280 8420 105290 8480
rect 105350 8420 105370 8480
rect 105430 8420 105450 8480
rect 105510 8420 105520 8480
rect 105280 8410 105520 8420
rect 105980 8640 106220 12220
rect 105980 8580 105990 8640
rect 106050 8580 106070 8640
rect 106130 8580 106150 8640
rect 106210 8580 106220 8640
rect 105980 8560 106220 8580
rect 105980 8500 105990 8560
rect 106050 8500 106070 8560
rect 106130 8500 106150 8560
rect 106210 8500 106220 8560
rect 105980 8480 106220 8500
rect 105980 8420 105990 8480
rect 106050 8420 106070 8480
rect 106130 8420 106150 8480
rect 106210 8420 106220 8480
rect 105980 8410 106220 8420
rect 106680 8640 106920 12220
rect 106680 8580 106690 8640
rect 106750 8580 106770 8640
rect 106830 8580 106850 8640
rect 106910 8580 106920 8640
rect 106680 8560 106920 8580
rect 106680 8500 106690 8560
rect 106750 8500 106770 8560
rect 106830 8500 106850 8560
rect 106910 8500 106920 8560
rect 106680 8480 106920 8500
rect 106680 8420 106690 8480
rect 106750 8420 106770 8480
rect 106830 8420 106850 8480
rect 106910 8420 106920 8480
rect 106680 8410 106920 8420
rect 108080 8640 108320 12220
rect 112410 10130 112490 10140
rect 112410 10070 112420 10130
rect 112480 10070 112490 10130
rect 112170 9860 112250 9870
rect 112170 9800 112180 9860
rect 112240 9800 112250 9860
rect 112170 9790 112250 9800
rect 112410 9860 112490 10070
rect 113350 10130 113430 10140
rect 113350 10070 113360 10130
rect 113420 10070 113430 10130
rect 113350 10060 113430 10070
rect 114170 10130 114250 10140
rect 114170 10070 114180 10130
rect 114240 10070 114250 10130
rect 114170 10060 114250 10070
rect 115110 10130 115190 10140
rect 115110 10070 115120 10130
rect 115180 10070 115190 10130
rect 112410 9800 112420 9860
rect 112480 9800 112490 9860
rect 112410 9790 112490 9800
rect 112530 9860 112610 9870
rect 112530 9800 112540 9860
rect 112600 9800 112610 9860
rect 112530 9790 112610 9800
rect 112180 9730 112240 9790
rect 112180 9090 112190 9730
rect 112230 9090 112240 9730
rect 112180 9070 112240 9090
rect 112300 9730 112360 9750
rect 112300 9090 112310 9730
rect 112350 9090 112360 9730
rect 112300 8970 112360 9090
rect 112420 9730 112480 9790
rect 112420 9090 112430 9730
rect 112470 9090 112480 9730
rect 112420 9060 112480 9090
rect 112540 9730 112600 9790
rect 112540 9090 112550 9730
rect 112590 9090 112600 9730
rect 113110 9680 113190 9690
rect 113110 9620 113120 9680
rect 113180 9620 113190 9680
rect 113110 9600 113190 9620
rect 113110 9540 113120 9600
rect 113180 9540 113190 9600
rect 113110 9520 113190 9540
rect 113110 9460 113120 9520
rect 113180 9460 113190 9520
rect 113110 9450 113190 9460
rect 113230 9680 113310 9690
rect 113230 9620 113240 9680
rect 113300 9620 113310 9680
rect 113230 9600 113310 9620
rect 113230 9540 113240 9600
rect 113300 9540 113310 9600
rect 113230 9520 113310 9540
rect 113230 9460 113240 9520
rect 113300 9460 113310 9520
rect 113230 9450 113310 9460
rect 112540 9070 112600 9090
rect 113120 9390 113180 9450
rect 113120 9090 113130 9390
rect 113170 9090 113180 9390
rect 113120 9070 113180 9090
rect 113240 9390 113300 9450
rect 113240 9090 113250 9390
rect 113290 9090 113300 9390
rect 113240 9070 113300 9090
rect 113360 9390 113420 10060
rect 113760 10020 113840 10030
rect 113760 9960 113770 10020
rect 113830 9960 113840 10020
rect 113760 9940 113840 9960
rect 113760 9880 113770 9940
rect 113830 9880 113840 9940
rect 113760 9860 113840 9880
rect 113760 9800 113770 9860
rect 113830 9800 113840 9860
rect 113470 9680 113550 9690
rect 113470 9620 113480 9680
rect 113540 9620 113550 9680
rect 113470 9600 113550 9620
rect 113470 9540 113480 9600
rect 113540 9540 113550 9600
rect 113470 9520 113550 9540
rect 113470 9460 113480 9520
rect 113540 9460 113550 9520
rect 113470 9450 113550 9460
rect 113760 9680 113840 9800
rect 114050 10020 114130 10030
rect 114050 9960 114060 10020
rect 114120 9960 114130 10020
rect 114050 9940 114130 9960
rect 114050 9880 114060 9940
rect 114120 9880 114130 9940
rect 114050 9860 114130 9880
rect 114050 9800 114060 9860
rect 114120 9800 114130 9860
rect 114050 9790 114130 9800
rect 113760 9620 113770 9680
rect 113830 9620 113840 9680
rect 113760 9600 113840 9620
rect 113760 9540 113770 9600
rect 113830 9540 113840 9600
rect 113760 9520 113840 9540
rect 113760 9460 113770 9520
rect 113830 9460 113840 9520
rect 113360 9090 113370 9390
rect 113410 9090 113420 9390
rect 113360 9060 113420 9090
rect 113480 9390 113540 9450
rect 113480 9090 113490 9390
rect 113530 9090 113540 9390
rect 113480 9070 113540 9090
rect 112410 9050 112490 9060
rect 112410 8990 112420 9050
rect 112480 8990 112490 9050
rect 112410 8980 112490 8990
rect 113350 9050 113430 9060
rect 113350 8990 113360 9050
rect 113420 8990 113430 9050
rect 113350 8980 113430 8990
rect 112300 8960 112380 8970
rect 112300 8900 112310 8960
rect 112370 8900 112380 8960
rect 112300 8890 112380 8900
rect 113260 8960 113320 8970
rect 113260 8890 113320 8900
rect 113650 8960 113730 8970
rect 113650 8900 113660 8960
rect 113720 8900 113730 8960
rect 113650 8890 113730 8900
rect 108080 8580 108090 8640
rect 108150 8580 108170 8640
rect 108230 8580 108250 8640
rect 108310 8580 108320 8640
rect 108080 8560 108320 8580
rect 108080 8500 108090 8560
rect 108150 8500 108170 8560
rect 108230 8500 108250 8560
rect 108310 8500 108320 8560
rect 108080 8480 108320 8500
rect 108080 8420 108090 8480
rect 108150 8420 108170 8480
rect 108230 8420 108250 8480
rect 108310 8420 108320 8480
rect 108080 8410 108320 8420
rect 109180 8640 109260 8650
rect 109180 8580 109190 8640
rect 109250 8580 109260 8640
rect 109180 8560 109260 8580
rect 109180 8500 109190 8560
rect 109250 8500 109260 8560
rect 109180 8480 109260 8500
rect 109180 8420 109190 8480
rect 109250 8420 109260 8480
rect 109180 7860 109260 8420
rect 109900 8640 109980 8650
rect 109900 8580 109910 8640
rect 109970 8580 109980 8640
rect 109900 8560 109980 8580
rect 109900 8500 109910 8560
rect 109970 8500 109980 8560
rect 109900 8480 109980 8500
rect 109900 8420 109910 8480
rect 109970 8420 109980 8480
rect 109300 8370 109380 8380
rect 109300 8310 109310 8370
rect 109370 8310 109380 8370
rect 109300 8290 109380 8310
rect 109300 8230 109310 8290
rect 109370 8230 109380 8290
rect 109300 8210 109380 8230
rect 109300 8150 109310 8210
rect 109370 8150 109380 8210
rect 109300 8130 109380 8150
rect 109300 8070 109310 8130
rect 109370 8070 109380 8130
rect 109300 8050 109380 8070
rect 109300 7990 109310 8050
rect 109370 7990 109380 8050
rect 109300 7970 109380 7990
rect 109300 7910 109310 7970
rect 109370 7910 109380 7970
rect 109300 7900 109380 7910
rect 109540 8370 109620 8380
rect 109540 8310 109550 8370
rect 109610 8310 109620 8370
rect 109540 8290 109620 8310
rect 109540 8230 109550 8290
rect 109610 8230 109620 8290
rect 109540 8210 109620 8230
rect 109540 8150 109550 8210
rect 109610 8150 109620 8210
rect 109540 8130 109620 8150
rect 109540 8070 109550 8130
rect 109610 8070 109620 8130
rect 109540 8050 109620 8070
rect 109540 7990 109550 8050
rect 109610 7990 109620 8050
rect 109540 7970 109620 7990
rect 109540 7910 109550 7970
rect 109610 7910 109620 7970
rect 109540 7900 109620 7910
rect 109780 8370 109860 8380
rect 109780 8310 109790 8370
rect 109850 8310 109860 8370
rect 109780 8290 109860 8310
rect 109780 8230 109790 8290
rect 109850 8230 109860 8290
rect 109780 8210 109860 8230
rect 109780 8150 109790 8210
rect 109850 8150 109860 8210
rect 109780 8130 109860 8150
rect 109780 8070 109790 8130
rect 109850 8070 109860 8130
rect 109780 8050 109860 8070
rect 109780 7990 109790 8050
rect 109850 7990 109860 8050
rect 109780 7970 109860 7990
rect 109780 7910 109790 7970
rect 109850 7910 109860 7970
rect 109780 7900 109860 7910
rect 109180 7800 109190 7860
rect 109250 7800 109260 7860
rect 109180 7790 109260 7800
rect 109190 7730 109250 7790
rect 109190 7090 109200 7730
rect 109240 7090 109250 7730
rect 109190 7070 109250 7090
rect 109310 7730 109370 7900
rect 109420 7860 109500 7870
rect 109420 7800 109430 7860
rect 109490 7800 109500 7860
rect 109420 7790 109500 7800
rect 109310 7090 109320 7730
rect 109360 7090 109370 7730
rect 109310 7060 109370 7090
rect 109430 7730 109490 7790
rect 109430 7090 109440 7730
rect 109480 7090 109490 7730
rect 109430 7070 109490 7090
rect 109550 7730 109610 7900
rect 109660 7860 109740 7870
rect 109660 7800 109670 7860
rect 109730 7800 109740 7860
rect 109660 7790 109740 7800
rect 109550 7090 109560 7730
rect 109600 7090 109610 7730
rect 109550 7060 109610 7090
rect 109670 7730 109730 7790
rect 109670 7090 109680 7730
rect 109720 7090 109730 7730
rect 109670 7070 109730 7090
rect 109790 7730 109850 7900
rect 109900 7860 109980 8420
rect 110620 8640 110700 8650
rect 110620 8580 110630 8640
rect 110690 8580 110700 8640
rect 110620 8560 110700 8580
rect 110620 8500 110630 8560
rect 110690 8500 110700 8560
rect 110620 8480 110700 8500
rect 110620 8420 110630 8480
rect 110690 8420 110700 8480
rect 110020 8370 110100 8380
rect 110020 8310 110030 8370
rect 110090 8310 110100 8370
rect 110020 8290 110100 8310
rect 110020 8230 110030 8290
rect 110090 8230 110100 8290
rect 110020 8210 110100 8230
rect 110020 8150 110030 8210
rect 110090 8150 110100 8210
rect 110020 8130 110100 8150
rect 110020 8070 110030 8130
rect 110090 8070 110100 8130
rect 110020 8050 110100 8070
rect 110020 7990 110030 8050
rect 110090 7990 110100 8050
rect 110020 7970 110100 7990
rect 110020 7910 110030 7970
rect 110090 7910 110100 7970
rect 110020 7900 110100 7910
rect 110260 8370 110340 8380
rect 110260 8310 110270 8370
rect 110330 8310 110340 8370
rect 110260 8290 110340 8310
rect 110260 8230 110270 8290
rect 110330 8230 110340 8290
rect 110260 8210 110340 8230
rect 110260 8150 110270 8210
rect 110330 8150 110340 8210
rect 110260 8130 110340 8150
rect 110260 8070 110270 8130
rect 110330 8070 110340 8130
rect 110260 8050 110340 8070
rect 110260 7990 110270 8050
rect 110330 7990 110340 8050
rect 110260 7970 110340 7990
rect 110260 7910 110270 7970
rect 110330 7910 110340 7970
rect 110260 7900 110340 7910
rect 110500 8370 110580 8380
rect 110500 8310 110510 8370
rect 110570 8310 110580 8370
rect 110500 8290 110580 8310
rect 110500 8230 110510 8290
rect 110570 8230 110580 8290
rect 110500 8210 110580 8230
rect 110500 8150 110510 8210
rect 110570 8150 110580 8210
rect 110500 8130 110580 8150
rect 110500 8070 110510 8130
rect 110570 8070 110580 8130
rect 110500 8050 110580 8070
rect 110500 7990 110510 8050
rect 110570 7990 110580 8050
rect 110500 7970 110580 7990
rect 110500 7910 110510 7970
rect 110570 7910 110580 7970
rect 110500 7900 110580 7910
rect 109900 7800 109910 7860
rect 109970 7800 109980 7860
rect 109900 7790 109980 7800
rect 109790 7090 109800 7730
rect 109840 7090 109850 7730
rect 109790 7060 109850 7090
rect 109910 7730 109970 7790
rect 109910 7090 109920 7730
rect 109960 7090 109970 7730
rect 109910 7070 109970 7090
rect 110030 7730 110090 7900
rect 110140 7860 110220 7870
rect 110140 7800 110150 7860
rect 110210 7800 110220 7860
rect 110140 7790 110220 7800
rect 110030 7090 110040 7730
rect 110080 7090 110090 7730
rect 110030 7060 110090 7090
rect 110150 7730 110210 7790
rect 110150 7090 110160 7730
rect 110200 7090 110210 7730
rect 110150 7070 110210 7090
rect 110270 7730 110330 7900
rect 110380 7860 110460 7870
rect 110380 7800 110390 7860
rect 110450 7800 110460 7860
rect 110380 7790 110460 7800
rect 110270 7090 110280 7730
rect 110320 7090 110330 7730
rect 110270 7060 110330 7090
rect 110390 7730 110450 7790
rect 110390 7090 110400 7730
rect 110440 7090 110450 7730
rect 110390 7070 110450 7090
rect 110510 7730 110570 7900
rect 110620 7860 110700 8420
rect 110620 7800 110630 7860
rect 110690 7800 110700 7860
rect 110620 7790 110700 7800
rect 111070 8640 111310 8650
rect 111070 8580 111080 8640
rect 111140 8580 111160 8640
rect 111220 8580 111240 8640
rect 111300 8580 111310 8640
rect 111070 8560 111310 8580
rect 111070 8500 111080 8560
rect 111140 8500 111160 8560
rect 111220 8500 111240 8560
rect 111300 8500 111310 8560
rect 111070 8480 111310 8500
rect 111070 8420 111080 8480
rect 111140 8420 111160 8480
rect 111220 8420 111240 8480
rect 111300 8420 111310 8480
rect 110510 7090 110520 7730
rect 110560 7090 110570 7730
rect 110510 7060 110570 7090
rect 110630 7730 110690 7790
rect 110630 7090 110640 7730
rect 110680 7090 110690 7730
rect 110630 7070 110690 7090
rect 109300 7050 109380 7060
rect 109300 6990 109310 7050
rect 109370 6990 109380 7050
rect 109300 6980 109380 6990
rect 109540 7050 109620 7060
rect 109540 6990 109550 7050
rect 109610 6990 109620 7050
rect 109540 6980 109620 6990
rect 109780 7050 109860 7060
rect 109780 6990 109790 7050
rect 109850 6990 109860 7050
rect 109780 6980 109860 6990
rect 110020 7050 110100 7060
rect 110020 6990 110030 7050
rect 110090 6990 110100 7050
rect 110020 6980 110100 6990
rect 110260 7050 110340 7060
rect 110260 6990 110270 7050
rect 110330 6990 110340 7050
rect 110260 6980 110340 6990
rect 110500 7050 110580 7060
rect 110500 6990 110510 7050
rect 110570 6990 110580 7050
rect 110500 6980 110580 6990
rect 110800 7050 111040 7060
rect 110800 6990 110810 7050
rect 110870 6990 110890 7050
rect 110950 6990 110970 7050
rect 111030 6990 111040 7050
rect 109370 6940 109430 6950
rect 109370 6870 109430 6880
rect 109490 6940 109550 6950
rect 109490 6870 109550 6880
rect 109610 6940 109670 6950
rect 109610 6870 109670 6880
rect 109730 6940 109790 6950
rect 109730 6870 109790 6880
rect 109850 6940 110030 6950
rect 109910 6880 109970 6940
rect 109850 6870 110030 6880
rect 110090 6940 110150 6950
rect 110090 6870 110150 6880
rect 110210 6940 110270 6950
rect 110210 6870 110270 6880
rect 110330 6940 110390 6950
rect 110330 6870 110390 6880
rect 110450 6940 110510 6950
rect 110450 6870 110510 6880
rect 109900 6820 109980 6870
rect 109900 6760 109910 6820
rect 109970 6760 109980 6820
rect 108510 6750 108590 6760
rect 109900 6750 109980 6760
rect 108510 6690 108520 6750
rect 108580 6690 108590 6750
rect 108510 6400 108590 6690
rect 109240 6710 109320 6720
rect 109240 6650 109250 6710
rect 109310 6650 109320 6710
rect 109240 6630 109320 6650
rect 109240 6570 109250 6630
rect 109310 6570 109320 6630
rect 109240 6550 109320 6570
rect 109240 6490 109250 6550
rect 109310 6490 109320 6550
rect 109240 6480 109320 6490
rect 109460 6710 109540 6720
rect 109460 6650 109470 6710
rect 109530 6650 109540 6710
rect 109460 6630 109540 6650
rect 109460 6570 109470 6630
rect 109530 6570 109540 6630
rect 109460 6550 109540 6570
rect 109460 6490 109470 6550
rect 109530 6490 109540 6550
rect 109460 6480 109540 6490
rect 109680 6710 109760 6720
rect 109680 6650 109690 6710
rect 109750 6650 109760 6710
rect 109680 6630 109760 6650
rect 109680 6570 109690 6630
rect 109750 6570 109760 6630
rect 109680 6550 109760 6570
rect 109680 6490 109690 6550
rect 109750 6490 109760 6550
rect 109680 6480 109760 6490
rect 109900 6710 109980 6720
rect 109900 6650 109910 6710
rect 109970 6650 109980 6710
rect 109900 6630 109980 6650
rect 109900 6570 109910 6630
rect 109970 6570 109980 6630
rect 109900 6550 109980 6570
rect 109900 6490 109910 6550
rect 109970 6490 109980 6550
rect 109900 6480 109980 6490
rect 110120 6710 110200 6720
rect 110120 6650 110130 6710
rect 110190 6650 110200 6710
rect 110120 6630 110200 6650
rect 110120 6570 110130 6630
rect 110190 6570 110200 6630
rect 110120 6550 110200 6570
rect 110120 6490 110130 6550
rect 110190 6490 110200 6550
rect 110120 6480 110200 6490
rect 110340 6710 110420 6720
rect 110340 6650 110350 6710
rect 110410 6650 110420 6710
rect 110340 6630 110420 6650
rect 110340 6570 110350 6630
rect 110410 6570 110420 6630
rect 110340 6550 110420 6570
rect 110340 6490 110350 6550
rect 110410 6490 110420 6550
rect 110340 6480 110420 6490
rect 110560 6710 110640 6720
rect 110560 6650 110570 6710
rect 110630 6650 110640 6710
rect 110560 6630 110640 6650
rect 110560 6570 110570 6630
rect 110630 6570 110640 6630
rect 110560 6550 110640 6570
rect 110560 6490 110570 6550
rect 110630 6490 110640 6550
rect 110560 6480 110640 6490
rect 109250 6400 109310 6480
rect 108408 6380 108690 6400
rect 108408 6340 108420 6380
rect 108460 6340 108530 6380
rect 108570 6340 108640 6380
rect 108680 6340 108690 6380
rect 108408 6320 108690 6340
rect 109250 6360 109260 6400
rect 109300 6360 109310 6400
rect 109250 6280 109310 6360
rect 109350 6380 109430 6390
rect 109350 6320 109360 6380
rect 109420 6320 109430 6380
rect 109350 6310 109430 6320
rect 108408 5170 108690 5190
rect 108408 5130 108420 5170
rect 108460 5130 108530 5170
rect 108570 5130 108640 5170
rect 108680 5130 108690 5170
rect 108408 5110 108690 5130
rect 109250 5140 109260 6280
rect 109300 5140 109310 6280
rect 109250 5120 109310 5140
rect 109360 6280 109420 6310
rect 109360 5140 109370 6280
rect 109410 5140 109420 6280
rect 109360 5110 109420 5140
rect 109470 6280 109530 6480
rect 109570 6380 109650 6390
rect 109570 6320 109580 6380
rect 109640 6320 109650 6380
rect 109570 6310 109650 6320
rect 109470 5140 109480 6280
rect 109520 5140 109530 6280
rect 109470 5120 109530 5140
rect 109580 6280 109640 6310
rect 109580 5140 109590 6280
rect 109630 5140 109640 6280
rect 109580 5110 109640 5140
rect 109690 6280 109750 6480
rect 109790 6380 109870 6390
rect 109790 6320 109800 6380
rect 109860 6320 109870 6380
rect 109790 6310 109870 6320
rect 109690 5140 109700 6280
rect 109740 5140 109750 6280
rect 109690 5120 109750 5140
rect 109800 6280 109860 6310
rect 109800 5140 109810 6280
rect 109850 5140 109860 6280
rect 109800 5110 109860 5140
rect 109910 6280 109970 6480
rect 110010 6380 110090 6390
rect 110010 6320 110020 6380
rect 110080 6320 110090 6380
rect 110010 6310 110090 6320
rect 109910 5140 109920 6280
rect 109960 5140 109970 6280
rect 109910 5120 109970 5140
rect 110020 6280 110080 6310
rect 110020 5140 110030 6280
rect 110070 5140 110080 6280
rect 110020 5110 110080 5140
rect 110130 6280 110190 6480
rect 110230 6380 110310 6390
rect 110230 6320 110240 6380
rect 110300 6320 110310 6380
rect 110230 6310 110310 6320
rect 110130 5140 110140 6280
rect 110180 5140 110190 6280
rect 110130 5120 110190 5140
rect 110240 6280 110300 6310
rect 110240 5140 110250 6280
rect 110290 5140 110300 6280
rect 110240 5110 110300 5140
rect 110350 6280 110410 6480
rect 110570 6400 110630 6480
rect 110450 6380 110530 6390
rect 110450 6320 110460 6380
rect 110520 6320 110530 6380
rect 110450 6310 110530 6320
rect 110570 6360 110580 6400
rect 110620 6360 110630 6400
rect 110350 5140 110360 6280
rect 110400 5140 110410 6280
rect 110350 5120 110410 5140
rect 110460 6280 110520 6310
rect 110460 5140 110470 6280
rect 110510 5140 110520 6280
rect 110460 5110 110520 5140
rect 110570 6280 110630 6360
rect 110570 5140 110580 6280
rect 110620 5140 110630 6280
rect 110570 5120 110630 5140
rect 108430 4940 108670 5110
rect 108430 4880 108440 4940
rect 108500 4880 108520 4940
rect 108580 4880 108600 4940
rect 108660 4880 108670 4940
rect 108430 4860 108670 4880
rect 108430 4800 108440 4860
rect 108500 4800 108520 4860
rect 108580 4800 108600 4860
rect 108660 4800 108670 4860
rect 108430 4780 108670 4800
rect 108430 4720 108440 4780
rect 108500 4720 108520 4780
rect 108580 4720 108600 4780
rect 108660 4720 108670 4780
rect 108430 4710 108670 4720
rect 109350 5100 109430 5110
rect 109350 5040 109360 5100
rect 109420 5040 109430 5100
rect 109350 4650 109430 5040
rect 109570 5100 109650 5110
rect 109570 5040 109580 5100
rect 109640 5040 109650 5100
rect 109570 4650 109650 5040
rect 109790 5100 109870 5110
rect 109790 5040 109800 5100
rect 109860 5040 109870 5100
rect 109790 4650 109870 5040
rect 110010 5100 110090 5110
rect 110010 5040 110020 5100
rect 110080 5040 110090 5100
rect 109900 4940 109980 4950
rect 109900 4880 109910 4940
rect 109970 4880 109980 4940
rect 109900 4860 109980 4880
rect 109900 4800 109910 4860
rect 109970 4800 109980 4860
rect 109900 4780 109980 4800
rect 109900 4720 109910 4780
rect 109970 4720 109980 4780
rect 109900 4710 109980 4720
rect 110010 4650 110090 5040
rect 110230 5100 110310 5110
rect 110230 5040 110240 5100
rect 110300 5040 110310 5100
rect 110230 4650 110310 5040
rect 110450 5100 110530 5110
rect 110450 5040 110460 5100
rect 110520 5040 110530 5100
rect 110450 4650 110530 5040
rect 107980 4640 108480 4650
rect 107980 4580 107990 4640
rect 108050 4580 108070 4640
rect 108130 4580 108160 4640
rect 108220 4580 108240 4640
rect 108300 4580 108330 4640
rect 108390 4580 108410 4640
rect 108470 4580 108480 4640
rect 107980 4560 108480 4580
rect 107980 4500 107990 4560
rect 108050 4500 108070 4560
rect 108130 4500 108160 4560
rect 108220 4500 108240 4560
rect 108300 4500 108330 4560
rect 108390 4500 108410 4560
rect 108470 4500 108480 4560
rect 107980 4480 108480 4500
rect 107980 4420 107990 4480
rect 108050 4420 108070 4480
rect 108130 4420 108160 4480
rect 108220 4420 108240 4480
rect 108300 4420 108330 4480
rect 108390 4420 108410 4480
rect 108470 4420 108480 4480
rect 107680 4100 107920 4110
rect 107680 4040 107690 4100
rect 107750 4040 107770 4100
rect 107830 4040 107850 4100
rect 107910 4040 107920 4100
rect 107680 4020 107920 4040
rect 107680 3960 107690 4020
rect 107750 3960 107770 4020
rect 107830 3960 107850 4020
rect 107910 3960 107920 4020
rect 107680 3940 107920 3960
rect 107680 3880 107690 3940
rect 107750 3880 107770 3940
rect 107830 3880 107850 3940
rect 107910 3880 107920 3940
rect 107680 1880 107920 3880
rect 107680 1820 107690 1880
rect 107750 1820 107770 1880
rect 107830 1820 107850 1880
rect 107910 1820 107920 1880
rect 107680 1800 107920 1820
rect 107680 1740 107690 1800
rect 107750 1740 107770 1800
rect 107830 1740 107850 1800
rect 107910 1740 107920 1800
rect 107680 1720 107920 1740
rect 107680 1660 107690 1720
rect 107750 1660 107770 1720
rect 107830 1660 107850 1720
rect 107910 1660 107920 1720
rect 104580 -1160 104820 -1150
rect 104580 -1220 104590 -1160
rect 104650 -1220 104670 -1160
rect 104730 -1220 104750 -1160
rect 104810 -1220 104820 -1160
rect 104580 -1240 104820 -1220
rect 104580 -1300 104590 -1240
rect 104650 -1300 104670 -1240
rect 104730 -1300 104750 -1240
rect 104810 -1300 104820 -1240
rect 104580 -1320 104820 -1300
rect 104580 -1380 104590 -1320
rect 104650 -1380 104670 -1320
rect 104730 -1380 104750 -1320
rect 104810 -1380 104820 -1320
rect 104580 -3000 104820 -1380
rect 105280 -1160 105520 -1150
rect 105280 -1220 105290 -1160
rect 105350 -1220 105370 -1160
rect 105430 -1220 105450 -1160
rect 105510 -1220 105520 -1160
rect 105280 -1240 105520 -1220
rect 105280 -1300 105290 -1240
rect 105350 -1300 105370 -1240
rect 105430 -1300 105450 -1240
rect 105510 -1300 105520 -1240
rect 105280 -1320 105520 -1300
rect 105280 -1380 105290 -1320
rect 105350 -1380 105370 -1320
rect 105430 -1380 105450 -1320
rect 105510 -1380 105520 -1320
rect 105280 -3000 105520 -1380
rect 105980 -1160 106220 -1150
rect 105980 -1220 105990 -1160
rect 106050 -1220 106070 -1160
rect 106130 -1220 106150 -1160
rect 106210 -1220 106220 -1160
rect 105980 -1240 106220 -1220
rect 105980 -1300 105990 -1240
rect 106050 -1300 106070 -1240
rect 106130 -1300 106150 -1240
rect 106210 -1300 106220 -1240
rect 105980 -1320 106220 -1300
rect 105980 -1380 105990 -1320
rect 106050 -1380 106070 -1320
rect 106130 -1380 106150 -1320
rect 106210 -1380 106220 -1320
rect 105980 -3000 106220 -1380
rect 106680 -1160 106920 -1150
rect 106680 -1220 106690 -1160
rect 106750 -1220 106770 -1160
rect 106830 -1220 106850 -1160
rect 106910 -1220 106920 -1160
rect 106680 -1240 106920 -1220
rect 106680 -1300 106690 -1240
rect 106750 -1300 106770 -1240
rect 106830 -1300 106850 -1240
rect 106910 -1300 106920 -1240
rect 106680 -1320 106920 -1300
rect 106680 -1380 106690 -1320
rect 106750 -1380 106770 -1320
rect 106830 -1380 106850 -1320
rect 106910 -1380 106920 -1320
rect 106680 -3000 106920 -1380
rect 107380 -1160 107620 -1150
rect 107380 -1220 107390 -1160
rect 107450 -1220 107470 -1160
rect 107530 -1220 107550 -1160
rect 107610 -1220 107620 -1160
rect 107380 -1240 107620 -1220
rect 107380 -1300 107390 -1240
rect 107450 -1300 107470 -1240
rect 107530 -1300 107550 -1240
rect 107610 -1300 107620 -1240
rect 107380 -1320 107620 -1300
rect 107380 -1380 107390 -1320
rect 107450 -1380 107470 -1320
rect 107530 -1380 107550 -1320
rect 107610 -1380 107620 -1320
rect 107380 -3000 107620 -1380
rect 107680 -1160 107920 1660
rect 107980 3420 108480 4420
rect 109350 4640 110530 4650
rect 109350 4580 109360 4640
rect 109420 4580 109470 4640
rect 109530 4580 109580 4640
rect 109640 4580 109690 4640
rect 109750 4580 109800 4640
rect 109860 4580 109910 4640
rect 109970 4580 110020 4640
rect 110080 4580 110130 4640
rect 110190 4580 110240 4640
rect 110300 4580 110350 4640
rect 110410 4580 110460 4640
rect 110520 4580 110530 4640
rect 109350 4560 110530 4580
rect 109350 4500 109360 4560
rect 109420 4500 109470 4560
rect 109530 4500 109580 4560
rect 109640 4500 109690 4560
rect 109750 4500 109800 4560
rect 109860 4500 109910 4560
rect 109970 4500 110020 4560
rect 110080 4500 110130 4560
rect 110190 4500 110240 4560
rect 110300 4500 110350 4560
rect 110410 4500 110460 4560
rect 110520 4500 110530 4560
rect 109350 4480 110530 4500
rect 109350 4420 109360 4480
rect 109420 4420 109470 4480
rect 109530 4420 109580 4480
rect 109640 4420 109690 4480
rect 109750 4420 109800 4480
rect 109860 4420 109910 4480
rect 109970 4420 110020 4480
rect 110080 4420 110130 4480
rect 110190 4420 110240 4480
rect 110300 4420 110350 4480
rect 110410 4420 110460 4480
rect 110520 4420 110530 4480
rect 109350 4410 110530 4420
rect 110800 4940 111040 6990
rect 110800 4880 110810 4940
rect 110870 4880 110890 4940
rect 110950 4880 110970 4940
rect 111030 4880 111040 4940
rect 110800 4860 111040 4880
rect 110800 4800 110810 4860
rect 110870 4800 110890 4860
rect 110950 4800 110970 4860
rect 111030 4800 111040 4860
rect 110800 4780 111040 4800
rect 110800 4720 110810 4780
rect 110870 4720 110890 4780
rect 110950 4720 110970 4780
rect 111030 4720 111040 4780
rect 109240 4370 109320 4380
rect 109240 4310 109250 4370
rect 109310 4310 109320 4370
rect 109240 4290 109320 4310
rect 109240 4230 109250 4290
rect 109310 4230 109320 4290
rect 109240 4210 109320 4230
rect 109240 4150 109250 4210
rect 109310 4150 109320 4210
rect 109240 4140 109320 4150
rect 110560 4370 110640 4380
rect 110560 4310 110570 4370
rect 110630 4310 110640 4370
rect 110560 4290 110640 4310
rect 110560 4230 110570 4290
rect 110630 4230 110640 4290
rect 110560 4210 110640 4230
rect 110560 4150 110570 4210
rect 110630 4150 110640 4210
rect 110560 4140 110640 4150
rect 107980 3360 108000 3420
rect 108060 3360 108100 3420
rect 108160 3360 108200 3420
rect 108260 3360 108300 3420
rect 108360 3360 108400 3420
rect 108460 3360 108480 3420
rect 109250 3850 109310 4140
rect 109350 4100 109430 4110
rect 109350 4040 109360 4100
rect 109420 4040 109430 4100
rect 109350 4020 109430 4040
rect 109350 3960 109360 4020
rect 109420 3960 109430 4020
rect 109350 3940 109430 3960
rect 109350 3880 109360 3940
rect 109420 3880 109430 3940
rect 109350 3870 109430 3880
rect 109570 4100 109650 4110
rect 109570 4040 109580 4100
rect 109640 4040 109650 4100
rect 109570 4020 109650 4040
rect 109570 3960 109580 4020
rect 109640 3960 109650 4020
rect 109570 3940 109650 3960
rect 109570 3880 109580 3940
rect 109640 3880 109650 3940
rect 109570 3870 109650 3880
rect 109790 4100 109870 4110
rect 109790 4040 109800 4100
rect 109860 4040 109870 4100
rect 109790 4020 109870 4040
rect 109790 3960 109800 4020
rect 109860 3960 109870 4020
rect 109790 3940 109870 3960
rect 109790 3880 109800 3940
rect 109860 3880 109870 3940
rect 109790 3870 109870 3880
rect 110010 4100 110090 4110
rect 110010 4040 110020 4100
rect 110080 4040 110090 4100
rect 110010 4020 110090 4040
rect 110010 3960 110020 4020
rect 110080 3960 110090 4020
rect 110010 3940 110090 3960
rect 110010 3880 110020 3940
rect 110080 3880 110090 3940
rect 110010 3870 110090 3880
rect 110230 4100 110310 4110
rect 110230 4040 110240 4100
rect 110300 4040 110310 4100
rect 110230 4020 110310 4040
rect 110230 3960 110240 4020
rect 110300 3960 110310 4020
rect 110230 3940 110310 3960
rect 110230 3880 110240 3940
rect 110300 3880 110310 3940
rect 110230 3870 110310 3880
rect 110450 4100 110530 4110
rect 110450 4040 110460 4100
rect 110520 4040 110530 4100
rect 110450 4020 110530 4040
rect 110450 3960 110460 4020
rect 110520 3960 110530 4020
rect 110450 3940 110530 3960
rect 110450 3880 110460 3940
rect 110520 3880 110530 3940
rect 110450 3870 110530 3880
rect 109250 3810 109260 3850
rect 109300 3810 109310 3850
rect 109250 3730 109310 3810
rect 109250 3390 109260 3730
rect 109300 3390 109310 3730
rect 109250 3370 109310 3390
rect 109360 3730 109420 3870
rect 109460 3830 109540 3840
rect 109460 3770 109470 3830
rect 109530 3770 109540 3830
rect 109460 3760 109540 3770
rect 109360 3390 109370 3730
rect 109410 3390 109420 3730
rect 109360 3370 109420 3390
rect 109470 3730 109530 3760
rect 109470 3390 109480 3730
rect 109520 3390 109530 3730
rect 107980 3320 108480 3360
rect 109470 3330 109530 3390
rect 109580 3730 109640 3870
rect 109680 3830 109760 3840
rect 109680 3770 109690 3830
rect 109750 3770 109760 3830
rect 109680 3760 109760 3770
rect 109580 3390 109590 3730
rect 109630 3390 109640 3730
rect 109580 3370 109640 3390
rect 109690 3730 109750 3760
rect 109690 3390 109700 3730
rect 109740 3390 109750 3730
rect 109690 3330 109750 3390
rect 109800 3730 109860 3870
rect 109900 3830 109980 3840
rect 109900 3770 109910 3830
rect 109970 3770 109980 3830
rect 109900 3760 109980 3770
rect 109800 3390 109810 3730
rect 109850 3390 109860 3730
rect 109800 3370 109860 3390
rect 109910 3730 109970 3760
rect 109910 3390 109920 3730
rect 109960 3390 109970 3730
rect 109910 3330 109970 3390
rect 110020 3730 110080 3870
rect 110120 3830 110200 3840
rect 110120 3770 110130 3830
rect 110190 3770 110200 3830
rect 110120 3760 110200 3770
rect 110020 3390 110030 3730
rect 110070 3390 110080 3730
rect 110020 3370 110080 3390
rect 110130 3730 110190 3760
rect 110130 3390 110140 3730
rect 110180 3390 110190 3730
rect 110130 3330 110190 3390
rect 110240 3730 110300 3870
rect 110340 3830 110420 3840
rect 110340 3770 110350 3830
rect 110410 3770 110420 3830
rect 110340 3760 110420 3770
rect 110240 3390 110250 3730
rect 110290 3390 110300 3730
rect 110240 3370 110300 3390
rect 110350 3730 110410 3760
rect 110350 3390 110360 3730
rect 110400 3390 110410 3730
rect 110350 3330 110410 3390
rect 110460 3730 110520 3870
rect 110460 3390 110470 3730
rect 110510 3390 110520 3730
rect 110460 3370 110520 3390
rect 110570 3850 110630 4140
rect 110570 3810 110580 3850
rect 110620 3810 110630 3850
rect 110570 3730 110630 3810
rect 110570 3390 110580 3730
rect 110620 3390 110630 3730
rect 110570 3370 110630 3390
rect 107980 3260 108000 3320
rect 108060 3260 108100 3320
rect 108160 3260 108200 3320
rect 108260 3260 108300 3320
rect 108360 3260 108400 3320
rect 108460 3260 108480 3320
rect 107980 3220 108480 3260
rect 108970 3320 109050 3330
rect 108970 3260 108980 3320
rect 109040 3260 109050 3320
rect 108970 3250 109050 3260
rect 109460 3320 109540 3330
rect 109460 3260 109470 3320
rect 109530 3260 109540 3320
rect 109460 3250 109540 3260
rect 109680 3320 109760 3330
rect 109680 3260 109690 3320
rect 109750 3260 109760 3320
rect 109680 3250 109760 3260
rect 109900 3320 109980 3330
rect 109900 3260 109910 3320
rect 109970 3260 109980 3320
rect 109900 3250 109980 3260
rect 110120 3320 110200 3330
rect 110120 3260 110130 3320
rect 110190 3260 110200 3320
rect 110120 3250 110200 3260
rect 110340 3320 110420 3330
rect 110340 3260 110350 3320
rect 110410 3260 110420 3320
rect 110340 3250 110420 3260
rect 107980 3160 108000 3220
rect 108060 3160 108100 3220
rect 108160 3160 108200 3220
rect 108260 3160 108300 3220
rect 108360 3160 108400 3220
rect 108460 3160 108480 3220
rect 107980 1040 108480 3160
rect 108510 2320 108580 2332
rect 108510 2240 108580 2250
rect 108630 2320 108700 2330
rect 108630 2240 108700 2250
rect 108750 2320 108820 2330
rect 108750 2240 108820 2250
rect 108870 2320 108940 2330
rect 108870 2240 108940 2250
rect 108530 1620 108570 2240
rect 108770 2180 108810 2240
rect 108990 2180 109030 3250
rect 110230 3190 110310 3200
rect 110230 3130 110240 3190
rect 110300 3130 110310 3190
rect 110230 3110 110310 3130
rect 110230 3050 110240 3110
rect 110300 3050 110310 3110
rect 110230 3040 110310 3050
rect 110800 3190 111040 4720
rect 110800 3130 110810 3190
rect 110870 3130 110890 3190
rect 110950 3130 110970 3190
rect 111030 3130 111040 3190
rect 110800 3110 111040 3130
rect 110800 3050 110810 3110
rect 110870 3050 110890 3110
rect 110950 3050 110970 3110
rect 111030 3050 111040 3110
rect 110800 3040 111040 3050
rect 111070 6710 111310 8420
rect 112010 8370 112090 8380
rect 112010 8310 112020 8370
rect 112080 8310 112090 8370
rect 112010 8290 112090 8310
rect 112010 8230 112020 8290
rect 112080 8230 112090 8290
rect 112010 8210 112090 8230
rect 112010 8150 112020 8210
rect 112080 8150 112090 8210
rect 112010 8130 112090 8150
rect 112010 8070 112020 8130
rect 112080 8070 112090 8130
rect 112010 8050 112090 8070
rect 112010 7990 112020 8050
rect 112080 7990 112090 8050
rect 112010 7970 112090 7990
rect 112010 7910 112020 7970
rect 112080 7910 112090 7970
rect 112010 7900 112090 7910
rect 112250 8370 112330 8380
rect 112250 8310 112260 8370
rect 112320 8310 112330 8370
rect 112250 8290 112330 8310
rect 112250 8230 112260 8290
rect 112320 8230 112330 8290
rect 112250 8210 112330 8230
rect 112250 8150 112260 8210
rect 112320 8150 112330 8210
rect 112250 8130 112330 8150
rect 112250 8070 112260 8130
rect 112320 8070 112330 8130
rect 112250 8050 112330 8070
rect 112250 7990 112260 8050
rect 112320 7990 112330 8050
rect 112250 7970 112330 7990
rect 112250 7910 112260 7970
rect 112320 7910 112330 7970
rect 112250 7900 112330 7910
rect 112490 8370 112570 8380
rect 112490 8310 112500 8370
rect 112560 8310 112570 8370
rect 112490 8290 112570 8310
rect 112490 8230 112500 8290
rect 112560 8230 112570 8290
rect 112490 8210 112570 8230
rect 112490 8150 112500 8210
rect 112560 8150 112570 8210
rect 112490 8130 112570 8150
rect 112490 8070 112500 8130
rect 112560 8070 112570 8130
rect 112490 8050 112570 8070
rect 112490 7990 112500 8050
rect 112560 7990 112570 8050
rect 112490 7970 112570 7990
rect 112490 7910 112500 7970
rect 112560 7910 112570 7970
rect 112490 7900 112570 7910
rect 112730 8370 112810 8380
rect 112730 8310 112740 8370
rect 112800 8310 112810 8370
rect 112730 8290 112810 8310
rect 112730 8230 112740 8290
rect 112800 8230 112810 8290
rect 112730 8210 112810 8230
rect 112730 8150 112740 8210
rect 112800 8150 112810 8210
rect 112730 8130 112810 8150
rect 112730 8070 112740 8130
rect 112800 8070 112810 8130
rect 112730 8050 112810 8070
rect 112730 7990 112740 8050
rect 112800 7990 112810 8050
rect 112730 7970 112810 7990
rect 112730 7910 112740 7970
rect 112800 7910 112810 7970
rect 112730 7900 112810 7910
rect 112970 8370 113050 8380
rect 112970 8310 112980 8370
rect 113040 8310 113050 8370
rect 112970 8290 113050 8310
rect 112970 8230 112980 8290
rect 113040 8230 113050 8290
rect 112970 8210 113050 8230
rect 112970 8150 112980 8210
rect 113040 8150 113050 8210
rect 112970 8130 113050 8150
rect 112970 8070 112980 8130
rect 113040 8070 113050 8130
rect 112970 8050 113050 8070
rect 112970 7990 112980 8050
rect 113040 7990 113050 8050
rect 112970 7970 113050 7990
rect 112970 7910 112980 7970
rect 113040 7910 113050 7970
rect 112970 7900 113050 7910
rect 113210 8370 113290 8380
rect 113210 8310 113220 8370
rect 113280 8310 113290 8370
rect 113210 8290 113290 8310
rect 113210 8230 113220 8290
rect 113280 8230 113290 8290
rect 113210 8210 113290 8230
rect 113210 8150 113220 8210
rect 113280 8150 113290 8210
rect 113210 8130 113290 8150
rect 113210 8070 113220 8130
rect 113280 8070 113290 8130
rect 113210 8050 113290 8070
rect 113210 7990 113220 8050
rect 113280 7990 113290 8050
rect 113210 7970 113290 7990
rect 113210 7910 113220 7970
rect 113280 7910 113290 7970
rect 113210 7900 113290 7910
rect 113450 8370 113530 8380
rect 113450 8310 113460 8370
rect 113520 8310 113530 8370
rect 113450 8290 113530 8310
rect 113450 8230 113460 8290
rect 113520 8230 113530 8290
rect 113450 8210 113530 8230
rect 113450 8150 113460 8210
rect 113520 8150 113530 8210
rect 113450 8130 113530 8150
rect 113450 8070 113460 8130
rect 113520 8070 113530 8130
rect 113450 8050 113530 8070
rect 113450 7990 113460 8050
rect 113520 7990 113530 8050
rect 113450 7970 113530 7990
rect 113450 7910 113460 7970
rect 113520 7910 113530 7970
rect 113450 7900 113530 7910
rect 112020 7850 112080 7900
rect 112020 7810 112030 7850
rect 112070 7810 112080 7850
rect 112020 7730 112080 7810
rect 112130 7830 112210 7840
rect 112130 7770 112140 7830
rect 112200 7770 112210 7830
rect 112130 7760 112210 7770
rect 112020 7090 112030 7730
rect 112070 7090 112080 7730
rect 112020 7070 112080 7090
rect 112140 7730 112200 7760
rect 112140 7090 112150 7730
rect 112190 7090 112200 7730
rect 112140 7060 112200 7090
rect 112260 7730 112320 7900
rect 112370 7830 112450 7840
rect 112370 7770 112380 7830
rect 112440 7770 112450 7830
rect 112370 7760 112450 7770
rect 112260 7090 112270 7730
rect 112310 7090 112320 7730
rect 112260 7070 112320 7090
rect 112380 7730 112440 7760
rect 112380 7090 112390 7730
rect 112430 7090 112440 7730
rect 112380 7060 112440 7090
rect 112500 7730 112560 7900
rect 112610 7830 112690 7840
rect 112610 7770 112620 7830
rect 112680 7770 112690 7830
rect 112610 7760 112690 7770
rect 112500 7090 112510 7730
rect 112550 7090 112560 7730
rect 112500 7070 112560 7090
rect 112620 7730 112680 7760
rect 112620 7090 112630 7730
rect 112670 7090 112680 7730
rect 112620 7060 112680 7090
rect 112740 7730 112800 7900
rect 112850 7830 112930 7840
rect 112850 7770 112860 7830
rect 112920 7770 112930 7830
rect 112850 7760 112930 7770
rect 112740 7090 112750 7730
rect 112790 7090 112800 7730
rect 112740 7070 112800 7090
rect 112860 7730 112920 7760
rect 112860 7090 112870 7730
rect 112910 7090 112920 7730
rect 112860 7060 112920 7090
rect 112980 7730 113040 7900
rect 113090 7830 113170 7840
rect 113090 7770 113100 7830
rect 113160 7770 113170 7830
rect 113090 7760 113170 7770
rect 112980 7090 112990 7730
rect 113030 7090 113040 7730
rect 112980 7070 113040 7090
rect 113100 7730 113160 7760
rect 113100 7090 113110 7730
rect 113150 7090 113160 7730
rect 113100 7060 113160 7090
rect 113220 7730 113280 7900
rect 113460 7850 113520 7900
rect 113330 7830 113410 7840
rect 113330 7770 113340 7830
rect 113400 7770 113410 7830
rect 113330 7760 113410 7770
rect 113460 7810 113470 7850
rect 113510 7810 113520 7850
rect 113220 7090 113230 7730
rect 113270 7090 113280 7730
rect 113220 7070 113280 7090
rect 113340 7730 113400 7760
rect 113340 7090 113350 7730
rect 113390 7090 113400 7730
rect 113340 7060 113400 7090
rect 113460 7730 113520 7810
rect 113460 7090 113470 7730
rect 113510 7090 113520 7730
rect 113460 7070 113520 7090
rect 112130 7050 112210 7060
rect 112130 6990 112140 7050
rect 112200 6990 112210 7050
rect 112130 6980 112210 6990
rect 112370 7050 112450 7060
rect 112370 6990 112380 7050
rect 112440 6990 112450 7050
rect 112370 6980 112450 6990
rect 112610 7050 112690 7060
rect 112610 6990 112620 7050
rect 112680 6990 112690 7050
rect 112610 6980 112690 6990
rect 112850 7050 112930 7060
rect 112850 6990 112860 7050
rect 112920 6990 112930 7050
rect 112850 6980 112930 6990
rect 113090 7050 113170 7060
rect 113090 6990 113100 7050
rect 113160 6990 113170 7050
rect 113090 6980 113170 6990
rect 113330 7050 113410 7060
rect 113330 6990 113340 7050
rect 113400 6990 113410 7050
rect 113330 6980 113410 6990
rect 113690 6950 113730 8890
rect 113760 8640 113840 9460
rect 114060 9730 114120 9790
rect 114060 9090 114070 9730
rect 114110 9090 114120 9730
rect 114060 9070 114120 9090
rect 114180 9730 114240 10060
rect 114290 10020 114370 10030
rect 114290 9960 114300 10020
rect 114360 9960 114370 10020
rect 114290 9940 114370 9960
rect 114290 9880 114300 9940
rect 114360 9880 114370 9940
rect 114290 9860 114370 9880
rect 114290 9800 114300 9860
rect 114360 9800 114370 9860
rect 114290 9790 114370 9800
rect 114410 10020 114490 10030
rect 114410 9960 114420 10020
rect 114480 9960 114490 10020
rect 114410 9940 114490 9960
rect 114410 9880 114420 9940
rect 114480 9880 114490 9940
rect 114410 9860 114490 9880
rect 114410 9800 114420 9860
rect 114480 9800 114490 9860
rect 114410 9790 114490 9800
rect 114990 9860 115070 9870
rect 114990 9800 115000 9860
rect 115060 9800 115070 9860
rect 114990 9790 115070 9800
rect 115110 9860 115190 10070
rect 115110 9800 115120 9860
rect 115180 9800 115190 9860
rect 115110 9790 115190 9800
rect 115350 9860 115430 9870
rect 115350 9800 115360 9860
rect 115420 9800 115430 9860
rect 115350 9790 115430 9800
rect 114180 9090 114190 9730
rect 114230 9090 114240 9730
rect 114180 9060 114240 9090
rect 114300 9730 114360 9790
rect 114300 9090 114310 9730
rect 114350 9090 114360 9730
rect 114300 9070 114360 9090
rect 114420 9730 114480 9790
rect 114420 9090 114430 9730
rect 114470 9090 114480 9730
rect 114420 9070 114480 9090
rect 115000 9730 115060 9790
rect 115000 9090 115010 9730
rect 115050 9090 115060 9730
rect 115000 9070 115060 9090
rect 115120 9730 115180 9790
rect 115120 9090 115130 9730
rect 115170 9090 115180 9730
rect 115120 9060 115180 9090
rect 115240 9730 115300 9750
rect 115240 9090 115250 9730
rect 115290 9090 115300 9730
rect 114170 9050 114250 9060
rect 114170 8990 114180 9050
rect 114240 8990 114250 9050
rect 114170 8980 114250 8990
rect 115110 9050 115190 9060
rect 115110 8990 115120 9050
rect 115180 8990 115190 9050
rect 115110 8980 115190 8990
rect 114280 8950 114340 8970
rect 114280 8910 114290 8950
rect 114330 8910 114340 8950
rect 113760 8580 113770 8640
rect 113830 8580 113840 8640
rect 113760 8560 113840 8580
rect 113760 8500 113770 8560
rect 113830 8500 113840 8560
rect 113760 8480 113840 8500
rect 113760 8420 113770 8480
rect 113830 8420 113840 8480
rect 113760 8410 113840 8420
rect 113870 8850 113950 8860
rect 113870 8790 113880 8850
rect 113940 8790 113950 8850
rect 114280 8840 114340 8910
rect 115152 8940 115212 8950
rect 115152 8870 115212 8880
rect 115240 8840 115300 9090
rect 115360 9730 115420 9790
rect 115360 9090 115370 9730
rect 115410 9090 115420 9730
rect 115360 9070 115420 9090
rect 113870 8780 113950 8790
rect 114270 8830 114350 8840
rect 112200 6940 112260 6950
rect 112200 6870 112260 6880
rect 112320 6940 112380 6950
rect 112320 6870 112380 6880
rect 112440 6940 112500 6950
rect 112440 6870 112500 6880
rect 112560 6940 112620 6950
rect 112560 6870 112620 6880
rect 112680 6940 112740 6950
rect 112680 6870 112740 6880
rect 112800 6940 112860 6950
rect 112800 6870 112860 6880
rect 112920 6940 112980 6950
rect 112920 6870 112980 6880
rect 113040 6940 113100 6950
rect 113040 6870 113100 6880
rect 113160 6940 113220 6950
rect 113160 6870 113220 6880
rect 113280 6940 113340 6950
rect 113280 6870 113340 6880
rect 113670 6940 113750 6950
rect 113670 6880 113680 6940
rect 113740 6880 113750 6940
rect 113670 6870 113750 6880
rect 113870 6830 113910 8780
rect 114270 8770 114280 8830
rect 114340 8770 114350 8830
rect 114270 8760 114350 8770
rect 115230 8830 115310 8840
rect 115230 8770 115240 8830
rect 115300 8770 115310 8830
rect 115230 8760 115310 8770
rect 116290 8640 116530 8650
rect 116290 8580 116300 8640
rect 116360 8580 116380 8640
rect 116440 8580 116460 8640
rect 116520 8580 116530 8640
rect 116290 8560 116530 8580
rect 116290 8500 116300 8560
rect 116360 8500 116380 8560
rect 116440 8500 116460 8560
rect 116520 8500 116530 8560
rect 116290 8480 116530 8500
rect 116290 8420 116300 8480
rect 116360 8420 116380 8480
rect 116440 8420 116460 8480
rect 116520 8420 116530 8480
rect 114070 8370 114150 8380
rect 114070 8310 114080 8370
rect 114140 8310 114150 8370
rect 114070 8290 114150 8310
rect 114070 8230 114080 8290
rect 114140 8230 114150 8290
rect 114070 8210 114150 8230
rect 114070 8150 114080 8210
rect 114140 8150 114150 8210
rect 114070 8130 114150 8150
rect 114070 8070 114080 8130
rect 114140 8070 114150 8130
rect 114070 8050 114150 8070
rect 114070 7990 114080 8050
rect 114140 7990 114150 8050
rect 114070 7970 114150 7990
rect 114070 7910 114080 7970
rect 114140 7910 114150 7970
rect 114070 7900 114150 7910
rect 114310 8370 114390 8380
rect 114310 8310 114320 8370
rect 114380 8310 114390 8370
rect 114310 8290 114390 8310
rect 114310 8230 114320 8290
rect 114380 8230 114390 8290
rect 114310 8210 114390 8230
rect 114310 8150 114320 8210
rect 114380 8150 114390 8210
rect 114310 8130 114390 8150
rect 114310 8070 114320 8130
rect 114380 8070 114390 8130
rect 114310 8050 114390 8070
rect 114310 7990 114320 8050
rect 114380 7990 114390 8050
rect 114310 7970 114390 7990
rect 114310 7910 114320 7970
rect 114380 7910 114390 7970
rect 114310 7900 114390 7910
rect 114550 8370 114630 8380
rect 114550 8310 114560 8370
rect 114620 8310 114630 8370
rect 114550 8290 114630 8310
rect 114550 8230 114560 8290
rect 114620 8230 114630 8290
rect 114550 8210 114630 8230
rect 114550 8150 114560 8210
rect 114620 8150 114630 8210
rect 114550 8130 114630 8150
rect 114550 8070 114560 8130
rect 114620 8070 114630 8130
rect 114550 8050 114630 8070
rect 114550 7990 114560 8050
rect 114620 7990 114630 8050
rect 114550 7970 114630 7990
rect 114550 7910 114560 7970
rect 114620 7910 114630 7970
rect 114550 7900 114630 7910
rect 114790 8370 114870 8380
rect 114790 8310 114800 8370
rect 114860 8310 114870 8370
rect 114790 8290 114870 8310
rect 114790 8230 114800 8290
rect 114860 8230 114870 8290
rect 114790 8210 114870 8230
rect 114790 8150 114800 8210
rect 114860 8150 114870 8210
rect 114790 8130 114870 8150
rect 114790 8070 114800 8130
rect 114860 8070 114870 8130
rect 114790 8050 114870 8070
rect 114790 7990 114800 8050
rect 114860 7990 114870 8050
rect 114790 7970 114870 7990
rect 114790 7910 114800 7970
rect 114860 7910 114870 7970
rect 114790 7900 114870 7910
rect 115030 8370 115110 8380
rect 115030 8310 115040 8370
rect 115100 8310 115110 8370
rect 115030 8290 115110 8310
rect 115030 8230 115040 8290
rect 115100 8230 115110 8290
rect 115030 8210 115110 8230
rect 115030 8150 115040 8210
rect 115100 8150 115110 8210
rect 115030 8130 115110 8150
rect 115030 8070 115040 8130
rect 115100 8070 115110 8130
rect 115030 8050 115110 8070
rect 115030 7990 115040 8050
rect 115100 7990 115110 8050
rect 115030 7970 115110 7990
rect 115030 7910 115040 7970
rect 115100 7910 115110 7970
rect 115030 7900 115110 7910
rect 115270 8370 115350 8380
rect 115270 8310 115280 8370
rect 115340 8310 115350 8370
rect 115270 8290 115350 8310
rect 115270 8230 115280 8290
rect 115340 8230 115350 8290
rect 115270 8210 115350 8230
rect 115270 8150 115280 8210
rect 115340 8150 115350 8210
rect 115270 8130 115350 8150
rect 115270 8070 115280 8130
rect 115340 8070 115350 8130
rect 115270 8050 115350 8070
rect 115270 7990 115280 8050
rect 115340 7990 115350 8050
rect 115270 7970 115350 7990
rect 115270 7910 115280 7970
rect 115340 7910 115350 7970
rect 115270 7900 115350 7910
rect 115510 8370 115590 8380
rect 115510 8310 115520 8370
rect 115580 8310 115590 8370
rect 115510 8290 115590 8310
rect 115510 8230 115520 8290
rect 115580 8230 115590 8290
rect 115510 8210 115590 8230
rect 115510 8150 115520 8210
rect 115580 8150 115590 8210
rect 115510 8130 115590 8150
rect 115510 8070 115520 8130
rect 115580 8070 115590 8130
rect 115510 8050 115590 8070
rect 115510 7990 115520 8050
rect 115580 7990 115590 8050
rect 115510 7970 115590 7990
rect 115510 7910 115520 7970
rect 115580 7910 115590 7970
rect 115510 7900 115590 7910
rect 114080 7850 114140 7900
rect 114080 7810 114090 7850
rect 114130 7810 114140 7850
rect 114080 7730 114140 7810
rect 114190 7830 114270 7840
rect 114190 7770 114200 7830
rect 114260 7770 114270 7830
rect 114190 7760 114270 7770
rect 114080 7090 114090 7730
rect 114130 7090 114140 7730
rect 114080 7070 114140 7090
rect 114200 7730 114260 7760
rect 114200 7090 114210 7730
rect 114250 7090 114260 7730
rect 114200 7060 114260 7090
rect 114320 7730 114380 7900
rect 114430 7830 114510 7840
rect 114430 7770 114440 7830
rect 114500 7770 114510 7830
rect 114430 7760 114510 7770
rect 114320 7090 114330 7730
rect 114370 7090 114380 7730
rect 114320 7070 114380 7090
rect 114440 7730 114500 7760
rect 114440 7090 114450 7730
rect 114490 7090 114500 7730
rect 114440 7060 114500 7090
rect 114560 7730 114620 7900
rect 114670 7830 114750 7840
rect 114670 7770 114680 7830
rect 114740 7770 114750 7830
rect 114670 7760 114750 7770
rect 114560 7090 114570 7730
rect 114610 7090 114620 7730
rect 114560 7070 114620 7090
rect 114680 7730 114740 7760
rect 114680 7090 114690 7730
rect 114730 7090 114740 7730
rect 114680 7060 114740 7090
rect 114800 7730 114860 7900
rect 114910 7830 114990 7840
rect 114910 7770 114920 7830
rect 114980 7770 114990 7830
rect 114910 7760 114990 7770
rect 114800 7090 114810 7730
rect 114850 7090 114860 7730
rect 114800 7070 114860 7090
rect 114920 7730 114980 7760
rect 114920 7090 114930 7730
rect 114970 7090 114980 7730
rect 114920 7060 114980 7090
rect 115040 7730 115100 7900
rect 115150 7830 115230 7840
rect 115150 7770 115160 7830
rect 115220 7770 115230 7830
rect 115150 7760 115230 7770
rect 115040 7090 115050 7730
rect 115090 7090 115100 7730
rect 115040 7070 115100 7090
rect 115160 7730 115220 7760
rect 115160 7090 115170 7730
rect 115210 7090 115220 7730
rect 115160 7060 115220 7090
rect 115280 7730 115340 7900
rect 115520 7850 115580 7900
rect 115390 7830 115470 7840
rect 115390 7770 115400 7830
rect 115460 7770 115470 7830
rect 115390 7760 115470 7770
rect 115520 7810 115530 7850
rect 115570 7810 115580 7850
rect 115280 7090 115290 7730
rect 115330 7090 115340 7730
rect 115280 7070 115340 7090
rect 115400 7730 115460 7760
rect 115400 7090 115410 7730
rect 115450 7090 115460 7730
rect 115400 7060 115460 7090
rect 115520 7730 115580 7810
rect 115520 7090 115530 7730
rect 115570 7090 115580 7730
rect 115520 7070 115580 7090
rect 114190 7050 114270 7060
rect 114190 6990 114200 7050
rect 114260 6990 114270 7050
rect 114190 6980 114270 6990
rect 114430 7050 114510 7060
rect 114430 6990 114440 7050
rect 114500 6990 114510 7050
rect 114430 6980 114510 6990
rect 114670 7050 114750 7060
rect 114670 6990 114680 7050
rect 114740 6990 114750 7050
rect 114670 6980 114750 6990
rect 114910 7050 114990 7060
rect 114910 6990 114920 7050
rect 114980 6990 114990 7050
rect 114910 6980 114990 6990
rect 115150 7050 115230 7060
rect 115150 6990 115160 7050
rect 115220 6990 115230 7050
rect 115150 6980 115230 6990
rect 115390 7050 115470 7060
rect 115390 6990 115400 7050
rect 115460 6990 115470 7050
rect 115390 6980 115470 6990
rect 114260 6940 114320 6950
rect 114260 6870 114320 6880
rect 114380 6940 114440 6950
rect 114380 6870 114440 6880
rect 114500 6940 114560 6950
rect 114500 6870 114560 6880
rect 114620 6940 114680 6950
rect 114620 6870 114680 6880
rect 114740 6940 114800 6950
rect 114740 6870 114800 6880
rect 114860 6940 114920 6950
rect 114860 6870 114920 6880
rect 114980 6940 115040 6950
rect 114980 6870 115040 6880
rect 115100 6940 115160 6950
rect 115100 6870 115160 6880
rect 115220 6940 115280 6950
rect 115220 6870 115280 6880
rect 115340 6940 115400 6950
rect 115340 6870 115400 6880
rect 113850 6820 113930 6830
rect 113850 6760 113860 6820
rect 113920 6760 113930 6820
rect 113850 6750 113930 6760
rect 111070 6650 111080 6710
rect 111140 6650 111160 6710
rect 111220 6650 111240 6710
rect 111300 6650 111310 6710
rect 111070 6630 111310 6650
rect 111070 6570 111080 6630
rect 111140 6570 111160 6630
rect 111220 6570 111240 6630
rect 111300 6570 111310 6630
rect 111070 6550 111310 6570
rect 111070 6490 111080 6550
rect 111140 6490 111160 6550
rect 111220 6490 111240 6550
rect 111300 6490 111310 6550
rect 111070 4370 111310 6490
rect 113020 6710 113100 6720
rect 113020 6650 113030 6710
rect 113090 6650 113100 6710
rect 113020 6630 113100 6650
rect 113020 6570 113030 6630
rect 113090 6570 113100 6630
rect 113020 6550 113100 6570
rect 113020 6490 113030 6550
rect 113090 6490 113100 6550
rect 113020 6480 113100 6490
rect 113360 6710 113420 6720
rect 113360 6630 113420 6650
rect 113360 6550 113420 6570
rect 113360 6480 113420 6490
rect 113680 6710 113760 6720
rect 113680 6650 113690 6710
rect 113750 6650 113760 6710
rect 113680 6630 113760 6650
rect 113680 6570 113690 6630
rect 113750 6570 113760 6630
rect 113680 6550 113760 6570
rect 113680 6490 113690 6550
rect 113750 6490 113760 6550
rect 113680 6480 113760 6490
rect 113840 6710 113920 6720
rect 113840 6650 113850 6710
rect 113910 6650 113920 6710
rect 113840 6630 113920 6650
rect 113840 6570 113850 6630
rect 113910 6570 113920 6630
rect 113840 6550 113920 6570
rect 113840 6490 113850 6550
rect 113910 6490 113920 6550
rect 113840 6480 113920 6490
rect 114180 6710 114240 6720
rect 114180 6630 114240 6650
rect 114180 6550 114240 6570
rect 114180 6480 114240 6490
rect 114500 6710 114580 6720
rect 114500 6650 114510 6710
rect 114570 6650 114580 6710
rect 114500 6630 114580 6650
rect 114500 6570 114510 6630
rect 114570 6570 114580 6630
rect 114500 6550 114580 6570
rect 114500 6490 114510 6550
rect 114570 6490 114580 6550
rect 114500 6480 114580 6490
rect 116290 6710 116530 8420
rect 116900 8640 116980 8650
rect 116900 8580 116910 8640
rect 116970 8580 116980 8640
rect 116900 8560 116980 8580
rect 116900 8500 116910 8560
rect 116970 8500 116980 8560
rect 116900 8480 116980 8500
rect 116900 8420 116910 8480
rect 116970 8420 116980 8480
rect 116900 7860 116980 8420
rect 117620 8640 117700 8650
rect 117620 8580 117630 8640
rect 117690 8580 117700 8640
rect 117620 8560 117700 8580
rect 117620 8500 117630 8560
rect 117690 8500 117700 8560
rect 117620 8480 117700 8500
rect 117620 8420 117630 8480
rect 117690 8420 117700 8480
rect 117020 8370 117100 8380
rect 117020 8310 117030 8370
rect 117090 8310 117100 8370
rect 117020 8290 117100 8310
rect 117020 8230 117030 8290
rect 117090 8230 117100 8290
rect 117020 8210 117100 8230
rect 117020 8150 117030 8210
rect 117090 8150 117100 8210
rect 117020 8130 117100 8150
rect 117020 8070 117030 8130
rect 117090 8070 117100 8130
rect 117020 8050 117100 8070
rect 117020 7990 117030 8050
rect 117090 7990 117100 8050
rect 117020 7970 117100 7990
rect 117020 7910 117030 7970
rect 117090 7910 117100 7970
rect 117020 7900 117100 7910
rect 117260 8370 117340 8380
rect 117260 8310 117270 8370
rect 117330 8310 117340 8370
rect 117260 8290 117340 8310
rect 117260 8230 117270 8290
rect 117330 8230 117340 8290
rect 117260 8210 117340 8230
rect 117260 8150 117270 8210
rect 117330 8150 117340 8210
rect 117260 8130 117340 8150
rect 117260 8070 117270 8130
rect 117330 8070 117340 8130
rect 117260 8050 117340 8070
rect 117260 7990 117270 8050
rect 117330 7990 117340 8050
rect 117260 7970 117340 7990
rect 117260 7910 117270 7970
rect 117330 7910 117340 7970
rect 117260 7900 117340 7910
rect 117500 8370 117580 8380
rect 117500 8310 117510 8370
rect 117570 8310 117580 8370
rect 117500 8290 117580 8310
rect 117500 8230 117510 8290
rect 117570 8230 117580 8290
rect 117500 8210 117580 8230
rect 117500 8150 117510 8210
rect 117570 8150 117580 8210
rect 117500 8130 117580 8150
rect 117500 8070 117510 8130
rect 117570 8070 117580 8130
rect 117500 8050 117580 8070
rect 117500 7990 117510 8050
rect 117570 7990 117580 8050
rect 117500 7970 117580 7990
rect 117500 7910 117510 7970
rect 117570 7910 117580 7970
rect 117500 7900 117580 7910
rect 116900 7800 116910 7860
rect 116970 7800 116980 7860
rect 116900 7790 116980 7800
rect 116910 7730 116970 7790
rect 116910 7090 116920 7730
rect 116960 7090 116970 7730
rect 116290 6650 116300 6710
rect 116360 6650 116380 6710
rect 116440 6650 116460 6710
rect 116520 6650 116530 6710
rect 116290 6630 116530 6650
rect 116290 6570 116300 6630
rect 116360 6570 116380 6630
rect 116440 6570 116460 6630
rect 116520 6570 116530 6630
rect 116290 6550 116530 6570
rect 116290 6490 116300 6550
rect 116360 6490 116380 6550
rect 116440 6490 116460 6550
rect 116520 6490 116530 6550
rect 113240 6440 113320 6450
rect 113240 6380 113250 6440
rect 113310 6380 113320 6440
rect 113240 6370 113320 6380
rect 113460 6440 113540 6450
rect 113460 6380 113470 6440
rect 113530 6380 113540 6440
rect 113460 6370 113540 6380
rect 114060 6440 114140 6450
rect 114060 6380 114070 6440
rect 114130 6380 114140 6440
rect 114060 6370 114140 6380
rect 114280 6440 114360 6450
rect 114280 6380 114290 6440
rect 114350 6380 114360 6440
rect 114280 6370 114360 6380
rect 113120 5820 113180 5830
rect 113600 5820 113660 5830
rect 113120 5750 113180 5760
rect 113214 5790 113274 5810
rect 113214 5750 113224 5790
rect 113264 5750 113274 5790
rect 113214 5730 113274 5750
rect 113350 5800 113430 5810
rect 113350 5740 113360 5800
rect 113420 5740 113430 5800
rect 113350 5730 113430 5740
rect 113506 5790 113566 5810
rect 113506 5750 113516 5790
rect 113556 5750 113566 5790
rect 113600 5750 113660 5760
rect 113940 5810 114000 5830
rect 114420 5810 114480 5830
rect 113940 5770 113950 5810
rect 113990 5770 114000 5810
rect 113940 5750 114000 5770
rect 114034 5790 114094 5810
rect 114034 5750 114044 5790
rect 114084 5750 114094 5790
rect 113506 5730 113566 5750
rect 113220 5670 113260 5730
rect 113200 5660 113280 5670
rect 113200 5600 113210 5660
rect 113270 5600 113280 5660
rect 113200 5590 113280 5600
rect 113520 5570 113560 5730
rect 111900 5560 111980 5570
rect 111900 5500 111910 5560
rect 111970 5500 111980 5560
rect 111900 5490 111980 5500
rect 113490 5560 113570 5570
rect 113490 5500 113500 5560
rect 113560 5500 113570 5560
rect 113490 5490 113570 5500
rect 111070 4310 111080 4370
rect 111140 4310 111160 4370
rect 111220 4310 111240 4370
rect 111300 4310 111310 4370
rect 111070 4290 111310 4310
rect 111070 4230 111080 4290
rect 111140 4230 111160 4290
rect 111220 4230 111240 4290
rect 111300 4230 111310 4290
rect 111070 4210 111310 4230
rect 111070 4150 111080 4210
rect 111140 4150 111160 4210
rect 111220 4150 111240 4210
rect 111300 4150 111310 4210
rect 109060 2950 109140 2960
rect 109060 2890 109070 2950
rect 109130 2890 109140 2950
rect 109060 2880 109140 2890
rect 109460 2950 109540 2960
rect 109460 2890 109470 2950
rect 109530 2890 109540 2950
rect 109460 2880 109540 2890
rect 109680 2950 109760 2960
rect 109680 2890 109690 2950
rect 109750 2890 109760 2950
rect 109680 2880 109760 2890
rect 109900 2950 109980 2960
rect 109900 2890 109910 2950
rect 109970 2890 109980 2950
rect 109900 2880 109980 2890
rect 110120 2950 110200 2960
rect 110120 2890 110130 2950
rect 110190 2890 110200 2950
rect 110120 2880 110200 2890
rect 110340 2950 110420 2960
rect 110340 2890 110350 2950
rect 110410 2890 110420 2950
rect 110340 2880 110420 2890
rect 109080 2320 109120 2880
rect 109250 2850 109310 2870
rect 109060 2310 109140 2320
rect 109060 2250 109070 2310
rect 109130 2250 109140 2310
rect 109060 2240 109140 2250
rect 109250 2310 109260 2850
rect 109300 2310 109310 2850
rect 109250 2230 109310 2310
rect 109250 2190 109260 2230
rect 109300 2190 109310 2230
rect 108750 2170 108830 2180
rect 108750 2110 108760 2170
rect 108820 2110 108830 2170
rect 108750 2100 108830 2110
rect 108970 2170 109050 2180
rect 108970 2110 108980 2170
rect 109040 2110 109050 2170
rect 108970 2100 109050 2110
rect 109250 1890 109310 2190
rect 109360 2850 109420 2870
rect 109360 2310 109370 2850
rect 109410 2310 109420 2850
rect 109360 2160 109420 2310
rect 109470 2850 109530 2880
rect 109470 2310 109480 2850
rect 109520 2310 109530 2850
rect 109470 2280 109530 2310
rect 109580 2850 109640 2870
rect 109580 2310 109590 2850
rect 109630 2310 109640 2850
rect 109460 2270 109540 2280
rect 109460 2210 109470 2270
rect 109530 2210 109540 2270
rect 109460 2200 109540 2210
rect 109580 2160 109640 2310
rect 109690 2850 109750 2880
rect 109690 2310 109700 2850
rect 109740 2310 109750 2850
rect 109690 2280 109750 2310
rect 109800 2850 109860 2870
rect 109800 2310 109810 2850
rect 109850 2310 109860 2850
rect 109680 2270 109760 2280
rect 109680 2210 109690 2270
rect 109750 2210 109760 2270
rect 109680 2200 109760 2210
rect 109800 2160 109860 2310
rect 109910 2850 109970 2880
rect 109910 2310 109920 2850
rect 109960 2310 109970 2850
rect 109910 2280 109970 2310
rect 110020 2850 110080 2870
rect 110020 2310 110030 2850
rect 110070 2310 110080 2850
rect 109900 2270 109980 2280
rect 109900 2210 109910 2270
rect 109970 2210 109980 2270
rect 109900 2200 109980 2210
rect 110020 2160 110080 2310
rect 110130 2850 110190 2880
rect 110130 2310 110140 2850
rect 110180 2310 110190 2850
rect 110130 2280 110190 2310
rect 110240 2850 110300 2870
rect 110240 2310 110250 2850
rect 110290 2310 110300 2850
rect 110120 2270 110200 2280
rect 110120 2210 110130 2270
rect 110190 2210 110200 2270
rect 110120 2200 110200 2210
rect 110240 2160 110300 2310
rect 110350 2850 110410 2880
rect 110350 2310 110360 2850
rect 110400 2310 110410 2850
rect 110350 2280 110410 2310
rect 110460 2850 110520 2870
rect 110460 2310 110470 2850
rect 110510 2310 110520 2850
rect 110340 2270 110420 2280
rect 110340 2210 110350 2270
rect 110410 2210 110420 2270
rect 110340 2200 110420 2210
rect 110460 2160 110520 2310
rect 110570 2850 110630 2870
rect 110570 2310 110580 2850
rect 110620 2310 110630 2850
rect 110570 2230 110630 2310
rect 110570 2190 110580 2230
rect 110620 2190 110630 2230
rect 109350 2150 109430 2160
rect 109350 2090 109360 2150
rect 109420 2090 109430 2150
rect 109350 2070 109430 2090
rect 109350 2010 109360 2070
rect 109420 2010 109430 2070
rect 109350 1990 109430 2010
rect 109350 1930 109360 1990
rect 109420 1930 109430 1990
rect 109350 1920 109430 1930
rect 109570 2150 109650 2160
rect 109570 2090 109580 2150
rect 109640 2090 109650 2150
rect 109570 2070 109650 2090
rect 109570 2010 109580 2070
rect 109640 2010 109650 2070
rect 109570 1990 109650 2010
rect 109570 1930 109580 1990
rect 109640 1930 109650 1990
rect 109570 1920 109650 1930
rect 109790 2150 109870 2160
rect 109790 2090 109800 2150
rect 109860 2090 109870 2150
rect 109790 2070 109870 2090
rect 109790 2010 109800 2070
rect 109860 2010 109870 2070
rect 109790 1990 109870 2010
rect 109790 1930 109800 1990
rect 109860 1930 109870 1990
rect 109790 1920 109870 1930
rect 110010 2150 110090 2160
rect 110010 2090 110020 2150
rect 110080 2090 110090 2150
rect 110010 2070 110090 2090
rect 110010 2010 110020 2070
rect 110080 2010 110090 2070
rect 110010 1990 110090 2010
rect 110010 1930 110020 1990
rect 110080 1930 110090 1990
rect 110010 1920 110090 1930
rect 110230 2150 110310 2160
rect 110230 2090 110240 2150
rect 110300 2090 110310 2150
rect 110230 2070 110310 2090
rect 110230 2010 110240 2070
rect 110300 2010 110310 2070
rect 110230 1990 110310 2010
rect 110230 1930 110240 1990
rect 110300 1930 110310 1990
rect 110230 1920 110310 1930
rect 110450 2150 110530 2160
rect 110450 2090 110460 2150
rect 110520 2090 110530 2150
rect 110450 2070 110530 2090
rect 110450 2010 110460 2070
rect 110520 2010 110530 2070
rect 110450 1990 110530 2010
rect 110450 1930 110460 1990
rect 110520 1930 110530 1990
rect 110450 1920 110530 1930
rect 110570 1890 110630 2190
rect 111070 2150 111310 4150
rect 111340 4590 111580 4600
rect 111340 4530 111350 4590
rect 111410 4530 111430 4590
rect 111490 4530 111510 4590
rect 111570 4530 111580 4590
rect 111340 4510 111580 4530
rect 111340 4450 111350 4510
rect 111410 4450 111430 4510
rect 111490 4450 111510 4510
rect 111570 4450 111580 4510
rect 111340 4430 111580 4450
rect 111340 4370 111350 4430
rect 111410 4370 111430 4430
rect 111490 4370 111510 4430
rect 111570 4370 111580 4430
rect 111340 4100 111580 4370
rect 111340 4040 111350 4100
rect 111410 4040 111430 4100
rect 111490 4040 111510 4100
rect 111570 4040 111580 4100
rect 111340 4020 111580 4040
rect 111340 3960 111350 4020
rect 111410 3960 111430 4020
rect 111490 3960 111510 4020
rect 111570 3960 111580 4020
rect 111340 3940 111580 3960
rect 111340 3880 111350 3940
rect 111410 3880 111430 3940
rect 111490 3880 111510 3940
rect 111570 3880 111580 3940
rect 111340 3280 111580 3880
rect 111340 3220 111350 3280
rect 111410 3220 111430 3280
rect 111490 3220 111510 3280
rect 111570 3220 111580 3280
rect 111340 3200 111580 3220
rect 111340 3140 111350 3200
rect 111410 3140 111430 3200
rect 111490 3140 111510 3200
rect 111570 3140 111580 3200
rect 111340 3120 111580 3140
rect 111340 3060 111350 3120
rect 111410 3060 111430 3120
rect 111490 3060 111510 3120
rect 111570 3060 111580 3120
rect 111340 3050 111580 3060
rect 111690 3910 111850 3920
rect 111690 3850 111700 3910
rect 111760 3850 111780 3910
rect 111840 3850 111850 3910
rect 111070 2090 111080 2150
rect 111140 2090 111160 2150
rect 111220 2090 111240 2150
rect 111300 2090 111310 2150
rect 111070 2070 111310 2090
rect 111070 2010 111080 2070
rect 111140 2010 111160 2070
rect 111220 2010 111240 2070
rect 111300 2010 111310 2070
rect 111070 1990 111310 2010
rect 111070 1930 111080 1990
rect 111140 1930 111160 1990
rect 111220 1930 111240 1990
rect 111300 1930 111310 1990
rect 111070 1920 111310 1930
rect 111340 2970 111580 2980
rect 111340 2910 111350 2970
rect 111410 2910 111430 2970
rect 111490 2910 111510 2970
rect 111570 2910 111580 2970
rect 111340 2890 111580 2910
rect 111340 2830 111350 2890
rect 111410 2830 111430 2890
rect 111490 2830 111510 2890
rect 111570 2830 111580 2890
rect 111340 2810 111580 2830
rect 111340 2750 111350 2810
rect 111410 2750 111430 2810
rect 111490 2750 111510 2810
rect 111570 2750 111580 2810
rect 109240 1880 109320 1890
rect 109240 1820 109250 1880
rect 109310 1820 109320 1880
rect 109240 1800 109320 1820
rect 109240 1740 109250 1800
rect 109310 1740 109320 1800
rect 109240 1720 109320 1740
rect 109240 1660 109250 1720
rect 109310 1660 109320 1720
rect 109240 1650 109320 1660
rect 110560 1880 110640 1890
rect 110560 1820 110570 1880
rect 110630 1820 110640 1880
rect 110560 1800 110640 1820
rect 110560 1740 110570 1800
rect 110630 1740 110640 1800
rect 110560 1720 110640 1740
rect 110560 1660 110570 1720
rect 110630 1660 110640 1720
rect 110560 1650 110640 1660
rect 108510 1610 108590 1620
rect 108510 1550 108520 1610
rect 108580 1550 108590 1610
rect 108510 1540 108590 1550
rect 107980 980 107990 1040
rect 108050 980 108070 1040
rect 108130 980 108160 1040
rect 108220 980 108240 1040
rect 108300 980 108330 1040
rect 108390 980 108410 1040
rect 108470 980 108480 1040
rect 107980 960 108480 980
rect 107980 900 107990 960
rect 108050 900 108070 960
rect 108130 900 108160 960
rect 108220 900 108240 960
rect 108300 900 108330 960
rect 108390 900 108410 960
rect 108470 900 108480 960
rect 107980 880 108480 900
rect 107980 820 107990 880
rect 108050 820 108070 880
rect 108130 820 108160 880
rect 108220 820 108240 880
rect 108300 820 108330 880
rect 108390 820 108410 880
rect 108470 820 108480 880
rect 107980 810 108480 820
rect 108640 1150 108720 1160
rect 108640 1090 108650 1150
rect 108710 1090 108720 1150
rect 108640 770 108720 1090
rect 108640 710 108650 770
rect 108710 710 108720 770
rect 108640 670 108720 710
rect 108650 660 108720 670
rect 108650 580 108720 590
rect 108770 1040 108850 1050
rect 108770 980 108780 1040
rect 108840 980 108850 1040
rect 108770 960 108850 980
rect 108770 900 108780 960
rect 108840 900 108850 960
rect 108770 880 108850 900
rect 108770 820 108780 880
rect 108840 820 108850 880
rect 108770 810 108850 820
rect 109500 1040 110380 1050
rect 109500 980 109510 1040
rect 109570 980 109590 1040
rect 109650 980 109670 1040
rect 109730 980 109750 1040
rect 109810 980 109830 1040
rect 109890 980 109910 1040
rect 109970 980 109990 1040
rect 110050 980 110070 1040
rect 110130 980 110150 1040
rect 110210 980 110230 1040
rect 110290 980 110310 1040
rect 110370 980 110380 1040
rect 109500 960 110380 980
rect 109500 900 109510 960
rect 109570 900 109590 960
rect 109650 900 109670 960
rect 109730 900 109750 960
rect 109810 900 109830 960
rect 109890 900 109910 960
rect 109970 900 109990 960
rect 110050 900 110070 960
rect 110130 900 110150 960
rect 110210 900 110230 960
rect 110290 900 110310 960
rect 110370 900 110380 960
rect 109500 880 110380 900
rect 109500 820 109510 880
rect 109570 820 109590 880
rect 109650 820 109670 880
rect 109730 820 109750 880
rect 109810 820 109830 880
rect 109890 820 109910 880
rect 109970 820 109990 880
rect 110050 820 110070 880
rect 110130 820 110150 880
rect 110210 820 110230 880
rect 110290 820 110310 880
rect 110370 820 110380 880
rect 109500 810 110380 820
rect 108770 660 108840 810
rect 108770 580 108840 590
rect 109310 650 109370 670
rect 109310 -690 109320 650
rect 109360 -690 109370 650
rect 109310 -770 109370 -690
rect 109510 650 109570 810
rect 109600 770 109680 780
rect 109600 710 109610 770
rect 109670 710 109680 770
rect 109600 700 109680 710
rect 109800 770 109880 780
rect 109800 710 109810 770
rect 109870 710 109880 770
rect 109800 700 109880 710
rect 109510 -690 109520 650
rect 109560 -690 109570 650
rect 109510 -720 109570 -690
rect 109710 650 109770 670
rect 109710 -690 109720 650
rect 109760 -690 109770 650
rect 109310 -810 109320 -770
rect 109360 -810 109370 -770
rect 109500 -730 109580 -720
rect 109500 -790 109510 -730
rect 109570 -790 109580 -730
rect 109500 -800 109580 -790
rect 109310 -1150 109370 -810
rect 109710 -1150 109770 -690
rect 109910 650 109970 810
rect 110000 770 110080 780
rect 110000 710 110010 770
rect 110070 710 110080 770
rect 110000 700 110080 710
rect 110200 770 110280 780
rect 110200 710 110210 770
rect 110270 710 110280 770
rect 110200 700 110280 710
rect 109910 -690 109920 650
rect 109960 -690 109970 650
rect 109910 -720 109970 -690
rect 110110 650 110170 670
rect 110110 -690 110120 650
rect 110160 -690 110170 650
rect 109900 -730 109980 -720
rect 109900 -790 109910 -730
rect 109970 -790 109980 -730
rect 109900 -800 109980 -790
rect 107680 -1220 107690 -1160
rect 107750 -1220 107770 -1160
rect 107830 -1220 107850 -1160
rect 107910 -1220 107920 -1160
rect 107680 -1240 107920 -1220
rect 107680 -1300 107690 -1240
rect 107750 -1300 107770 -1240
rect 107830 -1300 107850 -1240
rect 107910 -1300 107920 -1240
rect 107680 -1320 107920 -1300
rect 107680 -1380 107690 -1320
rect 107750 -1380 107770 -1320
rect 107830 -1380 107850 -1320
rect 107910 -1380 107920 -1320
rect 107680 -1390 107920 -1380
rect 108080 -1160 108320 -1150
rect 108080 -1220 108090 -1160
rect 108150 -1220 108170 -1160
rect 108230 -1220 108250 -1160
rect 108310 -1220 108320 -1160
rect 108080 -1240 108320 -1220
rect 108080 -1300 108090 -1240
rect 108150 -1300 108170 -1240
rect 108230 -1300 108250 -1240
rect 108310 -1300 108320 -1240
rect 108080 -1320 108320 -1300
rect 108080 -1380 108090 -1320
rect 108150 -1380 108170 -1320
rect 108230 -1380 108250 -1320
rect 108310 -1380 108320 -1320
rect 108080 -3000 108320 -1380
rect 108780 -1160 109020 -1150
rect 108780 -1220 108790 -1160
rect 108850 -1220 108870 -1160
rect 108930 -1220 108950 -1160
rect 109010 -1220 109020 -1160
rect 108780 -1240 109020 -1220
rect 108780 -1300 108790 -1240
rect 108850 -1300 108870 -1240
rect 108930 -1300 108950 -1240
rect 109010 -1300 109020 -1240
rect 108780 -1320 109020 -1300
rect 108780 -1380 108790 -1320
rect 108850 -1380 108870 -1320
rect 108930 -1380 108950 -1320
rect 109010 -1380 109020 -1320
rect 108780 -3000 109020 -1380
rect 109300 -1160 109380 -1150
rect 109300 -1220 109310 -1160
rect 109370 -1220 109380 -1160
rect 109300 -1240 109380 -1220
rect 109300 -1300 109310 -1240
rect 109370 -1300 109380 -1240
rect 109300 -1320 109380 -1300
rect 109300 -1380 109310 -1320
rect 109370 -1380 109380 -1320
rect 109300 -1390 109380 -1380
rect 109480 -1160 109770 -1150
rect 109480 -1220 109490 -1160
rect 109550 -1220 109570 -1160
rect 109630 -1220 109650 -1160
rect 109710 -1220 109770 -1160
rect 109480 -1240 109770 -1220
rect 109480 -1300 109490 -1240
rect 109550 -1300 109570 -1240
rect 109630 -1300 109650 -1240
rect 109710 -1300 109770 -1240
rect 109480 -1320 109770 -1300
rect 109480 -1380 109490 -1320
rect 109550 -1380 109570 -1320
rect 109630 -1380 109650 -1320
rect 109710 -1380 109770 -1320
rect 109480 -1390 109770 -1380
rect 110110 -1150 110170 -690
rect 110310 650 110370 810
rect 110310 -690 110320 650
rect 110360 -690 110370 650
rect 110310 -720 110370 -690
rect 110510 650 110570 670
rect 110510 -690 110520 650
rect 110560 -690 110570 650
rect 111340 -120 111580 2750
rect 111340 -180 111350 -120
rect 111410 -180 111430 -120
rect 111490 -180 111510 -120
rect 111570 -180 111580 -120
rect 111340 -200 111580 -180
rect 111340 -260 111350 -200
rect 111410 -260 111430 -200
rect 111490 -260 111510 -200
rect 111570 -260 111580 -200
rect 111340 -280 111580 -260
rect 111340 -340 111350 -280
rect 111410 -340 111430 -280
rect 111490 -340 111510 -280
rect 111570 -340 111580 -280
rect 111340 -350 111580 -340
rect 110300 -730 110380 -720
rect 110300 -790 110310 -730
rect 110370 -790 110380 -730
rect 110300 -800 110380 -790
rect 110510 -770 110570 -690
rect 110510 -810 110520 -770
rect 110560 -810 110570 -770
rect 110510 -1150 110570 -810
rect 111690 -500 111850 3850
rect 111900 1620 111940 5490
rect 113940 5460 113980 5750
rect 114034 5730 114094 5750
rect 114170 5800 114250 5810
rect 114170 5740 114180 5800
rect 114240 5740 114250 5800
rect 114170 5730 114250 5740
rect 114326 5790 114386 5810
rect 114326 5750 114336 5790
rect 114376 5750 114386 5790
rect 114420 5770 114430 5810
rect 114470 5770 114480 5810
rect 114420 5750 114480 5770
rect 114326 5730 114386 5750
rect 114040 5570 114080 5730
rect 114340 5670 114380 5730
rect 114320 5660 114400 5670
rect 114320 5600 114330 5660
rect 114390 5600 114400 5660
rect 114320 5590 114400 5600
rect 114030 5560 114110 5570
rect 114030 5500 114040 5560
rect 114100 5500 114110 5560
rect 114030 5490 114110 5500
rect 113700 5450 113780 5460
rect 113700 5390 113710 5450
rect 113770 5390 113780 5450
rect 113700 5380 113780 5390
rect 113920 5450 114000 5460
rect 113920 5390 113930 5450
rect 113990 5390 114000 5450
rect 113920 5380 114000 5390
rect 113720 5240 113760 5380
rect 114440 5350 114480 5750
rect 115620 5560 115700 5570
rect 115620 5500 115630 5560
rect 115690 5500 115700 5560
rect 115620 5490 115700 5500
rect 113870 5340 113950 5350
rect 113870 5280 113880 5340
rect 113940 5280 113950 5340
rect 113870 5270 113950 5280
rect 114420 5340 114500 5350
rect 114420 5280 114430 5340
rect 114490 5280 114500 5340
rect 114420 5270 114500 5280
rect 113890 5240 113930 5270
rect 113660 5230 113780 5240
rect 113660 5170 113710 5230
rect 113770 5170 113780 5230
rect 113660 5160 113780 5170
rect 113870 5220 113950 5240
rect 113870 5180 113890 5220
rect 113930 5180 113950 5220
rect 113870 5160 113950 5180
rect 113550 5100 113610 5120
rect 112170 4940 113350 4950
rect 112170 4880 112180 4940
rect 112240 4880 112290 4940
rect 112350 4880 112400 4940
rect 112460 4880 112510 4940
rect 112570 4880 112620 4940
rect 112680 4880 112730 4940
rect 112790 4880 112840 4940
rect 112900 4880 112950 4940
rect 113010 4880 113060 4940
rect 113120 4880 113170 4940
rect 113230 4880 113280 4940
rect 113340 4880 113350 4940
rect 112170 4860 113350 4880
rect 112170 4800 112180 4860
rect 112240 4800 112290 4860
rect 112350 4800 112400 4860
rect 112460 4800 112510 4860
rect 112570 4800 112620 4860
rect 112680 4800 112730 4860
rect 112790 4800 112840 4860
rect 112900 4800 112950 4860
rect 113010 4800 113060 4860
rect 113120 4800 113170 4860
rect 113230 4800 113280 4860
rect 113340 4800 113350 4860
rect 112170 4780 113350 4800
rect 112170 4720 112180 4780
rect 112240 4720 112290 4780
rect 112350 4720 112400 4780
rect 112460 4720 112510 4780
rect 112570 4720 112620 4780
rect 112680 4720 112730 4780
rect 112790 4720 112840 4780
rect 112900 4720 112950 4780
rect 113010 4720 113060 4780
rect 113120 4720 113170 4780
rect 113230 4720 113280 4780
rect 113340 4720 113350 4780
rect 112170 4710 113350 4720
rect 112170 4020 112250 4710
rect 112170 3960 112180 4020
rect 112240 3960 112250 4020
rect 112170 3950 112250 3960
rect 112390 4020 112470 4710
rect 112390 3960 112400 4020
rect 112460 3960 112470 4020
rect 112390 3950 112470 3960
rect 112610 4020 112690 4710
rect 112610 3960 112620 4020
rect 112680 3960 112690 4020
rect 112610 3950 112690 3960
rect 112830 4020 112910 4710
rect 112830 3960 112840 4020
rect 112900 3960 112910 4020
rect 112830 3950 112910 3960
rect 113050 4020 113130 4710
rect 113050 3960 113060 4020
rect 113120 3960 113130 4020
rect 113050 3950 113130 3960
rect 113270 4020 113350 4710
rect 113550 4660 113560 5100
rect 113600 4660 113610 5100
rect 113550 4600 113610 4660
rect 113660 5100 113720 5160
rect 113660 4660 113670 5100
rect 113710 4660 113720 5100
rect 113660 4640 113720 4660
rect 113770 5100 113830 5120
rect 113770 4660 113780 5100
rect 113820 4660 113830 5100
rect 113770 4600 113830 4660
rect 113880 5100 113940 5160
rect 113880 4660 113890 5100
rect 113930 4660 113940 5100
rect 113880 4640 113940 4660
rect 113990 5100 114050 5120
rect 113990 4660 114000 5100
rect 114040 4660 114050 5100
rect 113990 4600 114050 4660
rect 114250 4940 115430 4950
rect 114250 4880 114260 4940
rect 114320 4880 114370 4940
rect 114430 4880 114480 4940
rect 114540 4880 114590 4940
rect 114650 4880 114700 4940
rect 114760 4880 114810 4940
rect 114870 4880 114920 4940
rect 114980 4880 115030 4940
rect 115090 4880 115140 4940
rect 115200 4880 115250 4940
rect 115310 4880 115360 4940
rect 115420 4880 115430 4940
rect 114250 4860 115430 4880
rect 114250 4800 114260 4860
rect 114320 4800 114370 4860
rect 114430 4800 114480 4860
rect 114540 4800 114590 4860
rect 114650 4800 114700 4860
rect 114760 4800 114810 4860
rect 114870 4800 114920 4860
rect 114980 4800 115030 4860
rect 115090 4800 115140 4860
rect 115200 4800 115250 4860
rect 115310 4800 115360 4860
rect 115420 4800 115430 4860
rect 114250 4780 115430 4800
rect 114250 4720 114260 4780
rect 114320 4720 114370 4780
rect 114430 4720 114480 4780
rect 114540 4720 114590 4780
rect 114650 4720 114700 4780
rect 114760 4720 114810 4780
rect 114870 4720 114920 4780
rect 114980 4720 115030 4780
rect 115090 4720 115140 4780
rect 115200 4720 115250 4780
rect 115310 4720 115360 4780
rect 115420 4720 115430 4780
rect 114250 4710 115430 4720
rect 113540 4590 113620 4600
rect 113540 4530 113550 4590
rect 113610 4530 113620 4590
rect 113540 4510 113620 4530
rect 113540 4450 113550 4510
rect 113610 4450 113620 4510
rect 113540 4430 113620 4450
rect 113540 4370 113550 4430
rect 113610 4370 113620 4430
rect 113540 4360 113620 4370
rect 113760 4590 113840 4600
rect 113760 4530 113770 4590
rect 113830 4530 113840 4590
rect 113760 4510 113840 4530
rect 113760 4450 113770 4510
rect 113830 4450 113840 4510
rect 113760 4430 113840 4450
rect 113760 4370 113770 4430
rect 113830 4370 113840 4430
rect 113760 4360 113840 4370
rect 113980 4590 114060 4600
rect 113980 4530 113990 4590
rect 114050 4530 114060 4590
rect 113980 4510 114060 4530
rect 113980 4450 113990 4510
rect 114050 4450 114060 4510
rect 113980 4430 114060 4450
rect 113980 4370 113990 4430
rect 114050 4370 114060 4430
rect 113980 4360 114060 4370
rect 113270 3960 113280 4020
rect 113340 3960 113350 4020
rect 113270 3950 113350 3960
rect 113570 4020 113650 4030
rect 113570 3960 113580 4020
rect 113640 3960 113650 4020
rect 112232 3910 112298 3920
rect 112232 3850 112238 3910
rect 112292 3850 112298 3910
rect 112232 3840 112298 3850
rect 112342 3910 112408 3920
rect 112342 3850 112348 3910
rect 112402 3850 112408 3910
rect 112342 3840 112408 3850
rect 112452 3910 112518 3920
rect 112452 3850 112458 3910
rect 112512 3850 112518 3910
rect 112452 3840 112518 3850
rect 112562 3910 112628 3920
rect 112562 3850 112568 3910
rect 112622 3850 112628 3910
rect 112562 3840 112628 3850
rect 112672 3910 112738 3920
rect 112672 3850 112678 3910
rect 112732 3850 112738 3910
rect 112672 3840 112738 3850
rect 112782 3910 112848 3920
rect 112782 3850 112788 3910
rect 112842 3850 112848 3910
rect 112782 3840 112848 3850
rect 112892 3910 112958 3920
rect 112892 3850 112898 3910
rect 112952 3850 112958 3910
rect 112892 3840 112958 3850
rect 113002 3910 113068 3920
rect 113002 3850 113008 3910
rect 113062 3850 113068 3910
rect 113002 3840 113068 3850
rect 113112 3910 113178 3920
rect 113112 3850 113118 3910
rect 113172 3850 113178 3910
rect 113112 3840 113178 3850
rect 113222 3910 113288 3920
rect 113222 3850 113228 3910
rect 113282 3850 113288 3910
rect 113222 3840 113288 3850
rect 112060 3780 112130 3800
rect 112060 3540 112080 3780
rect 112120 3540 112130 3780
rect 112060 3520 112130 3540
rect 112070 3510 112130 3520
rect 112180 3780 112240 3810
rect 112180 3540 112190 3780
rect 112230 3540 112240 3780
rect 112070 3460 112130 3480
rect 112070 3420 112080 3460
rect 112120 3420 112130 3460
rect 112070 3290 112130 3420
rect 112180 3400 112240 3540
rect 112290 3780 112350 3810
rect 112290 3540 112300 3780
rect 112340 3540 112350 3780
rect 112290 3510 112350 3540
rect 112400 3780 112460 3810
rect 112400 3540 112410 3780
rect 112450 3540 112460 3780
rect 112280 3500 112360 3510
rect 112280 3440 112290 3500
rect 112350 3440 112360 3500
rect 112280 3430 112360 3440
rect 112170 3390 112250 3400
rect 112170 3330 112180 3390
rect 112240 3330 112250 3390
rect 112170 3320 112250 3330
rect 112060 3280 112140 3290
rect 112060 3220 112070 3280
rect 112130 3220 112140 3280
rect 112060 3200 112140 3220
rect 112060 3140 112070 3200
rect 112130 3140 112140 3200
rect 112060 3120 112140 3140
rect 112060 3060 112070 3120
rect 112130 3060 112140 3120
rect 112060 3050 112140 3060
rect 112290 2630 112350 3430
rect 112400 3400 112460 3540
rect 112510 3780 112570 3810
rect 112510 3540 112520 3780
rect 112560 3540 112570 3780
rect 112510 3510 112570 3540
rect 112620 3780 112680 3810
rect 112620 3540 112630 3780
rect 112670 3540 112680 3780
rect 112500 3500 112580 3510
rect 112500 3440 112510 3500
rect 112570 3440 112580 3500
rect 112500 3430 112580 3440
rect 112390 3390 112470 3400
rect 112390 3330 112400 3390
rect 112460 3330 112470 3390
rect 112390 3320 112470 3330
rect 112170 2610 112250 2620
rect 112080 2590 112140 2600
rect 112170 2550 112180 2610
rect 112240 2550 112250 2610
rect 112510 2630 112570 3430
rect 112620 3400 112680 3540
rect 112730 3780 112790 3810
rect 112730 3540 112740 3780
rect 112780 3540 112790 3780
rect 112730 3510 112790 3540
rect 112840 3780 112900 3810
rect 112840 3540 112850 3780
rect 112890 3540 112900 3780
rect 112720 3500 112800 3510
rect 112720 3440 112730 3500
rect 112790 3440 112800 3500
rect 112720 3430 112800 3440
rect 112610 3390 112690 3400
rect 112610 3330 112620 3390
rect 112680 3330 112690 3390
rect 112610 3320 112690 3330
rect 112290 2560 112350 2570
rect 112390 2610 112470 2620
rect 112170 2540 112250 2550
rect 112390 2550 112400 2610
rect 112460 2550 112470 2610
rect 112730 2630 112790 3430
rect 112840 3400 112900 3540
rect 112950 3780 113010 3810
rect 112950 3540 112960 3780
rect 113000 3540 113010 3780
rect 112950 3510 113010 3540
rect 113060 3780 113120 3810
rect 113060 3540 113070 3780
rect 113110 3540 113120 3780
rect 112940 3500 113020 3510
rect 112940 3440 112950 3500
rect 113010 3440 113020 3500
rect 112940 3430 113020 3440
rect 112830 3390 112910 3400
rect 112830 3330 112840 3390
rect 112900 3330 112910 3390
rect 112830 3320 112910 3330
rect 112510 2560 112570 2570
rect 112610 2610 112690 2620
rect 112390 2540 112470 2550
rect 112610 2550 112620 2610
rect 112680 2550 112690 2610
rect 112950 2630 113010 3430
rect 113060 3400 113120 3540
rect 113170 3780 113230 3810
rect 113170 3540 113180 3780
rect 113220 3540 113230 3780
rect 113170 3510 113230 3540
rect 113280 3780 113340 3810
rect 113280 3540 113290 3780
rect 113330 3540 113340 3780
rect 113160 3500 113240 3510
rect 113160 3440 113170 3500
rect 113230 3440 113240 3500
rect 113160 3430 113240 3440
rect 113050 3390 113130 3400
rect 113050 3330 113060 3390
rect 113120 3330 113130 3390
rect 113050 3320 113130 3330
rect 112730 2560 112790 2570
rect 112830 2610 112910 2620
rect 112610 2540 112690 2550
rect 112830 2550 112840 2610
rect 112900 2550 112910 2610
rect 113170 2630 113230 3430
rect 113280 3400 113340 3540
rect 113390 3780 113530 3800
rect 113390 3540 113400 3780
rect 113440 3540 113530 3780
rect 113390 3520 113530 3540
rect 113390 3460 113450 3520
rect 113390 3420 113400 3460
rect 113440 3420 113450 3460
rect 113270 3390 113350 3400
rect 113270 3330 113280 3390
rect 113340 3330 113350 3390
rect 113270 3320 113350 3330
rect 113390 3290 113450 3420
rect 113570 3390 113650 3960
rect 113570 3330 113580 3390
rect 113640 3330 113650 3390
rect 113570 3320 113650 3330
rect 113950 4020 114030 4030
rect 113950 3960 113960 4020
rect 114020 3960 114030 4020
rect 113950 3390 114030 3960
rect 114250 4020 114330 4710
rect 114250 3960 114260 4020
rect 114320 3960 114330 4020
rect 114250 3950 114330 3960
rect 114470 4020 114550 4710
rect 114470 3960 114480 4020
rect 114540 3960 114550 4020
rect 114470 3950 114550 3960
rect 114690 4020 114770 4710
rect 114690 3960 114700 4020
rect 114760 3960 114770 4020
rect 114690 3950 114770 3960
rect 114910 4020 114990 4710
rect 114910 3960 114920 4020
rect 114980 3960 114990 4020
rect 114910 3950 114990 3960
rect 115130 4020 115210 4710
rect 115130 3960 115140 4020
rect 115200 3960 115210 4020
rect 115130 3950 115210 3960
rect 115350 4020 115430 4710
rect 115350 3960 115360 4020
rect 115420 3960 115430 4020
rect 115350 3950 115430 3960
rect 114312 3910 114378 3920
rect 114312 3850 114318 3910
rect 114372 3850 114378 3910
rect 114312 3840 114378 3850
rect 114422 3910 114488 3920
rect 114422 3850 114428 3910
rect 114482 3850 114488 3910
rect 114422 3840 114488 3850
rect 114532 3910 114598 3920
rect 114532 3850 114538 3910
rect 114592 3850 114598 3910
rect 114532 3840 114598 3850
rect 114642 3910 114708 3920
rect 114642 3850 114648 3910
rect 114702 3850 114708 3910
rect 114642 3840 114708 3850
rect 114752 3910 114818 3920
rect 114752 3850 114758 3910
rect 114812 3850 114818 3910
rect 114752 3840 114818 3850
rect 114862 3910 114928 3920
rect 114862 3850 114868 3910
rect 114922 3850 114928 3910
rect 114862 3840 114928 3850
rect 114972 3910 115038 3920
rect 114972 3850 114978 3910
rect 115032 3850 115038 3910
rect 114972 3840 115038 3850
rect 115082 3910 115148 3920
rect 115082 3850 115088 3910
rect 115142 3850 115148 3910
rect 115082 3840 115148 3850
rect 115192 3910 115258 3920
rect 115192 3850 115198 3910
rect 115252 3850 115258 3910
rect 115192 3840 115258 3850
rect 115302 3910 115368 3920
rect 115302 3850 115308 3910
rect 115362 3850 115368 3910
rect 115302 3840 115368 3850
rect 114070 3780 114210 3800
rect 114070 3540 114160 3780
rect 114200 3540 114210 3780
rect 114070 3520 114210 3540
rect 113950 3330 113960 3390
rect 114020 3330 114030 3390
rect 113950 3320 114030 3330
rect 114150 3460 114210 3520
rect 114150 3420 114160 3460
rect 114200 3420 114210 3460
rect 114150 3290 114210 3420
rect 114260 3780 114320 3810
rect 114260 3540 114270 3780
rect 114310 3540 114320 3780
rect 114260 3400 114320 3540
rect 114370 3780 114430 3810
rect 114370 3540 114380 3780
rect 114420 3540 114430 3780
rect 114370 3510 114430 3540
rect 114480 3780 114540 3810
rect 114480 3540 114490 3780
rect 114530 3540 114540 3780
rect 114360 3500 114440 3510
rect 114360 3440 114370 3500
rect 114430 3440 114440 3500
rect 114360 3430 114440 3440
rect 114250 3390 114330 3400
rect 114250 3330 114260 3390
rect 114320 3330 114330 3390
rect 114250 3320 114330 3330
rect 113380 3280 113460 3290
rect 113380 3220 113390 3280
rect 113450 3220 113460 3280
rect 113380 3200 113460 3220
rect 113380 3140 113390 3200
rect 113450 3140 113460 3200
rect 113380 3120 113460 3140
rect 113380 3060 113390 3120
rect 113450 3060 113460 3120
rect 113380 3050 113460 3060
rect 114140 3280 114220 3290
rect 114140 3220 114150 3280
rect 114210 3220 114220 3280
rect 114140 3200 114220 3220
rect 114140 3140 114150 3200
rect 114210 3140 114220 3200
rect 114140 3120 114220 3140
rect 114140 3060 114150 3120
rect 114210 3060 114220 3120
rect 114140 3050 114220 3060
rect 113760 2970 113840 2980
rect 113760 2910 113770 2970
rect 113830 2910 113840 2970
rect 113760 2890 113840 2910
rect 113760 2830 113770 2890
rect 113830 2830 113840 2890
rect 113760 2810 113840 2830
rect 113760 2750 113770 2810
rect 113830 2750 113840 2810
rect 113760 2740 113840 2750
rect 112950 2560 113010 2570
rect 113050 2610 113130 2620
rect 112830 2540 112910 2550
rect 113050 2550 113060 2610
rect 113120 2550 113130 2610
rect 113170 2560 113230 2570
rect 113270 2610 113350 2620
rect 113050 2540 113130 2550
rect 113270 2550 113280 2610
rect 113340 2550 113350 2610
rect 113270 2540 113350 2550
rect 113380 2610 113440 2620
rect 113380 2540 113440 2550
rect 113680 2610 113740 2620
rect 113680 2540 113740 2550
rect 112080 2520 112140 2530
rect 112070 2410 112130 2430
rect 112070 2170 112080 2410
rect 112120 2170 112130 2410
rect 112070 2150 112130 2170
rect 112180 2410 112240 2540
rect 112280 2520 112360 2530
rect 112280 2460 112290 2520
rect 112350 2460 112360 2520
rect 112280 2450 112360 2460
rect 112180 2170 112190 2410
rect 112230 2170 112240 2410
rect 112180 2140 112240 2170
rect 112290 2410 112350 2450
rect 112290 2170 112300 2410
rect 112340 2170 112350 2410
rect 112170 2130 112250 2140
rect 112070 2090 112130 2110
rect 112070 2050 112080 2090
rect 112120 2050 112130 2090
rect 112170 2070 112180 2130
rect 112240 2070 112250 2130
rect 112170 2060 112250 2070
rect 112070 2030 112130 2050
rect 112080 1890 112120 2030
rect 112290 2000 112350 2170
rect 112400 2410 112460 2540
rect 112500 2520 112580 2530
rect 112500 2460 112510 2520
rect 112570 2460 112580 2520
rect 112500 2450 112580 2460
rect 112400 2170 112410 2410
rect 112450 2170 112460 2410
rect 112400 2140 112460 2170
rect 112510 2410 112570 2450
rect 112510 2170 112520 2410
rect 112560 2170 112570 2410
rect 112390 2130 112470 2140
rect 112390 2070 112400 2130
rect 112460 2070 112470 2130
rect 112390 2060 112470 2070
rect 112510 2000 112570 2170
rect 112620 2410 112680 2540
rect 112720 2520 112800 2530
rect 112720 2460 112730 2520
rect 112790 2460 112800 2520
rect 112720 2450 112800 2460
rect 112620 2170 112630 2410
rect 112670 2170 112680 2410
rect 112620 2140 112680 2170
rect 112730 2410 112790 2450
rect 112730 2170 112740 2410
rect 112780 2170 112790 2410
rect 112610 2130 112690 2140
rect 112610 2070 112620 2130
rect 112680 2070 112690 2130
rect 112610 2060 112690 2070
rect 112730 2000 112790 2170
rect 112840 2410 112900 2540
rect 112940 2520 113020 2530
rect 112940 2460 112950 2520
rect 113010 2460 113020 2520
rect 112940 2450 113020 2460
rect 112840 2170 112850 2410
rect 112890 2170 112900 2410
rect 112840 2140 112900 2170
rect 112950 2410 113010 2450
rect 112950 2170 112960 2410
rect 113000 2170 113010 2410
rect 112830 2130 112910 2140
rect 112830 2070 112840 2130
rect 112900 2070 112910 2130
rect 112830 2060 112910 2070
rect 112950 2000 113010 2170
rect 113060 2410 113120 2540
rect 113160 2520 113240 2530
rect 113160 2460 113170 2520
rect 113230 2460 113240 2520
rect 113160 2450 113240 2460
rect 113060 2170 113070 2410
rect 113110 2170 113120 2410
rect 113060 2140 113120 2170
rect 113170 2410 113230 2450
rect 113170 2170 113180 2410
rect 113220 2170 113230 2410
rect 113050 2130 113130 2140
rect 113050 2070 113060 2130
rect 113120 2070 113130 2130
rect 113050 2060 113130 2070
rect 113170 2000 113230 2170
rect 113280 2410 113340 2540
rect 113280 2170 113290 2410
rect 113330 2170 113340 2410
rect 113280 2140 113340 2170
rect 113390 2410 113610 2430
rect 113390 2170 113400 2410
rect 113440 2170 113560 2410
rect 113600 2170 113610 2410
rect 113390 2150 113610 2170
rect 113660 2410 113720 2430
rect 113660 2170 113670 2410
rect 113710 2170 113720 2410
rect 113270 2130 113350 2140
rect 113270 2070 113280 2130
rect 113340 2070 113350 2130
rect 113480 2110 113520 2150
rect 113660 2140 113720 2170
rect 113770 2410 113830 2740
rect 114370 2630 114430 3430
rect 114480 3400 114540 3540
rect 114590 3780 114650 3810
rect 114590 3540 114600 3780
rect 114640 3540 114650 3780
rect 114590 3510 114650 3540
rect 114700 3780 114760 3810
rect 114700 3540 114710 3780
rect 114750 3540 114760 3780
rect 114580 3500 114660 3510
rect 114580 3440 114590 3500
rect 114650 3440 114660 3500
rect 114580 3430 114660 3440
rect 114470 3390 114550 3400
rect 114470 3330 114480 3390
rect 114540 3330 114550 3390
rect 114470 3320 114550 3330
rect 113860 2610 113920 2620
rect 113860 2540 113920 2550
rect 114160 2610 114220 2620
rect 114160 2540 114220 2550
rect 114250 2610 114330 2620
rect 114250 2550 114260 2610
rect 114320 2550 114330 2610
rect 114590 2630 114650 3430
rect 114700 3400 114760 3540
rect 114810 3780 114870 3810
rect 114810 3540 114820 3780
rect 114860 3540 114870 3780
rect 114810 3510 114870 3540
rect 114920 3780 114980 3810
rect 114920 3540 114930 3780
rect 114970 3540 114980 3780
rect 114800 3500 114880 3510
rect 114800 3440 114810 3500
rect 114870 3440 114880 3500
rect 114800 3430 114880 3440
rect 114690 3390 114770 3400
rect 114690 3330 114700 3390
rect 114760 3330 114770 3390
rect 114690 3320 114770 3330
rect 114370 2560 114430 2570
rect 114470 2610 114550 2620
rect 114250 2540 114330 2550
rect 114470 2550 114480 2610
rect 114540 2550 114550 2610
rect 114810 2630 114870 3430
rect 114920 3400 114980 3540
rect 115030 3780 115090 3810
rect 115030 3540 115040 3780
rect 115080 3540 115090 3780
rect 115030 3510 115090 3540
rect 115140 3780 115200 3810
rect 115140 3540 115150 3780
rect 115190 3540 115200 3780
rect 115020 3500 115100 3510
rect 115020 3440 115030 3500
rect 115090 3440 115100 3500
rect 115020 3430 115100 3440
rect 114910 3390 114990 3400
rect 114910 3330 114920 3390
rect 114980 3330 114990 3390
rect 114910 3320 114990 3330
rect 114590 2560 114650 2570
rect 114690 2610 114770 2620
rect 114470 2540 114550 2550
rect 114690 2550 114700 2610
rect 114760 2550 114770 2610
rect 115030 2630 115090 3430
rect 115140 3400 115200 3540
rect 115250 3780 115310 3810
rect 115250 3540 115260 3780
rect 115300 3540 115310 3780
rect 115250 3510 115310 3540
rect 115360 3780 115420 3810
rect 115360 3540 115370 3780
rect 115410 3540 115420 3780
rect 115240 3500 115320 3510
rect 115240 3440 115250 3500
rect 115310 3440 115320 3500
rect 115240 3430 115320 3440
rect 115130 3390 115210 3400
rect 115130 3330 115140 3390
rect 115200 3330 115210 3390
rect 115130 3320 115210 3330
rect 114810 2560 114870 2570
rect 114910 2610 114990 2620
rect 114690 2540 114770 2550
rect 114910 2550 114920 2610
rect 114980 2550 114990 2610
rect 115250 2630 115310 3430
rect 115360 3400 115420 3540
rect 115470 3780 115530 3800
rect 115470 3540 115480 3780
rect 115520 3540 115530 3780
rect 115470 3520 115530 3540
rect 115470 3460 115530 3480
rect 115470 3420 115480 3460
rect 115520 3420 115530 3460
rect 115350 3390 115430 3400
rect 115350 3330 115360 3390
rect 115420 3330 115430 3390
rect 115350 3320 115430 3330
rect 115470 3290 115530 3420
rect 115460 3280 115540 3290
rect 115460 3220 115470 3280
rect 115530 3220 115540 3280
rect 115460 3200 115540 3220
rect 115460 3140 115470 3200
rect 115530 3140 115540 3200
rect 115460 3120 115540 3140
rect 115460 3060 115470 3120
rect 115530 3060 115540 3120
rect 115460 3050 115540 3060
rect 115030 2560 115090 2570
rect 115130 2610 115210 2620
rect 114910 2540 114990 2550
rect 115130 2550 115140 2610
rect 115200 2550 115210 2610
rect 115250 2560 115310 2570
rect 115350 2610 115430 2620
rect 115130 2540 115210 2550
rect 115350 2550 115360 2610
rect 115420 2550 115430 2610
rect 115350 2540 115430 2550
rect 115460 2590 115520 2600
rect 113770 2170 113780 2410
rect 113820 2170 113830 2410
rect 113770 2150 113830 2170
rect 113880 2410 113940 2430
rect 113880 2170 113890 2410
rect 113930 2170 113940 2410
rect 113880 2140 113940 2170
rect 113990 2410 114210 2430
rect 113990 2170 114000 2410
rect 114040 2170 114160 2410
rect 114200 2170 114210 2410
rect 113990 2150 114210 2170
rect 114260 2410 114320 2540
rect 114360 2520 114440 2530
rect 114360 2460 114370 2520
rect 114430 2460 114440 2520
rect 114360 2450 114440 2460
rect 114260 2170 114270 2410
rect 114310 2170 114320 2410
rect 113650 2130 113730 2140
rect 113270 2060 113350 2070
rect 113470 2090 113530 2110
rect 113470 2050 113480 2090
rect 113520 2050 113530 2090
rect 113470 2030 113530 2050
rect 113650 2070 113660 2130
rect 113720 2070 113730 2130
rect 112280 1990 112360 2000
rect 112280 1930 112290 1990
rect 112350 1930 112360 1990
rect 112280 1920 112360 1930
rect 112500 1990 112580 2000
rect 112500 1930 112510 1990
rect 112570 1930 112580 1990
rect 112500 1920 112580 1930
rect 112720 1990 112800 2000
rect 112720 1930 112730 1990
rect 112790 1930 112800 1990
rect 112720 1920 112800 1930
rect 112880 1990 113400 2000
rect 112880 1930 112950 1990
rect 113010 1930 113170 1990
rect 113230 1930 113400 1990
rect 112060 1880 112140 1890
rect 112060 1820 112070 1880
rect 112130 1820 112140 1880
rect 112060 1800 112140 1820
rect 112060 1740 112070 1800
rect 112130 1740 112140 1800
rect 112060 1720 112140 1740
rect 112060 1660 112070 1720
rect 112130 1660 112140 1720
rect 112060 1650 112140 1660
rect 111880 1610 111960 1620
rect 111880 1550 111890 1610
rect 111950 1550 111960 1610
rect 111880 1540 111960 1550
rect 112880 1030 113400 1930
rect 113480 1890 113520 2030
rect 113460 1880 113540 1890
rect 113460 1820 113470 1880
rect 113530 1820 113540 1880
rect 113460 1800 113540 1820
rect 113460 1740 113470 1800
rect 113530 1740 113540 1800
rect 113460 1720 113540 1740
rect 113460 1660 113470 1720
rect 113530 1660 113540 1720
rect 113460 1650 113540 1660
rect 112880 970 112890 1030
rect 112950 970 113110 1030
rect 113170 970 113330 1030
rect 113390 970 113400 1030
rect 112880 960 113400 970
rect 113540 1030 113620 1040
rect 113540 970 113550 1030
rect 113610 970 113620 1030
rect 113540 960 113620 970
rect 113650 1000 113730 2070
rect 113870 2130 113950 2140
rect 113870 2070 113880 2130
rect 113940 2070 113950 2130
rect 114080 2110 114120 2150
rect 114260 2140 114320 2170
rect 114370 2410 114430 2450
rect 114370 2170 114380 2410
rect 114420 2170 114430 2410
rect 114250 2130 114330 2140
rect 113650 960 113670 1000
rect 113710 960 113730 1000
rect 113760 1030 113840 1040
rect 113760 970 113770 1030
rect 113830 970 113840 1030
rect 113760 960 113840 970
rect 113870 1000 113950 2070
rect 114070 2090 114130 2110
rect 114070 2050 114080 2090
rect 114120 2050 114130 2090
rect 114250 2070 114260 2130
rect 114320 2070 114330 2130
rect 114250 2060 114330 2070
rect 114070 2030 114130 2050
rect 114080 1890 114120 2030
rect 114370 2000 114430 2170
rect 114480 2410 114540 2540
rect 114580 2520 114660 2530
rect 114580 2460 114590 2520
rect 114650 2460 114660 2520
rect 114580 2450 114660 2460
rect 114480 2170 114490 2410
rect 114530 2170 114540 2410
rect 114480 2140 114540 2170
rect 114590 2410 114650 2450
rect 114590 2170 114600 2410
rect 114640 2170 114650 2410
rect 114470 2130 114550 2140
rect 114470 2070 114480 2130
rect 114540 2070 114550 2130
rect 114470 2060 114550 2070
rect 114590 2000 114650 2170
rect 114700 2410 114760 2540
rect 114800 2520 114880 2530
rect 114800 2460 114810 2520
rect 114870 2460 114880 2520
rect 114800 2450 114880 2460
rect 114700 2170 114710 2410
rect 114750 2170 114760 2410
rect 114700 2140 114760 2170
rect 114810 2410 114870 2450
rect 114810 2170 114820 2410
rect 114860 2170 114870 2410
rect 114690 2130 114770 2140
rect 114690 2070 114700 2130
rect 114760 2070 114770 2130
rect 114690 2060 114770 2070
rect 114810 2000 114870 2170
rect 114920 2410 114980 2540
rect 115020 2520 115100 2530
rect 115020 2460 115030 2520
rect 115090 2460 115100 2520
rect 115020 2450 115100 2460
rect 114920 2170 114930 2410
rect 114970 2170 114980 2410
rect 114920 2140 114980 2170
rect 115030 2410 115090 2450
rect 115030 2170 115040 2410
rect 115080 2170 115090 2410
rect 114910 2130 114990 2140
rect 114910 2070 114920 2130
rect 114980 2070 114990 2130
rect 114910 2060 114990 2070
rect 115030 2000 115090 2170
rect 115140 2410 115200 2540
rect 115240 2520 115320 2530
rect 115240 2460 115250 2520
rect 115310 2460 115320 2520
rect 115240 2450 115320 2460
rect 115140 2170 115150 2410
rect 115190 2170 115200 2410
rect 115140 2140 115200 2170
rect 115250 2410 115310 2450
rect 115250 2170 115260 2410
rect 115300 2170 115310 2410
rect 115130 2130 115210 2140
rect 115130 2070 115140 2130
rect 115200 2070 115210 2130
rect 115130 2060 115210 2070
rect 115250 2000 115310 2170
rect 115360 2410 115420 2540
rect 115460 2520 115520 2530
rect 115360 2170 115370 2410
rect 115410 2170 115420 2410
rect 115360 2140 115420 2170
rect 115470 2410 115530 2430
rect 115470 2170 115480 2410
rect 115520 2170 115530 2410
rect 115470 2150 115530 2170
rect 115350 2130 115430 2140
rect 115350 2070 115360 2130
rect 115420 2070 115430 2130
rect 115350 2060 115430 2070
rect 115470 2090 115530 2110
rect 115470 2050 115480 2090
rect 115520 2050 115530 2090
rect 115470 2030 115530 2050
rect 114200 1990 114720 2000
rect 114200 1930 114370 1990
rect 114430 1930 114590 1990
rect 114650 1930 114720 1990
rect 114060 1880 114140 1890
rect 114060 1820 114070 1880
rect 114130 1820 114140 1880
rect 114060 1800 114140 1820
rect 114060 1740 114070 1800
rect 114130 1740 114140 1800
rect 114060 1720 114140 1740
rect 114060 1660 114070 1720
rect 114130 1660 114140 1720
rect 114060 1650 114140 1660
rect 113870 960 113890 1000
rect 113930 960 113950 1000
rect 113980 1030 114060 1040
rect 113980 970 113990 1030
rect 114050 970 114060 1030
rect 113980 960 114060 970
rect 114200 1030 114720 1930
rect 114800 1990 114880 2000
rect 114800 1930 114810 1990
rect 114870 1930 114880 1990
rect 114800 1920 114880 1930
rect 115020 1990 115100 2000
rect 115020 1930 115030 1990
rect 115090 1930 115100 1990
rect 115020 1920 115100 1930
rect 115240 1990 115320 2000
rect 115240 1930 115250 1990
rect 115310 1930 115320 1990
rect 115240 1920 115320 1930
rect 115480 1890 115520 2030
rect 115460 1880 115540 1890
rect 115460 1820 115470 1880
rect 115530 1820 115540 1880
rect 115460 1800 115540 1820
rect 115460 1740 115470 1800
rect 115530 1740 115540 1800
rect 115460 1720 115540 1740
rect 115460 1660 115470 1720
rect 115530 1660 115540 1720
rect 115460 1650 115540 1660
rect 115660 1620 115700 5490
rect 115730 5340 115810 5350
rect 115730 5280 115740 5340
rect 115800 5280 115810 5340
rect 115730 5270 115810 5280
rect 115640 1610 115720 1620
rect 115640 1550 115650 1610
rect 115710 1550 115720 1610
rect 115640 1540 115720 1550
rect 114200 970 114210 1030
rect 114270 970 114430 1030
rect 114490 970 114650 1030
rect 114710 970 114720 1030
rect 114200 960 114720 970
rect 114860 1030 114940 1040
rect 114860 970 114870 1030
rect 114930 970 114940 1030
rect 114860 960 114940 970
rect 112370 880 112510 900
rect 112370 440 112460 880
rect 112500 440 112510 880
rect 112370 420 112510 440
rect 112450 380 112510 420
rect 112560 880 112620 900
rect 112560 440 112570 880
rect 112610 440 112620 880
rect 112560 380 112620 440
rect 112670 880 112730 900
rect 112670 440 112680 880
rect 112720 440 112730 880
rect 111690 -560 111700 -500
rect 111760 -560 111780 -500
rect 111840 -560 111850 -500
rect 111690 -940 111850 -560
rect 111690 -1000 111700 -940
rect 111760 -1000 111780 -940
rect 111840 -1000 111850 -940
rect 111690 -1010 111850 -1000
rect 112440 370 112520 380
rect 112440 310 112450 370
rect 112510 310 112520 370
rect 112440 -1150 112520 310
rect 112550 370 112630 380
rect 112550 310 112560 370
rect 112620 310 112630 370
rect 112550 300 112630 310
rect 112670 -110 112730 440
rect 112780 880 112840 900
rect 112780 440 112790 880
rect 112830 440 112840 880
rect 112780 380 112840 440
rect 112890 880 112950 960
rect 112890 440 112900 880
rect 112940 440 112950 880
rect 112770 370 112850 380
rect 112770 310 112780 370
rect 112840 310 112850 370
rect 112770 300 112850 310
rect 112890 270 112950 440
rect 113000 880 113060 900
rect 113000 440 113010 880
rect 113050 440 113060 880
rect 113000 380 113060 440
rect 113110 880 113170 960
rect 113110 440 113120 880
rect 113160 440 113170 880
rect 112990 370 113070 380
rect 112990 310 113000 370
rect 113060 310 113070 370
rect 112990 300 113070 310
rect 113110 270 113170 440
rect 113220 880 113280 900
rect 113220 440 113230 880
rect 113270 440 113280 880
rect 113220 380 113280 440
rect 113330 880 113390 960
rect 113330 440 113340 880
rect 113380 440 113390 880
rect 113210 370 113290 380
rect 113210 310 113220 370
rect 113280 310 113290 370
rect 113210 300 113290 310
rect 113330 270 113390 440
rect 113440 880 113500 900
rect 113440 440 113450 880
rect 113490 440 113500 880
rect 113440 380 113500 440
rect 113550 880 113610 960
rect 113650 940 113730 960
rect 113550 440 113560 880
rect 113600 440 113610 880
rect 113430 370 113510 380
rect 113430 310 113440 370
rect 113500 310 113510 370
rect 113430 300 113510 310
rect 113550 270 113610 440
rect 113660 880 113720 900
rect 113660 440 113670 880
rect 113710 440 113720 880
rect 113660 380 113720 440
rect 113770 880 113830 960
rect 113870 940 113950 960
rect 113770 440 113780 880
rect 113820 440 113830 880
rect 113650 370 113730 380
rect 113650 310 113660 370
rect 113720 310 113730 370
rect 113650 300 113730 310
rect 113770 270 113830 440
rect 113880 880 113940 900
rect 113880 440 113890 880
rect 113930 440 113940 880
rect 113880 380 113940 440
rect 113990 880 114050 960
rect 113990 440 114000 880
rect 114040 440 114050 880
rect 113870 370 113950 380
rect 113870 310 113880 370
rect 113940 310 113950 370
rect 113870 300 113950 310
rect 113990 270 114050 440
rect 114100 880 114160 900
rect 114100 440 114110 880
rect 114150 440 114160 880
rect 114100 380 114160 440
rect 114210 880 114270 960
rect 114210 440 114220 880
rect 114260 440 114270 880
rect 114090 370 114170 380
rect 114090 310 114100 370
rect 114160 310 114170 370
rect 114090 300 114170 310
rect 114210 270 114270 440
rect 114320 880 114380 900
rect 114320 440 114330 880
rect 114370 440 114380 880
rect 114320 380 114380 440
rect 114430 880 114490 960
rect 114430 440 114440 880
rect 114480 440 114490 880
rect 114310 370 114390 380
rect 114310 310 114320 370
rect 114380 310 114390 370
rect 114310 300 114390 310
rect 114430 270 114490 440
rect 114540 880 114600 900
rect 114540 440 114550 880
rect 114590 440 114600 880
rect 114540 380 114600 440
rect 114650 880 114710 960
rect 114650 440 114660 880
rect 114700 440 114710 880
rect 114530 370 114610 380
rect 114530 310 114540 370
rect 114600 310 114610 370
rect 114530 300 114610 310
rect 114650 270 114710 440
rect 114760 880 114820 900
rect 114760 440 114770 880
rect 114810 440 114820 880
rect 114760 380 114820 440
rect 114870 880 114930 960
rect 114870 440 114880 880
rect 114920 440 114930 880
rect 114750 370 114830 380
rect 114750 310 114760 370
rect 114820 310 114830 370
rect 114750 300 114830 310
rect 114870 270 114930 440
rect 114980 880 115040 900
rect 114980 440 114990 880
rect 115030 440 115040 880
rect 114980 380 115040 440
rect 114970 370 115050 380
rect 114970 310 114980 370
rect 115040 310 115050 370
rect 112880 260 112960 270
rect 112880 200 112890 260
rect 112950 200 112960 260
rect 112880 180 112960 200
rect 112880 120 112890 180
rect 112950 120 112960 180
rect 112880 100 112960 120
rect 112880 40 112890 100
rect 112950 40 112960 100
rect 112880 30 112960 40
rect 113100 260 113180 270
rect 113100 200 113110 260
rect 113170 200 113180 260
rect 113100 180 113180 200
rect 113100 120 113110 180
rect 113170 120 113180 180
rect 113100 100 113180 120
rect 113100 40 113110 100
rect 113170 40 113180 100
rect 113100 30 113180 40
rect 113320 260 113400 270
rect 113320 200 113330 260
rect 113390 200 113400 260
rect 113320 180 113400 200
rect 113320 120 113330 180
rect 113390 120 113400 180
rect 113320 100 113400 120
rect 113320 40 113330 100
rect 113390 40 113400 100
rect 113320 30 113400 40
rect 113540 260 113620 270
rect 113540 200 113550 260
rect 113610 200 113620 260
rect 113540 180 113620 200
rect 113540 120 113550 180
rect 113610 120 113620 180
rect 113540 100 113620 120
rect 113540 40 113550 100
rect 113610 40 113620 100
rect 113540 30 113620 40
rect 113760 260 113840 270
rect 113760 200 113770 260
rect 113830 200 113840 260
rect 113760 180 113840 200
rect 113760 120 113770 180
rect 113830 120 113840 180
rect 113760 100 113840 120
rect 113760 40 113770 100
rect 113830 40 113840 100
rect 113760 30 113840 40
rect 113980 260 114060 270
rect 113980 200 113990 260
rect 114050 200 114060 260
rect 113980 180 114060 200
rect 113980 120 113990 180
rect 114050 120 114060 180
rect 113980 100 114060 120
rect 113980 40 113990 100
rect 114050 40 114060 100
rect 113980 30 114060 40
rect 114200 260 114280 270
rect 114200 200 114210 260
rect 114270 200 114280 260
rect 114200 180 114280 200
rect 114200 120 114210 180
rect 114270 120 114280 180
rect 114200 100 114280 120
rect 114200 40 114210 100
rect 114270 40 114280 100
rect 114200 30 114280 40
rect 114420 260 114500 270
rect 114420 200 114430 260
rect 114490 200 114500 260
rect 114420 180 114500 200
rect 114420 120 114430 180
rect 114490 120 114500 180
rect 114420 100 114500 120
rect 114420 40 114430 100
rect 114490 40 114500 100
rect 114420 30 114500 40
rect 114640 260 114720 270
rect 114640 200 114650 260
rect 114710 200 114720 260
rect 114640 180 114720 200
rect 114640 120 114650 180
rect 114710 120 114720 180
rect 114640 100 114720 120
rect 114640 40 114650 100
rect 114710 40 114720 100
rect 114640 30 114720 40
rect 114860 260 114940 270
rect 114860 200 114870 260
rect 114930 200 114940 260
rect 114860 180 114940 200
rect 114860 120 114870 180
rect 114930 120 114940 180
rect 114860 100 114940 120
rect 114860 40 114870 100
rect 114930 40 114940 100
rect 114860 30 114940 40
rect 114830 -10 114910 0
rect 114830 -70 114840 -10
rect 114900 -70 114910 -10
rect 114830 -80 114910 -70
rect 112660 -120 112740 -110
rect 112660 -180 112670 -120
rect 112730 -180 112740 -120
rect 112660 -200 112740 -180
rect 112660 -260 112670 -200
rect 112730 -260 112740 -200
rect 112660 -280 112740 -260
rect 112660 -340 112670 -280
rect 112730 -340 112740 -280
rect 112660 -350 112740 -340
rect 113080 -390 113160 -380
rect 113080 -450 113090 -390
rect 113150 -450 113160 -390
rect 113080 -460 113160 -450
rect 113300 -390 113380 -380
rect 113300 -450 113310 -390
rect 113370 -450 113380 -390
rect 113300 -460 113380 -450
rect 113740 -390 113820 -380
rect 113740 -450 113750 -390
rect 113810 -450 113820 -390
rect 113740 -460 113820 -450
rect 112970 -500 113050 -490
rect 112970 -560 112980 -500
rect 113040 -560 113050 -500
rect 112970 -570 113050 -560
rect 112790 -630 112930 -610
rect 112790 -870 112880 -630
rect 112920 -870 112930 -630
rect 112790 -890 112930 -870
rect 112870 -950 112930 -890
rect 112980 -630 113040 -570
rect 112980 -870 112990 -630
rect 113030 -870 113040 -630
rect 112980 -930 113040 -870
rect 113090 -630 113150 -460
rect 113190 -500 113270 -490
rect 113190 -560 113200 -500
rect 113260 -560 113270 -500
rect 113190 -570 113270 -560
rect 113090 -870 113100 -630
rect 113140 -870 113150 -630
rect 112870 -990 112880 -950
rect 112920 -990 112930 -950
rect 112870 -1150 112930 -990
rect 112970 -940 113050 -930
rect 112970 -1000 112980 -940
rect 113040 -1000 113050 -940
rect 112970 -1010 113050 -1000
rect 113090 -1040 113150 -870
rect 113200 -630 113260 -570
rect 113200 -870 113210 -630
rect 113250 -870 113260 -630
rect 113200 -930 113260 -870
rect 113310 -630 113370 -460
rect 113410 -500 113490 -490
rect 113410 -560 113420 -500
rect 113480 -560 113490 -500
rect 113410 -570 113490 -560
rect 113310 -870 113320 -630
rect 113360 -870 113370 -630
rect 113190 -940 113270 -930
rect 113190 -1000 113200 -940
rect 113260 -1000 113270 -940
rect 113190 -1010 113270 -1000
rect 113310 -1040 113370 -870
rect 113420 -630 113480 -570
rect 113420 -870 113430 -630
rect 113470 -870 113480 -630
rect 113420 -930 113480 -870
rect 113530 -630 113670 -610
rect 113530 -870 113540 -630
rect 113580 -870 113670 -630
rect 113530 -890 113670 -870
rect 113750 -630 113810 -460
rect 114080 -500 114160 -490
rect 114080 -560 114090 -500
rect 114150 -560 114160 -500
rect 114080 -570 114160 -560
rect 113750 -870 113760 -630
rect 113800 -870 113810 -630
rect 114430 -650 114490 -630
rect 114430 -870 114490 -850
rect 113410 -940 113490 -930
rect 113410 -1000 113420 -940
rect 113480 -1000 113490 -940
rect 113410 -1010 113490 -1000
rect 113530 -950 113590 -890
rect 113530 -990 113540 -950
rect 113580 -990 113590 -950
rect 113080 -1050 113160 -1040
rect 113080 -1110 113090 -1050
rect 113150 -1110 113160 -1050
rect 113080 -1120 113160 -1110
rect 113300 -1050 113380 -1040
rect 113300 -1110 113310 -1050
rect 113370 -1110 113380 -1050
rect 113300 -1120 113380 -1110
rect 113530 -1150 113590 -990
rect 113750 -1040 113810 -870
rect 114080 -940 114160 -930
rect 114080 -1000 114090 -940
rect 114150 -1000 114160 -940
rect 114080 -1010 114160 -1000
rect 113740 -1050 113820 -1040
rect 113740 -1110 113750 -1050
rect 113810 -1110 113820 -1050
rect 113740 -1120 113820 -1110
rect 110110 -1160 110420 -1150
rect 110110 -1220 110190 -1160
rect 110250 -1220 110270 -1160
rect 110330 -1220 110350 -1160
rect 110410 -1220 110420 -1160
rect 110110 -1240 110420 -1220
rect 110110 -1300 110190 -1240
rect 110250 -1300 110270 -1240
rect 110330 -1300 110350 -1240
rect 110410 -1300 110420 -1240
rect 110110 -1320 110420 -1300
rect 110110 -1380 110190 -1320
rect 110250 -1380 110270 -1320
rect 110330 -1380 110350 -1320
rect 110410 -1380 110420 -1320
rect 110110 -1390 110420 -1380
rect 110500 -1160 110580 -1150
rect 110500 -1220 110510 -1160
rect 110570 -1220 110580 -1160
rect 110500 -1240 110580 -1220
rect 110500 -1300 110510 -1240
rect 110570 -1300 110580 -1240
rect 110500 -1320 110580 -1300
rect 110500 -1380 110510 -1320
rect 110570 -1380 110580 -1320
rect 110500 -1390 110580 -1380
rect 110880 -1160 111120 -1150
rect 110880 -1220 110890 -1160
rect 110950 -1220 110970 -1160
rect 111030 -1220 111050 -1160
rect 111110 -1220 111120 -1160
rect 110880 -1240 111120 -1220
rect 110880 -1300 110890 -1240
rect 110950 -1300 110970 -1240
rect 111030 -1300 111050 -1240
rect 111110 -1300 111120 -1240
rect 110880 -1320 111120 -1300
rect 110880 -1380 110890 -1320
rect 110950 -1380 110970 -1320
rect 111030 -1380 111050 -1320
rect 111110 -1380 111120 -1320
rect 109480 -3000 109720 -1390
rect 110180 -3000 110420 -1390
rect 110880 -3000 111120 -1380
rect 111580 -1160 111820 -1150
rect 111580 -1220 111590 -1160
rect 111650 -1220 111670 -1160
rect 111730 -1220 111750 -1160
rect 111810 -1220 111820 -1160
rect 111580 -1240 111820 -1220
rect 111580 -1300 111590 -1240
rect 111650 -1300 111670 -1240
rect 111730 -1300 111750 -1240
rect 111810 -1300 111820 -1240
rect 111580 -1320 111820 -1300
rect 111580 -1380 111590 -1320
rect 111650 -1380 111670 -1320
rect 111730 -1380 111750 -1320
rect 111810 -1380 111820 -1320
rect 111580 -3000 111820 -1380
rect 112280 -1160 112520 -1150
rect 112280 -1220 112290 -1160
rect 112350 -1220 112370 -1160
rect 112430 -1220 112450 -1160
rect 112510 -1220 112520 -1160
rect 112280 -1240 112520 -1220
rect 112280 -1300 112290 -1240
rect 112350 -1300 112370 -1240
rect 112430 -1300 112450 -1240
rect 112510 -1300 112520 -1240
rect 112280 -1320 112520 -1300
rect 112280 -1380 112290 -1320
rect 112350 -1380 112370 -1320
rect 112430 -1380 112450 -1320
rect 112510 -1380 112520 -1320
rect 112280 -3000 112520 -1380
rect 112860 -1160 112940 -1150
rect 112860 -1220 112870 -1160
rect 112930 -1220 112940 -1160
rect 112860 -1240 112940 -1220
rect 112860 -1300 112870 -1240
rect 112930 -1300 112940 -1240
rect 112860 -1320 112940 -1300
rect 112860 -1380 112870 -1320
rect 112930 -1380 112940 -1320
rect 112860 -1390 112940 -1380
rect 112980 -1160 113220 -1150
rect 112980 -1220 112990 -1160
rect 113050 -1220 113070 -1160
rect 113130 -1220 113150 -1160
rect 113210 -1220 113220 -1160
rect 112980 -1240 113220 -1220
rect 112980 -1300 112990 -1240
rect 113050 -1300 113070 -1240
rect 113130 -1300 113150 -1240
rect 113210 -1300 113220 -1240
rect 112980 -1320 113220 -1300
rect 112980 -1380 112990 -1320
rect 113050 -1380 113070 -1320
rect 113130 -1380 113150 -1320
rect 113210 -1380 113220 -1320
rect 112980 -3000 113220 -1380
rect 113520 -1160 113600 -1150
rect 113520 -1220 113530 -1160
rect 113590 -1220 113600 -1160
rect 113520 -1240 113600 -1220
rect 113520 -1300 113530 -1240
rect 113590 -1300 113600 -1240
rect 113520 -1320 113600 -1300
rect 113520 -1380 113530 -1320
rect 113590 -1380 113600 -1320
rect 113520 -1390 113600 -1380
rect 113680 -1160 113920 -1150
rect 113680 -1220 113690 -1160
rect 113750 -1220 113770 -1160
rect 113830 -1220 113850 -1160
rect 113910 -1220 113920 -1160
rect 113680 -1240 113920 -1220
rect 113680 -1300 113690 -1240
rect 113750 -1300 113770 -1240
rect 113830 -1300 113850 -1240
rect 113910 -1300 113920 -1240
rect 113680 -1320 113920 -1300
rect 113680 -1380 113690 -1320
rect 113750 -1380 113770 -1320
rect 113830 -1380 113850 -1320
rect 113910 -1380 113920 -1320
rect 113680 -3000 113920 -1380
rect 114380 -1160 114620 -1150
rect 114380 -1220 114390 -1160
rect 114450 -1220 114470 -1160
rect 114530 -1220 114550 -1160
rect 114610 -1220 114620 -1160
rect 114380 -1240 114620 -1220
rect 114380 -1300 114390 -1240
rect 114450 -1300 114470 -1240
rect 114530 -1300 114550 -1240
rect 114610 -1300 114620 -1240
rect 114380 -1320 114620 -1300
rect 114380 -1380 114390 -1320
rect 114450 -1380 114470 -1320
rect 114530 -1380 114550 -1320
rect 114610 -1380 114620 -1320
rect 114380 -3000 114620 -1380
rect 114970 -1160 115050 310
rect 115420 260 115660 270
rect 115420 200 115430 260
rect 115490 200 115510 260
rect 115570 200 115590 260
rect 115650 200 115660 260
rect 115420 180 115660 200
rect 115420 120 115430 180
rect 115490 120 115510 180
rect 115570 120 115590 180
rect 115650 120 115660 180
rect 115420 100 115660 120
rect 115420 40 115430 100
rect 115490 40 115510 100
rect 115570 40 115590 100
rect 115650 40 115660 100
rect 115420 -640 115660 40
rect 115750 0 115790 5270
rect 116020 4590 116260 4600
rect 116020 4530 116030 4590
rect 116090 4530 116110 4590
rect 116170 4530 116190 4590
rect 116250 4530 116260 4590
rect 116020 4510 116260 4530
rect 116020 4450 116030 4510
rect 116090 4450 116110 4510
rect 116170 4450 116190 4510
rect 116250 4450 116260 4510
rect 116020 4430 116260 4450
rect 116020 4370 116030 4430
rect 116090 4370 116110 4430
rect 116170 4370 116190 4430
rect 116250 4370 116260 4430
rect 116020 4100 116260 4370
rect 116020 4040 116030 4100
rect 116090 4040 116110 4100
rect 116170 4040 116190 4100
rect 116250 4040 116260 4100
rect 116020 4020 116260 4040
rect 116020 3960 116030 4020
rect 116090 3960 116110 4020
rect 116170 3960 116190 4020
rect 116250 3960 116260 4020
rect 116020 3940 116260 3960
rect 116020 3880 116030 3940
rect 116090 3880 116110 3940
rect 116170 3880 116190 3940
rect 116250 3880 116260 3940
rect 116020 3280 116260 3880
rect 116020 3220 116030 3280
rect 116090 3220 116110 3280
rect 116170 3220 116190 3280
rect 116250 3220 116260 3280
rect 116020 3200 116260 3220
rect 116020 3140 116030 3200
rect 116090 3140 116110 3200
rect 116170 3140 116190 3200
rect 116250 3140 116260 3200
rect 116020 3120 116260 3140
rect 116020 3060 116030 3120
rect 116090 3060 116110 3120
rect 116170 3060 116190 3120
rect 116250 3060 116260 3120
rect 116020 3050 116260 3060
rect 116290 4370 116530 6490
rect 116290 4310 116300 4370
rect 116360 4310 116380 4370
rect 116440 4310 116460 4370
rect 116520 4310 116530 4370
rect 116290 4290 116530 4310
rect 116290 4230 116300 4290
rect 116360 4230 116380 4290
rect 116440 4230 116460 4290
rect 116520 4230 116530 4290
rect 116290 4210 116530 4230
rect 116290 4150 116300 4210
rect 116360 4150 116380 4210
rect 116440 4150 116460 4210
rect 116520 4150 116530 4210
rect 116020 2970 116260 2980
rect 116020 2910 116030 2970
rect 116090 2910 116110 2970
rect 116170 2910 116190 2970
rect 116250 2910 116260 2970
rect 116020 2890 116260 2910
rect 116020 2830 116030 2890
rect 116090 2830 116110 2890
rect 116170 2830 116190 2890
rect 116250 2830 116260 2890
rect 116020 2810 116260 2830
rect 116020 2750 116030 2810
rect 116090 2750 116110 2810
rect 116170 2750 116190 2810
rect 116250 2750 116260 2810
rect 115730 -10 115810 0
rect 115730 -70 115740 -10
rect 115800 -70 115810 -10
rect 115730 -80 115810 -70
rect 116020 -120 116260 2750
rect 116290 2160 116530 4150
rect 116560 7050 116800 7060
rect 116560 6990 116570 7050
rect 116630 6990 116650 7050
rect 116710 6990 116730 7050
rect 116790 6990 116800 7050
rect 116560 4940 116800 6990
rect 116910 7010 116970 7090
rect 117030 7730 117090 7900
rect 117140 7860 117220 7870
rect 117140 7800 117150 7860
rect 117210 7800 117220 7860
rect 117140 7790 117220 7800
rect 117030 7090 117040 7730
rect 117080 7090 117090 7730
rect 117030 7060 117090 7090
rect 117150 7730 117210 7790
rect 117150 7090 117160 7730
rect 117200 7090 117210 7730
rect 117150 7070 117210 7090
rect 117270 7730 117330 7900
rect 117380 7860 117460 7870
rect 117380 7800 117390 7860
rect 117450 7800 117460 7860
rect 117380 7790 117460 7800
rect 117270 7090 117280 7730
rect 117320 7090 117330 7730
rect 117270 7060 117330 7090
rect 117390 7730 117450 7790
rect 117390 7090 117400 7730
rect 117440 7090 117450 7730
rect 117390 7070 117450 7090
rect 117510 7730 117570 7900
rect 117620 7860 117700 8420
rect 118340 8640 118420 8650
rect 118340 8580 118350 8640
rect 118410 8580 118420 8640
rect 118340 8560 118420 8580
rect 118340 8500 118350 8560
rect 118410 8500 118420 8560
rect 118340 8480 118420 8500
rect 118340 8420 118350 8480
rect 118410 8420 118420 8480
rect 117740 8370 117820 8380
rect 117740 8310 117750 8370
rect 117810 8310 117820 8370
rect 117740 8290 117820 8310
rect 117740 8230 117750 8290
rect 117810 8230 117820 8290
rect 117740 8210 117820 8230
rect 117740 8150 117750 8210
rect 117810 8150 117820 8210
rect 117740 8130 117820 8150
rect 117740 8070 117750 8130
rect 117810 8070 117820 8130
rect 117740 8050 117820 8070
rect 117740 7990 117750 8050
rect 117810 7990 117820 8050
rect 117740 7970 117820 7990
rect 117740 7910 117750 7970
rect 117810 7910 117820 7970
rect 117740 7900 117820 7910
rect 117980 8370 118060 8380
rect 117980 8310 117990 8370
rect 118050 8310 118060 8370
rect 117980 8290 118060 8310
rect 117980 8230 117990 8290
rect 118050 8230 118060 8290
rect 117980 8210 118060 8230
rect 117980 8150 117990 8210
rect 118050 8150 118060 8210
rect 117980 8130 118060 8150
rect 117980 8070 117990 8130
rect 118050 8070 118060 8130
rect 117980 8050 118060 8070
rect 117980 7990 117990 8050
rect 118050 7990 118060 8050
rect 117980 7970 118060 7990
rect 117980 7910 117990 7970
rect 118050 7910 118060 7970
rect 117980 7900 118060 7910
rect 118220 8370 118300 8380
rect 118220 8310 118230 8370
rect 118290 8310 118300 8370
rect 118220 8290 118300 8310
rect 118220 8230 118230 8290
rect 118290 8230 118300 8290
rect 118220 8210 118300 8230
rect 118220 8150 118230 8210
rect 118290 8150 118300 8210
rect 118220 8130 118300 8150
rect 118220 8070 118230 8130
rect 118290 8070 118300 8130
rect 118220 8050 118300 8070
rect 118220 7990 118230 8050
rect 118290 7990 118300 8050
rect 118220 7970 118300 7990
rect 118220 7910 118230 7970
rect 118290 7910 118300 7970
rect 118220 7900 118300 7910
rect 117620 7800 117630 7860
rect 117690 7800 117700 7860
rect 117620 7790 117700 7800
rect 117510 7090 117520 7730
rect 117560 7090 117570 7730
rect 117510 7060 117570 7090
rect 117630 7730 117690 7790
rect 117630 7090 117640 7730
rect 117680 7090 117690 7730
rect 117630 7070 117690 7090
rect 117750 7730 117810 7900
rect 117860 7860 117940 7870
rect 117860 7800 117870 7860
rect 117930 7800 117940 7860
rect 117860 7790 117940 7800
rect 117750 7090 117760 7730
rect 117800 7090 117810 7730
rect 117750 7060 117810 7090
rect 117870 7730 117930 7790
rect 117870 7090 117880 7730
rect 117920 7090 117930 7730
rect 117870 7070 117930 7090
rect 117990 7730 118050 7900
rect 118100 7860 118180 7870
rect 118100 7800 118110 7860
rect 118170 7800 118180 7860
rect 118100 7790 118180 7800
rect 117990 7090 118000 7730
rect 118040 7090 118050 7730
rect 117990 7060 118050 7090
rect 118110 7730 118170 7790
rect 118110 7090 118120 7730
rect 118160 7090 118170 7730
rect 118110 7070 118170 7090
rect 118230 7730 118290 7900
rect 118340 7860 118420 8420
rect 119280 8640 119520 12220
rect 119280 8580 119290 8640
rect 119350 8580 119370 8640
rect 119430 8580 119450 8640
rect 119510 8580 119520 8640
rect 119280 8560 119520 8580
rect 119280 8500 119290 8560
rect 119350 8500 119370 8560
rect 119430 8500 119450 8560
rect 119510 8500 119520 8560
rect 119280 8480 119520 8500
rect 119280 8420 119290 8480
rect 119350 8420 119370 8480
rect 119430 8420 119450 8480
rect 119510 8420 119520 8480
rect 119280 8410 119520 8420
rect 120680 8640 120920 12220
rect 120680 8580 120690 8640
rect 120750 8580 120770 8640
rect 120830 8580 120850 8640
rect 120910 8580 120920 8640
rect 120680 8560 120920 8580
rect 120680 8500 120690 8560
rect 120750 8500 120770 8560
rect 120830 8500 120850 8560
rect 120910 8500 120920 8560
rect 120680 8480 120920 8500
rect 120680 8420 120690 8480
rect 120750 8420 120770 8480
rect 120830 8420 120850 8480
rect 120910 8420 120920 8480
rect 120680 8410 120920 8420
rect 121380 8640 121620 12220
rect 121380 8580 121390 8640
rect 121450 8580 121470 8640
rect 121530 8580 121550 8640
rect 121610 8580 121620 8640
rect 121380 8560 121620 8580
rect 121380 8500 121390 8560
rect 121450 8500 121470 8560
rect 121530 8500 121550 8560
rect 121610 8500 121620 8560
rect 121380 8480 121620 8500
rect 121380 8420 121390 8480
rect 121450 8420 121470 8480
rect 121530 8420 121550 8480
rect 121610 8420 121620 8480
rect 121380 8410 121620 8420
rect 122080 8640 122320 12220
rect 122080 8580 122090 8640
rect 122150 8580 122170 8640
rect 122230 8580 122250 8640
rect 122310 8580 122320 8640
rect 122080 8560 122320 8580
rect 122080 8500 122090 8560
rect 122150 8500 122170 8560
rect 122230 8500 122250 8560
rect 122310 8500 122320 8560
rect 122080 8480 122320 8500
rect 122080 8420 122090 8480
rect 122150 8420 122170 8480
rect 122230 8420 122250 8480
rect 122310 8420 122320 8480
rect 122080 8410 122320 8420
rect 122780 8640 123020 12220
rect 122780 8580 122790 8640
rect 122850 8580 122870 8640
rect 122930 8580 122950 8640
rect 123010 8580 123020 8640
rect 122780 8560 123020 8580
rect 122780 8500 122790 8560
rect 122850 8500 122870 8560
rect 122930 8500 122950 8560
rect 123010 8500 123020 8560
rect 122780 8480 123020 8500
rect 122780 8420 122790 8480
rect 122850 8420 122870 8480
rect 122930 8420 122950 8480
rect 123010 8420 123020 8480
rect 122780 8410 123020 8420
rect 118340 7800 118350 7860
rect 118410 7800 118420 7860
rect 118340 7790 118420 7800
rect 118230 7090 118240 7730
rect 118280 7090 118290 7730
rect 118230 7060 118290 7090
rect 118350 7730 118410 7790
rect 118350 7090 118360 7730
rect 118400 7090 118410 7730
rect 116910 6970 116920 7010
rect 116960 6970 116970 7010
rect 117020 7050 117100 7060
rect 117020 6990 117030 7050
rect 117090 6990 117100 7050
rect 117020 6980 117100 6990
rect 117260 7050 117340 7060
rect 117260 6990 117270 7050
rect 117330 6990 117340 7050
rect 117260 6980 117340 6990
rect 117500 7050 117580 7060
rect 117500 6990 117510 7050
rect 117570 6990 117580 7050
rect 117500 6980 117580 6990
rect 117740 7050 117820 7060
rect 117740 6990 117750 7050
rect 117810 6990 117820 7050
rect 117740 6980 117820 6990
rect 117980 7050 118060 7060
rect 117980 6990 117990 7050
rect 118050 6990 118060 7050
rect 117980 6980 118060 6990
rect 118220 7050 118300 7060
rect 118220 6990 118230 7050
rect 118290 6990 118300 7050
rect 118220 6980 118300 6990
rect 118350 7010 118410 7090
rect 116910 6950 116970 6970
rect 118350 6970 118360 7010
rect 118400 6970 118410 7010
rect 118350 6950 118410 6970
rect 117090 6940 117150 6950
rect 117090 6870 117150 6880
rect 117210 6940 117270 6950
rect 117210 6870 117270 6880
rect 117330 6940 117390 6950
rect 117330 6870 117390 6880
rect 117450 6940 117510 6950
rect 117450 6870 117510 6880
rect 117570 6940 117750 6950
rect 117630 6880 117690 6940
rect 117570 6870 117750 6880
rect 117810 6940 117870 6950
rect 117810 6870 117870 6880
rect 117930 6940 117990 6950
rect 117930 6870 117990 6880
rect 118050 6940 118110 6950
rect 118050 6870 118110 6880
rect 118170 6940 118230 6950
rect 118170 6870 118230 6880
rect 117620 6820 117700 6870
rect 117620 6760 117630 6820
rect 117690 6760 117700 6820
rect 117620 6750 117700 6760
rect 119010 6750 119090 6760
rect 116960 6710 117040 6720
rect 116960 6650 116970 6710
rect 117030 6650 117040 6710
rect 116960 6630 117040 6650
rect 116960 6570 116970 6630
rect 117030 6570 117040 6630
rect 116960 6550 117040 6570
rect 116960 6490 116970 6550
rect 117030 6490 117040 6550
rect 116960 6480 117040 6490
rect 117180 6710 117260 6720
rect 117180 6650 117190 6710
rect 117250 6650 117260 6710
rect 117180 6630 117260 6650
rect 117180 6570 117190 6630
rect 117250 6570 117260 6630
rect 117180 6550 117260 6570
rect 117180 6490 117190 6550
rect 117250 6490 117260 6550
rect 117180 6480 117260 6490
rect 117400 6710 117480 6720
rect 117400 6650 117410 6710
rect 117470 6650 117480 6710
rect 117400 6630 117480 6650
rect 117400 6570 117410 6630
rect 117470 6570 117480 6630
rect 117400 6550 117480 6570
rect 117400 6490 117410 6550
rect 117470 6490 117480 6550
rect 117400 6480 117480 6490
rect 117620 6710 117700 6720
rect 117620 6650 117630 6710
rect 117690 6650 117700 6710
rect 117620 6630 117700 6650
rect 117620 6570 117630 6630
rect 117690 6570 117700 6630
rect 117620 6550 117700 6570
rect 117620 6490 117630 6550
rect 117690 6490 117700 6550
rect 117620 6480 117700 6490
rect 117840 6710 117920 6720
rect 117840 6650 117850 6710
rect 117910 6650 117920 6710
rect 117840 6630 117920 6650
rect 117840 6570 117850 6630
rect 117910 6570 117920 6630
rect 117840 6550 117920 6570
rect 117840 6490 117850 6550
rect 117910 6490 117920 6550
rect 117840 6480 117920 6490
rect 118060 6710 118140 6720
rect 118060 6650 118070 6710
rect 118130 6650 118140 6710
rect 118060 6630 118140 6650
rect 118060 6570 118070 6630
rect 118130 6570 118140 6630
rect 118060 6550 118140 6570
rect 118060 6490 118070 6550
rect 118130 6490 118140 6550
rect 118060 6480 118140 6490
rect 118280 6710 118360 6720
rect 118280 6650 118290 6710
rect 118350 6650 118360 6710
rect 118280 6630 118360 6650
rect 118280 6570 118290 6630
rect 118350 6570 118360 6630
rect 118280 6550 118360 6570
rect 118280 6490 118290 6550
rect 118350 6490 118360 6550
rect 118280 6480 118360 6490
rect 119010 6690 119020 6750
rect 119080 6690 119090 6750
rect 116970 6400 117030 6480
rect 116970 6360 116980 6400
rect 117020 6360 117030 6400
rect 116970 6280 117030 6360
rect 117070 6380 117150 6390
rect 117070 6320 117080 6380
rect 117140 6320 117150 6380
rect 117070 6310 117150 6320
rect 116970 5140 116980 6280
rect 117020 5140 117030 6280
rect 116970 5120 117030 5140
rect 117080 6280 117140 6310
rect 117080 5140 117090 6280
rect 117130 5140 117140 6280
rect 117080 5110 117140 5140
rect 117190 6280 117250 6480
rect 117290 6380 117370 6390
rect 117290 6320 117300 6380
rect 117360 6320 117370 6380
rect 117290 6310 117370 6320
rect 117190 5140 117200 6280
rect 117240 5140 117250 6280
rect 117190 5120 117250 5140
rect 117300 6280 117360 6310
rect 117300 5140 117310 6280
rect 117350 5140 117360 6280
rect 117300 5110 117360 5140
rect 117410 6280 117470 6480
rect 117510 6380 117590 6390
rect 117510 6320 117520 6380
rect 117580 6320 117590 6380
rect 117510 6310 117590 6320
rect 117410 5140 117420 6280
rect 117460 5140 117470 6280
rect 117410 5120 117470 5140
rect 117520 6280 117580 6310
rect 117520 5140 117530 6280
rect 117570 5140 117580 6280
rect 117520 5110 117580 5140
rect 117630 6280 117690 6480
rect 117730 6380 117810 6390
rect 117730 6320 117740 6380
rect 117800 6320 117810 6380
rect 117730 6310 117810 6320
rect 117630 5140 117640 6280
rect 117680 5140 117690 6280
rect 117630 5120 117690 5140
rect 117740 6280 117800 6310
rect 117740 5140 117750 6280
rect 117790 5140 117800 6280
rect 117740 5110 117800 5140
rect 117850 6280 117910 6480
rect 117950 6380 118030 6390
rect 117950 6320 117960 6380
rect 118020 6320 118030 6380
rect 117950 6310 118030 6320
rect 117850 5140 117860 6280
rect 117900 5140 117910 6280
rect 117850 5120 117910 5140
rect 117960 6280 118020 6310
rect 117960 5140 117970 6280
rect 118010 5140 118020 6280
rect 117960 5110 118020 5140
rect 118070 6280 118130 6480
rect 118290 6400 118350 6480
rect 119010 6400 119090 6690
rect 118170 6380 118250 6390
rect 118170 6320 118180 6380
rect 118240 6320 118250 6380
rect 118170 6310 118250 6320
rect 118290 6360 118300 6400
rect 118340 6360 118350 6400
rect 118070 5140 118080 6280
rect 118120 5140 118130 6280
rect 118070 5120 118130 5140
rect 118180 6280 118240 6310
rect 118180 5140 118190 6280
rect 118230 5140 118240 6280
rect 118180 5110 118240 5140
rect 118290 6280 118350 6360
rect 118910 6380 119192 6400
rect 118910 6340 118920 6380
rect 118960 6340 119030 6380
rect 119070 6340 119140 6380
rect 119180 6340 119192 6380
rect 118910 6320 119192 6340
rect 118290 5140 118300 6280
rect 118340 5140 118350 6280
rect 118290 5120 118350 5140
rect 118910 5170 119192 5190
rect 118910 5130 118920 5170
rect 118960 5130 119030 5170
rect 119070 5130 119140 5170
rect 119180 5130 119192 5170
rect 118910 5110 119192 5130
rect 116560 4880 116570 4940
rect 116630 4880 116650 4940
rect 116710 4880 116730 4940
rect 116790 4880 116800 4940
rect 116560 4860 116800 4880
rect 116560 4800 116570 4860
rect 116630 4800 116650 4860
rect 116710 4800 116730 4860
rect 116790 4800 116800 4860
rect 116560 4780 116800 4800
rect 116560 4720 116570 4780
rect 116630 4720 116650 4780
rect 116710 4720 116730 4780
rect 116790 4720 116800 4780
rect 116560 3190 116800 4720
rect 117070 5100 117150 5110
rect 117070 5040 117080 5100
rect 117140 5040 117150 5100
rect 117070 4650 117150 5040
rect 117290 5100 117370 5110
rect 117290 5040 117300 5100
rect 117360 5040 117370 5100
rect 117290 4650 117370 5040
rect 117510 5100 117590 5110
rect 117510 5040 117520 5100
rect 117580 5040 117590 5100
rect 117510 4650 117590 5040
rect 117730 5100 117810 5110
rect 117730 5040 117740 5100
rect 117800 5040 117810 5100
rect 117620 4940 117700 4950
rect 117620 4880 117630 4940
rect 117690 4880 117700 4940
rect 117620 4860 117700 4880
rect 117620 4800 117630 4860
rect 117690 4800 117700 4860
rect 117620 4780 117700 4800
rect 117620 4720 117630 4780
rect 117690 4720 117700 4780
rect 117620 4710 117700 4720
rect 117730 4650 117810 5040
rect 117950 5100 118030 5110
rect 117950 5040 117960 5100
rect 118020 5040 118030 5100
rect 117950 4650 118030 5040
rect 118170 5100 118250 5110
rect 118170 5040 118180 5100
rect 118240 5040 118250 5100
rect 118170 4650 118250 5040
rect 118930 4940 119170 5110
rect 118930 4880 118940 4940
rect 119000 4880 119020 4940
rect 119080 4880 119100 4940
rect 119160 4880 119170 4940
rect 118930 4860 119170 4880
rect 118930 4800 118940 4860
rect 119000 4800 119020 4860
rect 119080 4800 119100 4860
rect 119160 4800 119170 4860
rect 118930 4780 119170 4800
rect 118930 4720 118940 4780
rect 119000 4720 119020 4780
rect 119080 4720 119100 4780
rect 119160 4720 119170 4780
rect 118930 4710 119170 4720
rect 117070 4640 118250 4650
rect 117070 4580 117080 4640
rect 117140 4580 117190 4640
rect 117250 4580 117300 4640
rect 117360 4580 117410 4640
rect 117470 4580 117520 4640
rect 117580 4580 117630 4640
rect 117690 4580 117740 4640
rect 117800 4580 117850 4640
rect 117910 4580 117960 4640
rect 118020 4580 118070 4640
rect 118130 4580 118180 4640
rect 118240 4580 118250 4640
rect 117070 4560 118250 4580
rect 117070 4500 117080 4560
rect 117140 4500 117190 4560
rect 117250 4500 117300 4560
rect 117360 4500 117410 4560
rect 117470 4500 117520 4560
rect 117580 4500 117630 4560
rect 117690 4500 117740 4560
rect 117800 4500 117850 4560
rect 117910 4500 117960 4560
rect 118020 4500 118070 4560
rect 118130 4500 118180 4560
rect 118240 4500 118250 4560
rect 117070 4480 118250 4500
rect 117070 4420 117080 4480
rect 117140 4420 117190 4480
rect 117250 4420 117300 4480
rect 117360 4420 117410 4480
rect 117470 4420 117520 4480
rect 117580 4420 117630 4480
rect 117690 4420 117740 4480
rect 117800 4420 117850 4480
rect 117910 4420 117960 4480
rect 118020 4420 118070 4480
rect 118130 4420 118180 4480
rect 118240 4420 118250 4480
rect 117070 4410 118250 4420
rect 119120 4640 119620 4650
rect 119120 4580 119130 4640
rect 119190 4580 119210 4640
rect 119270 4580 119300 4640
rect 119360 4580 119380 4640
rect 119440 4580 119470 4640
rect 119530 4580 119550 4640
rect 119610 4580 119620 4640
rect 119120 4560 119620 4580
rect 119120 4500 119130 4560
rect 119190 4500 119210 4560
rect 119270 4500 119300 4560
rect 119360 4500 119380 4560
rect 119440 4500 119470 4560
rect 119530 4500 119550 4560
rect 119610 4500 119620 4560
rect 119120 4480 119620 4500
rect 119120 4420 119130 4480
rect 119190 4420 119210 4480
rect 119270 4420 119300 4480
rect 119360 4420 119380 4480
rect 119440 4420 119470 4480
rect 119530 4420 119550 4480
rect 119610 4420 119620 4480
rect 116960 4370 117040 4380
rect 116960 4310 116970 4370
rect 117030 4310 117040 4370
rect 116960 4290 117040 4310
rect 116960 4230 116970 4290
rect 117030 4230 117040 4290
rect 116960 4210 117040 4230
rect 116960 4150 116970 4210
rect 117030 4150 117040 4210
rect 116960 4140 117040 4150
rect 118280 4370 118360 4380
rect 118280 4310 118290 4370
rect 118350 4310 118360 4370
rect 118280 4290 118360 4310
rect 118280 4230 118290 4290
rect 118350 4230 118360 4290
rect 118280 4210 118360 4230
rect 118280 4150 118290 4210
rect 118350 4150 118360 4210
rect 118280 4140 118360 4150
rect 116970 3850 117030 4140
rect 117070 4100 117150 4110
rect 117070 4040 117080 4100
rect 117140 4040 117150 4100
rect 117070 4020 117150 4040
rect 117070 3960 117080 4020
rect 117140 3960 117150 4020
rect 117070 3940 117150 3960
rect 117070 3880 117080 3940
rect 117140 3880 117150 3940
rect 117070 3870 117150 3880
rect 117290 4100 117370 4110
rect 117290 4040 117300 4100
rect 117360 4040 117370 4100
rect 117290 4020 117370 4040
rect 117290 3960 117300 4020
rect 117360 3960 117370 4020
rect 117290 3940 117370 3960
rect 117290 3880 117300 3940
rect 117360 3880 117370 3940
rect 117290 3870 117370 3880
rect 117510 4100 117590 4110
rect 117510 4040 117520 4100
rect 117580 4040 117590 4100
rect 117510 4020 117590 4040
rect 117510 3960 117520 4020
rect 117580 3960 117590 4020
rect 117510 3940 117590 3960
rect 117510 3880 117520 3940
rect 117580 3880 117590 3940
rect 117510 3870 117590 3880
rect 117730 4100 117810 4110
rect 117730 4040 117740 4100
rect 117800 4040 117810 4100
rect 117730 4020 117810 4040
rect 117730 3960 117740 4020
rect 117800 3960 117810 4020
rect 117730 3940 117810 3960
rect 117730 3880 117740 3940
rect 117800 3880 117810 3940
rect 117730 3870 117810 3880
rect 117950 4100 118030 4110
rect 117950 4040 117960 4100
rect 118020 4040 118030 4100
rect 117950 4020 118030 4040
rect 117950 3960 117960 4020
rect 118020 3960 118030 4020
rect 117950 3940 118030 3960
rect 117950 3880 117960 3940
rect 118020 3880 118030 3940
rect 117950 3870 118030 3880
rect 118170 4100 118250 4110
rect 118170 4040 118180 4100
rect 118240 4040 118250 4100
rect 118170 4020 118250 4040
rect 118170 3960 118180 4020
rect 118240 3960 118250 4020
rect 118170 3940 118250 3960
rect 118170 3880 118180 3940
rect 118240 3880 118250 3940
rect 118170 3870 118250 3880
rect 116970 3810 116980 3850
rect 117020 3810 117030 3850
rect 116970 3730 117030 3810
rect 116970 3390 116980 3730
rect 117020 3390 117030 3730
rect 116970 3370 117030 3390
rect 117080 3730 117140 3870
rect 117180 3830 117260 3840
rect 117180 3770 117190 3830
rect 117250 3770 117260 3830
rect 117180 3760 117260 3770
rect 117080 3390 117090 3730
rect 117130 3390 117140 3730
rect 117080 3370 117140 3390
rect 117190 3730 117250 3760
rect 117190 3390 117200 3730
rect 117240 3390 117250 3730
rect 117190 3330 117250 3390
rect 117300 3730 117360 3870
rect 117400 3830 117480 3840
rect 117400 3770 117410 3830
rect 117470 3770 117480 3830
rect 117400 3760 117480 3770
rect 117300 3390 117310 3730
rect 117350 3390 117360 3730
rect 117300 3370 117360 3390
rect 117410 3730 117470 3760
rect 117410 3390 117420 3730
rect 117460 3390 117470 3730
rect 117410 3330 117470 3390
rect 117520 3730 117580 3870
rect 117620 3830 117700 3840
rect 117620 3770 117630 3830
rect 117690 3770 117700 3830
rect 117620 3760 117700 3770
rect 117520 3390 117530 3730
rect 117570 3390 117580 3730
rect 117520 3370 117580 3390
rect 117630 3730 117690 3760
rect 117630 3390 117640 3730
rect 117680 3390 117690 3730
rect 117630 3330 117690 3390
rect 117740 3730 117800 3870
rect 117840 3830 117920 3840
rect 117840 3770 117850 3830
rect 117910 3770 117920 3830
rect 117840 3760 117920 3770
rect 117740 3390 117750 3730
rect 117790 3390 117800 3730
rect 117740 3370 117800 3390
rect 117850 3730 117910 3760
rect 117850 3390 117860 3730
rect 117900 3390 117910 3730
rect 117850 3330 117910 3390
rect 117960 3730 118020 3870
rect 118060 3830 118140 3840
rect 118060 3770 118070 3830
rect 118130 3770 118140 3830
rect 118060 3760 118140 3770
rect 117960 3390 117970 3730
rect 118010 3390 118020 3730
rect 117960 3370 118020 3390
rect 118070 3730 118130 3760
rect 118070 3390 118080 3730
rect 118120 3390 118130 3730
rect 118070 3330 118130 3390
rect 118180 3730 118240 3870
rect 118180 3390 118190 3730
rect 118230 3390 118240 3730
rect 118180 3370 118240 3390
rect 118290 3850 118350 4140
rect 118290 3810 118300 3850
rect 118340 3810 118350 3850
rect 118290 3730 118350 3810
rect 118290 3390 118300 3730
rect 118340 3390 118350 3730
rect 118290 3370 118350 3390
rect 119120 3420 119620 4420
rect 119120 3360 119140 3420
rect 119200 3360 119240 3420
rect 119300 3360 119340 3420
rect 119400 3360 119440 3420
rect 119500 3360 119540 3420
rect 119600 3360 119620 3420
rect 117180 3320 117260 3330
rect 117180 3260 117190 3320
rect 117250 3260 117260 3320
rect 117180 3250 117260 3260
rect 117400 3320 117480 3330
rect 117400 3260 117410 3320
rect 117470 3260 117480 3320
rect 117400 3250 117480 3260
rect 117620 3320 117700 3330
rect 117620 3260 117630 3320
rect 117690 3260 117700 3320
rect 117620 3250 117700 3260
rect 117840 3320 117920 3330
rect 117840 3260 117850 3320
rect 117910 3260 117920 3320
rect 117840 3250 117920 3260
rect 118060 3320 118140 3330
rect 118060 3260 118070 3320
rect 118130 3260 118140 3320
rect 118060 3250 118140 3260
rect 118550 3320 118630 3330
rect 118550 3260 118560 3320
rect 118620 3260 118630 3320
rect 118550 3250 118630 3260
rect 119120 3320 119620 3360
rect 119120 3260 119140 3320
rect 119200 3260 119240 3320
rect 119300 3260 119340 3320
rect 119400 3260 119440 3320
rect 119500 3260 119540 3320
rect 119600 3260 119620 3320
rect 116560 3130 116570 3190
rect 116630 3130 116650 3190
rect 116710 3130 116730 3190
rect 116790 3130 116800 3190
rect 116560 3110 116800 3130
rect 116560 3050 116570 3110
rect 116630 3050 116650 3110
rect 116710 3050 116730 3110
rect 116790 3050 116800 3110
rect 116560 3040 116800 3050
rect 117290 3190 117370 3200
rect 117290 3130 117300 3190
rect 117360 3130 117370 3190
rect 117290 3110 117370 3130
rect 117290 3050 117300 3110
rect 117360 3050 117370 3110
rect 117290 3040 117370 3050
rect 117180 2950 117260 2960
rect 117180 2890 117190 2950
rect 117250 2890 117260 2950
rect 117180 2880 117260 2890
rect 117400 2950 117480 2960
rect 117400 2890 117410 2950
rect 117470 2890 117480 2950
rect 117400 2880 117480 2890
rect 117620 2950 117700 2960
rect 117620 2890 117630 2950
rect 117690 2890 117700 2950
rect 117620 2880 117700 2890
rect 117840 2950 117920 2960
rect 117840 2890 117850 2950
rect 117910 2890 117920 2950
rect 117840 2880 117920 2890
rect 118060 2950 118140 2960
rect 118060 2890 118070 2950
rect 118130 2890 118140 2950
rect 118060 2880 118140 2890
rect 118460 2950 118540 2960
rect 118460 2890 118470 2950
rect 118530 2890 118540 2950
rect 118460 2880 118540 2890
rect 116290 2100 116300 2160
rect 116360 2100 116380 2160
rect 116440 2100 116460 2160
rect 116520 2100 116530 2160
rect 116290 2080 116530 2100
rect 116290 2020 116300 2080
rect 116360 2020 116380 2080
rect 116440 2020 116460 2080
rect 116520 2020 116530 2080
rect 116290 2000 116530 2020
rect 116290 1940 116300 2000
rect 116360 1940 116380 2000
rect 116440 1940 116460 2000
rect 116520 1940 116530 2000
rect 116290 1930 116530 1940
rect 116970 2850 117030 2870
rect 116970 2310 116980 2850
rect 117020 2310 117030 2850
rect 116970 2230 117030 2310
rect 116970 2190 116980 2230
rect 117020 2190 117030 2230
rect 116970 1890 117030 2190
rect 117080 2850 117140 2870
rect 117080 2310 117090 2850
rect 117130 2310 117140 2850
rect 117080 2170 117140 2310
rect 117190 2850 117250 2880
rect 117190 2310 117200 2850
rect 117240 2310 117250 2850
rect 117190 2280 117250 2310
rect 117300 2850 117360 2870
rect 117300 2310 117310 2850
rect 117350 2310 117360 2850
rect 117180 2270 117260 2280
rect 117180 2210 117190 2270
rect 117250 2210 117260 2270
rect 117180 2200 117260 2210
rect 117300 2170 117360 2310
rect 117410 2850 117470 2880
rect 117410 2310 117420 2850
rect 117460 2310 117470 2850
rect 117410 2280 117470 2310
rect 117520 2850 117580 2870
rect 117520 2310 117530 2850
rect 117570 2310 117580 2850
rect 117400 2270 117480 2280
rect 117400 2210 117410 2270
rect 117470 2210 117480 2270
rect 117400 2200 117480 2210
rect 117520 2170 117580 2310
rect 117630 2850 117690 2880
rect 117630 2310 117640 2850
rect 117680 2310 117690 2850
rect 117630 2280 117690 2310
rect 117740 2850 117800 2870
rect 117740 2310 117750 2850
rect 117790 2310 117800 2850
rect 117620 2270 117700 2280
rect 117620 2210 117630 2270
rect 117690 2210 117700 2270
rect 117620 2200 117700 2210
rect 117740 2170 117800 2310
rect 117850 2850 117910 2880
rect 117850 2310 117860 2850
rect 117900 2310 117910 2850
rect 117850 2280 117910 2310
rect 117960 2850 118020 2870
rect 117960 2310 117970 2850
rect 118010 2310 118020 2850
rect 117840 2270 117920 2280
rect 117840 2210 117850 2270
rect 117910 2210 117920 2270
rect 117840 2200 117920 2210
rect 117960 2170 118020 2310
rect 118070 2850 118130 2880
rect 118070 2310 118080 2850
rect 118120 2310 118130 2850
rect 118070 2280 118130 2310
rect 118180 2850 118240 2870
rect 118180 2310 118190 2850
rect 118230 2310 118240 2850
rect 118060 2270 118140 2280
rect 118060 2210 118070 2270
rect 118130 2210 118140 2270
rect 118060 2200 118140 2210
rect 118180 2170 118240 2310
rect 118290 2850 118350 2870
rect 118290 2310 118300 2850
rect 118340 2310 118350 2850
rect 118480 2320 118520 2880
rect 118290 2230 118350 2310
rect 118460 2310 118540 2320
rect 118460 2250 118470 2310
rect 118530 2250 118540 2310
rect 118460 2240 118540 2250
rect 118290 2190 118300 2230
rect 118340 2190 118350 2230
rect 117070 2160 117150 2170
rect 117070 2100 117080 2160
rect 117140 2100 117150 2160
rect 117070 2080 117150 2100
rect 117070 2020 117080 2080
rect 117140 2020 117150 2080
rect 117070 2000 117150 2020
rect 117070 1940 117080 2000
rect 117140 1940 117150 2000
rect 117070 1930 117150 1940
rect 117290 2160 117370 2170
rect 117290 2100 117300 2160
rect 117360 2100 117370 2160
rect 117290 2080 117370 2100
rect 117290 2020 117300 2080
rect 117360 2020 117370 2080
rect 117290 2000 117370 2020
rect 117290 1940 117300 2000
rect 117360 1940 117370 2000
rect 117290 1930 117370 1940
rect 117510 2160 117590 2170
rect 117510 2100 117520 2160
rect 117580 2100 117590 2160
rect 117510 2080 117590 2100
rect 117510 2020 117520 2080
rect 117580 2020 117590 2080
rect 117510 2000 117590 2020
rect 117510 1940 117520 2000
rect 117580 1940 117590 2000
rect 117510 1930 117590 1940
rect 117730 2160 117810 2170
rect 117730 2100 117740 2160
rect 117800 2100 117810 2160
rect 117730 2080 117810 2100
rect 117730 2020 117740 2080
rect 117800 2020 117810 2080
rect 117730 2000 117810 2020
rect 117730 1940 117740 2000
rect 117800 1940 117810 2000
rect 117730 1930 117810 1940
rect 117950 2160 118030 2170
rect 117950 2100 117960 2160
rect 118020 2100 118030 2160
rect 117950 2080 118030 2100
rect 117950 2020 117960 2080
rect 118020 2020 118030 2080
rect 117950 2000 118030 2020
rect 117950 1940 117960 2000
rect 118020 1940 118030 2000
rect 117950 1930 118030 1940
rect 118170 2160 118250 2170
rect 118170 2100 118180 2160
rect 118240 2100 118250 2160
rect 118170 2080 118250 2100
rect 118170 2020 118180 2080
rect 118240 2020 118250 2080
rect 118170 2000 118250 2020
rect 118170 1940 118180 2000
rect 118240 1940 118250 2000
rect 118170 1930 118250 1940
rect 118290 1890 118350 2190
rect 118570 2180 118610 3250
rect 119120 3220 119620 3260
rect 119120 3160 119140 3220
rect 119200 3160 119240 3220
rect 119300 3160 119340 3220
rect 119400 3160 119440 3220
rect 119500 3160 119540 3220
rect 119600 3160 119620 3220
rect 118660 2320 118730 2330
rect 118660 2240 118730 2250
rect 118780 2320 118850 2330
rect 118780 2240 118850 2250
rect 118900 2320 118970 2330
rect 118900 2240 118970 2250
rect 119020 2320 119090 2332
rect 119020 2240 119090 2250
rect 118790 2180 118830 2240
rect 118550 2170 118630 2180
rect 118550 2110 118560 2170
rect 118620 2110 118630 2170
rect 118550 2100 118630 2110
rect 118770 2170 118850 2180
rect 118770 2110 118780 2170
rect 118840 2110 118850 2170
rect 118770 2100 118850 2110
rect 116960 1880 117040 1890
rect 116960 1820 116970 1880
rect 117030 1820 117040 1880
rect 116960 1800 117040 1820
rect 116960 1740 116970 1800
rect 117030 1740 117040 1800
rect 116960 1720 117040 1740
rect 116960 1660 116970 1720
rect 117030 1660 117040 1720
rect 116960 1650 117040 1660
rect 118280 1880 118360 1890
rect 118280 1820 118290 1880
rect 118350 1820 118360 1880
rect 118280 1800 118360 1820
rect 118280 1740 118290 1800
rect 118350 1740 118360 1800
rect 118280 1720 118360 1740
rect 118280 1660 118290 1720
rect 118350 1660 118360 1720
rect 118280 1650 118360 1660
rect 119030 1620 119070 2240
rect 119010 1610 119090 1620
rect 119010 1550 119020 1610
rect 119080 1550 119090 1610
rect 119010 1540 119090 1550
rect 118880 1150 118960 1160
rect 118880 1090 118890 1150
rect 118950 1090 118960 1150
rect 117220 1040 118100 1050
rect 117220 980 117230 1040
rect 117290 980 117310 1040
rect 117370 980 117390 1040
rect 117450 980 117470 1040
rect 117530 980 117550 1040
rect 117610 980 117630 1040
rect 117690 980 117710 1040
rect 117770 980 117790 1040
rect 117850 980 117870 1040
rect 117930 980 117950 1040
rect 118010 980 118030 1040
rect 118090 980 118100 1040
rect 117220 960 118100 980
rect 117220 900 117230 960
rect 117290 900 117310 960
rect 117370 900 117390 960
rect 117450 900 117470 960
rect 117530 900 117550 960
rect 117610 900 117630 960
rect 117690 900 117710 960
rect 117770 900 117790 960
rect 117850 900 117870 960
rect 117930 900 117950 960
rect 118010 900 118030 960
rect 118090 900 118100 960
rect 117220 880 118100 900
rect 117220 820 117230 880
rect 117290 820 117310 880
rect 117370 820 117390 880
rect 117450 820 117470 880
rect 117530 820 117550 880
rect 117610 820 117630 880
rect 117690 820 117710 880
rect 117770 820 117790 880
rect 117850 820 117870 880
rect 117930 820 117950 880
rect 118010 820 118030 880
rect 118090 820 118100 880
rect 117220 810 118100 820
rect 118750 1040 118830 1050
rect 118750 980 118760 1040
rect 118820 980 118830 1040
rect 118750 960 118830 980
rect 118750 900 118760 960
rect 118820 900 118830 960
rect 118750 880 118830 900
rect 118750 820 118760 880
rect 118820 820 118830 880
rect 118750 810 118830 820
rect 116020 -180 116030 -120
rect 116090 -180 116110 -120
rect 116170 -180 116190 -120
rect 116250 -180 116260 -120
rect 116020 -200 116260 -180
rect 116020 -260 116030 -200
rect 116090 -260 116110 -200
rect 116170 -260 116190 -200
rect 116250 -260 116260 -200
rect 116020 -280 116260 -260
rect 116020 -340 116030 -280
rect 116090 -340 116110 -280
rect 116170 -340 116190 -280
rect 116250 -340 116260 -280
rect 116020 -350 116260 -340
rect 117030 650 117090 670
rect 115420 -700 115430 -640
rect 115490 -700 115510 -640
rect 115570 -700 115590 -640
rect 115650 -700 115660 -640
rect 115420 -720 115660 -700
rect 115420 -780 115430 -720
rect 115490 -780 115510 -720
rect 115570 -780 115590 -720
rect 115650 -780 115660 -720
rect 115420 -800 115660 -780
rect 115420 -860 115430 -800
rect 115490 -860 115510 -800
rect 115570 -860 115590 -800
rect 115650 -860 115660 -800
rect 115420 -870 115660 -860
rect 117030 -690 117040 650
rect 117080 -690 117090 650
rect 117030 -770 117090 -690
rect 117230 650 117290 810
rect 117320 770 117400 780
rect 117320 710 117330 770
rect 117390 710 117400 770
rect 117320 700 117400 710
rect 117520 770 117600 780
rect 117520 710 117530 770
rect 117590 710 117600 770
rect 117520 700 117600 710
rect 117230 -690 117240 650
rect 117280 -690 117290 650
rect 117230 -720 117290 -690
rect 117430 650 117490 670
rect 117430 -690 117440 650
rect 117480 -690 117490 650
rect 117030 -810 117040 -770
rect 117080 -810 117090 -770
rect 117220 -730 117300 -720
rect 117220 -790 117230 -730
rect 117290 -790 117300 -730
rect 117220 -800 117300 -790
rect 117030 -1150 117090 -810
rect 117430 -1150 117490 -690
rect 117630 650 117690 810
rect 117720 770 117800 780
rect 117720 710 117730 770
rect 117790 710 117800 770
rect 117720 700 117800 710
rect 117920 770 118000 780
rect 117920 710 117930 770
rect 117990 710 118000 770
rect 117920 700 118000 710
rect 117630 -690 117640 650
rect 117680 -690 117690 650
rect 117630 -720 117690 -690
rect 117830 650 117890 670
rect 117830 -690 117840 650
rect 117880 -690 117890 650
rect 117620 -730 117700 -720
rect 117620 -790 117630 -730
rect 117690 -790 117700 -730
rect 117620 -800 117700 -790
rect 114970 -1220 114980 -1160
rect 115040 -1220 115050 -1160
rect 114970 -1240 115050 -1220
rect 114970 -1300 114980 -1240
rect 115040 -1300 115050 -1240
rect 114970 -1320 115050 -1300
rect 114970 -1380 114980 -1320
rect 115040 -1380 115050 -1320
rect 114970 -1390 115050 -1380
rect 115080 -1160 115320 -1150
rect 115080 -1220 115090 -1160
rect 115150 -1220 115170 -1160
rect 115230 -1220 115250 -1160
rect 115310 -1220 115320 -1160
rect 115080 -1240 115320 -1220
rect 115080 -1300 115090 -1240
rect 115150 -1300 115170 -1240
rect 115230 -1300 115250 -1240
rect 115310 -1300 115320 -1240
rect 115080 -1320 115320 -1300
rect 115080 -1380 115090 -1320
rect 115150 -1380 115170 -1320
rect 115230 -1380 115250 -1320
rect 115310 -1380 115320 -1320
rect 115080 -3000 115320 -1380
rect 115780 -1160 116020 -1150
rect 115780 -1220 115790 -1160
rect 115850 -1220 115870 -1160
rect 115930 -1220 115950 -1160
rect 116010 -1220 116020 -1160
rect 115780 -1240 116020 -1220
rect 115780 -1300 115790 -1240
rect 115850 -1300 115870 -1240
rect 115930 -1300 115950 -1240
rect 116010 -1300 116020 -1240
rect 115780 -1320 116020 -1300
rect 115780 -1380 115790 -1320
rect 115850 -1380 115870 -1320
rect 115930 -1380 115950 -1320
rect 116010 -1380 116020 -1320
rect 115780 -3000 116020 -1380
rect 116480 -1160 116720 -1150
rect 116480 -1220 116490 -1160
rect 116550 -1220 116570 -1160
rect 116630 -1220 116650 -1160
rect 116710 -1220 116720 -1160
rect 116480 -1240 116720 -1220
rect 116480 -1300 116490 -1240
rect 116550 -1300 116570 -1240
rect 116630 -1300 116650 -1240
rect 116710 -1300 116720 -1240
rect 116480 -1320 116720 -1300
rect 116480 -1380 116490 -1320
rect 116550 -1380 116570 -1320
rect 116630 -1380 116650 -1320
rect 116710 -1380 116720 -1320
rect 116480 -3000 116720 -1380
rect 117020 -1160 117100 -1150
rect 117020 -1220 117030 -1160
rect 117090 -1220 117100 -1160
rect 117020 -1240 117100 -1220
rect 117020 -1300 117030 -1240
rect 117090 -1300 117100 -1240
rect 117020 -1320 117100 -1300
rect 117020 -1380 117030 -1320
rect 117090 -1380 117100 -1320
rect 117020 -1390 117100 -1380
rect 117180 -1160 117490 -1150
rect 117180 -1220 117190 -1160
rect 117250 -1220 117270 -1160
rect 117330 -1220 117350 -1160
rect 117410 -1220 117490 -1160
rect 117180 -1240 117490 -1220
rect 117180 -1300 117190 -1240
rect 117250 -1300 117270 -1240
rect 117330 -1300 117350 -1240
rect 117410 -1300 117490 -1240
rect 117180 -1320 117490 -1300
rect 117180 -1380 117190 -1320
rect 117250 -1380 117270 -1320
rect 117330 -1380 117350 -1320
rect 117410 -1380 117490 -1320
rect 117180 -1390 117490 -1380
rect 117830 -1150 117890 -690
rect 118030 650 118090 810
rect 118030 -690 118040 650
rect 118080 -690 118090 650
rect 118030 -720 118090 -690
rect 118230 650 118290 670
rect 118230 -690 118240 650
rect 118280 -690 118290 650
rect 118760 660 118830 810
rect 118760 580 118830 590
rect 118880 770 118960 1090
rect 119120 1040 119620 3160
rect 119120 980 119130 1040
rect 119190 980 119210 1040
rect 119270 980 119300 1040
rect 119360 980 119380 1040
rect 119440 980 119470 1040
rect 119530 980 119550 1040
rect 119610 980 119620 1040
rect 119120 960 119620 980
rect 119120 900 119130 960
rect 119190 900 119210 960
rect 119270 900 119300 960
rect 119360 900 119380 960
rect 119440 900 119470 960
rect 119530 900 119550 960
rect 119610 900 119620 960
rect 119120 880 119620 900
rect 119120 820 119130 880
rect 119190 820 119210 880
rect 119270 820 119300 880
rect 119360 820 119380 880
rect 119440 820 119470 880
rect 119530 820 119550 880
rect 119610 820 119620 880
rect 119120 810 119620 820
rect 119680 4100 119920 4110
rect 119680 4040 119690 4100
rect 119750 4040 119770 4100
rect 119830 4040 119850 4100
rect 119910 4040 119920 4100
rect 119680 4020 119920 4040
rect 119680 3960 119690 4020
rect 119750 3960 119770 4020
rect 119830 3960 119850 4020
rect 119910 3960 119920 4020
rect 119680 3940 119920 3960
rect 119680 3880 119690 3940
rect 119750 3880 119770 3940
rect 119830 3880 119850 3940
rect 119910 3880 119920 3940
rect 119680 1880 119920 3880
rect 119680 1820 119690 1880
rect 119750 1820 119770 1880
rect 119830 1820 119850 1880
rect 119910 1820 119920 1880
rect 119680 1800 119920 1820
rect 119680 1740 119690 1800
rect 119750 1740 119770 1800
rect 119830 1740 119850 1800
rect 119910 1740 119920 1800
rect 119680 1720 119920 1740
rect 119680 1660 119690 1720
rect 119750 1660 119770 1720
rect 119830 1660 119850 1720
rect 119910 1660 119920 1720
rect 118880 710 118890 770
rect 118950 710 118960 770
rect 118880 670 118960 710
rect 118880 660 118950 670
rect 118880 580 118950 590
rect 118020 -730 118100 -720
rect 118020 -790 118030 -730
rect 118090 -790 118100 -730
rect 118020 -800 118100 -790
rect 118230 -770 118290 -690
rect 118230 -810 118240 -770
rect 118280 -810 118290 -770
rect 118230 -1150 118290 -810
rect 117830 -1160 118120 -1150
rect 117830 -1220 117890 -1160
rect 117950 -1220 117970 -1160
rect 118030 -1220 118050 -1160
rect 118110 -1220 118120 -1160
rect 117830 -1240 118120 -1220
rect 117830 -1300 117890 -1240
rect 117950 -1300 117970 -1240
rect 118030 -1300 118050 -1240
rect 118110 -1300 118120 -1240
rect 117830 -1320 118120 -1300
rect 117830 -1380 117890 -1320
rect 117950 -1380 117970 -1320
rect 118030 -1380 118050 -1320
rect 118110 -1380 118120 -1320
rect 117830 -1390 118120 -1380
rect 118220 -1160 118300 -1150
rect 118220 -1220 118230 -1160
rect 118290 -1220 118300 -1160
rect 118220 -1240 118300 -1220
rect 118220 -1300 118230 -1240
rect 118290 -1300 118300 -1240
rect 118220 -1320 118300 -1300
rect 118220 -1380 118230 -1320
rect 118290 -1380 118300 -1320
rect 118220 -1390 118300 -1380
rect 118740 -1160 118980 -1150
rect 118740 -1220 118750 -1160
rect 118810 -1220 118830 -1160
rect 118890 -1220 118910 -1160
rect 118970 -1220 118980 -1160
rect 118740 -1240 118980 -1220
rect 118740 -1300 118750 -1240
rect 118810 -1300 118830 -1240
rect 118890 -1300 118910 -1240
rect 118970 -1300 118980 -1240
rect 118740 -1320 118980 -1300
rect 118740 -1380 118750 -1320
rect 118810 -1380 118830 -1320
rect 118890 -1380 118910 -1320
rect 118970 -1380 118980 -1320
rect 118740 -1390 118980 -1380
rect 119280 -1160 119520 -1150
rect 119280 -1220 119290 -1160
rect 119350 -1220 119370 -1160
rect 119430 -1220 119450 -1160
rect 119510 -1220 119520 -1160
rect 119280 -1240 119520 -1220
rect 119280 -1300 119290 -1240
rect 119350 -1300 119370 -1240
rect 119430 -1300 119450 -1240
rect 119510 -1300 119520 -1240
rect 119280 -1320 119520 -1300
rect 119280 -1380 119290 -1320
rect 119350 -1380 119370 -1320
rect 119430 -1380 119450 -1320
rect 119510 -1380 119520 -1320
rect 117180 -3000 117420 -1390
rect 117880 -3000 118120 -1390
rect 118580 -3000 118820 -1390
rect 119280 -3000 119520 -1380
rect 119680 -1160 119920 1660
rect 119680 -1220 119690 -1160
rect 119750 -1220 119770 -1160
rect 119830 -1220 119850 -1160
rect 119910 -1220 119920 -1160
rect 119680 -1240 119920 -1220
rect 119680 -1300 119690 -1240
rect 119750 -1300 119770 -1240
rect 119830 -1300 119850 -1240
rect 119910 -1300 119920 -1240
rect 119680 -1320 119920 -1300
rect 119680 -1380 119690 -1320
rect 119750 -1380 119770 -1320
rect 119830 -1380 119850 -1320
rect 119910 -1380 119920 -1320
rect 119680 -1390 119920 -1380
rect 119980 -1160 120220 -1150
rect 119980 -1220 119990 -1160
rect 120050 -1220 120070 -1160
rect 120130 -1220 120150 -1160
rect 120210 -1220 120220 -1160
rect 119980 -1240 120220 -1220
rect 119980 -1300 119990 -1240
rect 120050 -1300 120070 -1240
rect 120130 -1300 120150 -1240
rect 120210 -1300 120220 -1240
rect 119980 -1320 120220 -1300
rect 119980 -1380 119990 -1320
rect 120050 -1380 120070 -1320
rect 120130 -1380 120150 -1320
rect 120210 -1380 120220 -1320
rect 119980 -3000 120220 -1380
rect 120680 -1160 120920 -1150
rect 120680 -1220 120690 -1160
rect 120750 -1220 120770 -1160
rect 120830 -1220 120850 -1160
rect 120910 -1220 120920 -1160
rect 120680 -1240 120920 -1220
rect 120680 -1300 120690 -1240
rect 120750 -1300 120770 -1240
rect 120830 -1300 120850 -1240
rect 120910 -1300 120920 -1240
rect 120680 -1320 120920 -1300
rect 120680 -1380 120690 -1320
rect 120750 -1380 120770 -1320
rect 120830 -1380 120850 -1320
rect 120910 -1380 120920 -1320
rect 120680 -3000 120920 -1380
rect 121380 -1160 121620 -1150
rect 121380 -1220 121390 -1160
rect 121450 -1220 121470 -1160
rect 121530 -1220 121550 -1160
rect 121610 -1220 121620 -1160
rect 121380 -1240 121620 -1220
rect 121380 -1300 121390 -1240
rect 121450 -1300 121470 -1240
rect 121530 -1300 121550 -1240
rect 121610 -1300 121620 -1240
rect 121380 -1320 121620 -1300
rect 121380 -1380 121390 -1320
rect 121450 -1380 121470 -1320
rect 121530 -1380 121550 -1320
rect 121610 -1380 121620 -1320
rect 121380 -3000 121620 -1380
rect 122080 -1160 122320 -1150
rect 122080 -1220 122090 -1160
rect 122150 -1220 122170 -1160
rect 122230 -1220 122250 -1160
rect 122310 -1220 122320 -1160
rect 122080 -1240 122320 -1220
rect 122080 -1300 122090 -1240
rect 122150 -1300 122170 -1240
rect 122230 -1300 122250 -1240
rect 122310 -1300 122320 -1240
rect 122080 -1320 122320 -1300
rect 122080 -1380 122090 -1320
rect 122150 -1380 122170 -1320
rect 122230 -1380 122250 -1320
rect 122310 -1380 122320 -1320
rect 122080 -3000 122320 -1380
rect 122780 -1160 123020 -1150
rect 122780 -1220 122790 -1160
rect 122850 -1220 122870 -1160
rect 122930 -1220 122950 -1160
rect 123010 -1220 123020 -1160
rect 122780 -1240 123020 -1220
rect 122780 -1300 122790 -1240
rect 122850 -1300 122870 -1240
rect 122930 -1300 122950 -1240
rect 123010 -1300 123020 -1240
rect 122780 -1320 123020 -1300
rect 122780 -1380 122790 -1320
rect 122850 -1380 122870 -1320
rect 122930 -1380 122950 -1320
rect 123010 -1380 123020 -1320
rect 122780 -3000 123020 -1380
<< via1 >>
rect 104590 8580 104650 8640
rect 104670 8580 104730 8640
rect 104750 8580 104810 8640
rect 104590 8500 104650 8560
rect 104670 8500 104730 8560
rect 104750 8500 104810 8560
rect 104590 8420 104650 8480
rect 104670 8420 104730 8480
rect 104750 8420 104810 8480
rect 105290 8580 105350 8640
rect 105370 8580 105430 8640
rect 105450 8580 105510 8640
rect 105290 8500 105350 8560
rect 105370 8500 105430 8560
rect 105450 8500 105510 8560
rect 105290 8420 105350 8480
rect 105370 8420 105430 8480
rect 105450 8420 105510 8480
rect 105990 8580 106050 8640
rect 106070 8580 106130 8640
rect 106150 8580 106210 8640
rect 105990 8500 106050 8560
rect 106070 8500 106130 8560
rect 106150 8500 106210 8560
rect 105990 8420 106050 8480
rect 106070 8420 106130 8480
rect 106150 8420 106210 8480
rect 106690 8580 106750 8640
rect 106770 8580 106830 8640
rect 106850 8580 106910 8640
rect 106690 8500 106750 8560
rect 106770 8500 106830 8560
rect 106850 8500 106910 8560
rect 106690 8420 106750 8480
rect 106770 8420 106830 8480
rect 106850 8420 106910 8480
rect 112420 10070 112480 10130
rect 112180 9850 112240 9860
rect 112180 9810 112190 9850
rect 112190 9810 112230 9850
rect 112230 9810 112240 9850
rect 112180 9800 112240 9810
rect 113360 10070 113420 10130
rect 114180 10070 114240 10130
rect 115120 10070 115180 10130
rect 112420 9800 112480 9860
rect 112540 9850 112600 9860
rect 112540 9810 112550 9850
rect 112550 9810 112590 9850
rect 112590 9810 112600 9850
rect 112540 9800 112600 9810
rect 113120 9620 113180 9680
rect 113120 9540 113180 9600
rect 113120 9510 113180 9520
rect 113120 9470 113130 9510
rect 113130 9470 113170 9510
rect 113170 9470 113180 9510
rect 113120 9460 113180 9470
rect 113240 9620 113300 9680
rect 113240 9540 113300 9600
rect 113240 9460 113300 9520
rect 113770 9960 113830 10020
rect 113770 9880 113830 9940
rect 113770 9800 113830 9860
rect 113480 9620 113540 9680
rect 113480 9540 113540 9600
rect 113480 9510 113540 9520
rect 113480 9470 113490 9510
rect 113490 9470 113530 9510
rect 113530 9470 113540 9510
rect 113480 9460 113540 9470
rect 114060 9960 114120 10020
rect 114060 9880 114120 9940
rect 114060 9850 114120 9860
rect 114060 9810 114070 9850
rect 114070 9810 114110 9850
rect 114110 9810 114120 9850
rect 114060 9800 114120 9810
rect 113770 9620 113830 9680
rect 113770 9540 113830 9600
rect 113770 9460 113830 9520
rect 112420 8990 112480 9050
rect 113360 8990 113420 9050
rect 112310 8950 112370 8960
rect 112310 8910 112320 8950
rect 112320 8910 112360 8950
rect 112360 8910 112370 8950
rect 112310 8900 112370 8910
rect 113260 8950 113320 8960
rect 113260 8910 113270 8950
rect 113270 8910 113310 8950
rect 113310 8910 113320 8950
rect 113260 8900 113320 8910
rect 113660 8900 113720 8960
rect 108090 8580 108150 8640
rect 108170 8580 108230 8640
rect 108250 8580 108310 8640
rect 108090 8500 108150 8560
rect 108170 8500 108230 8560
rect 108250 8500 108310 8560
rect 108090 8420 108150 8480
rect 108170 8420 108230 8480
rect 108250 8420 108310 8480
rect 109190 8580 109250 8640
rect 109190 8500 109250 8560
rect 109190 8420 109250 8480
rect 109910 8580 109970 8640
rect 109910 8500 109970 8560
rect 109910 8420 109970 8480
rect 109310 8310 109370 8370
rect 109310 8230 109370 8290
rect 109310 8150 109370 8210
rect 109310 8070 109370 8130
rect 109310 7990 109370 8050
rect 109310 7910 109370 7970
rect 109550 8310 109610 8370
rect 109550 8230 109610 8290
rect 109550 8150 109610 8210
rect 109550 8070 109610 8130
rect 109550 7990 109610 8050
rect 109550 7910 109610 7970
rect 109790 8310 109850 8370
rect 109790 8230 109850 8290
rect 109790 8150 109850 8210
rect 109790 8070 109850 8130
rect 109790 7990 109850 8050
rect 109790 7910 109850 7970
rect 109190 7800 109250 7860
rect 109430 7800 109490 7860
rect 109670 7800 109730 7860
rect 110630 8580 110690 8640
rect 110630 8500 110690 8560
rect 110630 8420 110690 8480
rect 110030 8310 110090 8370
rect 110030 8230 110090 8290
rect 110030 8150 110090 8210
rect 110030 8070 110090 8130
rect 110030 7990 110090 8050
rect 110030 7910 110090 7970
rect 110270 8310 110330 8370
rect 110270 8230 110330 8290
rect 110270 8150 110330 8210
rect 110270 8070 110330 8130
rect 110270 7990 110330 8050
rect 110270 7910 110330 7970
rect 110510 8310 110570 8370
rect 110510 8230 110570 8290
rect 110510 8150 110570 8210
rect 110510 8070 110570 8130
rect 110510 7990 110570 8050
rect 110510 7910 110570 7970
rect 109910 7800 109970 7860
rect 110150 7800 110210 7860
rect 110390 7800 110450 7860
rect 110630 7800 110690 7860
rect 111080 8580 111140 8640
rect 111160 8580 111220 8640
rect 111240 8580 111300 8640
rect 111080 8500 111140 8560
rect 111160 8500 111220 8560
rect 111240 8500 111300 8560
rect 111080 8420 111140 8480
rect 111160 8420 111220 8480
rect 111240 8420 111300 8480
rect 109310 6990 109370 7050
rect 109550 6990 109610 7050
rect 109790 6990 109850 7050
rect 110030 6990 110090 7050
rect 110270 6990 110330 7050
rect 110510 6990 110570 7050
rect 110810 6990 110870 7050
rect 110890 6990 110950 7050
rect 110970 6990 111030 7050
rect 109370 6930 109430 6940
rect 109370 6890 109380 6930
rect 109380 6890 109420 6930
rect 109420 6890 109430 6930
rect 109370 6880 109430 6890
rect 109490 6930 109550 6940
rect 109490 6890 109500 6930
rect 109500 6890 109540 6930
rect 109540 6890 109550 6930
rect 109490 6880 109550 6890
rect 109610 6930 109670 6940
rect 109610 6890 109620 6930
rect 109620 6890 109660 6930
rect 109660 6890 109670 6930
rect 109610 6880 109670 6890
rect 109730 6930 109790 6940
rect 109730 6890 109740 6930
rect 109740 6890 109780 6930
rect 109780 6890 109790 6930
rect 109730 6880 109790 6890
rect 109850 6930 109910 6940
rect 109850 6890 109860 6930
rect 109860 6890 109900 6930
rect 109900 6890 109910 6930
rect 109850 6880 109910 6890
rect 109970 6930 110030 6940
rect 109970 6890 109980 6930
rect 109980 6890 110020 6930
rect 110020 6890 110030 6930
rect 109970 6880 110030 6890
rect 110090 6930 110150 6940
rect 110090 6890 110100 6930
rect 110100 6890 110140 6930
rect 110140 6890 110150 6930
rect 110090 6880 110150 6890
rect 110210 6930 110270 6940
rect 110210 6890 110220 6930
rect 110220 6890 110260 6930
rect 110260 6890 110270 6930
rect 110210 6880 110270 6890
rect 110330 6930 110390 6940
rect 110330 6890 110340 6930
rect 110340 6890 110380 6930
rect 110380 6890 110390 6930
rect 110330 6880 110390 6890
rect 110450 6930 110510 6940
rect 110450 6890 110460 6930
rect 110460 6890 110500 6930
rect 110500 6890 110510 6930
rect 110450 6880 110510 6890
rect 109910 6760 109970 6820
rect 108520 6690 108580 6750
rect 109250 6650 109310 6710
rect 109250 6570 109310 6630
rect 109250 6490 109310 6550
rect 109470 6650 109530 6710
rect 109470 6570 109530 6630
rect 109470 6490 109530 6550
rect 109690 6650 109750 6710
rect 109690 6570 109750 6630
rect 109690 6490 109750 6550
rect 109910 6650 109970 6710
rect 109910 6570 109970 6630
rect 109910 6490 109970 6550
rect 110130 6650 110190 6710
rect 110130 6570 110190 6630
rect 110130 6490 110190 6550
rect 110350 6650 110410 6710
rect 110350 6570 110410 6630
rect 110350 6490 110410 6550
rect 110570 6650 110630 6710
rect 110570 6570 110630 6630
rect 110570 6490 110630 6550
rect 109360 6320 109420 6380
rect 109580 6320 109640 6380
rect 109800 6320 109860 6380
rect 110020 6320 110080 6380
rect 110240 6320 110300 6380
rect 110460 6320 110520 6380
rect 108440 4880 108500 4940
rect 108520 4880 108580 4940
rect 108600 4880 108660 4940
rect 108440 4800 108500 4860
rect 108520 4800 108580 4860
rect 108600 4800 108660 4860
rect 108440 4720 108500 4780
rect 108520 4720 108580 4780
rect 108600 4720 108660 4780
rect 109360 5040 109420 5100
rect 109580 5040 109640 5100
rect 109800 5040 109860 5100
rect 110020 5040 110080 5100
rect 109910 4930 109970 4940
rect 109910 4890 109920 4930
rect 109920 4890 109960 4930
rect 109960 4890 109970 4930
rect 109910 4880 109970 4890
rect 109910 4850 109970 4860
rect 109910 4810 109920 4850
rect 109920 4810 109960 4850
rect 109960 4810 109970 4850
rect 109910 4800 109970 4810
rect 109910 4770 109970 4780
rect 109910 4730 109920 4770
rect 109920 4730 109960 4770
rect 109960 4730 109970 4770
rect 109910 4720 109970 4730
rect 110240 5040 110300 5100
rect 110460 5040 110520 5100
rect 107990 4580 108050 4640
rect 108070 4580 108130 4640
rect 108160 4580 108220 4640
rect 108240 4580 108300 4640
rect 108330 4580 108390 4640
rect 108410 4580 108470 4640
rect 107990 4500 108050 4560
rect 108070 4500 108130 4560
rect 108160 4500 108220 4560
rect 108240 4500 108300 4560
rect 108330 4500 108390 4560
rect 108410 4500 108470 4560
rect 107990 4420 108050 4480
rect 108070 4420 108130 4480
rect 108160 4420 108220 4480
rect 108240 4420 108300 4480
rect 108330 4420 108390 4480
rect 108410 4420 108470 4480
rect 107690 4040 107750 4100
rect 107770 4040 107830 4100
rect 107850 4040 107910 4100
rect 107690 3960 107750 4020
rect 107770 3960 107830 4020
rect 107850 3960 107910 4020
rect 107690 3880 107750 3940
rect 107770 3880 107830 3940
rect 107850 3880 107910 3940
rect 107690 1820 107750 1880
rect 107770 1820 107830 1880
rect 107850 1820 107910 1880
rect 107690 1740 107750 1800
rect 107770 1740 107830 1800
rect 107850 1740 107910 1800
rect 107690 1660 107750 1720
rect 107770 1660 107830 1720
rect 107850 1660 107910 1720
rect 104590 -1220 104650 -1160
rect 104670 -1220 104730 -1160
rect 104750 -1220 104810 -1160
rect 104590 -1300 104650 -1240
rect 104670 -1300 104730 -1240
rect 104750 -1300 104810 -1240
rect 104590 -1380 104650 -1320
rect 104670 -1380 104730 -1320
rect 104750 -1380 104810 -1320
rect 105290 -1220 105350 -1160
rect 105370 -1220 105430 -1160
rect 105450 -1220 105510 -1160
rect 105290 -1300 105350 -1240
rect 105370 -1300 105430 -1240
rect 105450 -1300 105510 -1240
rect 105290 -1380 105350 -1320
rect 105370 -1380 105430 -1320
rect 105450 -1380 105510 -1320
rect 105990 -1220 106050 -1160
rect 106070 -1220 106130 -1160
rect 106150 -1220 106210 -1160
rect 105990 -1300 106050 -1240
rect 106070 -1300 106130 -1240
rect 106150 -1300 106210 -1240
rect 105990 -1380 106050 -1320
rect 106070 -1380 106130 -1320
rect 106150 -1380 106210 -1320
rect 106690 -1220 106750 -1160
rect 106770 -1220 106830 -1160
rect 106850 -1220 106910 -1160
rect 106690 -1300 106750 -1240
rect 106770 -1300 106830 -1240
rect 106850 -1300 106910 -1240
rect 106690 -1380 106750 -1320
rect 106770 -1380 106830 -1320
rect 106850 -1380 106910 -1320
rect 107390 -1220 107450 -1160
rect 107470 -1220 107530 -1160
rect 107550 -1220 107610 -1160
rect 107390 -1300 107450 -1240
rect 107470 -1300 107530 -1240
rect 107550 -1300 107610 -1240
rect 107390 -1380 107450 -1320
rect 107470 -1380 107530 -1320
rect 107550 -1380 107610 -1320
rect 109360 4580 109420 4640
rect 109470 4580 109530 4640
rect 109580 4580 109640 4640
rect 109690 4580 109750 4640
rect 109800 4580 109860 4640
rect 109910 4580 109970 4640
rect 110020 4580 110080 4640
rect 110130 4580 110190 4640
rect 110240 4580 110300 4640
rect 110350 4580 110410 4640
rect 110460 4580 110520 4640
rect 109360 4500 109420 4560
rect 109470 4500 109530 4560
rect 109580 4500 109640 4560
rect 109690 4500 109750 4560
rect 109800 4500 109860 4560
rect 109910 4500 109970 4560
rect 110020 4500 110080 4560
rect 110130 4500 110190 4560
rect 110240 4500 110300 4560
rect 110350 4500 110410 4560
rect 110460 4500 110520 4560
rect 109360 4420 109420 4480
rect 109470 4420 109530 4480
rect 109580 4420 109640 4480
rect 109690 4420 109750 4480
rect 109800 4420 109860 4480
rect 109910 4420 109970 4480
rect 110020 4420 110080 4480
rect 110130 4420 110190 4480
rect 110240 4420 110300 4480
rect 110350 4420 110410 4480
rect 110460 4420 110520 4480
rect 110810 4880 110870 4940
rect 110890 4880 110950 4940
rect 110970 4880 111030 4940
rect 110810 4800 110870 4860
rect 110890 4800 110950 4860
rect 110970 4800 111030 4860
rect 110810 4720 110870 4780
rect 110890 4720 110950 4780
rect 110970 4720 111030 4780
rect 109250 4310 109310 4370
rect 109250 4230 109310 4290
rect 109250 4150 109310 4210
rect 110570 4310 110630 4370
rect 110570 4230 110630 4290
rect 110570 4150 110630 4210
rect 108000 3360 108060 3420
rect 108100 3360 108160 3420
rect 108200 3360 108260 3420
rect 108300 3360 108360 3420
rect 108400 3360 108460 3420
rect 109360 4040 109420 4100
rect 109360 3960 109420 4020
rect 109360 3880 109420 3940
rect 109580 4040 109640 4100
rect 109580 3960 109640 4020
rect 109580 3880 109640 3940
rect 109800 4040 109860 4100
rect 109800 3960 109860 4020
rect 109800 3880 109860 3940
rect 110020 4040 110080 4100
rect 110020 3960 110080 4020
rect 110020 3880 110080 3940
rect 110240 4040 110300 4100
rect 110240 3960 110300 4020
rect 110240 3880 110300 3940
rect 110460 4040 110520 4100
rect 110460 3960 110520 4020
rect 110460 3880 110520 3940
rect 109470 3770 109530 3830
rect 109690 3770 109750 3830
rect 109910 3770 109970 3830
rect 110130 3770 110190 3830
rect 110350 3770 110410 3830
rect 108000 3260 108060 3320
rect 108100 3260 108160 3320
rect 108200 3260 108260 3320
rect 108300 3260 108360 3320
rect 108400 3260 108460 3320
rect 108980 3260 109040 3320
rect 109470 3310 109530 3320
rect 109470 3270 109480 3310
rect 109480 3270 109520 3310
rect 109520 3270 109530 3310
rect 109470 3260 109530 3270
rect 109690 3310 109750 3320
rect 109690 3270 109700 3310
rect 109700 3270 109740 3310
rect 109740 3270 109750 3310
rect 109690 3260 109750 3270
rect 109910 3310 109970 3320
rect 109910 3270 109920 3310
rect 109920 3270 109960 3310
rect 109960 3270 109970 3310
rect 109910 3260 109970 3270
rect 110130 3310 110190 3320
rect 110130 3270 110140 3310
rect 110140 3270 110180 3310
rect 110180 3270 110190 3310
rect 110130 3260 110190 3270
rect 110350 3310 110410 3320
rect 110350 3270 110360 3310
rect 110360 3270 110400 3310
rect 110400 3270 110410 3310
rect 110350 3260 110410 3270
rect 108000 3160 108060 3220
rect 108100 3160 108160 3220
rect 108200 3160 108260 3220
rect 108300 3160 108360 3220
rect 108400 3160 108460 3220
rect 108510 2310 108580 2320
rect 108510 2260 108520 2310
rect 108520 2260 108570 2310
rect 108570 2260 108580 2310
rect 108510 2250 108580 2260
rect 108630 2310 108700 2320
rect 108630 2260 108640 2310
rect 108640 2260 108690 2310
rect 108690 2260 108700 2310
rect 108630 2250 108700 2260
rect 108750 2310 108820 2320
rect 108750 2260 108760 2310
rect 108760 2260 108810 2310
rect 108810 2260 108820 2310
rect 108750 2250 108820 2260
rect 108870 2310 108940 2320
rect 108870 2260 108880 2310
rect 108880 2260 108930 2310
rect 108930 2260 108940 2310
rect 108870 2250 108940 2260
rect 110240 3180 110300 3190
rect 110240 3140 110250 3180
rect 110250 3140 110290 3180
rect 110290 3140 110300 3180
rect 110240 3130 110300 3140
rect 110240 3100 110300 3110
rect 110240 3060 110250 3100
rect 110250 3060 110290 3100
rect 110290 3060 110300 3100
rect 110240 3050 110300 3060
rect 110810 3130 110870 3190
rect 110890 3130 110950 3190
rect 110970 3130 111030 3190
rect 110810 3050 110870 3110
rect 110890 3050 110950 3110
rect 110970 3050 111030 3110
rect 112020 8310 112080 8370
rect 112020 8230 112080 8290
rect 112020 8150 112080 8210
rect 112020 8070 112080 8130
rect 112020 7990 112080 8050
rect 112020 7910 112080 7970
rect 112260 8310 112320 8370
rect 112260 8230 112320 8290
rect 112260 8150 112320 8210
rect 112260 8070 112320 8130
rect 112260 7990 112320 8050
rect 112260 7910 112320 7970
rect 112500 8310 112560 8370
rect 112500 8230 112560 8290
rect 112500 8150 112560 8210
rect 112500 8070 112560 8130
rect 112500 7990 112560 8050
rect 112500 7910 112560 7970
rect 112740 8310 112800 8370
rect 112740 8230 112800 8290
rect 112740 8150 112800 8210
rect 112740 8070 112800 8130
rect 112740 7990 112800 8050
rect 112740 7910 112800 7970
rect 112980 8310 113040 8370
rect 112980 8230 113040 8290
rect 112980 8150 113040 8210
rect 112980 8070 113040 8130
rect 112980 7990 113040 8050
rect 112980 7910 113040 7970
rect 113220 8310 113280 8370
rect 113220 8230 113280 8290
rect 113220 8150 113280 8210
rect 113220 8070 113280 8130
rect 113220 7990 113280 8050
rect 113220 7910 113280 7970
rect 113460 8310 113520 8370
rect 113460 8230 113520 8290
rect 113460 8150 113520 8210
rect 113460 8070 113520 8130
rect 113460 7990 113520 8050
rect 113460 7910 113520 7970
rect 112140 7770 112200 7830
rect 112380 7770 112440 7830
rect 112620 7770 112680 7830
rect 112860 7770 112920 7830
rect 113100 7770 113160 7830
rect 113340 7770 113400 7830
rect 112140 6990 112200 7050
rect 112380 6990 112440 7050
rect 112620 6990 112680 7050
rect 112860 6990 112920 7050
rect 113100 6990 113160 7050
rect 113340 6990 113400 7050
rect 114300 9960 114360 10020
rect 114300 9880 114360 9940
rect 114300 9800 114360 9860
rect 114420 9960 114480 10020
rect 114420 9880 114480 9940
rect 114420 9850 114480 9860
rect 114420 9810 114430 9850
rect 114430 9810 114470 9850
rect 114470 9810 114480 9850
rect 114420 9800 114480 9810
rect 115000 9850 115060 9860
rect 115000 9810 115010 9850
rect 115010 9810 115050 9850
rect 115050 9810 115060 9850
rect 115000 9800 115060 9810
rect 115120 9800 115180 9860
rect 115360 9850 115420 9860
rect 115360 9810 115370 9850
rect 115370 9810 115410 9850
rect 115410 9810 115420 9850
rect 115360 9800 115420 9810
rect 114180 8990 114240 9050
rect 115120 8990 115180 9050
rect 113770 8580 113830 8640
rect 113770 8500 113830 8560
rect 113770 8420 113830 8480
rect 113880 8790 113940 8850
rect 115152 8930 115212 8940
rect 115152 8890 115162 8930
rect 115162 8890 115202 8930
rect 115202 8890 115212 8930
rect 115152 8880 115212 8890
rect 112200 6930 112260 6940
rect 112200 6890 112210 6930
rect 112210 6890 112250 6930
rect 112250 6890 112260 6930
rect 112200 6880 112260 6890
rect 112320 6930 112380 6940
rect 112320 6890 112330 6930
rect 112330 6890 112370 6930
rect 112370 6890 112380 6930
rect 112320 6880 112380 6890
rect 112440 6930 112500 6940
rect 112440 6890 112450 6930
rect 112450 6890 112490 6930
rect 112490 6890 112500 6930
rect 112440 6880 112500 6890
rect 112560 6930 112620 6940
rect 112560 6890 112570 6930
rect 112570 6890 112610 6930
rect 112610 6890 112620 6930
rect 112560 6880 112620 6890
rect 112680 6930 112740 6940
rect 112680 6890 112690 6930
rect 112690 6890 112730 6930
rect 112730 6890 112740 6930
rect 112680 6880 112740 6890
rect 112800 6930 112860 6940
rect 112800 6890 112810 6930
rect 112810 6890 112850 6930
rect 112850 6890 112860 6930
rect 112800 6880 112860 6890
rect 112920 6930 112980 6940
rect 112920 6890 112930 6930
rect 112930 6890 112970 6930
rect 112970 6890 112980 6930
rect 112920 6880 112980 6890
rect 113040 6930 113100 6940
rect 113040 6890 113050 6930
rect 113050 6890 113090 6930
rect 113090 6890 113100 6930
rect 113040 6880 113100 6890
rect 113160 6930 113220 6940
rect 113160 6890 113170 6930
rect 113170 6890 113210 6930
rect 113210 6890 113220 6930
rect 113160 6880 113220 6890
rect 113280 6930 113340 6940
rect 113280 6890 113290 6930
rect 113290 6890 113330 6930
rect 113330 6890 113340 6930
rect 113280 6880 113340 6890
rect 113680 6880 113740 6940
rect 114280 8770 114340 8830
rect 115240 8770 115300 8830
rect 116300 8580 116360 8640
rect 116380 8580 116440 8640
rect 116460 8580 116520 8640
rect 116300 8500 116360 8560
rect 116380 8500 116440 8560
rect 116460 8500 116520 8560
rect 116300 8420 116360 8480
rect 116380 8420 116440 8480
rect 116460 8420 116520 8480
rect 114080 8310 114140 8370
rect 114080 8230 114140 8290
rect 114080 8150 114140 8210
rect 114080 8070 114140 8130
rect 114080 7990 114140 8050
rect 114080 7910 114140 7970
rect 114320 8310 114380 8370
rect 114320 8230 114380 8290
rect 114320 8150 114380 8210
rect 114320 8070 114380 8130
rect 114320 7990 114380 8050
rect 114320 7910 114380 7970
rect 114560 8310 114620 8370
rect 114560 8230 114620 8290
rect 114560 8150 114620 8210
rect 114560 8070 114620 8130
rect 114560 7990 114620 8050
rect 114560 7910 114620 7970
rect 114800 8310 114860 8370
rect 114800 8230 114860 8290
rect 114800 8150 114860 8210
rect 114800 8070 114860 8130
rect 114800 7990 114860 8050
rect 114800 7910 114860 7970
rect 115040 8310 115100 8370
rect 115040 8230 115100 8290
rect 115040 8150 115100 8210
rect 115040 8070 115100 8130
rect 115040 7990 115100 8050
rect 115040 7910 115100 7970
rect 115280 8310 115340 8370
rect 115280 8230 115340 8290
rect 115280 8150 115340 8210
rect 115280 8070 115340 8130
rect 115280 7990 115340 8050
rect 115280 7910 115340 7970
rect 115520 8310 115580 8370
rect 115520 8230 115580 8290
rect 115520 8150 115580 8210
rect 115520 8070 115580 8130
rect 115520 7990 115580 8050
rect 115520 7910 115580 7970
rect 114200 7770 114260 7830
rect 114440 7770 114500 7830
rect 114680 7770 114740 7830
rect 114920 7770 114980 7830
rect 115160 7770 115220 7830
rect 115400 7770 115460 7830
rect 114200 6990 114260 7050
rect 114440 6990 114500 7050
rect 114680 6990 114740 7050
rect 114920 6990 114980 7050
rect 115160 6990 115220 7050
rect 115400 6990 115460 7050
rect 114260 6930 114320 6940
rect 114260 6890 114270 6930
rect 114270 6890 114310 6930
rect 114310 6890 114320 6930
rect 114260 6880 114320 6890
rect 114380 6930 114440 6940
rect 114380 6890 114390 6930
rect 114390 6890 114430 6930
rect 114430 6890 114440 6930
rect 114380 6880 114440 6890
rect 114500 6930 114560 6940
rect 114500 6890 114510 6930
rect 114510 6890 114550 6930
rect 114550 6890 114560 6930
rect 114500 6880 114560 6890
rect 114620 6930 114680 6940
rect 114620 6890 114630 6930
rect 114630 6890 114670 6930
rect 114670 6890 114680 6930
rect 114620 6880 114680 6890
rect 114740 6930 114800 6940
rect 114740 6890 114750 6930
rect 114750 6890 114790 6930
rect 114790 6890 114800 6930
rect 114740 6880 114800 6890
rect 114860 6930 114920 6940
rect 114860 6890 114870 6930
rect 114870 6890 114910 6930
rect 114910 6890 114920 6930
rect 114860 6880 114920 6890
rect 114980 6930 115040 6940
rect 114980 6890 114990 6930
rect 114990 6890 115030 6930
rect 115030 6890 115040 6930
rect 114980 6880 115040 6890
rect 115100 6930 115160 6940
rect 115100 6890 115110 6930
rect 115110 6890 115150 6930
rect 115150 6890 115160 6930
rect 115100 6880 115160 6890
rect 115220 6930 115280 6940
rect 115220 6890 115230 6930
rect 115230 6890 115270 6930
rect 115270 6890 115280 6930
rect 115220 6880 115280 6890
rect 115340 6930 115400 6940
rect 115340 6890 115350 6930
rect 115350 6890 115390 6930
rect 115390 6890 115400 6930
rect 115340 6880 115400 6890
rect 113860 6760 113920 6820
rect 111080 6650 111140 6710
rect 111160 6650 111220 6710
rect 111240 6650 111300 6710
rect 111080 6570 111140 6630
rect 111160 6570 111220 6630
rect 111240 6570 111300 6630
rect 111080 6490 111140 6550
rect 111160 6490 111220 6550
rect 111240 6490 111300 6550
rect 113030 6650 113090 6710
rect 113030 6570 113090 6630
rect 113030 6540 113090 6550
rect 113030 6500 113040 6540
rect 113040 6500 113080 6540
rect 113080 6500 113090 6540
rect 113030 6490 113090 6500
rect 113360 6650 113420 6710
rect 113360 6570 113420 6630
rect 113360 6540 113420 6550
rect 113360 6500 113370 6540
rect 113370 6500 113410 6540
rect 113410 6500 113420 6540
rect 113360 6490 113420 6500
rect 113690 6650 113750 6710
rect 113690 6570 113750 6630
rect 113690 6540 113750 6550
rect 113690 6500 113700 6540
rect 113700 6500 113740 6540
rect 113740 6500 113750 6540
rect 113690 6490 113750 6500
rect 113850 6650 113910 6710
rect 113850 6570 113910 6630
rect 113850 6540 113910 6550
rect 113850 6500 113860 6540
rect 113860 6500 113900 6540
rect 113900 6500 113910 6540
rect 113850 6490 113910 6500
rect 114180 6650 114240 6710
rect 114180 6570 114240 6630
rect 114180 6540 114240 6550
rect 114180 6500 114190 6540
rect 114190 6500 114230 6540
rect 114230 6500 114240 6540
rect 114180 6490 114240 6500
rect 114510 6650 114570 6710
rect 114510 6570 114570 6630
rect 114510 6540 114570 6550
rect 114510 6500 114520 6540
rect 114520 6500 114560 6540
rect 114560 6500 114570 6540
rect 114510 6490 114570 6500
rect 116910 8580 116970 8640
rect 116910 8500 116970 8560
rect 116910 8420 116970 8480
rect 117630 8580 117690 8640
rect 117630 8500 117690 8560
rect 117630 8420 117690 8480
rect 117030 8310 117090 8370
rect 117030 8230 117090 8290
rect 117030 8150 117090 8210
rect 117030 8070 117090 8130
rect 117030 7990 117090 8050
rect 117030 7910 117090 7970
rect 117270 8310 117330 8370
rect 117270 8230 117330 8290
rect 117270 8150 117330 8210
rect 117270 8070 117330 8130
rect 117270 7990 117330 8050
rect 117270 7910 117330 7970
rect 117510 8310 117570 8370
rect 117510 8230 117570 8290
rect 117510 8150 117570 8210
rect 117510 8070 117570 8130
rect 117510 7990 117570 8050
rect 117510 7910 117570 7970
rect 116910 7850 116970 7860
rect 116910 7810 116920 7850
rect 116920 7810 116960 7850
rect 116960 7810 116970 7850
rect 116910 7800 116970 7810
rect 116300 6650 116360 6710
rect 116380 6650 116440 6710
rect 116460 6650 116520 6710
rect 116300 6570 116360 6630
rect 116380 6570 116440 6630
rect 116460 6570 116520 6630
rect 116300 6490 116360 6550
rect 116380 6490 116440 6550
rect 116460 6490 116520 6550
rect 113250 6430 113310 6440
rect 113250 6390 113260 6430
rect 113260 6390 113300 6430
rect 113300 6390 113310 6430
rect 113250 6380 113310 6390
rect 113470 6430 113530 6440
rect 113470 6390 113480 6430
rect 113480 6390 113520 6430
rect 113520 6390 113530 6430
rect 113470 6380 113530 6390
rect 114070 6430 114130 6440
rect 114070 6390 114080 6430
rect 114080 6390 114120 6430
rect 114120 6390 114130 6430
rect 114070 6380 114130 6390
rect 114290 6430 114350 6440
rect 114290 6390 114300 6430
rect 114300 6390 114340 6430
rect 114340 6390 114350 6430
rect 114290 6380 114350 6390
rect 113120 5810 113180 5820
rect 113600 5810 113660 5820
rect 113120 5770 113130 5810
rect 113130 5770 113170 5810
rect 113170 5770 113180 5810
rect 113120 5760 113180 5770
rect 113360 5790 113420 5800
rect 113360 5750 113370 5790
rect 113370 5750 113410 5790
rect 113410 5750 113420 5790
rect 113360 5740 113420 5750
rect 113600 5770 113610 5810
rect 113610 5770 113650 5810
rect 113650 5770 113660 5810
rect 113600 5760 113660 5770
rect 113210 5650 113270 5660
rect 113210 5610 113220 5650
rect 113220 5610 113260 5650
rect 113260 5610 113270 5650
rect 113210 5600 113270 5610
rect 111910 5500 111970 5560
rect 113500 5500 113560 5560
rect 111080 4310 111140 4370
rect 111160 4310 111220 4370
rect 111240 4310 111300 4370
rect 111080 4230 111140 4290
rect 111160 4230 111220 4290
rect 111240 4230 111300 4290
rect 111080 4150 111140 4210
rect 111160 4150 111220 4210
rect 111240 4150 111300 4210
rect 109070 2890 109130 2950
rect 109470 2890 109530 2950
rect 109690 2890 109750 2950
rect 109910 2890 109970 2950
rect 110130 2890 110190 2950
rect 110350 2890 110410 2950
rect 109070 2250 109130 2310
rect 108760 2110 108820 2170
rect 108980 2110 109040 2170
rect 109470 2210 109530 2270
rect 109690 2210 109750 2270
rect 109910 2210 109970 2270
rect 110130 2210 110190 2270
rect 110350 2210 110410 2270
rect 109360 2090 109420 2150
rect 109360 2010 109420 2070
rect 109360 1930 109420 1990
rect 109580 2090 109640 2150
rect 109580 2010 109640 2070
rect 109580 1930 109640 1990
rect 109800 2090 109860 2150
rect 109800 2010 109860 2070
rect 109800 1930 109860 1990
rect 110020 2090 110080 2150
rect 110020 2010 110080 2070
rect 110020 1930 110080 1990
rect 110240 2090 110300 2150
rect 110240 2010 110300 2070
rect 110240 1930 110300 1990
rect 110460 2090 110520 2150
rect 110460 2010 110520 2070
rect 110460 1930 110520 1990
rect 111350 4530 111410 4590
rect 111430 4530 111490 4590
rect 111510 4530 111570 4590
rect 111350 4450 111410 4510
rect 111430 4450 111490 4510
rect 111510 4450 111570 4510
rect 111350 4370 111410 4430
rect 111430 4370 111490 4430
rect 111510 4370 111570 4430
rect 111350 4040 111410 4100
rect 111430 4040 111490 4100
rect 111510 4040 111570 4100
rect 111350 3960 111410 4020
rect 111430 3960 111490 4020
rect 111510 3960 111570 4020
rect 111350 3880 111410 3940
rect 111430 3880 111490 3940
rect 111510 3880 111570 3940
rect 111350 3220 111410 3280
rect 111430 3220 111490 3280
rect 111510 3220 111570 3280
rect 111350 3140 111410 3200
rect 111430 3140 111490 3200
rect 111510 3140 111570 3200
rect 111350 3060 111410 3120
rect 111430 3060 111490 3120
rect 111510 3060 111570 3120
rect 111700 3850 111760 3910
rect 111780 3850 111840 3910
rect 111080 2090 111140 2150
rect 111160 2090 111220 2150
rect 111240 2090 111300 2150
rect 111080 2010 111140 2070
rect 111160 2010 111220 2070
rect 111240 2010 111300 2070
rect 111080 1930 111140 1990
rect 111160 1930 111220 1990
rect 111240 1930 111300 1990
rect 111350 2910 111410 2970
rect 111430 2910 111490 2970
rect 111510 2910 111570 2970
rect 111350 2830 111410 2890
rect 111430 2830 111490 2890
rect 111510 2830 111570 2890
rect 111350 2750 111410 2810
rect 111430 2750 111490 2810
rect 111510 2750 111570 2810
rect 109250 1820 109310 1880
rect 109250 1740 109310 1800
rect 109250 1660 109310 1720
rect 110570 1820 110630 1880
rect 110570 1740 110630 1800
rect 110570 1660 110630 1720
rect 108520 1550 108580 1610
rect 107990 980 108050 1040
rect 108070 980 108130 1040
rect 108160 980 108220 1040
rect 108240 980 108300 1040
rect 108330 980 108390 1040
rect 108410 980 108470 1040
rect 107990 900 108050 960
rect 108070 900 108130 960
rect 108160 900 108220 960
rect 108240 900 108300 960
rect 108330 900 108390 960
rect 108410 900 108470 960
rect 107990 820 108050 880
rect 108070 820 108130 880
rect 108160 820 108220 880
rect 108240 820 108300 880
rect 108330 820 108390 880
rect 108410 820 108470 880
rect 108650 1090 108710 1150
rect 108650 710 108710 770
rect 108650 650 108720 660
rect 108650 600 108660 650
rect 108660 600 108710 650
rect 108710 600 108720 650
rect 108650 590 108720 600
rect 108780 980 108840 1040
rect 108780 900 108840 960
rect 108780 820 108840 880
rect 109510 980 109570 1040
rect 109590 980 109650 1040
rect 109670 980 109730 1040
rect 109750 980 109810 1040
rect 109830 980 109890 1040
rect 109910 980 109970 1040
rect 109990 980 110050 1040
rect 110070 980 110130 1040
rect 110150 980 110210 1040
rect 110230 980 110290 1040
rect 110310 980 110370 1040
rect 109510 900 109570 960
rect 109590 900 109650 960
rect 109670 900 109730 960
rect 109750 900 109810 960
rect 109830 900 109890 960
rect 109910 900 109970 960
rect 109990 900 110050 960
rect 110070 900 110130 960
rect 110150 900 110210 960
rect 110230 900 110290 960
rect 110310 900 110370 960
rect 109510 820 109570 880
rect 109590 820 109650 880
rect 109670 820 109730 880
rect 109750 820 109810 880
rect 109830 820 109890 880
rect 109910 820 109970 880
rect 109990 820 110050 880
rect 110070 820 110130 880
rect 110150 820 110210 880
rect 110230 820 110290 880
rect 110310 820 110370 880
rect 108770 650 108840 660
rect 108770 600 108780 650
rect 108780 600 108830 650
rect 108830 600 108840 650
rect 108770 590 108840 600
rect 109610 760 109670 770
rect 109610 720 109620 760
rect 109620 720 109660 760
rect 109660 720 109670 760
rect 109610 710 109670 720
rect 109810 760 109870 770
rect 109810 720 109820 760
rect 109820 720 109860 760
rect 109860 720 109870 760
rect 109810 710 109870 720
rect 109510 -790 109570 -730
rect 110010 760 110070 770
rect 110010 720 110020 760
rect 110020 720 110060 760
rect 110060 720 110070 760
rect 110010 710 110070 720
rect 110210 760 110270 770
rect 110210 720 110220 760
rect 110220 720 110260 760
rect 110260 720 110270 760
rect 110210 710 110270 720
rect 109910 -790 109970 -730
rect 107690 -1220 107750 -1160
rect 107770 -1220 107830 -1160
rect 107850 -1220 107910 -1160
rect 107690 -1300 107750 -1240
rect 107770 -1300 107830 -1240
rect 107850 -1300 107910 -1240
rect 107690 -1380 107750 -1320
rect 107770 -1380 107830 -1320
rect 107850 -1380 107910 -1320
rect 108090 -1220 108150 -1160
rect 108170 -1220 108230 -1160
rect 108250 -1220 108310 -1160
rect 108090 -1300 108150 -1240
rect 108170 -1300 108230 -1240
rect 108250 -1300 108310 -1240
rect 108090 -1380 108150 -1320
rect 108170 -1380 108230 -1320
rect 108250 -1380 108310 -1320
rect 108790 -1220 108850 -1160
rect 108870 -1220 108930 -1160
rect 108950 -1220 109010 -1160
rect 108790 -1300 108850 -1240
rect 108870 -1300 108930 -1240
rect 108950 -1300 109010 -1240
rect 108790 -1380 108850 -1320
rect 108870 -1380 108930 -1320
rect 108950 -1380 109010 -1320
rect 109310 -1220 109370 -1160
rect 109310 -1300 109370 -1240
rect 109310 -1380 109370 -1320
rect 109490 -1220 109550 -1160
rect 109570 -1220 109630 -1160
rect 109650 -1220 109710 -1160
rect 109490 -1300 109550 -1240
rect 109570 -1300 109630 -1240
rect 109650 -1300 109710 -1240
rect 109490 -1380 109550 -1320
rect 109570 -1380 109630 -1320
rect 109650 -1380 109710 -1320
rect 111350 -180 111410 -120
rect 111430 -180 111490 -120
rect 111510 -180 111570 -120
rect 111350 -260 111410 -200
rect 111430 -260 111490 -200
rect 111510 -260 111570 -200
rect 111350 -340 111410 -280
rect 111430 -340 111490 -280
rect 111510 -340 111570 -280
rect 110310 -790 110370 -730
rect 114180 5790 114240 5800
rect 114180 5750 114190 5790
rect 114190 5750 114230 5790
rect 114230 5750 114240 5790
rect 114180 5740 114240 5750
rect 114330 5650 114390 5660
rect 114330 5610 114340 5650
rect 114340 5610 114380 5650
rect 114380 5610 114390 5650
rect 114330 5600 114390 5610
rect 114040 5500 114100 5560
rect 113710 5390 113770 5450
rect 113930 5390 113990 5450
rect 115630 5500 115690 5560
rect 113880 5280 113940 5340
rect 114430 5280 114490 5340
rect 113710 5220 113770 5230
rect 113710 5180 113720 5220
rect 113720 5180 113760 5220
rect 113760 5180 113770 5220
rect 113710 5170 113770 5180
rect 112180 4880 112240 4940
rect 112290 4880 112350 4940
rect 112400 4880 112460 4940
rect 112510 4880 112570 4940
rect 112620 4880 112680 4940
rect 112730 4880 112790 4940
rect 112840 4880 112900 4940
rect 112950 4880 113010 4940
rect 113060 4880 113120 4940
rect 113170 4880 113230 4940
rect 113280 4880 113340 4940
rect 112180 4800 112240 4860
rect 112290 4800 112350 4860
rect 112400 4800 112460 4860
rect 112510 4800 112570 4860
rect 112620 4800 112680 4860
rect 112730 4800 112790 4860
rect 112840 4800 112900 4860
rect 112950 4800 113010 4860
rect 113060 4800 113120 4860
rect 113170 4800 113230 4860
rect 113280 4800 113340 4860
rect 112180 4720 112240 4780
rect 112290 4720 112350 4780
rect 112400 4720 112460 4780
rect 112510 4720 112570 4780
rect 112620 4720 112680 4780
rect 112730 4720 112790 4780
rect 112840 4720 112900 4780
rect 112950 4720 113010 4780
rect 113060 4720 113120 4780
rect 113170 4720 113230 4780
rect 113280 4720 113340 4780
rect 112180 3960 112240 4020
rect 112400 3960 112460 4020
rect 112620 3960 112680 4020
rect 112840 3960 112900 4020
rect 113060 3960 113120 4020
rect 114260 4880 114320 4940
rect 114370 4880 114430 4940
rect 114480 4880 114540 4940
rect 114590 4880 114650 4940
rect 114700 4880 114760 4940
rect 114810 4880 114870 4940
rect 114920 4880 114980 4940
rect 115030 4880 115090 4940
rect 115140 4880 115200 4940
rect 115250 4880 115310 4940
rect 115360 4880 115420 4940
rect 114260 4800 114320 4860
rect 114370 4800 114430 4860
rect 114480 4800 114540 4860
rect 114590 4800 114650 4860
rect 114700 4800 114760 4860
rect 114810 4800 114870 4860
rect 114920 4800 114980 4860
rect 115030 4800 115090 4860
rect 115140 4800 115200 4860
rect 115250 4800 115310 4860
rect 115360 4800 115420 4860
rect 114260 4720 114320 4780
rect 114370 4720 114430 4780
rect 114480 4720 114540 4780
rect 114590 4720 114650 4780
rect 114700 4720 114760 4780
rect 114810 4720 114870 4780
rect 114920 4720 114980 4780
rect 115030 4720 115090 4780
rect 115140 4720 115200 4780
rect 115250 4720 115310 4780
rect 115360 4720 115420 4780
rect 113550 4580 113610 4590
rect 113550 4540 113560 4580
rect 113560 4540 113600 4580
rect 113600 4540 113610 4580
rect 113550 4530 113610 4540
rect 113550 4450 113610 4510
rect 113550 4370 113610 4430
rect 113770 4530 113830 4590
rect 113770 4450 113830 4510
rect 113770 4370 113830 4430
rect 113990 4580 114050 4590
rect 113990 4540 114000 4580
rect 114000 4540 114040 4580
rect 114040 4540 114050 4580
rect 113990 4530 114050 4540
rect 113990 4450 114050 4510
rect 113990 4370 114050 4430
rect 113280 3960 113340 4020
rect 113580 3960 113640 4020
rect 112238 3900 112292 3910
rect 112238 3860 112245 3900
rect 112245 3860 112285 3900
rect 112285 3860 112292 3900
rect 112238 3850 112292 3860
rect 112348 3900 112402 3910
rect 112348 3860 112355 3900
rect 112355 3860 112395 3900
rect 112395 3860 112402 3900
rect 112348 3850 112402 3860
rect 112458 3900 112512 3910
rect 112458 3860 112465 3900
rect 112465 3860 112505 3900
rect 112505 3860 112512 3900
rect 112458 3850 112512 3860
rect 112568 3900 112622 3910
rect 112568 3860 112575 3900
rect 112575 3860 112615 3900
rect 112615 3860 112622 3900
rect 112568 3850 112622 3860
rect 112678 3900 112732 3910
rect 112678 3860 112685 3900
rect 112685 3860 112725 3900
rect 112725 3860 112732 3900
rect 112678 3850 112732 3860
rect 112788 3900 112842 3910
rect 112788 3860 112795 3900
rect 112795 3860 112835 3900
rect 112835 3860 112842 3900
rect 112788 3850 112842 3860
rect 112898 3900 112952 3910
rect 112898 3860 112905 3900
rect 112905 3860 112945 3900
rect 112945 3860 112952 3900
rect 112898 3850 112952 3860
rect 113008 3900 113062 3910
rect 113008 3860 113015 3900
rect 113015 3860 113055 3900
rect 113055 3860 113062 3900
rect 113008 3850 113062 3860
rect 113118 3900 113172 3910
rect 113118 3860 113125 3900
rect 113125 3860 113165 3900
rect 113165 3860 113172 3900
rect 113118 3850 113172 3860
rect 113228 3900 113282 3910
rect 113228 3860 113235 3900
rect 113235 3860 113275 3900
rect 113275 3860 113282 3900
rect 113228 3850 113282 3860
rect 112290 3440 112350 3500
rect 112180 3330 112240 3390
rect 112070 3220 112130 3280
rect 112070 3140 112130 3200
rect 112070 3060 112130 3120
rect 112510 3440 112570 3500
rect 112400 3330 112460 3390
rect 112080 2580 112140 2590
rect 112080 2540 112090 2580
rect 112090 2540 112130 2580
rect 112130 2540 112140 2580
rect 112180 2550 112240 2610
rect 112290 2570 112350 2630
rect 112730 3440 112790 3500
rect 112620 3330 112680 3390
rect 112400 2550 112460 2610
rect 112510 2570 112570 2630
rect 112950 3440 113010 3500
rect 112840 3330 112900 3390
rect 112620 2550 112680 2610
rect 112730 2570 112790 2630
rect 113170 3440 113230 3500
rect 113060 3330 113120 3390
rect 112840 2550 112900 2610
rect 112950 2570 113010 2630
rect 113280 3330 113340 3390
rect 113580 3330 113640 3390
rect 113960 3960 114020 4020
rect 114260 3960 114320 4020
rect 114480 3960 114540 4020
rect 114700 3960 114760 4020
rect 114920 3960 114980 4020
rect 115140 3960 115200 4020
rect 115360 3960 115420 4020
rect 114318 3900 114372 3910
rect 114318 3860 114325 3900
rect 114325 3860 114365 3900
rect 114365 3860 114372 3900
rect 114318 3850 114372 3860
rect 114428 3900 114482 3910
rect 114428 3860 114435 3900
rect 114435 3860 114475 3900
rect 114475 3860 114482 3900
rect 114428 3850 114482 3860
rect 114538 3900 114592 3910
rect 114538 3860 114545 3900
rect 114545 3860 114585 3900
rect 114585 3860 114592 3900
rect 114538 3850 114592 3860
rect 114648 3900 114702 3910
rect 114648 3860 114655 3900
rect 114655 3860 114695 3900
rect 114695 3860 114702 3900
rect 114648 3850 114702 3860
rect 114758 3900 114812 3910
rect 114758 3860 114765 3900
rect 114765 3860 114805 3900
rect 114805 3860 114812 3900
rect 114758 3850 114812 3860
rect 114868 3900 114922 3910
rect 114868 3860 114875 3900
rect 114875 3860 114915 3900
rect 114915 3860 114922 3900
rect 114868 3850 114922 3860
rect 114978 3900 115032 3910
rect 114978 3860 114985 3900
rect 114985 3860 115025 3900
rect 115025 3860 115032 3900
rect 114978 3850 115032 3860
rect 115088 3900 115142 3910
rect 115088 3860 115095 3900
rect 115095 3860 115135 3900
rect 115135 3860 115142 3900
rect 115088 3850 115142 3860
rect 115198 3900 115252 3910
rect 115198 3860 115205 3900
rect 115205 3860 115245 3900
rect 115245 3860 115252 3900
rect 115198 3850 115252 3860
rect 115308 3900 115362 3910
rect 115308 3860 115315 3900
rect 115315 3860 115355 3900
rect 115355 3860 115362 3900
rect 115308 3850 115362 3860
rect 113960 3330 114020 3390
rect 114370 3440 114430 3500
rect 114260 3330 114320 3390
rect 113390 3220 113450 3280
rect 113390 3140 113450 3200
rect 113390 3060 113450 3120
rect 114150 3220 114210 3280
rect 114150 3140 114210 3200
rect 114150 3060 114210 3120
rect 113770 2910 113830 2970
rect 113770 2830 113830 2890
rect 113770 2750 113830 2810
rect 113060 2550 113120 2610
rect 113170 2570 113230 2630
rect 113280 2550 113340 2610
rect 113380 2600 113440 2610
rect 113380 2560 113390 2600
rect 113390 2560 113430 2600
rect 113430 2560 113440 2600
rect 113380 2550 113440 2560
rect 113680 2600 113740 2610
rect 113680 2560 113690 2600
rect 113690 2560 113730 2600
rect 113730 2560 113740 2600
rect 113680 2550 113740 2560
rect 112080 2530 112140 2540
rect 112290 2460 112350 2520
rect 112180 2070 112240 2130
rect 112510 2460 112570 2520
rect 112400 2070 112460 2130
rect 112730 2460 112790 2520
rect 112620 2070 112680 2130
rect 112950 2460 113010 2520
rect 112840 2070 112900 2130
rect 113170 2460 113230 2520
rect 113060 2070 113120 2130
rect 113280 2070 113340 2130
rect 114590 3440 114650 3500
rect 114480 3330 114540 3390
rect 113860 2600 113920 2610
rect 113860 2560 113870 2600
rect 113870 2560 113910 2600
rect 113910 2560 113920 2600
rect 113860 2550 113920 2560
rect 114160 2600 114220 2610
rect 114160 2560 114170 2600
rect 114170 2560 114210 2600
rect 114210 2560 114220 2600
rect 114160 2550 114220 2560
rect 114260 2550 114320 2610
rect 114370 2570 114430 2630
rect 114810 3440 114870 3500
rect 114700 3330 114760 3390
rect 114480 2550 114540 2610
rect 114590 2570 114650 2630
rect 115030 3440 115090 3500
rect 114920 3330 114980 3390
rect 114700 2550 114760 2610
rect 114810 2570 114870 2630
rect 115250 3440 115310 3500
rect 115140 3330 115200 3390
rect 114920 2550 114980 2610
rect 115030 2570 115090 2630
rect 115360 3330 115420 3390
rect 115470 3220 115530 3280
rect 115470 3140 115530 3200
rect 115470 3060 115530 3120
rect 115140 2550 115200 2610
rect 115250 2570 115310 2630
rect 115360 2550 115420 2610
rect 115460 2580 115520 2590
rect 115460 2540 115470 2580
rect 115470 2540 115510 2580
rect 115510 2540 115520 2580
rect 114370 2460 114430 2520
rect 113660 2070 113720 2130
rect 112290 1930 112350 1990
rect 112510 1930 112570 1990
rect 112730 1930 112790 1990
rect 112950 1930 113010 1990
rect 113170 1930 113230 1990
rect 112070 1820 112130 1880
rect 112070 1740 112130 1800
rect 112070 1660 112130 1720
rect 111890 1550 111950 1610
rect 113470 1820 113530 1880
rect 113470 1740 113530 1800
rect 113470 1660 113530 1720
rect 112890 970 112950 1030
rect 113110 970 113170 1030
rect 113330 970 113390 1030
rect 113550 970 113610 1030
rect 113880 2070 113940 2130
rect 113770 970 113830 1030
rect 114260 2070 114320 2130
rect 114590 2460 114650 2520
rect 114480 2070 114540 2130
rect 114810 2460 114870 2520
rect 114700 2070 114760 2130
rect 115030 2460 115090 2520
rect 114920 2070 114980 2130
rect 115250 2460 115310 2520
rect 115140 2070 115200 2130
rect 115460 2530 115520 2540
rect 115360 2070 115420 2130
rect 114370 1930 114430 1990
rect 114590 1930 114650 1990
rect 114070 1820 114130 1880
rect 114070 1740 114130 1800
rect 114070 1660 114130 1720
rect 113990 970 114050 1030
rect 114810 1930 114870 1990
rect 115030 1930 115090 1990
rect 115250 1930 115310 1990
rect 115470 1820 115530 1880
rect 115470 1740 115530 1800
rect 115470 1660 115530 1720
rect 115740 5280 115800 5340
rect 115650 1550 115710 1610
rect 114210 970 114270 1030
rect 114430 970 114490 1030
rect 114650 970 114710 1030
rect 114870 970 114930 1030
rect 111700 -560 111760 -500
rect 111780 -560 111840 -500
rect 111700 -1000 111760 -940
rect 111780 -1000 111840 -940
rect 112450 360 112510 370
rect 112450 320 112460 360
rect 112460 320 112500 360
rect 112500 320 112510 360
rect 112450 310 112510 320
rect 112560 310 112620 370
rect 112780 310 112840 370
rect 113000 310 113060 370
rect 113220 310 113280 370
rect 113440 310 113500 370
rect 113660 310 113720 370
rect 113880 310 113940 370
rect 114100 310 114160 370
rect 114320 310 114380 370
rect 114540 310 114600 370
rect 114760 310 114820 370
rect 114980 360 115040 370
rect 114980 320 114990 360
rect 114990 320 115030 360
rect 115030 320 115040 360
rect 114980 310 115040 320
rect 112890 200 112950 260
rect 112890 120 112950 180
rect 112890 40 112950 100
rect 113110 200 113170 260
rect 113110 120 113170 180
rect 113110 40 113170 100
rect 113330 200 113390 260
rect 113330 120 113390 180
rect 113330 40 113390 100
rect 113550 200 113610 260
rect 113550 120 113610 180
rect 113550 40 113610 100
rect 113770 200 113830 260
rect 113770 120 113830 180
rect 113770 40 113830 100
rect 113990 200 114050 260
rect 113990 120 114050 180
rect 113990 40 114050 100
rect 114210 200 114270 260
rect 114210 120 114270 180
rect 114210 40 114270 100
rect 114430 200 114490 260
rect 114430 120 114490 180
rect 114430 40 114490 100
rect 114650 200 114710 260
rect 114650 120 114710 180
rect 114650 40 114710 100
rect 114870 200 114930 260
rect 114870 120 114930 180
rect 114870 40 114930 100
rect 114840 -20 114900 -10
rect 114840 -60 114850 -20
rect 114850 -60 114890 -20
rect 114890 -60 114900 -20
rect 114840 -70 114900 -60
rect 112670 -180 112730 -120
rect 112670 -260 112730 -200
rect 112670 -340 112730 -280
rect 113090 -450 113150 -390
rect 113310 -450 113370 -390
rect 113750 -450 113810 -390
rect 112980 -560 113040 -500
rect 113200 -510 113260 -500
rect 113200 -550 113210 -510
rect 113210 -550 113250 -510
rect 113250 -550 113260 -510
rect 113200 -560 113260 -550
rect 112980 -1000 113040 -940
rect 113420 -560 113480 -500
rect 113200 -1000 113260 -940
rect 114090 -510 114150 -500
rect 114090 -550 114100 -510
rect 114100 -550 114140 -510
rect 114140 -550 114150 -510
rect 114090 -560 114150 -550
rect 114430 -850 114440 -650
rect 114440 -850 114480 -650
rect 114480 -850 114490 -650
rect 113420 -1000 113480 -940
rect 113090 -1110 113150 -1050
rect 113310 -1110 113370 -1050
rect 114090 -950 114150 -940
rect 114090 -990 114100 -950
rect 114100 -990 114140 -950
rect 114140 -990 114150 -950
rect 114090 -1000 114150 -990
rect 113750 -1110 113810 -1050
rect 110190 -1220 110250 -1160
rect 110270 -1220 110330 -1160
rect 110350 -1220 110410 -1160
rect 110190 -1300 110250 -1240
rect 110270 -1300 110330 -1240
rect 110350 -1300 110410 -1240
rect 110190 -1380 110250 -1320
rect 110270 -1380 110330 -1320
rect 110350 -1380 110410 -1320
rect 110510 -1220 110570 -1160
rect 110510 -1300 110570 -1240
rect 110510 -1380 110570 -1320
rect 110890 -1220 110950 -1160
rect 110970 -1220 111030 -1160
rect 111050 -1220 111110 -1160
rect 110890 -1300 110950 -1240
rect 110970 -1300 111030 -1240
rect 111050 -1300 111110 -1240
rect 110890 -1380 110950 -1320
rect 110970 -1380 111030 -1320
rect 111050 -1380 111110 -1320
rect 111590 -1220 111650 -1160
rect 111670 -1220 111730 -1160
rect 111750 -1220 111810 -1160
rect 111590 -1300 111650 -1240
rect 111670 -1300 111730 -1240
rect 111750 -1300 111810 -1240
rect 111590 -1380 111650 -1320
rect 111670 -1380 111730 -1320
rect 111750 -1380 111810 -1320
rect 112290 -1220 112350 -1160
rect 112370 -1220 112430 -1160
rect 112450 -1220 112510 -1160
rect 112290 -1300 112350 -1240
rect 112370 -1300 112430 -1240
rect 112450 -1300 112510 -1240
rect 112290 -1380 112350 -1320
rect 112370 -1380 112430 -1320
rect 112450 -1380 112510 -1320
rect 112870 -1220 112930 -1160
rect 112870 -1300 112930 -1240
rect 112870 -1380 112930 -1320
rect 112990 -1220 113050 -1160
rect 113070 -1220 113130 -1160
rect 113150 -1220 113210 -1160
rect 112990 -1300 113050 -1240
rect 113070 -1300 113130 -1240
rect 113150 -1300 113210 -1240
rect 112990 -1380 113050 -1320
rect 113070 -1380 113130 -1320
rect 113150 -1380 113210 -1320
rect 113530 -1220 113590 -1160
rect 113530 -1300 113590 -1240
rect 113530 -1380 113590 -1320
rect 113690 -1220 113750 -1160
rect 113770 -1220 113830 -1160
rect 113850 -1220 113910 -1160
rect 113690 -1300 113750 -1240
rect 113770 -1300 113830 -1240
rect 113850 -1300 113910 -1240
rect 113690 -1380 113750 -1320
rect 113770 -1380 113830 -1320
rect 113850 -1380 113910 -1320
rect 114390 -1220 114450 -1160
rect 114470 -1220 114530 -1160
rect 114550 -1220 114610 -1160
rect 114390 -1300 114450 -1240
rect 114470 -1300 114530 -1240
rect 114550 -1300 114610 -1240
rect 114390 -1380 114450 -1320
rect 114470 -1380 114530 -1320
rect 114550 -1380 114610 -1320
rect 115430 200 115490 260
rect 115510 200 115570 260
rect 115590 200 115650 260
rect 115430 120 115490 180
rect 115510 120 115570 180
rect 115590 120 115650 180
rect 115430 40 115490 100
rect 115510 40 115570 100
rect 115590 40 115650 100
rect 116030 4530 116090 4590
rect 116110 4530 116170 4590
rect 116190 4530 116250 4590
rect 116030 4450 116090 4510
rect 116110 4450 116170 4510
rect 116190 4450 116250 4510
rect 116030 4370 116090 4430
rect 116110 4370 116170 4430
rect 116190 4370 116250 4430
rect 116030 4040 116090 4100
rect 116110 4040 116170 4100
rect 116190 4040 116250 4100
rect 116030 3960 116090 4020
rect 116110 3960 116170 4020
rect 116190 3960 116250 4020
rect 116030 3880 116090 3940
rect 116110 3880 116170 3940
rect 116190 3880 116250 3940
rect 116030 3220 116090 3280
rect 116110 3220 116170 3280
rect 116190 3220 116250 3280
rect 116030 3140 116090 3200
rect 116110 3140 116170 3200
rect 116190 3140 116250 3200
rect 116030 3060 116090 3120
rect 116110 3060 116170 3120
rect 116190 3060 116250 3120
rect 116300 4310 116360 4370
rect 116380 4310 116440 4370
rect 116460 4310 116520 4370
rect 116300 4230 116360 4290
rect 116380 4230 116440 4290
rect 116460 4230 116520 4290
rect 116300 4150 116360 4210
rect 116380 4150 116440 4210
rect 116460 4150 116520 4210
rect 116030 2910 116090 2970
rect 116110 2910 116170 2970
rect 116190 2910 116250 2970
rect 116030 2830 116090 2890
rect 116110 2830 116170 2890
rect 116190 2830 116250 2890
rect 116030 2750 116090 2810
rect 116110 2750 116170 2810
rect 116190 2750 116250 2810
rect 115740 -70 115800 -10
rect 116570 6990 116630 7050
rect 116650 6990 116710 7050
rect 116730 6990 116790 7050
rect 117150 7800 117210 7860
rect 117390 7800 117450 7860
rect 118350 8580 118410 8640
rect 118350 8500 118410 8560
rect 118350 8420 118410 8480
rect 117750 8310 117810 8370
rect 117750 8230 117810 8290
rect 117750 8150 117810 8210
rect 117750 8070 117810 8130
rect 117750 7990 117810 8050
rect 117750 7910 117810 7970
rect 117990 8310 118050 8370
rect 117990 8230 118050 8290
rect 117990 8150 118050 8210
rect 117990 8070 118050 8130
rect 117990 7990 118050 8050
rect 117990 7910 118050 7970
rect 118230 8310 118290 8370
rect 118230 8230 118290 8290
rect 118230 8150 118290 8210
rect 118230 8070 118290 8130
rect 118230 7990 118290 8050
rect 118230 7910 118290 7970
rect 117630 7800 117690 7860
rect 117870 7800 117930 7860
rect 118110 7800 118170 7860
rect 119290 8580 119350 8640
rect 119370 8580 119430 8640
rect 119450 8580 119510 8640
rect 119290 8500 119350 8560
rect 119370 8500 119430 8560
rect 119450 8500 119510 8560
rect 119290 8420 119350 8480
rect 119370 8420 119430 8480
rect 119450 8420 119510 8480
rect 120690 8580 120750 8640
rect 120770 8580 120830 8640
rect 120850 8580 120910 8640
rect 120690 8500 120750 8560
rect 120770 8500 120830 8560
rect 120850 8500 120910 8560
rect 120690 8420 120750 8480
rect 120770 8420 120830 8480
rect 120850 8420 120910 8480
rect 121390 8580 121450 8640
rect 121470 8580 121530 8640
rect 121550 8580 121610 8640
rect 121390 8500 121450 8560
rect 121470 8500 121530 8560
rect 121550 8500 121610 8560
rect 121390 8420 121450 8480
rect 121470 8420 121530 8480
rect 121550 8420 121610 8480
rect 122090 8580 122150 8640
rect 122170 8580 122230 8640
rect 122250 8580 122310 8640
rect 122090 8500 122150 8560
rect 122170 8500 122230 8560
rect 122250 8500 122310 8560
rect 122090 8420 122150 8480
rect 122170 8420 122230 8480
rect 122250 8420 122310 8480
rect 122790 8580 122850 8640
rect 122870 8580 122930 8640
rect 122950 8580 123010 8640
rect 122790 8500 122850 8560
rect 122870 8500 122930 8560
rect 122950 8500 123010 8560
rect 122790 8420 122850 8480
rect 122870 8420 122930 8480
rect 122950 8420 123010 8480
rect 118350 7850 118410 7860
rect 118350 7810 118360 7850
rect 118360 7810 118400 7850
rect 118400 7810 118410 7850
rect 118350 7800 118410 7810
rect 117030 6990 117090 7050
rect 117270 6990 117330 7050
rect 117510 6990 117570 7050
rect 117750 6990 117810 7050
rect 117990 6990 118050 7050
rect 118230 6990 118290 7050
rect 117090 6930 117150 6940
rect 117090 6890 117100 6930
rect 117100 6890 117140 6930
rect 117140 6890 117150 6930
rect 117090 6880 117150 6890
rect 117210 6930 117270 6940
rect 117210 6890 117220 6930
rect 117220 6890 117260 6930
rect 117260 6890 117270 6930
rect 117210 6880 117270 6890
rect 117330 6930 117390 6940
rect 117330 6890 117340 6930
rect 117340 6890 117380 6930
rect 117380 6890 117390 6930
rect 117330 6880 117390 6890
rect 117450 6930 117510 6940
rect 117450 6890 117460 6930
rect 117460 6890 117500 6930
rect 117500 6890 117510 6930
rect 117450 6880 117510 6890
rect 117570 6930 117630 6940
rect 117570 6890 117580 6930
rect 117580 6890 117620 6930
rect 117620 6890 117630 6930
rect 117570 6880 117630 6890
rect 117690 6930 117750 6940
rect 117690 6890 117700 6930
rect 117700 6890 117740 6930
rect 117740 6890 117750 6930
rect 117690 6880 117750 6890
rect 117810 6930 117870 6940
rect 117810 6890 117820 6930
rect 117820 6890 117860 6930
rect 117860 6890 117870 6930
rect 117810 6880 117870 6890
rect 117930 6930 117990 6940
rect 117930 6890 117940 6930
rect 117940 6890 117980 6930
rect 117980 6890 117990 6930
rect 117930 6880 117990 6890
rect 118050 6930 118110 6940
rect 118050 6890 118060 6930
rect 118060 6890 118100 6930
rect 118100 6890 118110 6930
rect 118050 6880 118110 6890
rect 118170 6930 118230 6940
rect 118170 6890 118180 6930
rect 118180 6890 118220 6930
rect 118220 6890 118230 6930
rect 118170 6880 118230 6890
rect 117630 6760 117690 6820
rect 116970 6650 117030 6710
rect 116970 6570 117030 6630
rect 116970 6490 117030 6550
rect 117190 6650 117250 6710
rect 117190 6570 117250 6630
rect 117190 6490 117250 6550
rect 117410 6650 117470 6710
rect 117410 6570 117470 6630
rect 117410 6490 117470 6550
rect 117630 6650 117690 6710
rect 117630 6570 117690 6630
rect 117630 6490 117690 6550
rect 117850 6650 117910 6710
rect 117850 6570 117910 6630
rect 117850 6490 117910 6550
rect 118070 6650 118130 6710
rect 118070 6570 118130 6630
rect 118070 6490 118130 6550
rect 118290 6650 118350 6710
rect 118290 6570 118350 6630
rect 118290 6490 118350 6550
rect 119020 6690 119080 6750
rect 117080 6320 117140 6380
rect 117300 6320 117360 6380
rect 117520 6320 117580 6380
rect 117740 6320 117800 6380
rect 117960 6320 118020 6380
rect 118180 6320 118240 6380
rect 116570 4880 116630 4940
rect 116650 4880 116710 4940
rect 116730 4880 116790 4940
rect 116570 4800 116630 4860
rect 116650 4800 116710 4860
rect 116730 4800 116790 4860
rect 116570 4720 116630 4780
rect 116650 4720 116710 4780
rect 116730 4720 116790 4780
rect 117080 5040 117140 5100
rect 117300 5040 117360 5100
rect 117520 5040 117580 5100
rect 117740 5040 117800 5100
rect 117630 4930 117690 4940
rect 117630 4890 117640 4930
rect 117640 4890 117680 4930
rect 117680 4890 117690 4930
rect 117630 4880 117690 4890
rect 117630 4850 117690 4860
rect 117630 4810 117640 4850
rect 117640 4810 117680 4850
rect 117680 4810 117690 4850
rect 117630 4800 117690 4810
rect 117630 4770 117690 4780
rect 117630 4730 117640 4770
rect 117640 4730 117680 4770
rect 117680 4730 117690 4770
rect 117630 4720 117690 4730
rect 117960 5040 118020 5100
rect 118180 5040 118240 5100
rect 118940 4880 119000 4940
rect 119020 4880 119080 4940
rect 119100 4880 119160 4940
rect 118940 4800 119000 4860
rect 119020 4800 119080 4860
rect 119100 4800 119160 4860
rect 118940 4720 119000 4780
rect 119020 4720 119080 4780
rect 119100 4720 119160 4780
rect 117080 4580 117140 4640
rect 117190 4580 117250 4640
rect 117300 4580 117360 4640
rect 117410 4580 117470 4640
rect 117520 4580 117580 4640
rect 117630 4580 117690 4640
rect 117740 4580 117800 4640
rect 117850 4580 117910 4640
rect 117960 4580 118020 4640
rect 118070 4580 118130 4640
rect 118180 4580 118240 4640
rect 117080 4500 117140 4560
rect 117190 4500 117250 4560
rect 117300 4500 117360 4560
rect 117410 4500 117470 4560
rect 117520 4500 117580 4560
rect 117630 4500 117690 4560
rect 117740 4500 117800 4560
rect 117850 4500 117910 4560
rect 117960 4500 118020 4560
rect 118070 4500 118130 4560
rect 118180 4500 118240 4560
rect 117080 4420 117140 4480
rect 117190 4420 117250 4480
rect 117300 4420 117360 4480
rect 117410 4420 117470 4480
rect 117520 4420 117580 4480
rect 117630 4420 117690 4480
rect 117740 4420 117800 4480
rect 117850 4420 117910 4480
rect 117960 4420 118020 4480
rect 118070 4420 118130 4480
rect 118180 4420 118240 4480
rect 119130 4580 119190 4640
rect 119210 4580 119270 4640
rect 119300 4580 119360 4640
rect 119380 4580 119440 4640
rect 119470 4580 119530 4640
rect 119550 4580 119610 4640
rect 119130 4500 119190 4560
rect 119210 4500 119270 4560
rect 119300 4500 119360 4560
rect 119380 4500 119440 4560
rect 119470 4500 119530 4560
rect 119550 4500 119610 4560
rect 119130 4420 119190 4480
rect 119210 4420 119270 4480
rect 119300 4420 119360 4480
rect 119380 4420 119440 4480
rect 119470 4420 119530 4480
rect 119550 4420 119610 4480
rect 116970 4310 117030 4370
rect 116970 4230 117030 4290
rect 116970 4150 117030 4210
rect 118290 4310 118350 4370
rect 118290 4230 118350 4290
rect 118290 4150 118350 4210
rect 117080 4040 117140 4100
rect 117080 3960 117140 4020
rect 117080 3880 117140 3940
rect 117300 4040 117360 4100
rect 117300 3960 117360 4020
rect 117300 3880 117360 3940
rect 117520 4040 117580 4100
rect 117520 3960 117580 4020
rect 117520 3880 117580 3940
rect 117740 4040 117800 4100
rect 117740 3960 117800 4020
rect 117740 3880 117800 3940
rect 117960 4040 118020 4100
rect 117960 3960 118020 4020
rect 117960 3880 118020 3940
rect 118180 4040 118240 4100
rect 118180 3960 118240 4020
rect 118180 3880 118240 3940
rect 117190 3770 117250 3830
rect 117410 3770 117470 3830
rect 117630 3770 117690 3830
rect 117850 3770 117910 3830
rect 118070 3770 118130 3830
rect 119140 3360 119200 3420
rect 119240 3360 119300 3420
rect 119340 3360 119400 3420
rect 119440 3360 119500 3420
rect 119540 3360 119600 3420
rect 117190 3310 117250 3320
rect 117190 3270 117200 3310
rect 117200 3270 117240 3310
rect 117240 3270 117250 3310
rect 117190 3260 117250 3270
rect 117410 3310 117470 3320
rect 117410 3270 117420 3310
rect 117420 3270 117460 3310
rect 117460 3270 117470 3310
rect 117410 3260 117470 3270
rect 117630 3310 117690 3320
rect 117630 3270 117640 3310
rect 117640 3270 117680 3310
rect 117680 3270 117690 3310
rect 117630 3260 117690 3270
rect 117850 3310 117910 3320
rect 117850 3270 117860 3310
rect 117860 3270 117900 3310
rect 117900 3270 117910 3310
rect 117850 3260 117910 3270
rect 118070 3310 118130 3320
rect 118070 3270 118080 3310
rect 118080 3270 118120 3310
rect 118120 3270 118130 3310
rect 118070 3260 118130 3270
rect 118560 3260 118620 3320
rect 119140 3260 119200 3320
rect 119240 3260 119300 3320
rect 119340 3260 119400 3320
rect 119440 3260 119500 3320
rect 119540 3260 119600 3320
rect 116570 3130 116630 3190
rect 116650 3130 116710 3190
rect 116730 3130 116790 3190
rect 116570 3050 116630 3110
rect 116650 3050 116710 3110
rect 116730 3050 116790 3110
rect 117300 3180 117360 3190
rect 117300 3140 117310 3180
rect 117310 3140 117350 3180
rect 117350 3140 117360 3180
rect 117300 3130 117360 3140
rect 117300 3100 117360 3110
rect 117300 3060 117310 3100
rect 117310 3060 117350 3100
rect 117350 3060 117360 3100
rect 117300 3050 117360 3060
rect 117190 2890 117250 2950
rect 117410 2890 117470 2950
rect 117630 2890 117690 2950
rect 117850 2890 117910 2950
rect 118070 2890 118130 2950
rect 118470 2890 118530 2950
rect 116300 2100 116360 2160
rect 116380 2100 116440 2160
rect 116460 2100 116520 2160
rect 116300 2020 116360 2080
rect 116380 2020 116440 2080
rect 116460 2020 116520 2080
rect 116300 1940 116360 2000
rect 116380 1940 116440 2000
rect 116460 1940 116520 2000
rect 117190 2210 117250 2270
rect 117410 2210 117470 2270
rect 117630 2210 117690 2270
rect 117850 2210 117910 2270
rect 118070 2210 118130 2270
rect 118470 2250 118530 2310
rect 117080 2100 117140 2160
rect 117080 2020 117140 2080
rect 117080 1940 117140 2000
rect 117300 2100 117360 2160
rect 117300 2020 117360 2080
rect 117300 1940 117360 2000
rect 117520 2100 117580 2160
rect 117520 2020 117580 2080
rect 117520 1940 117580 2000
rect 117740 2100 117800 2160
rect 117740 2020 117800 2080
rect 117740 1940 117800 2000
rect 117960 2100 118020 2160
rect 117960 2020 118020 2080
rect 117960 1940 118020 2000
rect 118180 2100 118240 2160
rect 118180 2020 118240 2080
rect 118180 1940 118240 2000
rect 119140 3160 119200 3220
rect 119240 3160 119300 3220
rect 119340 3160 119400 3220
rect 119440 3160 119500 3220
rect 119540 3160 119600 3220
rect 118660 2310 118730 2320
rect 118660 2260 118670 2310
rect 118670 2260 118720 2310
rect 118720 2260 118730 2310
rect 118660 2250 118730 2260
rect 118780 2310 118850 2320
rect 118780 2260 118790 2310
rect 118790 2260 118840 2310
rect 118840 2260 118850 2310
rect 118780 2250 118850 2260
rect 118900 2310 118970 2320
rect 118900 2260 118910 2310
rect 118910 2260 118960 2310
rect 118960 2260 118970 2310
rect 118900 2250 118970 2260
rect 119020 2310 119090 2320
rect 119020 2260 119030 2310
rect 119030 2260 119080 2310
rect 119080 2260 119090 2310
rect 119020 2250 119090 2260
rect 118560 2110 118620 2170
rect 118780 2110 118840 2170
rect 116970 1820 117030 1880
rect 116970 1740 117030 1800
rect 116970 1660 117030 1720
rect 118290 1820 118350 1880
rect 118290 1740 118350 1800
rect 118290 1660 118350 1720
rect 119020 1550 119080 1610
rect 118890 1090 118950 1150
rect 117230 980 117290 1040
rect 117310 980 117370 1040
rect 117390 980 117450 1040
rect 117470 980 117530 1040
rect 117550 980 117610 1040
rect 117630 980 117690 1040
rect 117710 980 117770 1040
rect 117790 980 117850 1040
rect 117870 980 117930 1040
rect 117950 980 118010 1040
rect 118030 980 118090 1040
rect 117230 900 117290 960
rect 117310 900 117370 960
rect 117390 900 117450 960
rect 117470 900 117530 960
rect 117550 900 117610 960
rect 117630 900 117690 960
rect 117710 900 117770 960
rect 117790 900 117850 960
rect 117870 900 117930 960
rect 117950 900 118010 960
rect 118030 900 118090 960
rect 117230 820 117290 880
rect 117310 820 117370 880
rect 117390 820 117450 880
rect 117470 820 117530 880
rect 117550 820 117610 880
rect 117630 820 117690 880
rect 117710 820 117770 880
rect 117790 820 117850 880
rect 117870 820 117930 880
rect 117950 820 118010 880
rect 118030 820 118090 880
rect 118760 980 118820 1040
rect 118760 900 118820 960
rect 118760 820 118820 880
rect 116030 -180 116090 -120
rect 116110 -180 116170 -120
rect 116190 -180 116250 -120
rect 116030 -260 116090 -200
rect 116110 -260 116170 -200
rect 116190 -260 116250 -200
rect 116030 -340 116090 -280
rect 116110 -340 116170 -280
rect 116190 -340 116250 -280
rect 115430 -700 115490 -640
rect 115510 -700 115570 -640
rect 115590 -700 115650 -640
rect 115430 -780 115490 -720
rect 115510 -780 115570 -720
rect 115590 -780 115650 -720
rect 115430 -860 115490 -800
rect 115510 -860 115570 -800
rect 115590 -860 115650 -800
rect 117330 760 117390 770
rect 117330 720 117340 760
rect 117340 720 117380 760
rect 117380 720 117390 760
rect 117330 710 117390 720
rect 117530 760 117590 770
rect 117530 720 117540 760
rect 117540 720 117580 760
rect 117580 720 117590 760
rect 117530 710 117590 720
rect 117230 -790 117290 -730
rect 117730 760 117790 770
rect 117730 720 117740 760
rect 117740 720 117780 760
rect 117780 720 117790 760
rect 117730 710 117790 720
rect 117930 760 117990 770
rect 117930 720 117940 760
rect 117940 720 117980 760
rect 117980 720 117990 760
rect 117930 710 117990 720
rect 117630 -790 117690 -730
rect 114980 -1220 115040 -1160
rect 114980 -1300 115040 -1240
rect 114980 -1380 115040 -1320
rect 115090 -1220 115150 -1160
rect 115170 -1220 115230 -1160
rect 115250 -1220 115310 -1160
rect 115090 -1300 115150 -1240
rect 115170 -1300 115230 -1240
rect 115250 -1300 115310 -1240
rect 115090 -1380 115150 -1320
rect 115170 -1380 115230 -1320
rect 115250 -1380 115310 -1320
rect 115790 -1220 115850 -1160
rect 115870 -1220 115930 -1160
rect 115950 -1220 116010 -1160
rect 115790 -1300 115850 -1240
rect 115870 -1300 115930 -1240
rect 115950 -1300 116010 -1240
rect 115790 -1380 115850 -1320
rect 115870 -1380 115930 -1320
rect 115950 -1380 116010 -1320
rect 116490 -1220 116550 -1160
rect 116570 -1220 116630 -1160
rect 116650 -1220 116710 -1160
rect 116490 -1300 116550 -1240
rect 116570 -1300 116630 -1240
rect 116650 -1300 116710 -1240
rect 116490 -1380 116550 -1320
rect 116570 -1380 116630 -1320
rect 116650 -1380 116710 -1320
rect 117030 -1220 117090 -1160
rect 117030 -1300 117090 -1240
rect 117030 -1380 117090 -1320
rect 117190 -1220 117250 -1160
rect 117270 -1220 117330 -1160
rect 117350 -1220 117410 -1160
rect 117190 -1300 117250 -1240
rect 117270 -1300 117330 -1240
rect 117350 -1300 117410 -1240
rect 117190 -1380 117250 -1320
rect 117270 -1380 117330 -1320
rect 117350 -1380 117410 -1320
rect 118760 650 118830 660
rect 118760 600 118770 650
rect 118770 600 118820 650
rect 118820 600 118830 650
rect 118760 590 118830 600
rect 119130 980 119190 1040
rect 119210 980 119270 1040
rect 119300 980 119360 1040
rect 119380 980 119440 1040
rect 119470 980 119530 1040
rect 119550 980 119610 1040
rect 119130 900 119190 960
rect 119210 900 119270 960
rect 119300 900 119360 960
rect 119380 900 119440 960
rect 119470 900 119530 960
rect 119550 900 119610 960
rect 119130 820 119190 880
rect 119210 820 119270 880
rect 119300 820 119360 880
rect 119380 820 119440 880
rect 119470 820 119530 880
rect 119550 820 119610 880
rect 119690 4040 119750 4100
rect 119770 4040 119830 4100
rect 119850 4040 119910 4100
rect 119690 3960 119750 4020
rect 119770 3960 119830 4020
rect 119850 3960 119910 4020
rect 119690 3880 119750 3940
rect 119770 3880 119830 3940
rect 119850 3880 119910 3940
rect 119690 1820 119750 1880
rect 119770 1820 119830 1880
rect 119850 1820 119910 1880
rect 119690 1740 119750 1800
rect 119770 1740 119830 1800
rect 119850 1740 119910 1800
rect 119690 1660 119750 1720
rect 119770 1660 119830 1720
rect 119850 1660 119910 1720
rect 118890 710 118950 770
rect 118880 650 118950 660
rect 118880 600 118890 650
rect 118890 600 118940 650
rect 118940 600 118950 650
rect 118880 590 118950 600
rect 118030 -790 118090 -730
rect 117890 -1220 117950 -1160
rect 117970 -1220 118030 -1160
rect 118050 -1220 118110 -1160
rect 117890 -1300 117950 -1240
rect 117970 -1300 118030 -1240
rect 118050 -1300 118110 -1240
rect 117890 -1380 117950 -1320
rect 117970 -1380 118030 -1320
rect 118050 -1380 118110 -1320
rect 118230 -1220 118290 -1160
rect 118230 -1300 118290 -1240
rect 118230 -1380 118290 -1320
rect 118750 -1220 118810 -1160
rect 118830 -1220 118890 -1160
rect 118910 -1220 118970 -1160
rect 118750 -1300 118810 -1240
rect 118830 -1300 118890 -1240
rect 118910 -1300 118970 -1240
rect 118750 -1380 118810 -1320
rect 118830 -1380 118890 -1320
rect 118910 -1380 118970 -1320
rect 119290 -1220 119350 -1160
rect 119370 -1220 119430 -1160
rect 119450 -1220 119510 -1160
rect 119290 -1300 119350 -1240
rect 119370 -1300 119430 -1240
rect 119450 -1300 119510 -1240
rect 119290 -1380 119350 -1320
rect 119370 -1380 119430 -1320
rect 119450 -1380 119510 -1320
rect 119690 -1220 119750 -1160
rect 119770 -1220 119830 -1160
rect 119850 -1220 119910 -1160
rect 119690 -1300 119750 -1240
rect 119770 -1300 119830 -1240
rect 119850 -1300 119910 -1240
rect 119690 -1380 119750 -1320
rect 119770 -1380 119830 -1320
rect 119850 -1380 119910 -1320
rect 119990 -1220 120050 -1160
rect 120070 -1220 120130 -1160
rect 120150 -1220 120210 -1160
rect 119990 -1300 120050 -1240
rect 120070 -1300 120130 -1240
rect 120150 -1300 120210 -1240
rect 119990 -1380 120050 -1320
rect 120070 -1380 120130 -1320
rect 120150 -1380 120210 -1320
rect 120690 -1220 120750 -1160
rect 120770 -1220 120830 -1160
rect 120850 -1220 120910 -1160
rect 120690 -1300 120750 -1240
rect 120770 -1300 120830 -1240
rect 120850 -1300 120910 -1240
rect 120690 -1380 120750 -1320
rect 120770 -1380 120830 -1320
rect 120850 -1380 120910 -1320
rect 121390 -1220 121450 -1160
rect 121470 -1220 121530 -1160
rect 121550 -1220 121610 -1160
rect 121390 -1300 121450 -1240
rect 121470 -1300 121530 -1240
rect 121550 -1300 121610 -1240
rect 121390 -1380 121450 -1320
rect 121470 -1380 121530 -1320
rect 121550 -1380 121610 -1320
rect 122090 -1220 122150 -1160
rect 122170 -1220 122230 -1160
rect 122250 -1220 122310 -1160
rect 122090 -1300 122150 -1240
rect 122170 -1300 122230 -1240
rect 122250 -1300 122310 -1240
rect 122090 -1380 122150 -1320
rect 122170 -1380 122230 -1320
rect 122250 -1380 122310 -1320
rect 122790 -1220 122850 -1160
rect 122870 -1220 122930 -1160
rect 122950 -1220 123010 -1160
rect 122790 -1300 122850 -1240
rect 122870 -1300 122930 -1240
rect 122950 -1300 123010 -1240
rect 122790 -1380 122850 -1320
rect 122870 -1380 122930 -1320
rect 122950 -1380 123010 -1320
<< metal2 >>
rect 112410 10130 112490 10140
rect 112410 10070 112420 10130
rect 112480 10120 112490 10130
rect 113350 10130 113430 10140
rect 113350 10120 113360 10130
rect 112480 10080 113360 10120
rect 112480 10070 112490 10080
rect 112410 10060 112490 10070
rect 113350 10070 113360 10080
rect 113420 10070 113430 10130
rect 113350 10060 113430 10070
rect 114170 10130 114250 10140
rect 114170 10070 114180 10130
rect 114240 10120 114250 10130
rect 115110 10130 115190 10140
rect 115110 10120 115120 10130
rect 114240 10080 115120 10120
rect 114240 10070 114250 10080
rect 114170 10060 114250 10070
rect 115110 10070 115120 10080
rect 115180 10070 115190 10130
rect 115110 10060 115190 10070
rect 113760 10020 114490 10030
rect 113760 9960 113770 10020
rect 113830 9960 114060 10020
rect 114120 9960 114300 10020
rect 114360 9960 114420 10020
rect 114480 9960 114490 10020
rect 113760 9940 114490 9960
rect 113760 9880 113770 9940
rect 113830 9880 114060 9940
rect 114120 9880 114300 9940
rect 114360 9880 114420 9940
rect 114480 9880 114490 9940
rect 112170 9860 112250 9870
rect 112170 9800 112180 9860
rect 112240 9850 112250 9860
rect 112410 9860 112490 9870
rect 112410 9850 112420 9860
rect 112240 9810 112420 9850
rect 112240 9800 112250 9810
rect 112170 9790 112250 9800
rect 112410 9800 112420 9810
rect 112480 9850 112490 9860
rect 112530 9860 112610 9870
rect 112530 9850 112540 9860
rect 112480 9810 112540 9850
rect 112480 9800 112490 9810
rect 112410 9790 112490 9800
rect 112530 9800 112540 9810
rect 112600 9800 112610 9860
rect 112530 9790 112610 9800
rect 113760 9860 114490 9880
rect 113760 9800 113770 9860
rect 113830 9800 114060 9860
rect 114120 9800 114300 9860
rect 114360 9800 114420 9860
rect 114480 9800 114490 9860
rect 113760 9790 114490 9800
rect 114990 9860 115070 9870
rect 114990 9800 115000 9860
rect 115060 9850 115070 9860
rect 115110 9860 115190 9870
rect 115110 9850 115120 9860
rect 115060 9810 115120 9850
rect 115060 9800 115070 9810
rect 114990 9790 115070 9800
rect 115110 9800 115120 9810
rect 115180 9850 115190 9860
rect 115350 9860 115430 9870
rect 115350 9850 115360 9860
rect 115180 9810 115360 9850
rect 115180 9800 115190 9810
rect 115110 9790 115190 9800
rect 115350 9800 115360 9810
rect 115420 9800 115430 9860
rect 115350 9790 115430 9800
rect 113110 9680 113840 9690
rect 113110 9620 113120 9680
rect 113180 9620 113240 9680
rect 113300 9620 113480 9680
rect 113540 9620 113770 9680
rect 113830 9620 113840 9680
rect 113110 9600 113840 9620
rect 113110 9540 113120 9600
rect 113180 9540 113240 9600
rect 113300 9540 113480 9600
rect 113540 9540 113770 9600
rect 113830 9540 113840 9600
rect 113110 9520 113840 9540
rect 113110 9460 113120 9520
rect 113180 9460 113240 9520
rect 113300 9460 113480 9520
rect 113540 9460 113770 9520
rect 113830 9460 113840 9520
rect 113110 9450 113840 9460
rect 112410 9050 112490 9060
rect 112410 8990 112420 9050
rect 112480 9040 112490 9050
rect 113350 9050 113430 9060
rect 113350 9040 113360 9050
rect 112480 9000 113360 9040
rect 112480 8990 112490 9000
rect 112410 8980 112490 8990
rect 113350 8990 113360 9000
rect 113420 8990 113430 9050
rect 113350 8980 113430 8990
rect 114170 9050 114250 9060
rect 114170 8990 114180 9050
rect 114240 9040 114250 9050
rect 115110 9050 115190 9060
rect 115110 9040 115120 9050
rect 114240 9000 115120 9040
rect 114240 8990 114250 9000
rect 114170 8980 114250 8990
rect 115110 8990 115120 9000
rect 115180 8990 115190 9050
rect 115110 8980 115190 8990
rect 112300 8960 112380 8970
rect 112300 8900 112310 8960
rect 112370 8950 112380 8960
rect 113260 8960 113320 8970
rect 112370 8910 113260 8950
rect 112370 8900 112380 8910
rect 112300 8890 112380 8900
rect 113650 8960 113730 8970
rect 113650 8950 113660 8960
rect 113320 8910 113660 8950
rect 113260 8890 113320 8900
rect 113650 8900 113660 8910
rect 113720 8950 113730 8960
rect 113720 8940 115212 8950
rect 113720 8910 115152 8940
rect 113720 8900 113730 8910
rect 113650 8890 113730 8900
rect 115152 8870 115212 8880
rect 113870 8850 113950 8860
rect 113870 8790 113880 8850
rect 113940 8820 113950 8850
rect 114270 8830 114350 8840
rect 114270 8820 114280 8830
rect 113940 8790 114280 8820
rect 113870 8780 114280 8790
rect 114270 8770 114280 8780
rect 114340 8820 114350 8830
rect 115230 8830 115310 8840
rect 115230 8820 115240 8830
rect 114340 8780 115240 8820
rect 114340 8770 114350 8780
rect 114270 8760 114350 8770
rect 115230 8770 115240 8780
rect 115300 8770 115310 8830
rect 115230 8760 115310 8770
rect 104580 8640 123020 8650
rect 104580 8580 104590 8640
rect 104650 8580 104670 8640
rect 104730 8580 104750 8640
rect 104810 8580 105290 8640
rect 105350 8580 105370 8640
rect 105430 8580 105450 8640
rect 105510 8580 105990 8640
rect 106050 8580 106070 8640
rect 106130 8580 106150 8640
rect 106210 8580 106690 8640
rect 106750 8580 106770 8640
rect 106830 8580 106850 8640
rect 106910 8580 108090 8640
rect 108150 8580 108170 8640
rect 108230 8580 108250 8640
rect 108310 8580 109190 8640
rect 109250 8580 109910 8640
rect 109970 8580 110630 8640
rect 110690 8580 111080 8640
rect 111140 8580 111160 8640
rect 111220 8580 111240 8640
rect 111300 8580 113770 8640
rect 113830 8580 116300 8640
rect 116360 8580 116380 8640
rect 116440 8580 116460 8640
rect 116520 8580 116910 8640
rect 116970 8580 117630 8640
rect 117690 8580 118350 8640
rect 118410 8580 119290 8640
rect 119350 8580 119370 8640
rect 119430 8580 119450 8640
rect 119510 8580 120690 8640
rect 120750 8580 120770 8640
rect 120830 8580 120850 8640
rect 120910 8580 121390 8640
rect 121450 8580 121470 8640
rect 121530 8580 121550 8640
rect 121610 8580 122090 8640
rect 122150 8580 122170 8640
rect 122230 8580 122250 8640
rect 122310 8580 122790 8640
rect 122850 8580 122870 8640
rect 122930 8580 122950 8640
rect 123010 8580 123020 8640
rect 104580 8560 123020 8580
rect 104580 8500 104590 8560
rect 104650 8500 104670 8560
rect 104730 8500 104750 8560
rect 104810 8500 105290 8560
rect 105350 8500 105370 8560
rect 105430 8500 105450 8560
rect 105510 8500 105990 8560
rect 106050 8500 106070 8560
rect 106130 8500 106150 8560
rect 106210 8500 106690 8560
rect 106750 8500 106770 8560
rect 106830 8500 106850 8560
rect 106910 8500 108090 8560
rect 108150 8500 108170 8560
rect 108230 8500 108250 8560
rect 108310 8500 109190 8560
rect 109250 8500 109910 8560
rect 109970 8500 110630 8560
rect 110690 8500 111080 8560
rect 111140 8500 111160 8560
rect 111220 8500 111240 8560
rect 111300 8500 113770 8560
rect 113830 8500 116300 8560
rect 116360 8500 116380 8560
rect 116440 8500 116460 8560
rect 116520 8500 116910 8560
rect 116970 8500 117630 8560
rect 117690 8500 118350 8560
rect 118410 8500 119290 8560
rect 119350 8500 119370 8560
rect 119430 8500 119450 8560
rect 119510 8500 120690 8560
rect 120750 8500 120770 8560
rect 120830 8500 120850 8560
rect 120910 8500 121390 8560
rect 121450 8500 121470 8560
rect 121530 8500 121550 8560
rect 121610 8500 122090 8560
rect 122150 8500 122170 8560
rect 122230 8500 122250 8560
rect 122310 8500 122790 8560
rect 122850 8500 122870 8560
rect 122930 8500 122950 8560
rect 123010 8500 123020 8560
rect 104580 8480 123020 8500
rect 104580 8420 104590 8480
rect 104650 8420 104670 8480
rect 104730 8420 104750 8480
rect 104810 8420 105290 8480
rect 105350 8420 105370 8480
rect 105430 8420 105450 8480
rect 105510 8420 105990 8480
rect 106050 8420 106070 8480
rect 106130 8420 106150 8480
rect 106210 8420 106690 8480
rect 106750 8420 106770 8480
rect 106830 8420 106850 8480
rect 106910 8420 108090 8480
rect 108150 8420 108170 8480
rect 108230 8420 108250 8480
rect 108310 8420 109190 8480
rect 109250 8420 109910 8480
rect 109970 8420 110630 8480
rect 110690 8420 111080 8480
rect 111140 8420 111160 8480
rect 111220 8420 111240 8480
rect 111300 8420 113770 8480
rect 113830 8420 116300 8480
rect 116360 8420 116380 8480
rect 116440 8420 116460 8480
rect 116520 8420 116910 8480
rect 116970 8420 117630 8480
rect 117690 8420 118350 8480
rect 118410 8420 119290 8480
rect 119350 8420 119370 8480
rect 119430 8420 119450 8480
rect 119510 8420 120690 8480
rect 120750 8420 120770 8480
rect 120830 8420 120850 8480
rect 120910 8420 121390 8480
rect 121450 8420 121470 8480
rect 121530 8420 121550 8480
rect 121610 8420 122090 8480
rect 122150 8420 122170 8480
rect 122230 8420 122250 8480
rect 122310 8420 122790 8480
rect 122850 8420 122870 8480
rect 122930 8420 122950 8480
rect 123010 8420 123020 8480
rect 104580 8410 123020 8420
rect 109300 8370 113530 8380
rect 109300 8310 109310 8370
rect 109370 8310 109550 8370
rect 109610 8310 109790 8370
rect 109850 8310 110030 8370
rect 110090 8310 110270 8370
rect 110330 8310 110510 8370
rect 110570 8310 112020 8370
rect 112080 8310 112260 8370
rect 112320 8310 112500 8370
rect 112560 8310 112740 8370
rect 112800 8310 112980 8370
rect 113040 8310 113220 8370
rect 113280 8310 113460 8370
rect 113520 8310 113530 8370
rect 109300 8290 113530 8310
rect 109300 8230 109310 8290
rect 109370 8230 109550 8290
rect 109610 8230 109790 8290
rect 109850 8230 110030 8290
rect 110090 8230 110270 8290
rect 110330 8230 110510 8290
rect 110570 8230 112020 8290
rect 112080 8230 112260 8290
rect 112320 8230 112500 8290
rect 112560 8230 112740 8290
rect 112800 8230 112980 8290
rect 113040 8230 113220 8290
rect 113280 8230 113460 8290
rect 113520 8230 113530 8290
rect 109300 8210 113530 8230
rect 109300 8150 109310 8210
rect 109370 8150 109550 8210
rect 109610 8150 109790 8210
rect 109850 8150 110030 8210
rect 110090 8150 110270 8210
rect 110330 8150 110510 8210
rect 110570 8150 112020 8210
rect 112080 8150 112260 8210
rect 112320 8150 112500 8210
rect 112560 8150 112740 8210
rect 112800 8150 112980 8210
rect 113040 8150 113220 8210
rect 113280 8150 113460 8210
rect 113520 8150 113530 8210
rect 109300 8130 113530 8150
rect 109300 8070 109310 8130
rect 109370 8070 109550 8130
rect 109610 8070 109790 8130
rect 109850 8070 110030 8130
rect 110090 8070 110270 8130
rect 110330 8070 110510 8130
rect 110570 8070 112020 8130
rect 112080 8070 112260 8130
rect 112320 8070 112500 8130
rect 112560 8070 112740 8130
rect 112800 8070 112980 8130
rect 113040 8070 113220 8130
rect 113280 8070 113460 8130
rect 113520 8070 113530 8130
rect 109300 8050 113530 8070
rect 109300 7990 109310 8050
rect 109370 7990 109550 8050
rect 109610 7990 109790 8050
rect 109850 7990 110030 8050
rect 110090 7990 110270 8050
rect 110330 7990 110510 8050
rect 110570 7990 112020 8050
rect 112080 7990 112260 8050
rect 112320 7990 112500 8050
rect 112560 7990 112740 8050
rect 112800 7990 112980 8050
rect 113040 7990 113220 8050
rect 113280 7990 113460 8050
rect 113520 7990 113530 8050
rect 109300 7970 113530 7990
rect 109300 7910 109310 7970
rect 109370 7910 109550 7970
rect 109610 7910 109790 7970
rect 109850 7910 110030 7970
rect 110090 7910 110270 7970
rect 110330 7910 110510 7970
rect 110570 7910 112020 7970
rect 112080 7910 112260 7970
rect 112320 7910 112500 7970
rect 112560 7910 112740 7970
rect 112800 7910 112980 7970
rect 113040 7910 113220 7970
rect 113280 7910 113460 7970
rect 113520 7910 113530 7970
rect 109300 7900 113530 7910
rect 114070 8370 118300 8380
rect 114070 8310 114080 8370
rect 114140 8310 114320 8370
rect 114380 8310 114560 8370
rect 114620 8310 114800 8370
rect 114860 8310 115040 8370
rect 115100 8310 115280 8370
rect 115340 8310 115520 8370
rect 115580 8310 117030 8370
rect 117090 8310 117270 8370
rect 117330 8310 117510 8370
rect 117570 8310 117750 8370
rect 117810 8310 117990 8370
rect 118050 8310 118230 8370
rect 118290 8310 118300 8370
rect 114070 8290 118300 8310
rect 114070 8230 114080 8290
rect 114140 8230 114320 8290
rect 114380 8230 114560 8290
rect 114620 8230 114800 8290
rect 114860 8230 115040 8290
rect 115100 8230 115280 8290
rect 115340 8230 115520 8290
rect 115580 8230 117030 8290
rect 117090 8230 117270 8290
rect 117330 8230 117510 8290
rect 117570 8230 117750 8290
rect 117810 8230 117990 8290
rect 118050 8230 118230 8290
rect 118290 8230 118300 8290
rect 114070 8210 118300 8230
rect 114070 8150 114080 8210
rect 114140 8150 114320 8210
rect 114380 8150 114560 8210
rect 114620 8150 114800 8210
rect 114860 8150 115040 8210
rect 115100 8150 115280 8210
rect 115340 8150 115520 8210
rect 115580 8150 117030 8210
rect 117090 8150 117270 8210
rect 117330 8150 117510 8210
rect 117570 8150 117750 8210
rect 117810 8150 117990 8210
rect 118050 8150 118230 8210
rect 118290 8150 118300 8210
rect 114070 8130 118300 8150
rect 114070 8070 114080 8130
rect 114140 8070 114320 8130
rect 114380 8070 114560 8130
rect 114620 8070 114800 8130
rect 114860 8070 115040 8130
rect 115100 8070 115280 8130
rect 115340 8070 115520 8130
rect 115580 8070 117030 8130
rect 117090 8070 117270 8130
rect 117330 8070 117510 8130
rect 117570 8070 117750 8130
rect 117810 8070 117990 8130
rect 118050 8070 118230 8130
rect 118290 8070 118300 8130
rect 114070 8050 118300 8070
rect 114070 7990 114080 8050
rect 114140 7990 114320 8050
rect 114380 7990 114560 8050
rect 114620 7990 114800 8050
rect 114860 7990 115040 8050
rect 115100 7990 115280 8050
rect 115340 7990 115520 8050
rect 115580 7990 117030 8050
rect 117090 7990 117270 8050
rect 117330 7990 117510 8050
rect 117570 7990 117750 8050
rect 117810 7990 117990 8050
rect 118050 7990 118230 8050
rect 118290 7990 118300 8050
rect 114070 7970 118300 7990
rect 114070 7910 114080 7970
rect 114140 7910 114320 7970
rect 114380 7910 114560 7970
rect 114620 7910 114800 7970
rect 114860 7910 115040 7970
rect 115100 7910 115280 7970
rect 115340 7910 115520 7970
rect 115580 7910 117030 7970
rect 117090 7910 117270 7970
rect 117330 7910 117510 7970
rect 117570 7910 117750 7970
rect 117810 7910 117990 7970
rect 118050 7910 118230 7970
rect 118290 7910 118300 7970
rect 114070 7900 118300 7910
rect 109180 7860 109260 7870
rect 109180 7800 109190 7860
rect 109250 7850 109260 7860
rect 109420 7860 109500 7870
rect 109420 7850 109430 7860
rect 109250 7810 109430 7850
rect 109250 7800 109260 7810
rect 109180 7790 109260 7800
rect 109420 7800 109430 7810
rect 109490 7850 109500 7860
rect 109660 7860 109740 7870
rect 109660 7850 109670 7860
rect 109490 7810 109670 7850
rect 109490 7800 109500 7810
rect 109420 7790 109500 7800
rect 109660 7800 109670 7810
rect 109730 7850 109740 7860
rect 109900 7860 109980 7870
rect 109900 7850 109910 7860
rect 109730 7810 109910 7850
rect 109730 7800 109740 7810
rect 109660 7790 109740 7800
rect 109900 7800 109910 7810
rect 109970 7850 109980 7860
rect 110140 7860 110220 7870
rect 110140 7850 110150 7860
rect 109970 7810 110150 7850
rect 109970 7800 109980 7810
rect 109900 7790 109980 7800
rect 110140 7800 110150 7810
rect 110210 7850 110220 7860
rect 110380 7860 110460 7870
rect 110380 7850 110390 7860
rect 110210 7810 110390 7850
rect 110210 7800 110220 7810
rect 110140 7790 110220 7800
rect 110380 7800 110390 7810
rect 110450 7850 110460 7860
rect 110620 7860 110700 7870
rect 110620 7850 110630 7860
rect 110450 7810 110630 7850
rect 110450 7800 110460 7810
rect 110380 7790 110460 7800
rect 110620 7800 110630 7810
rect 110690 7800 110700 7860
rect 116900 7860 116980 7870
rect 110620 7790 110700 7800
rect 112130 7830 112210 7840
rect 112130 7770 112140 7830
rect 112200 7820 112210 7830
rect 112370 7830 112450 7840
rect 112370 7820 112380 7830
rect 112200 7780 112380 7820
rect 112200 7770 112210 7780
rect 112130 7760 112210 7770
rect 112370 7770 112380 7780
rect 112440 7820 112450 7830
rect 112610 7830 112690 7840
rect 112610 7820 112620 7830
rect 112440 7780 112620 7820
rect 112440 7770 112450 7780
rect 112370 7760 112450 7770
rect 112610 7770 112620 7780
rect 112680 7820 112690 7830
rect 112850 7830 112930 7840
rect 112850 7820 112860 7830
rect 112680 7780 112860 7820
rect 112680 7770 112690 7780
rect 112610 7760 112690 7770
rect 112850 7770 112860 7780
rect 112920 7820 112930 7830
rect 113090 7830 113170 7840
rect 113090 7820 113100 7830
rect 112920 7780 113100 7820
rect 112920 7770 112930 7780
rect 112850 7760 112930 7770
rect 113090 7770 113100 7780
rect 113160 7820 113170 7830
rect 113330 7830 113410 7840
rect 113330 7820 113340 7830
rect 113160 7780 113340 7820
rect 113160 7770 113170 7780
rect 113090 7760 113170 7770
rect 113330 7770 113340 7780
rect 113400 7770 113410 7830
rect 113330 7760 113410 7770
rect 114190 7830 114270 7840
rect 114190 7770 114200 7830
rect 114260 7820 114270 7830
rect 114430 7830 114510 7840
rect 114430 7820 114440 7830
rect 114260 7780 114440 7820
rect 114260 7770 114270 7780
rect 114190 7760 114270 7770
rect 114430 7770 114440 7780
rect 114500 7820 114510 7830
rect 114670 7830 114750 7840
rect 114670 7820 114680 7830
rect 114500 7780 114680 7820
rect 114500 7770 114510 7780
rect 114430 7760 114510 7770
rect 114670 7770 114680 7780
rect 114740 7820 114750 7830
rect 114910 7830 114990 7840
rect 114910 7820 114920 7830
rect 114740 7780 114920 7820
rect 114740 7770 114750 7780
rect 114670 7760 114750 7770
rect 114910 7770 114920 7780
rect 114980 7820 114990 7830
rect 115150 7830 115230 7840
rect 115150 7820 115160 7830
rect 114980 7780 115160 7820
rect 114980 7770 114990 7780
rect 114910 7760 114990 7770
rect 115150 7770 115160 7780
rect 115220 7820 115230 7830
rect 115390 7830 115470 7840
rect 115390 7820 115400 7830
rect 115220 7780 115400 7820
rect 115220 7770 115230 7780
rect 115150 7760 115230 7770
rect 115390 7770 115400 7780
rect 115460 7770 115470 7830
rect 116900 7800 116910 7860
rect 116970 7850 116980 7860
rect 117140 7860 117220 7870
rect 117140 7850 117150 7860
rect 116970 7810 117150 7850
rect 116970 7800 116980 7810
rect 116900 7790 116980 7800
rect 117140 7800 117150 7810
rect 117210 7850 117220 7860
rect 117380 7860 117460 7870
rect 117380 7850 117390 7860
rect 117210 7810 117390 7850
rect 117210 7800 117220 7810
rect 117140 7790 117220 7800
rect 117380 7800 117390 7810
rect 117450 7850 117460 7860
rect 117620 7860 117700 7870
rect 117620 7850 117630 7860
rect 117450 7810 117630 7850
rect 117450 7800 117460 7810
rect 117380 7790 117460 7800
rect 117620 7800 117630 7810
rect 117690 7850 117700 7860
rect 117860 7860 117940 7870
rect 117860 7850 117870 7860
rect 117690 7810 117870 7850
rect 117690 7800 117700 7810
rect 117620 7790 117700 7800
rect 117860 7800 117870 7810
rect 117930 7850 117940 7860
rect 118100 7860 118180 7870
rect 118100 7850 118110 7860
rect 117930 7810 118110 7850
rect 117930 7800 117940 7810
rect 117860 7790 117940 7800
rect 118100 7800 118110 7810
rect 118170 7850 118180 7860
rect 118340 7860 118420 7870
rect 118340 7850 118350 7860
rect 118170 7810 118350 7850
rect 118170 7800 118180 7810
rect 118100 7790 118180 7800
rect 118340 7800 118350 7810
rect 118410 7800 118420 7860
rect 118340 7790 118420 7800
rect 115390 7760 115470 7770
rect 109300 7050 109380 7060
rect 109300 6990 109310 7050
rect 109370 7040 109380 7050
rect 109540 7050 109620 7060
rect 109540 7040 109550 7050
rect 109370 7000 109550 7040
rect 109370 6990 109380 7000
rect 109300 6980 109380 6990
rect 109540 6990 109550 7000
rect 109610 7040 109620 7050
rect 109780 7050 109860 7060
rect 109780 7040 109790 7050
rect 109610 7000 109790 7040
rect 109610 6990 109620 7000
rect 109540 6980 109620 6990
rect 109780 6990 109790 7000
rect 109850 7040 109860 7050
rect 110020 7050 110100 7060
rect 110020 7040 110030 7050
rect 109850 7000 110030 7040
rect 109850 6990 109860 7000
rect 109780 6980 109860 6990
rect 110020 6990 110030 7000
rect 110090 7040 110100 7050
rect 110260 7050 110340 7060
rect 110260 7040 110270 7050
rect 110090 7000 110270 7040
rect 110090 6990 110100 7000
rect 110020 6980 110100 6990
rect 110260 6990 110270 7000
rect 110330 7040 110340 7050
rect 110500 7050 110580 7060
rect 110500 7040 110510 7050
rect 110330 7000 110510 7040
rect 110330 6990 110340 7000
rect 110260 6980 110340 6990
rect 110500 6990 110510 7000
rect 110570 6990 110580 7050
rect 110500 6980 110580 6990
rect 110800 7050 113410 7060
rect 110800 6990 110810 7050
rect 110870 6990 110890 7050
rect 110950 6990 110970 7050
rect 111030 6990 112140 7050
rect 112200 6990 112380 7050
rect 112440 6990 112620 7050
rect 112680 6990 112860 7050
rect 112920 6990 113100 7050
rect 113160 6990 113340 7050
rect 113400 6990 113410 7050
rect 110800 6980 113410 6990
rect 114190 7050 116800 7060
rect 114190 6990 114200 7050
rect 114260 6990 114440 7050
rect 114500 6990 114680 7050
rect 114740 6990 114920 7050
rect 114980 6990 115160 7050
rect 115220 6990 115400 7050
rect 115460 6990 116570 7050
rect 116630 6990 116650 7050
rect 116710 6990 116730 7050
rect 116790 6990 116800 7050
rect 114190 6980 116800 6990
rect 117020 7050 117100 7060
rect 117020 6990 117030 7050
rect 117090 7040 117100 7050
rect 117260 7050 117340 7060
rect 117260 7040 117270 7050
rect 117090 7000 117270 7040
rect 117090 6990 117100 7000
rect 117020 6980 117100 6990
rect 117260 6990 117270 7000
rect 117330 7040 117340 7050
rect 117500 7050 117580 7060
rect 117500 7040 117510 7050
rect 117330 7000 117510 7040
rect 117330 6990 117340 7000
rect 117260 6980 117340 6990
rect 117500 6990 117510 7000
rect 117570 7040 117580 7050
rect 117740 7050 117820 7060
rect 117740 7040 117750 7050
rect 117570 7000 117750 7040
rect 117570 6990 117580 7000
rect 117500 6980 117580 6990
rect 117740 6990 117750 7000
rect 117810 7040 117820 7050
rect 117980 7050 118060 7060
rect 117980 7040 117990 7050
rect 117810 7000 117990 7040
rect 117810 6990 117820 7000
rect 117740 6980 117820 6990
rect 117980 6990 117990 7000
rect 118050 7040 118060 7050
rect 118220 7050 118300 7060
rect 118220 7040 118230 7050
rect 118050 7000 118230 7040
rect 118050 6990 118060 7000
rect 117980 6980 118060 6990
rect 118220 6990 118230 7000
rect 118290 6990 118300 7050
rect 118220 6980 118300 6990
rect 109370 6940 110510 6950
rect 109430 6880 109490 6940
rect 109550 6880 109610 6940
rect 109670 6880 109730 6940
rect 109790 6880 109850 6940
rect 109910 6880 109970 6940
rect 110030 6880 110090 6940
rect 110150 6880 110210 6940
rect 110270 6880 110330 6940
rect 110390 6880 110450 6940
rect 109370 6870 110510 6880
rect 112200 6940 115400 6950
rect 112260 6880 112320 6940
rect 112380 6880 112440 6940
rect 112500 6880 112560 6940
rect 112620 6880 112680 6940
rect 112740 6880 112800 6940
rect 112860 6880 112920 6940
rect 112980 6880 113040 6940
rect 113100 6880 113160 6940
rect 113220 6880 113280 6940
rect 113340 6880 113680 6940
rect 113740 6880 114260 6940
rect 114320 6880 114380 6940
rect 114440 6880 114500 6940
rect 114560 6880 114620 6940
rect 114680 6880 114740 6940
rect 114800 6880 114860 6940
rect 114920 6880 114980 6940
rect 115040 6880 115100 6940
rect 115160 6880 115220 6940
rect 115280 6880 115340 6940
rect 112200 6870 115400 6880
rect 117090 6940 118230 6950
rect 117150 6880 117210 6940
rect 117270 6880 117330 6940
rect 117390 6880 117450 6940
rect 117510 6880 117570 6940
rect 117630 6880 117690 6940
rect 117750 6880 117810 6940
rect 117870 6880 117930 6940
rect 117990 6880 118050 6940
rect 118110 6880 118170 6940
rect 117090 6870 118230 6880
rect 109900 6820 117700 6830
rect 109900 6760 109910 6820
rect 109970 6760 113860 6820
rect 113920 6760 117630 6820
rect 117690 6760 117700 6820
rect 108510 6750 108590 6760
rect 109900 6750 117700 6760
rect 119010 6750 119090 6760
rect 108510 6690 108520 6750
rect 108580 6690 108590 6750
rect 108510 6680 108590 6690
rect 109240 6710 118360 6720
rect 109240 6650 109250 6710
rect 109310 6650 109470 6710
rect 109530 6650 109690 6710
rect 109750 6650 109910 6710
rect 109970 6650 110130 6710
rect 110190 6650 110350 6710
rect 110410 6650 110570 6710
rect 110630 6650 111080 6710
rect 111140 6650 111160 6710
rect 111220 6650 111240 6710
rect 111300 6650 113030 6710
rect 113090 6650 113360 6710
rect 113420 6650 113690 6710
rect 113750 6650 113850 6710
rect 113910 6650 114180 6710
rect 114240 6650 114510 6710
rect 114570 6650 116300 6710
rect 116360 6650 116380 6710
rect 116440 6650 116460 6710
rect 116520 6650 116970 6710
rect 117030 6650 117190 6710
rect 117250 6650 117410 6710
rect 117470 6650 117630 6710
rect 117690 6650 117850 6710
rect 117910 6650 118070 6710
rect 118130 6650 118290 6710
rect 118350 6650 118360 6710
rect 119010 6690 119020 6750
rect 119080 6690 119090 6750
rect 119010 6680 119090 6690
rect 109240 6630 118360 6650
rect 109240 6570 109250 6630
rect 109310 6570 109470 6630
rect 109530 6570 109690 6630
rect 109750 6570 109910 6630
rect 109970 6570 110130 6630
rect 110190 6570 110350 6630
rect 110410 6570 110570 6630
rect 110630 6570 111080 6630
rect 111140 6570 111160 6630
rect 111220 6570 111240 6630
rect 111300 6570 113030 6630
rect 113090 6570 113360 6630
rect 113420 6570 113690 6630
rect 113750 6570 113850 6630
rect 113910 6570 114180 6630
rect 114240 6570 114510 6630
rect 114570 6570 116300 6630
rect 116360 6570 116380 6630
rect 116440 6570 116460 6630
rect 116520 6570 116970 6630
rect 117030 6570 117190 6630
rect 117250 6570 117410 6630
rect 117470 6570 117630 6630
rect 117690 6570 117850 6630
rect 117910 6570 118070 6630
rect 118130 6570 118290 6630
rect 118350 6570 118360 6630
rect 109240 6550 118360 6570
rect 109240 6490 109250 6550
rect 109310 6490 109470 6550
rect 109530 6490 109690 6550
rect 109750 6490 109910 6550
rect 109970 6490 110130 6550
rect 110190 6490 110350 6550
rect 110410 6490 110570 6550
rect 110630 6490 111080 6550
rect 111140 6490 111160 6550
rect 111220 6490 111240 6550
rect 111300 6490 113030 6550
rect 113090 6490 113360 6550
rect 113420 6490 113690 6550
rect 113750 6490 113850 6550
rect 113910 6490 114180 6550
rect 114240 6490 114510 6550
rect 114570 6490 116300 6550
rect 116360 6490 116380 6550
rect 116440 6490 116460 6550
rect 116520 6490 116970 6550
rect 117030 6490 117190 6550
rect 117250 6490 117410 6550
rect 117470 6490 117630 6550
rect 117690 6490 117850 6550
rect 117910 6490 118070 6550
rect 118130 6490 118290 6550
rect 118350 6490 118360 6550
rect 109240 6480 118360 6490
rect 113240 6440 113320 6450
rect 109350 6380 109430 6390
rect 109350 6320 109360 6380
rect 109420 6370 109430 6380
rect 109570 6380 109650 6390
rect 109570 6370 109580 6380
rect 109420 6330 109580 6370
rect 109420 6320 109430 6330
rect 109350 6310 109430 6320
rect 109570 6320 109580 6330
rect 109640 6370 109650 6380
rect 109790 6380 109870 6390
rect 109790 6370 109800 6380
rect 109640 6330 109800 6370
rect 109640 6320 109650 6330
rect 109570 6310 109650 6320
rect 109790 6320 109800 6330
rect 109860 6370 109870 6380
rect 110010 6380 110090 6390
rect 110010 6370 110020 6380
rect 109860 6330 110020 6370
rect 109860 6320 109870 6330
rect 109790 6310 109870 6320
rect 110010 6320 110020 6330
rect 110080 6370 110090 6380
rect 110230 6380 110310 6390
rect 110230 6370 110240 6380
rect 110080 6330 110240 6370
rect 110080 6320 110090 6330
rect 110010 6310 110090 6320
rect 110230 6320 110240 6330
rect 110300 6370 110310 6380
rect 110450 6380 110530 6390
rect 110450 6370 110460 6380
rect 110300 6330 110460 6370
rect 110300 6320 110310 6330
rect 110230 6310 110310 6320
rect 110450 6320 110460 6330
rect 110520 6320 110530 6380
rect 113240 6380 113250 6440
rect 113310 6430 113320 6440
rect 113460 6440 113540 6450
rect 113460 6430 113470 6440
rect 113310 6390 113470 6430
rect 113310 6380 113320 6390
rect 113240 6370 113320 6380
rect 113460 6380 113470 6390
rect 113530 6380 113540 6440
rect 113460 6370 113540 6380
rect 114060 6440 114140 6450
rect 114060 6380 114070 6440
rect 114130 6430 114140 6440
rect 114280 6440 114360 6450
rect 114280 6430 114290 6440
rect 114130 6390 114290 6430
rect 114130 6380 114140 6390
rect 114060 6370 114140 6380
rect 114280 6380 114290 6390
rect 114350 6380 114360 6440
rect 114280 6370 114360 6380
rect 117070 6380 117150 6390
rect 110450 6310 110530 6320
rect 117070 6320 117080 6380
rect 117140 6370 117150 6380
rect 117290 6380 117370 6390
rect 117290 6370 117300 6380
rect 117140 6330 117300 6370
rect 117140 6320 117150 6330
rect 117070 6310 117150 6320
rect 117290 6320 117300 6330
rect 117360 6370 117370 6380
rect 117510 6380 117590 6390
rect 117510 6370 117520 6380
rect 117360 6330 117520 6370
rect 117360 6320 117370 6330
rect 117290 6310 117370 6320
rect 117510 6320 117520 6330
rect 117580 6370 117590 6380
rect 117730 6380 117810 6390
rect 117730 6370 117740 6380
rect 117580 6330 117740 6370
rect 117580 6320 117590 6330
rect 117510 6310 117590 6320
rect 117730 6320 117740 6330
rect 117800 6370 117810 6380
rect 117950 6380 118030 6390
rect 117950 6370 117960 6380
rect 117800 6330 117960 6370
rect 117800 6320 117810 6330
rect 117730 6310 117810 6320
rect 117950 6320 117960 6330
rect 118020 6370 118030 6380
rect 118170 6380 118250 6390
rect 118170 6370 118180 6380
rect 118020 6330 118180 6370
rect 118020 6320 118030 6330
rect 117950 6310 118030 6320
rect 118170 6320 118180 6330
rect 118240 6320 118250 6380
rect 118170 6310 118250 6320
rect 113120 5820 113180 5830
rect 113600 5820 113660 5830
rect 113350 5800 113430 5810
rect 113350 5790 113360 5800
rect 113180 5760 113360 5790
rect 113120 5750 113360 5760
rect 113350 5740 113360 5750
rect 113420 5790 113430 5800
rect 113420 5760 113600 5790
rect 114170 5800 114250 5810
rect 114170 5790 114180 5800
rect 113660 5760 114180 5790
rect 113420 5750 114180 5760
rect 113420 5740 113430 5750
rect 113350 5730 113430 5740
rect 114170 5740 114180 5750
rect 114240 5790 114250 5800
rect 114240 5750 114260 5790
rect 114240 5740 114250 5750
rect 114170 5730 114250 5740
rect 113200 5660 113280 5670
rect 113200 5650 113210 5660
rect 112730 5610 113210 5650
rect 113200 5600 113210 5610
rect 113270 5650 113280 5660
rect 114320 5660 114400 5670
rect 114320 5650 114330 5660
rect 113270 5610 114330 5650
rect 113270 5600 113280 5610
rect 113200 5590 113280 5600
rect 114320 5600 114330 5610
rect 114390 5600 114400 5660
rect 114320 5590 114400 5600
rect 111900 5560 111980 5570
rect 111900 5500 111910 5560
rect 111970 5550 111980 5560
rect 113490 5560 113570 5570
rect 113490 5550 113500 5560
rect 111970 5510 113500 5550
rect 111970 5500 111980 5510
rect 111900 5490 111980 5500
rect 113490 5500 113500 5510
rect 113560 5550 113570 5560
rect 114030 5560 114110 5570
rect 114030 5550 114040 5560
rect 113560 5510 114040 5550
rect 113560 5500 113570 5510
rect 113490 5490 113570 5500
rect 114030 5500 114040 5510
rect 114100 5550 114110 5560
rect 115620 5560 115700 5570
rect 115620 5550 115630 5560
rect 114100 5510 115630 5550
rect 114100 5500 114110 5510
rect 114030 5490 114110 5500
rect 115620 5500 115630 5510
rect 115690 5500 115700 5560
rect 115620 5490 115700 5500
rect 113700 5450 113780 5460
rect 113700 5390 113710 5450
rect 113770 5440 113780 5450
rect 113920 5450 114000 5460
rect 113920 5440 113930 5450
rect 113770 5400 113930 5440
rect 113770 5390 113780 5400
rect 113700 5380 113780 5390
rect 113920 5390 113930 5400
rect 113990 5390 114000 5450
rect 113920 5380 114000 5390
rect 113870 5340 113950 5350
rect 113870 5280 113880 5340
rect 113940 5330 113950 5340
rect 114420 5340 114500 5350
rect 114420 5330 114430 5340
rect 113940 5290 114430 5330
rect 113940 5280 113950 5290
rect 113870 5270 113950 5280
rect 114420 5280 114430 5290
rect 114490 5330 114500 5340
rect 115730 5340 115810 5350
rect 115730 5330 115740 5340
rect 114490 5290 115740 5330
rect 114490 5280 114500 5290
rect 114420 5270 114500 5280
rect 115730 5280 115740 5290
rect 115800 5280 115810 5340
rect 115730 5270 115810 5280
rect 113700 5230 113780 5240
rect 113700 5170 113710 5230
rect 113770 5170 113780 5230
rect 113700 5160 113780 5170
rect 109350 5100 109430 5110
rect 109350 5040 109360 5100
rect 109420 5090 109430 5100
rect 109570 5100 109650 5110
rect 109570 5090 109580 5100
rect 109420 5050 109580 5090
rect 109420 5040 109430 5050
rect 109350 5030 109430 5040
rect 109570 5040 109580 5050
rect 109640 5090 109650 5100
rect 109790 5100 109870 5110
rect 109790 5090 109800 5100
rect 109640 5050 109800 5090
rect 109640 5040 109650 5050
rect 109570 5030 109650 5040
rect 109790 5040 109800 5050
rect 109860 5090 109870 5100
rect 110010 5100 110090 5110
rect 110010 5090 110020 5100
rect 109860 5050 110020 5090
rect 109860 5040 109870 5050
rect 109790 5030 109870 5040
rect 110010 5040 110020 5050
rect 110080 5090 110090 5100
rect 110230 5100 110310 5110
rect 110230 5090 110240 5100
rect 110080 5050 110240 5090
rect 110080 5040 110090 5050
rect 110010 5030 110090 5040
rect 110230 5040 110240 5050
rect 110300 5090 110310 5100
rect 110450 5100 110530 5110
rect 110450 5090 110460 5100
rect 110300 5050 110460 5090
rect 110300 5040 110310 5050
rect 110230 5030 110310 5040
rect 110450 5040 110460 5050
rect 110520 5040 110530 5100
rect 110450 5030 110530 5040
rect 117070 5100 117150 5110
rect 117070 5040 117080 5100
rect 117140 5090 117150 5100
rect 117290 5100 117370 5110
rect 117290 5090 117300 5100
rect 117140 5050 117300 5090
rect 117140 5040 117150 5050
rect 117070 5030 117150 5040
rect 117290 5040 117300 5050
rect 117360 5090 117370 5100
rect 117510 5100 117590 5110
rect 117510 5090 117520 5100
rect 117360 5050 117520 5090
rect 117360 5040 117370 5050
rect 117290 5030 117370 5040
rect 117510 5040 117520 5050
rect 117580 5090 117590 5100
rect 117730 5100 117810 5110
rect 117730 5090 117740 5100
rect 117580 5050 117740 5090
rect 117580 5040 117590 5050
rect 117510 5030 117590 5040
rect 117730 5040 117740 5050
rect 117800 5090 117810 5100
rect 117950 5100 118030 5110
rect 117950 5090 117960 5100
rect 117800 5050 117960 5090
rect 117800 5040 117810 5050
rect 117730 5030 117810 5040
rect 117950 5040 117960 5050
rect 118020 5090 118030 5100
rect 118170 5100 118250 5110
rect 118170 5090 118180 5100
rect 118020 5050 118180 5090
rect 118020 5040 118030 5050
rect 117950 5030 118030 5040
rect 118170 5040 118180 5050
rect 118240 5040 118250 5100
rect 118170 5030 118250 5040
rect 108430 4940 113350 4950
rect 108430 4880 108440 4940
rect 108500 4880 108520 4940
rect 108580 4880 108600 4940
rect 108660 4880 109910 4940
rect 109970 4880 110810 4940
rect 110870 4880 110890 4940
rect 110950 4880 110970 4940
rect 111030 4880 112180 4940
rect 112240 4880 112290 4940
rect 112350 4880 112400 4940
rect 112460 4880 112510 4940
rect 112570 4880 112620 4940
rect 112680 4880 112730 4940
rect 112790 4880 112840 4940
rect 112900 4880 112950 4940
rect 113010 4880 113060 4940
rect 113120 4880 113170 4940
rect 113230 4880 113280 4940
rect 113340 4880 113350 4940
rect 108430 4860 113350 4880
rect 108430 4800 108440 4860
rect 108500 4800 108520 4860
rect 108580 4800 108600 4860
rect 108660 4800 109910 4860
rect 109970 4800 110810 4860
rect 110870 4800 110890 4860
rect 110950 4800 110970 4860
rect 111030 4800 112180 4860
rect 112240 4800 112290 4860
rect 112350 4800 112400 4860
rect 112460 4800 112510 4860
rect 112570 4800 112620 4860
rect 112680 4800 112730 4860
rect 112790 4800 112840 4860
rect 112900 4800 112950 4860
rect 113010 4800 113060 4860
rect 113120 4800 113170 4860
rect 113230 4800 113280 4860
rect 113340 4800 113350 4860
rect 108430 4780 113350 4800
rect 108430 4720 108440 4780
rect 108500 4720 108520 4780
rect 108580 4720 108600 4780
rect 108660 4720 109910 4780
rect 109970 4720 110810 4780
rect 110870 4720 110890 4780
rect 110950 4720 110970 4780
rect 111030 4720 112180 4780
rect 112240 4720 112290 4780
rect 112350 4720 112400 4780
rect 112460 4720 112510 4780
rect 112570 4720 112620 4780
rect 112680 4720 112730 4780
rect 112790 4720 112840 4780
rect 112900 4720 112950 4780
rect 113010 4720 113060 4780
rect 113120 4720 113170 4780
rect 113230 4720 113280 4780
rect 113340 4720 113350 4780
rect 108430 4710 113350 4720
rect 114250 4940 119170 4950
rect 114250 4880 114260 4940
rect 114320 4880 114370 4940
rect 114430 4880 114480 4940
rect 114540 4880 114590 4940
rect 114650 4880 114700 4940
rect 114760 4880 114810 4940
rect 114870 4880 114920 4940
rect 114980 4880 115030 4940
rect 115090 4880 115140 4940
rect 115200 4880 115250 4940
rect 115310 4880 115360 4940
rect 115420 4880 116570 4940
rect 116630 4880 116650 4940
rect 116710 4880 116730 4940
rect 116790 4880 117630 4940
rect 117690 4880 118940 4940
rect 119000 4880 119020 4940
rect 119080 4880 119100 4940
rect 119160 4880 119170 4940
rect 114250 4860 119170 4880
rect 114250 4800 114260 4860
rect 114320 4800 114370 4860
rect 114430 4800 114480 4860
rect 114540 4800 114590 4860
rect 114650 4800 114700 4860
rect 114760 4800 114810 4860
rect 114870 4800 114920 4860
rect 114980 4800 115030 4860
rect 115090 4800 115140 4860
rect 115200 4800 115250 4860
rect 115310 4800 115360 4860
rect 115420 4800 116570 4860
rect 116630 4800 116650 4860
rect 116710 4800 116730 4860
rect 116790 4800 117630 4860
rect 117690 4800 118940 4860
rect 119000 4800 119020 4860
rect 119080 4800 119100 4860
rect 119160 4800 119170 4860
rect 114250 4780 119170 4800
rect 114250 4720 114260 4780
rect 114320 4720 114370 4780
rect 114430 4720 114480 4780
rect 114540 4720 114590 4780
rect 114650 4720 114700 4780
rect 114760 4720 114810 4780
rect 114870 4720 114920 4780
rect 114980 4720 115030 4780
rect 115090 4720 115140 4780
rect 115200 4720 115250 4780
rect 115310 4720 115360 4780
rect 115420 4720 116570 4780
rect 116630 4720 116650 4780
rect 116710 4720 116730 4780
rect 116790 4720 117630 4780
rect 117690 4720 118940 4780
rect 119000 4720 119020 4780
rect 119080 4720 119100 4780
rect 119160 4720 119170 4780
rect 114250 4710 119170 4720
rect 107980 4640 110530 4650
rect 107980 4580 107990 4640
rect 108050 4580 108070 4640
rect 108130 4580 108160 4640
rect 108220 4580 108240 4640
rect 108300 4580 108330 4640
rect 108390 4580 108410 4640
rect 108470 4580 109360 4640
rect 109420 4580 109470 4640
rect 109530 4580 109580 4640
rect 109640 4580 109690 4640
rect 109750 4580 109800 4640
rect 109860 4580 109910 4640
rect 109970 4580 110020 4640
rect 110080 4580 110130 4640
rect 110190 4580 110240 4640
rect 110300 4580 110350 4640
rect 110410 4580 110460 4640
rect 110520 4580 110530 4640
rect 117070 4640 119620 4650
rect 107980 4560 110530 4580
rect 107980 4500 107990 4560
rect 108050 4500 108070 4560
rect 108130 4500 108160 4560
rect 108220 4500 108240 4560
rect 108300 4500 108330 4560
rect 108390 4500 108410 4560
rect 108470 4500 109360 4560
rect 109420 4500 109470 4560
rect 109530 4500 109580 4560
rect 109640 4500 109690 4560
rect 109750 4500 109800 4560
rect 109860 4500 109910 4560
rect 109970 4500 110020 4560
rect 110080 4500 110130 4560
rect 110190 4500 110240 4560
rect 110300 4500 110350 4560
rect 110410 4500 110460 4560
rect 110520 4500 110530 4560
rect 107980 4480 110530 4500
rect 107980 4420 107990 4480
rect 108050 4420 108070 4480
rect 108130 4420 108160 4480
rect 108220 4420 108240 4480
rect 108300 4420 108330 4480
rect 108390 4420 108410 4480
rect 108470 4420 109360 4480
rect 109420 4420 109470 4480
rect 109530 4420 109580 4480
rect 109640 4420 109690 4480
rect 109750 4420 109800 4480
rect 109860 4420 109910 4480
rect 109970 4420 110020 4480
rect 110080 4420 110130 4480
rect 110190 4420 110240 4480
rect 110300 4420 110350 4480
rect 110410 4420 110460 4480
rect 110520 4420 110530 4480
rect 107980 4410 110530 4420
rect 111340 4590 116260 4600
rect 111340 4530 111350 4590
rect 111410 4530 111430 4590
rect 111490 4530 111510 4590
rect 111570 4530 113550 4590
rect 113610 4530 113770 4590
rect 113830 4530 113990 4590
rect 114050 4530 116030 4590
rect 116090 4530 116110 4590
rect 116170 4530 116190 4590
rect 116250 4530 116260 4590
rect 111340 4510 116260 4530
rect 111340 4450 111350 4510
rect 111410 4450 111430 4510
rect 111490 4450 111510 4510
rect 111570 4450 113550 4510
rect 113610 4450 113770 4510
rect 113830 4450 113990 4510
rect 114050 4450 116030 4510
rect 116090 4450 116110 4510
rect 116170 4450 116190 4510
rect 116250 4450 116260 4510
rect 111340 4430 116260 4450
rect 109240 4370 111310 4380
rect 109240 4310 109250 4370
rect 109310 4310 110570 4370
rect 110630 4310 111080 4370
rect 111140 4310 111160 4370
rect 111220 4310 111240 4370
rect 111300 4310 111310 4370
rect 111340 4370 111350 4430
rect 111410 4370 111430 4430
rect 111490 4370 111510 4430
rect 111570 4370 113550 4430
rect 113610 4370 113770 4430
rect 113830 4370 113990 4430
rect 114050 4370 116030 4430
rect 116090 4370 116110 4430
rect 116170 4370 116190 4430
rect 116250 4370 116260 4430
rect 117070 4580 117080 4640
rect 117140 4580 117190 4640
rect 117250 4580 117300 4640
rect 117360 4580 117410 4640
rect 117470 4580 117520 4640
rect 117580 4580 117630 4640
rect 117690 4580 117740 4640
rect 117800 4580 117850 4640
rect 117910 4580 117960 4640
rect 118020 4580 118070 4640
rect 118130 4580 118180 4640
rect 118240 4580 119130 4640
rect 119190 4580 119210 4640
rect 119270 4580 119300 4640
rect 119360 4580 119380 4640
rect 119440 4580 119470 4640
rect 119530 4580 119550 4640
rect 119610 4580 119620 4640
rect 117070 4560 119620 4580
rect 117070 4500 117080 4560
rect 117140 4500 117190 4560
rect 117250 4500 117300 4560
rect 117360 4500 117410 4560
rect 117470 4500 117520 4560
rect 117580 4500 117630 4560
rect 117690 4500 117740 4560
rect 117800 4500 117850 4560
rect 117910 4500 117960 4560
rect 118020 4500 118070 4560
rect 118130 4500 118180 4560
rect 118240 4500 119130 4560
rect 119190 4500 119210 4560
rect 119270 4500 119300 4560
rect 119360 4500 119380 4560
rect 119440 4500 119470 4560
rect 119530 4500 119550 4560
rect 119610 4500 119620 4560
rect 117070 4480 119620 4500
rect 117070 4420 117080 4480
rect 117140 4420 117190 4480
rect 117250 4420 117300 4480
rect 117360 4420 117410 4480
rect 117470 4420 117520 4480
rect 117580 4420 117630 4480
rect 117690 4420 117740 4480
rect 117800 4420 117850 4480
rect 117910 4420 117960 4480
rect 118020 4420 118070 4480
rect 118130 4420 118180 4480
rect 118240 4420 119130 4480
rect 119190 4420 119210 4480
rect 119270 4420 119300 4480
rect 119360 4420 119380 4480
rect 119440 4420 119470 4480
rect 119530 4420 119550 4480
rect 119610 4420 119620 4480
rect 117070 4410 119620 4420
rect 111340 4360 116260 4370
rect 116290 4370 118360 4380
rect 109240 4290 111310 4310
rect 109240 4230 109250 4290
rect 109310 4230 110570 4290
rect 110630 4230 111080 4290
rect 111140 4230 111160 4290
rect 111220 4230 111240 4290
rect 111300 4230 111310 4290
rect 109240 4210 111310 4230
rect 109240 4150 109250 4210
rect 109310 4150 110570 4210
rect 110630 4150 111080 4210
rect 111140 4150 111160 4210
rect 111220 4150 111240 4210
rect 111300 4150 111310 4210
rect 109240 4140 111310 4150
rect 116290 4310 116300 4370
rect 116360 4310 116380 4370
rect 116440 4310 116460 4370
rect 116520 4310 116970 4370
rect 117030 4310 118290 4370
rect 118350 4310 118360 4370
rect 116290 4290 118360 4310
rect 116290 4230 116300 4290
rect 116360 4230 116380 4290
rect 116440 4230 116460 4290
rect 116520 4230 116970 4290
rect 117030 4230 118290 4290
rect 118350 4230 118360 4290
rect 116290 4210 118360 4230
rect 116290 4150 116300 4210
rect 116360 4150 116380 4210
rect 116440 4150 116460 4210
rect 116520 4150 116970 4210
rect 117030 4150 118290 4210
rect 118350 4150 118360 4210
rect 116290 4140 118360 4150
rect 107680 4100 110530 4110
rect 107680 4040 107690 4100
rect 107750 4040 107770 4100
rect 107830 4040 107850 4100
rect 107910 4040 109360 4100
rect 109420 4040 109580 4100
rect 109640 4040 109800 4100
rect 109860 4040 110020 4100
rect 110080 4040 110240 4100
rect 110300 4040 110460 4100
rect 110520 4040 110530 4100
rect 107680 4020 110530 4040
rect 107680 3960 107690 4020
rect 107750 3960 107770 4020
rect 107830 3960 107850 4020
rect 107910 3960 109360 4020
rect 109420 3960 109580 4020
rect 109640 3960 109800 4020
rect 109860 3960 110020 4020
rect 110080 3960 110240 4020
rect 110300 3960 110460 4020
rect 110520 3960 110530 4020
rect 107680 3940 110530 3960
rect 107680 3880 107690 3940
rect 107750 3880 107770 3940
rect 107830 3880 107850 3940
rect 107910 3880 109360 3940
rect 109420 3880 109580 3940
rect 109640 3880 109800 3940
rect 109860 3880 110020 3940
rect 110080 3880 110240 3940
rect 110300 3880 110460 3940
rect 110520 3880 110530 3940
rect 107680 3870 110530 3880
rect 111340 4100 111580 4110
rect 111340 4040 111350 4100
rect 111410 4040 111430 4100
rect 111490 4040 111510 4100
rect 111570 4040 111580 4100
rect 111340 4020 111580 4040
rect 116020 4100 119920 4110
rect 116020 4040 116030 4100
rect 116090 4040 116110 4100
rect 116170 4040 116190 4100
rect 116250 4040 117080 4100
rect 117140 4040 117300 4100
rect 117360 4040 117520 4100
rect 117580 4040 117740 4100
rect 117800 4040 117960 4100
rect 118020 4040 118180 4100
rect 118240 4040 119690 4100
rect 119750 4040 119770 4100
rect 119830 4040 119850 4100
rect 119910 4040 119920 4100
rect 111340 3960 111350 4020
rect 111410 3960 111430 4020
rect 111490 3960 111510 4020
rect 111570 3960 111580 4020
rect 111340 3940 111580 3960
rect 112170 4020 113650 4030
rect 112170 3960 112180 4020
rect 112240 3960 112400 4020
rect 112460 3960 112620 4020
rect 112680 3960 112840 4020
rect 112900 3960 113060 4020
rect 113120 3960 113280 4020
rect 113340 3960 113580 4020
rect 113640 3960 113650 4020
rect 112170 3950 113650 3960
rect 113950 4020 115430 4030
rect 113950 3960 113960 4020
rect 114020 3960 114260 4020
rect 114320 3960 114480 4020
rect 114540 3960 114700 4020
rect 114760 3960 114920 4020
rect 114980 3960 115140 4020
rect 115200 3960 115360 4020
rect 115420 3960 115430 4020
rect 113950 3950 115430 3960
rect 116020 4020 119920 4040
rect 116020 3960 116030 4020
rect 116090 3960 116110 4020
rect 116170 3960 116190 4020
rect 116250 3960 117080 4020
rect 117140 3960 117300 4020
rect 117360 3960 117520 4020
rect 117580 3960 117740 4020
rect 117800 3960 117960 4020
rect 118020 3960 118180 4020
rect 118240 3960 119690 4020
rect 119750 3960 119770 4020
rect 119830 3960 119850 4020
rect 119910 3960 119920 4020
rect 111340 3880 111350 3940
rect 111410 3880 111430 3940
rect 111490 3880 111510 3940
rect 111570 3880 111580 3940
rect 116020 3940 119920 3960
rect 111340 3870 111580 3880
rect 111690 3910 115368 3920
rect 109250 3860 109310 3870
rect 111690 3850 111700 3910
rect 111760 3850 111780 3910
rect 111840 3850 112238 3910
rect 112292 3850 112348 3910
rect 112402 3850 112458 3910
rect 112512 3850 112568 3910
rect 112622 3850 112678 3910
rect 112732 3850 112788 3910
rect 112842 3850 112898 3910
rect 112952 3850 113008 3910
rect 113062 3850 113118 3910
rect 113172 3850 113228 3910
rect 113282 3850 114318 3910
rect 114372 3850 114428 3910
rect 114482 3850 114538 3910
rect 114592 3850 114648 3910
rect 114702 3850 114758 3910
rect 114812 3850 114868 3910
rect 114922 3850 114978 3910
rect 115032 3850 115088 3910
rect 115142 3850 115198 3910
rect 115252 3850 115308 3910
rect 115362 3850 115368 3910
rect 116020 3880 116030 3940
rect 116090 3880 116110 3940
rect 116170 3880 116190 3940
rect 116250 3880 117080 3940
rect 117140 3880 117300 3940
rect 117360 3880 117520 3940
rect 117580 3880 117740 3940
rect 117800 3880 117960 3940
rect 118020 3880 118180 3940
rect 118240 3880 119690 3940
rect 119750 3880 119770 3940
rect 119830 3880 119850 3940
rect 119910 3880 119920 3940
rect 116020 3870 119920 3880
rect 116970 3860 117030 3870
rect 118290 3860 118350 3870
rect 111690 3840 115368 3850
rect 109460 3830 109540 3840
rect 109460 3770 109470 3830
rect 109530 3820 109540 3830
rect 109680 3830 109760 3840
rect 109680 3820 109690 3830
rect 109530 3780 109690 3820
rect 109530 3770 109540 3780
rect 109460 3760 109540 3770
rect 109680 3770 109690 3780
rect 109750 3820 109760 3830
rect 109900 3830 109980 3840
rect 109900 3820 109910 3830
rect 109750 3780 109910 3820
rect 109750 3770 109760 3780
rect 109680 3760 109760 3770
rect 109900 3770 109910 3780
rect 109970 3820 109980 3830
rect 110120 3830 110200 3840
rect 110120 3820 110130 3830
rect 109970 3780 110130 3820
rect 109970 3770 109980 3780
rect 109900 3760 109980 3770
rect 110120 3770 110130 3780
rect 110190 3820 110200 3830
rect 110340 3830 110420 3840
rect 110340 3820 110350 3830
rect 110190 3780 110350 3820
rect 110190 3770 110200 3780
rect 110120 3760 110200 3770
rect 110340 3770 110350 3780
rect 110410 3770 110420 3830
rect 110340 3760 110420 3770
rect 117180 3830 117260 3840
rect 117180 3770 117190 3830
rect 117250 3820 117260 3830
rect 117400 3830 117480 3840
rect 117400 3820 117410 3830
rect 117250 3780 117410 3820
rect 117250 3770 117260 3780
rect 117180 3760 117260 3770
rect 117400 3770 117410 3780
rect 117470 3820 117480 3830
rect 117620 3830 117700 3840
rect 117620 3820 117630 3830
rect 117470 3780 117630 3820
rect 117470 3770 117480 3780
rect 117400 3760 117480 3770
rect 117620 3770 117630 3780
rect 117690 3820 117700 3830
rect 117840 3830 117920 3840
rect 117840 3820 117850 3830
rect 117690 3780 117850 3820
rect 117690 3770 117700 3780
rect 117620 3760 117700 3770
rect 117840 3770 117850 3780
rect 117910 3820 117920 3830
rect 118060 3830 118140 3840
rect 118060 3820 118070 3830
rect 117910 3780 118070 3820
rect 117910 3770 117920 3780
rect 117840 3760 117920 3770
rect 118060 3770 118070 3780
rect 118130 3770 118140 3830
rect 118060 3760 118140 3770
rect 112280 3500 112360 3510
rect 112280 3440 112290 3500
rect 112350 3490 112360 3500
rect 112500 3500 112580 3510
rect 112500 3490 112510 3500
rect 112350 3450 112510 3490
rect 112350 3440 112360 3450
rect 107980 3420 108480 3440
rect 112280 3430 112360 3440
rect 112500 3440 112510 3450
rect 112570 3490 112580 3500
rect 112720 3500 112800 3510
rect 112720 3490 112730 3500
rect 112570 3450 112730 3490
rect 112570 3440 112580 3450
rect 112500 3430 112580 3440
rect 112720 3440 112730 3450
rect 112790 3490 112800 3500
rect 112940 3500 113020 3510
rect 112940 3490 112950 3500
rect 112790 3450 112950 3490
rect 112790 3440 112800 3450
rect 112720 3430 112800 3440
rect 112940 3440 112950 3450
rect 113010 3490 113020 3500
rect 113160 3500 113240 3510
rect 113160 3490 113170 3500
rect 113010 3450 113170 3490
rect 113010 3440 113020 3450
rect 112940 3430 113020 3440
rect 113160 3440 113170 3450
rect 113230 3440 113240 3500
rect 113160 3430 113240 3440
rect 114360 3500 114440 3510
rect 114360 3440 114370 3500
rect 114430 3490 114440 3500
rect 114580 3500 114660 3510
rect 114580 3490 114590 3500
rect 114430 3450 114590 3490
rect 114430 3440 114440 3450
rect 114360 3430 114440 3440
rect 114580 3440 114590 3450
rect 114650 3490 114660 3500
rect 114800 3500 114880 3510
rect 114800 3490 114810 3500
rect 114650 3450 114810 3490
rect 114650 3440 114660 3450
rect 114580 3430 114660 3440
rect 114800 3440 114810 3450
rect 114870 3490 114880 3500
rect 115020 3500 115100 3510
rect 115020 3490 115030 3500
rect 114870 3450 115030 3490
rect 114870 3440 114880 3450
rect 114800 3430 114880 3440
rect 115020 3440 115030 3450
rect 115090 3490 115100 3500
rect 115240 3500 115320 3510
rect 115240 3490 115250 3500
rect 115090 3450 115250 3490
rect 115090 3440 115100 3450
rect 115020 3430 115100 3440
rect 115240 3440 115250 3450
rect 115310 3440 115320 3500
rect 115240 3430 115320 3440
rect 107980 3360 108000 3420
rect 108060 3360 108100 3420
rect 108160 3360 108200 3420
rect 108260 3360 108300 3420
rect 108360 3360 108400 3420
rect 108460 3360 108480 3420
rect 119120 3420 119620 3440
rect 107980 3320 108480 3360
rect 112170 3390 113650 3400
rect 112170 3330 112180 3390
rect 112240 3330 112400 3390
rect 112460 3330 112620 3390
rect 112680 3330 112840 3390
rect 112900 3330 113060 3390
rect 113120 3330 113280 3390
rect 113340 3330 113580 3390
rect 113640 3330 113650 3390
rect 107980 3260 108000 3320
rect 108060 3260 108100 3320
rect 108160 3260 108200 3320
rect 108260 3260 108300 3320
rect 108360 3260 108400 3320
rect 108460 3260 108480 3320
rect 107980 3220 108480 3260
rect 108970 3320 109050 3330
rect 108970 3260 108980 3320
rect 109040 3310 109050 3320
rect 109460 3320 109540 3330
rect 109460 3310 109470 3320
rect 109040 3270 109470 3310
rect 109040 3260 109050 3270
rect 108970 3250 109050 3260
rect 109460 3260 109470 3270
rect 109530 3310 109540 3320
rect 109680 3320 109760 3330
rect 109680 3310 109690 3320
rect 109530 3270 109690 3310
rect 109530 3260 109540 3270
rect 109460 3250 109540 3260
rect 109680 3260 109690 3270
rect 109750 3310 109760 3320
rect 109900 3320 109980 3330
rect 109900 3310 109910 3320
rect 109750 3270 109910 3310
rect 109750 3260 109760 3270
rect 109680 3250 109760 3260
rect 109900 3260 109910 3270
rect 109970 3310 109980 3320
rect 110120 3320 110200 3330
rect 110120 3310 110130 3320
rect 109970 3270 110130 3310
rect 109970 3260 109980 3270
rect 109900 3250 109980 3260
rect 110120 3260 110130 3270
rect 110190 3310 110200 3320
rect 110340 3320 110420 3330
rect 112170 3320 113650 3330
rect 113950 3390 115430 3400
rect 113950 3330 113960 3390
rect 114020 3330 114260 3390
rect 114320 3330 114480 3390
rect 114540 3330 114700 3390
rect 114760 3330 114920 3390
rect 114980 3330 115140 3390
rect 115200 3330 115360 3390
rect 115420 3330 115430 3390
rect 119120 3360 119140 3420
rect 119200 3360 119240 3420
rect 119300 3360 119340 3420
rect 119400 3360 119440 3420
rect 119500 3360 119540 3420
rect 119600 3360 119620 3420
rect 113950 3320 115430 3330
rect 117180 3320 117260 3330
rect 110340 3310 110350 3320
rect 110190 3270 110350 3310
rect 110190 3260 110200 3270
rect 110120 3250 110200 3260
rect 110340 3260 110350 3270
rect 110410 3260 110420 3320
rect 110340 3250 110420 3260
rect 111340 3280 116260 3290
rect 107980 3160 108000 3220
rect 108060 3160 108100 3220
rect 108160 3160 108200 3220
rect 108260 3160 108300 3220
rect 108360 3160 108400 3220
rect 108460 3160 108480 3220
rect 111340 3220 111350 3280
rect 111410 3220 111430 3280
rect 111490 3220 111510 3280
rect 111570 3220 112070 3280
rect 112130 3220 113390 3280
rect 113450 3220 114150 3280
rect 114210 3220 115470 3280
rect 115530 3220 116030 3280
rect 116090 3220 116110 3280
rect 116170 3220 116190 3280
rect 116250 3220 116260 3280
rect 117180 3260 117190 3320
rect 117250 3310 117260 3320
rect 117400 3320 117480 3330
rect 117400 3310 117410 3320
rect 117250 3270 117410 3310
rect 117250 3260 117260 3270
rect 117180 3250 117260 3260
rect 117400 3260 117410 3270
rect 117470 3310 117480 3320
rect 117620 3320 117700 3330
rect 117620 3310 117630 3320
rect 117470 3270 117630 3310
rect 117470 3260 117480 3270
rect 117400 3250 117480 3260
rect 117620 3260 117630 3270
rect 117690 3310 117700 3320
rect 117840 3320 117920 3330
rect 117840 3310 117850 3320
rect 117690 3270 117850 3310
rect 117690 3260 117700 3270
rect 117620 3250 117700 3260
rect 117840 3260 117850 3270
rect 117910 3310 117920 3320
rect 118060 3320 118140 3330
rect 118060 3310 118070 3320
rect 117910 3270 118070 3310
rect 117910 3260 117920 3270
rect 117840 3250 117920 3260
rect 118060 3260 118070 3270
rect 118130 3310 118140 3320
rect 118550 3320 118630 3330
rect 118550 3310 118560 3320
rect 118130 3270 118560 3310
rect 118130 3260 118140 3270
rect 118060 3250 118140 3260
rect 118550 3260 118560 3270
rect 118620 3260 118630 3320
rect 118550 3250 118630 3260
rect 119120 3320 119620 3360
rect 119120 3260 119140 3320
rect 119200 3260 119240 3320
rect 119300 3260 119340 3320
rect 119400 3260 119440 3320
rect 119500 3260 119540 3320
rect 119600 3260 119620 3320
rect 111340 3200 116260 3220
rect 119120 3220 119620 3260
rect 107980 3140 108480 3160
rect 110230 3190 111040 3200
rect 110230 3130 110240 3190
rect 110300 3130 110810 3190
rect 110870 3130 110890 3190
rect 110950 3130 110970 3190
rect 111030 3130 111040 3190
rect 110230 3110 111040 3130
rect 110230 3050 110240 3110
rect 110300 3050 110810 3110
rect 110870 3050 110890 3110
rect 110950 3050 110970 3110
rect 111030 3050 111040 3110
rect 111340 3140 111350 3200
rect 111410 3140 111430 3200
rect 111490 3140 111510 3200
rect 111570 3140 112070 3200
rect 112130 3140 113390 3200
rect 113450 3140 114150 3200
rect 114210 3140 115470 3200
rect 115530 3140 116030 3200
rect 116090 3140 116110 3200
rect 116170 3140 116190 3200
rect 116250 3140 116260 3200
rect 111340 3120 116260 3140
rect 111340 3060 111350 3120
rect 111410 3060 111430 3120
rect 111490 3060 111510 3120
rect 111570 3060 112070 3120
rect 112130 3060 113390 3120
rect 113450 3060 114150 3120
rect 114210 3060 115470 3120
rect 115530 3060 116030 3120
rect 116090 3060 116110 3120
rect 116170 3060 116190 3120
rect 116250 3060 116260 3120
rect 111340 3050 116260 3060
rect 116560 3190 117370 3200
rect 116560 3130 116570 3190
rect 116630 3130 116650 3190
rect 116710 3130 116730 3190
rect 116790 3130 117300 3190
rect 117360 3130 117370 3190
rect 119120 3160 119140 3220
rect 119200 3160 119240 3220
rect 119300 3160 119340 3220
rect 119400 3160 119440 3220
rect 119500 3160 119540 3220
rect 119600 3160 119620 3220
rect 119120 3140 119620 3160
rect 116560 3110 117370 3130
rect 116560 3050 116570 3110
rect 116630 3050 116650 3110
rect 116710 3050 116730 3110
rect 116790 3050 117300 3110
rect 117360 3050 117370 3110
rect 110230 3040 111040 3050
rect 116560 3040 117370 3050
rect 111340 2970 116260 2980
rect 109060 2950 109140 2960
rect 109060 2890 109070 2950
rect 109130 2940 109140 2950
rect 109460 2950 109540 2960
rect 109460 2940 109470 2950
rect 109130 2900 109470 2940
rect 109130 2890 109140 2900
rect 109060 2880 109140 2890
rect 109460 2890 109470 2900
rect 109530 2940 109540 2950
rect 109680 2950 109760 2960
rect 109680 2940 109690 2950
rect 109530 2900 109690 2940
rect 109530 2890 109540 2900
rect 109460 2880 109540 2890
rect 109680 2890 109690 2900
rect 109750 2940 109760 2950
rect 109900 2950 109980 2960
rect 109900 2940 109910 2950
rect 109750 2900 109910 2940
rect 109750 2890 109760 2900
rect 109680 2880 109760 2890
rect 109900 2890 109910 2900
rect 109970 2940 109980 2950
rect 110120 2950 110200 2960
rect 110120 2940 110130 2950
rect 109970 2900 110130 2940
rect 109970 2890 109980 2900
rect 109900 2880 109980 2890
rect 110120 2890 110130 2900
rect 110190 2940 110200 2950
rect 110340 2950 110420 2960
rect 110340 2940 110350 2950
rect 110190 2900 110350 2940
rect 110190 2890 110200 2900
rect 110120 2880 110200 2890
rect 110340 2890 110350 2900
rect 110410 2890 110420 2950
rect 110340 2880 110420 2890
rect 111340 2910 111350 2970
rect 111410 2910 111430 2970
rect 111490 2910 111510 2970
rect 111570 2910 113770 2970
rect 113830 2910 116030 2970
rect 116090 2910 116110 2970
rect 116170 2910 116190 2970
rect 116250 2910 116260 2970
rect 111340 2890 116260 2910
rect 111340 2830 111350 2890
rect 111410 2830 111430 2890
rect 111490 2830 111510 2890
rect 111570 2830 113770 2890
rect 113830 2830 116030 2890
rect 116090 2830 116110 2890
rect 116170 2830 116190 2890
rect 116250 2830 116260 2890
rect 117180 2950 117260 2960
rect 117180 2890 117190 2950
rect 117250 2940 117260 2950
rect 117400 2950 117480 2960
rect 117400 2940 117410 2950
rect 117250 2900 117410 2940
rect 117250 2890 117260 2900
rect 117180 2880 117260 2890
rect 117400 2890 117410 2900
rect 117470 2940 117480 2950
rect 117620 2950 117700 2960
rect 117620 2940 117630 2950
rect 117470 2900 117630 2940
rect 117470 2890 117480 2900
rect 117400 2880 117480 2890
rect 117620 2890 117630 2900
rect 117690 2940 117700 2950
rect 117840 2950 117920 2960
rect 117840 2940 117850 2950
rect 117690 2900 117850 2940
rect 117690 2890 117700 2900
rect 117620 2880 117700 2890
rect 117840 2890 117850 2900
rect 117910 2940 117920 2950
rect 118060 2950 118140 2960
rect 118060 2940 118070 2950
rect 117910 2900 118070 2940
rect 117910 2890 117920 2900
rect 117840 2880 117920 2890
rect 118060 2890 118070 2900
rect 118130 2940 118140 2950
rect 118460 2950 118540 2960
rect 118460 2940 118470 2950
rect 118130 2900 118470 2940
rect 118130 2890 118140 2900
rect 118060 2880 118140 2890
rect 118460 2890 118470 2900
rect 118530 2890 118540 2950
rect 118460 2880 118540 2890
rect 111340 2810 116260 2830
rect 111340 2750 111350 2810
rect 111410 2750 111430 2810
rect 111490 2750 111510 2810
rect 111570 2750 113770 2810
rect 113830 2750 116030 2810
rect 116090 2750 116110 2810
rect 116170 2750 116190 2810
rect 116250 2750 116260 2810
rect 111340 2740 116260 2750
rect 112290 2630 112350 2640
rect 112170 2610 112250 2620
rect 112080 2590 112140 2600
rect 112060 2540 112080 2580
rect 112170 2550 112180 2610
rect 112240 2600 112250 2610
rect 112240 2570 112290 2600
rect 112510 2630 112570 2640
rect 112390 2610 112470 2620
rect 112390 2600 112400 2610
rect 112350 2570 112400 2600
rect 112240 2560 112400 2570
rect 112240 2550 112250 2560
rect 112170 2540 112250 2550
rect 112390 2550 112400 2560
rect 112460 2600 112470 2610
rect 112460 2570 112510 2600
rect 112730 2630 112790 2640
rect 112610 2610 112690 2620
rect 112610 2600 112620 2610
rect 112570 2570 112620 2600
rect 112460 2560 112620 2570
rect 112460 2550 112470 2560
rect 112390 2540 112470 2550
rect 112610 2550 112620 2560
rect 112680 2600 112690 2610
rect 112680 2570 112730 2600
rect 112950 2630 113010 2640
rect 112830 2610 112910 2620
rect 112830 2600 112840 2610
rect 112790 2570 112840 2600
rect 112680 2560 112840 2570
rect 112680 2550 112690 2560
rect 112610 2540 112690 2550
rect 112830 2550 112840 2560
rect 112900 2600 112910 2610
rect 112900 2570 112950 2600
rect 113170 2630 113230 2640
rect 113050 2610 113130 2620
rect 113050 2600 113060 2610
rect 113010 2570 113060 2600
rect 112900 2560 113060 2570
rect 112900 2550 112910 2560
rect 112830 2540 112910 2550
rect 113050 2550 113060 2560
rect 113120 2600 113130 2610
rect 113120 2570 113170 2600
rect 114370 2630 114430 2640
rect 113270 2610 113350 2620
rect 113270 2600 113280 2610
rect 113230 2570 113280 2600
rect 113120 2560 113280 2570
rect 113120 2550 113130 2560
rect 113050 2540 113130 2550
rect 113270 2550 113280 2560
rect 113340 2550 113350 2610
rect 113270 2540 113350 2550
rect 113380 2610 113440 2620
rect 113680 2610 113740 2620
rect 113440 2560 113680 2600
rect 113380 2540 113440 2550
rect 113680 2540 113740 2550
rect 113860 2610 113920 2620
rect 114160 2610 114220 2620
rect 113920 2560 114160 2600
rect 113860 2540 113920 2550
rect 114160 2540 114220 2550
rect 114250 2610 114330 2620
rect 114250 2550 114260 2610
rect 114320 2600 114330 2610
rect 114320 2570 114370 2600
rect 114590 2630 114650 2640
rect 114470 2610 114550 2620
rect 114470 2600 114480 2610
rect 114430 2570 114480 2600
rect 114320 2560 114480 2570
rect 114320 2550 114330 2560
rect 114250 2540 114330 2550
rect 114470 2550 114480 2560
rect 114540 2600 114550 2610
rect 114540 2570 114590 2600
rect 114810 2630 114870 2640
rect 114690 2610 114770 2620
rect 114690 2600 114700 2610
rect 114650 2570 114700 2600
rect 114540 2560 114700 2570
rect 114540 2550 114550 2560
rect 114470 2540 114550 2550
rect 114690 2550 114700 2560
rect 114760 2600 114770 2610
rect 114760 2570 114810 2600
rect 115030 2630 115090 2640
rect 114910 2610 114990 2620
rect 114910 2600 114920 2610
rect 114870 2570 114920 2600
rect 114760 2560 114920 2570
rect 114760 2550 114770 2560
rect 114690 2540 114770 2550
rect 114910 2550 114920 2560
rect 114980 2600 114990 2610
rect 114980 2570 115030 2600
rect 115250 2630 115310 2640
rect 115130 2610 115210 2620
rect 115130 2600 115140 2610
rect 115090 2570 115140 2600
rect 114980 2560 115140 2570
rect 114980 2550 114990 2560
rect 114910 2540 114990 2550
rect 115130 2550 115140 2560
rect 115200 2600 115210 2610
rect 115200 2570 115250 2600
rect 115350 2610 115430 2620
rect 115350 2600 115360 2610
rect 115310 2570 115360 2600
rect 115200 2560 115360 2570
rect 115200 2550 115210 2560
rect 115130 2540 115210 2550
rect 115350 2550 115360 2560
rect 115420 2550 115430 2610
rect 115350 2540 115430 2550
rect 115460 2590 115520 2600
rect 115520 2540 115540 2580
rect 112080 2520 112140 2530
rect 112280 2520 112360 2530
rect 112280 2460 112290 2520
rect 112350 2510 112360 2520
rect 112500 2520 112580 2530
rect 112500 2510 112510 2520
rect 112350 2470 112510 2510
rect 112350 2460 112360 2470
rect 112280 2450 112360 2460
rect 112500 2460 112510 2470
rect 112570 2510 112580 2520
rect 112720 2520 112800 2530
rect 112720 2510 112730 2520
rect 112570 2470 112730 2510
rect 112570 2460 112580 2470
rect 112500 2450 112580 2460
rect 112720 2460 112730 2470
rect 112790 2510 112800 2520
rect 112940 2520 113020 2530
rect 112940 2510 112950 2520
rect 112790 2470 112950 2510
rect 112790 2460 112800 2470
rect 112720 2450 112800 2460
rect 112940 2460 112950 2470
rect 113010 2510 113020 2520
rect 113160 2520 113240 2530
rect 113160 2510 113170 2520
rect 113010 2470 113170 2510
rect 113010 2460 113020 2470
rect 112940 2450 113020 2460
rect 113160 2460 113170 2470
rect 113230 2510 113240 2520
rect 114360 2520 114440 2530
rect 114360 2510 114370 2520
rect 113230 2470 114370 2510
rect 113230 2460 113240 2470
rect 113160 2450 113240 2460
rect 114360 2460 114370 2470
rect 114430 2510 114440 2520
rect 114580 2520 114660 2530
rect 114580 2510 114590 2520
rect 114430 2470 114590 2510
rect 114430 2460 114440 2470
rect 114360 2450 114440 2460
rect 114580 2460 114590 2470
rect 114650 2510 114660 2520
rect 114800 2520 114880 2530
rect 114800 2510 114810 2520
rect 114650 2470 114810 2510
rect 114650 2460 114660 2470
rect 114580 2450 114660 2460
rect 114800 2460 114810 2470
rect 114870 2510 114880 2520
rect 115020 2520 115100 2530
rect 115020 2510 115030 2520
rect 114870 2470 115030 2510
rect 114870 2460 114880 2470
rect 114800 2450 114880 2460
rect 115020 2460 115030 2470
rect 115090 2510 115100 2520
rect 115240 2520 115320 2530
rect 115460 2520 115520 2530
rect 115240 2510 115250 2520
rect 115090 2470 115250 2510
rect 115090 2460 115100 2470
rect 115020 2450 115100 2460
rect 115240 2460 115250 2470
rect 115310 2460 115320 2520
rect 115240 2450 115320 2460
rect 108510 2330 108580 2332
rect 119020 2330 119090 2332
rect 108510 2320 108700 2330
rect 108580 2250 108630 2320
rect 108510 2240 108700 2250
rect 108750 2320 108820 2330
rect 108750 2240 108820 2250
rect 108870 2320 108940 2330
rect 118660 2320 118730 2330
rect 109060 2310 109140 2320
rect 109060 2300 109070 2310
rect 108940 2260 109070 2300
rect 108870 2240 108940 2250
rect 109060 2250 109070 2260
rect 109130 2250 109140 2310
rect 118460 2310 118540 2320
rect 109060 2240 109140 2250
rect 109460 2270 109540 2280
rect 109460 2210 109470 2270
rect 109530 2260 109540 2270
rect 109680 2270 109760 2280
rect 109680 2260 109690 2270
rect 109530 2220 109690 2260
rect 109530 2210 109540 2220
rect 109460 2200 109540 2210
rect 109680 2210 109690 2220
rect 109750 2260 109760 2270
rect 109900 2270 109980 2280
rect 109900 2260 109910 2270
rect 109750 2220 109910 2260
rect 109750 2210 109760 2220
rect 109680 2200 109760 2210
rect 109900 2210 109910 2220
rect 109970 2260 109980 2270
rect 110120 2270 110200 2280
rect 110120 2260 110130 2270
rect 109970 2220 110130 2260
rect 109970 2210 109980 2220
rect 109900 2200 109980 2210
rect 110120 2210 110130 2220
rect 110190 2260 110200 2270
rect 110340 2270 110420 2280
rect 110340 2260 110350 2270
rect 110190 2220 110350 2260
rect 110190 2210 110200 2220
rect 110120 2200 110200 2210
rect 110340 2210 110350 2220
rect 110410 2210 110420 2270
rect 110340 2200 110420 2210
rect 117180 2270 117260 2280
rect 117180 2210 117190 2270
rect 117250 2260 117260 2270
rect 117400 2270 117480 2280
rect 117400 2260 117410 2270
rect 117250 2220 117410 2260
rect 117250 2210 117260 2220
rect 117180 2200 117260 2210
rect 117400 2210 117410 2220
rect 117470 2260 117480 2270
rect 117620 2270 117700 2280
rect 117620 2260 117630 2270
rect 117470 2220 117630 2260
rect 117470 2210 117480 2220
rect 117400 2200 117480 2210
rect 117620 2210 117630 2220
rect 117690 2260 117700 2270
rect 117840 2270 117920 2280
rect 117840 2260 117850 2270
rect 117690 2220 117850 2260
rect 117690 2210 117700 2220
rect 117620 2200 117700 2210
rect 117840 2210 117850 2220
rect 117910 2260 117920 2270
rect 118060 2270 118140 2280
rect 118060 2260 118070 2270
rect 117910 2220 118070 2260
rect 117910 2210 117920 2220
rect 117840 2200 117920 2210
rect 118060 2210 118070 2220
rect 118130 2210 118140 2270
rect 118460 2250 118470 2310
rect 118530 2300 118540 2310
rect 118530 2260 118660 2300
rect 118530 2250 118540 2260
rect 118460 2240 118540 2250
rect 118660 2240 118730 2250
rect 118780 2320 118850 2330
rect 118780 2240 118850 2250
rect 118900 2320 119090 2330
rect 118970 2250 119020 2320
rect 118900 2240 119090 2250
rect 118060 2200 118140 2210
rect 108750 2170 108830 2180
rect 108750 2110 108760 2170
rect 108820 2150 108830 2170
rect 108970 2170 109050 2180
rect 118550 2170 118630 2180
rect 108970 2150 108980 2170
rect 108820 2120 108980 2150
rect 108820 2110 108830 2120
rect 108750 2100 108830 2110
rect 108970 2110 108980 2120
rect 109040 2110 109050 2170
rect 116290 2160 118250 2170
rect 108970 2100 109050 2110
rect 109350 2150 111310 2160
rect 109350 2090 109360 2150
rect 109420 2090 109580 2150
rect 109640 2090 109800 2150
rect 109860 2090 110020 2150
rect 110080 2090 110240 2150
rect 110300 2090 110460 2150
rect 110520 2090 111080 2150
rect 111140 2090 111160 2150
rect 111220 2090 111240 2150
rect 111300 2090 111310 2150
rect 109350 2070 111310 2090
rect 109350 2010 109360 2070
rect 109420 2010 109580 2070
rect 109640 2010 109800 2070
rect 109860 2010 110020 2070
rect 110080 2010 110240 2070
rect 110300 2010 110460 2070
rect 110520 2010 111080 2070
rect 111140 2010 111160 2070
rect 111220 2010 111240 2070
rect 111300 2010 111310 2070
rect 112170 2130 112250 2140
rect 112170 2070 112180 2130
rect 112240 2120 112250 2130
rect 112390 2130 112470 2140
rect 112390 2120 112400 2130
rect 112240 2080 112400 2120
rect 112240 2070 112250 2080
rect 112170 2060 112250 2070
rect 112390 2070 112400 2080
rect 112460 2120 112470 2130
rect 112610 2130 112690 2140
rect 112610 2120 112620 2130
rect 112460 2080 112620 2120
rect 112460 2070 112470 2080
rect 112390 2060 112470 2070
rect 112610 2070 112620 2080
rect 112680 2120 112690 2130
rect 112830 2130 112910 2140
rect 112830 2120 112840 2130
rect 112680 2080 112840 2120
rect 112680 2070 112690 2080
rect 112610 2060 112690 2070
rect 112830 2070 112840 2080
rect 112900 2120 112910 2130
rect 113050 2130 113130 2140
rect 113050 2120 113060 2130
rect 112900 2080 113060 2120
rect 112900 2070 112910 2080
rect 112830 2060 112910 2070
rect 113050 2070 113060 2080
rect 113120 2120 113130 2130
rect 113270 2130 113350 2140
rect 113270 2120 113280 2130
rect 113120 2080 113280 2120
rect 113120 2070 113130 2080
rect 113050 2060 113130 2070
rect 113270 2070 113280 2080
rect 113340 2070 113350 2130
rect 113270 2060 113350 2070
rect 113650 2130 113730 2140
rect 113650 2070 113660 2130
rect 113720 2120 113730 2130
rect 113870 2130 113950 2140
rect 113870 2120 113880 2130
rect 113720 2080 113880 2120
rect 113720 2070 113730 2080
rect 113650 2060 113730 2070
rect 113870 2070 113880 2080
rect 113940 2070 113950 2130
rect 113870 2060 113950 2070
rect 114250 2130 114330 2140
rect 114250 2070 114260 2130
rect 114320 2120 114330 2130
rect 114470 2130 114550 2140
rect 114470 2120 114480 2130
rect 114320 2080 114480 2120
rect 114320 2070 114330 2080
rect 114250 2060 114330 2070
rect 114470 2070 114480 2080
rect 114540 2120 114550 2130
rect 114690 2130 114770 2140
rect 114690 2120 114700 2130
rect 114540 2080 114700 2120
rect 114540 2070 114550 2080
rect 114470 2060 114550 2070
rect 114690 2070 114700 2080
rect 114760 2120 114770 2130
rect 114910 2130 114990 2140
rect 114910 2120 114920 2130
rect 114760 2080 114920 2120
rect 114760 2070 114770 2080
rect 114690 2060 114770 2070
rect 114910 2070 114920 2080
rect 114980 2120 114990 2130
rect 115130 2130 115210 2140
rect 115130 2120 115140 2130
rect 114980 2080 115140 2120
rect 114980 2070 114990 2080
rect 114910 2060 114990 2070
rect 115130 2070 115140 2080
rect 115200 2120 115210 2130
rect 115350 2130 115430 2140
rect 115350 2120 115360 2130
rect 115200 2080 115360 2120
rect 115200 2070 115210 2080
rect 115130 2060 115210 2070
rect 115350 2070 115360 2080
rect 115420 2070 115430 2130
rect 115350 2060 115430 2070
rect 116290 2100 116300 2160
rect 116360 2100 116380 2160
rect 116440 2100 116460 2160
rect 116520 2100 117080 2160
rect 117140 2100 117300 2160
rect 117360 2100 117520 2160
rect 117580 2100 117740 2160
rect 117800 2100 117960 2160
rect 118020 2100 118180 2160
rect 118240 2100 118250 2160
rect 118550 2110 118560 2170
rect 118620 2160 118630 2170
rect 118770 2170 118850 2180
rect 118770 2160 118780 2170
rect 118620 2120 118780 2160
rect 118620 2110 118630 2120
rect 118550 2100 118630 2110
rect 118770 2110 118780 2120
rect 118840 2110 118850 2170
rect 118770 2100 118850 2110
rect 116290 2080 118250 2100
rect 109350 1990 111310 2010
rect 116290 2020 116300 2080
rect 116360 2020 116380 2080
rect 116440 2020 116460 2080
rect 116520 2020 117080 2080
rect 117140 2020 117300 2080
rect 117360 2020 117520 2080
rect 117580 2020 117740 2080
rect 117800 2020 117960 2080
rect 118020 2020 118180 2080
rect 118240 2020 118250 2080
rect 116290 2000 118250 2020
rect 109350 1930 109360 1990
rect 109420 1930 109580 1990
rect 109640 1930 109800 1990
rect 109860 1930 110020 1990
rect 110080 1930 110240 1990
rect 110300 1930 110460 1990
rect 110520 1930 111080 1990
rect 111140 1930 111160 1990
rect 111220 1930 111240 1990
rect 111300 1930 111310 1990
rect 109350 1920 111310 1930
rect 112280 1990 115320 2000
rect 112280 1930 112290 1990
rect 112350 1930 112510 1990
rect 112570 1930 112730 1990
rect 112790 1930 112950 1990
rect 113010 1930 113170 1990
rect 113230 1930 114370 1990
rect 114430 1930 114590 1990
rect 114650 1930 114810 1990
rect 114870 1930 115030 1990
rect 115090 1930 115250 1990
rect 115310 1930 115320 1990
rect 116290 1940 116300 2000
rect 116360 1940 116380 2000
rect 116440 1940 116460 2000
rect 116520 1940 117080 2000
rect 117140 1940 117300 2000
rect 117360 1940 117520 2000
rect 117580 1940 117740 2000
rect 117800 1940 117960 2000
rect 118020 1940 118180 2000
rect 118240 1940 118250 2000
rect 116290 1930 118250 1940
rect 112280 1920 115320 1930
rect 107680 1880 119920 1890
rect 107680 1820 107690 1880
rect 107750 1820 107770 1880
rect 107830 1820 107850 1880
rect 107910 1820 109250 1880
rect 109310 1820 110570 1880
rect 110630 1820 112070 1880
rect 112130 1820 113470 1880
rect 113530 1820 114070 1880
rect 114130 1820 115470 1880
rect 115530 1820 116970 1880
rect 117030 1820 118290 1880
rect 118350 1820 119690 1880
rect 119750 1820 119770 1880
rect 119830 1820 119850 1880
rect 119910 1820 119920 1880
rect 107680 1800 119920 1820
rect 107680 1740 107690 1800
rect 107750 1740 107770 1800
rect 107830 1740 107850 1800
rect 107910 1740 109250 1800
rect 109310 1740 110570 1800
rect 110630 1740 112070 1800
rect 112130 1740 113470 1800
rect 113530 1740 114070 1800
rect 114130 1740 115470 1800
rect 115530 1740 116970 1800
rect 117030 1740 118290 1800
rect 118350 1740 119690 1800
rect 119750 1740 119770 1800
rect 119830 1740 119850 1800
rect 119910 1740 119920 1800
rect 107680 1720 119920 1740
rect 107680 1660 107690 1720
rect 107750 1660 107770 1720
rect 107830 1660 107850 1720
rect 107910 1660 109250 1720
rect 109310 1660 110570 1720
rect 110630 1660 112070 1720
rect 112130 1660 113470 1720
rect 113530 1660 114070 1720
rect 114130 1660 115470 1720
rect 115530 1660 116970 1720
rect 117030 1660 118290 1720
rect 118350 1660 119690 1720
rect 119750 1660 119770 1720
rect 119830 1660 119850 1720
rect 119910 1660 119920 1720
rect 107680 1650 119920 1660
rect 108510 1610 108590 1620
rect 108510 1550 108520 1610
rect 108580 1600 108590 1610
rect 111880 1610 111960 1620
rect 111880 1600 111890 1610
rect 108580 1560 111890 1600
rect 108580 1550 108590 1560
rect 108510 1540 108590 1550
rect 111880 1550 111890 1560
rect 111950 1550 111960 1610
rect 111880 1540 111960 1550
rect 115640 1610 115720 1620
rect 115640 1550 115650 1610
rect 115710 1600 115720 1610
rect 119010 1610 119090 1620
rect 119010 1600 119020 1610
rect 115710 1560 119020 1600
rect 115710 1550 115720 1560
rect 115640 1540 115720 1550
rect 119010 1550 119020 1560
rect 119080 1550 119090 1610
rect 119010 1540 119090 1550
rect 108640 1150 118960 1160
rect 108640 1090 108650 1150
rect 108710 1090 118890 1150
rect 118950 1090 118960 1150
rect 108640 1080 118960 1090
rect 107980 1040 110380 1050
rect 117220 1040 119620 1050
rect 107980 980 107990 1040
rect 108050 980 108070 1040
rect 108130 980 108160 1040
rect 108220 980 108240 1040
rect 108300 980 108330 1040
rect 108390 980 108410 1040
rect 108470 980 108780 1040
rect 108840 980 109510 1040
rect 109570 980 109590 1040
rect 109650 980 109670 1040
rect 109730 980 109750 1040
rect 109810 980 109830 1040
rect 109890 980 109910 1040
rect 109970 980 109990 1040
rect 110050 980 110070 1040
rect 110130 980 110150 1040
rect 110210 980 110230 1040
rect 110290 980 110310 1040
rect 110370 980 110380 1040
rect 107980 960 110380 980
rect 112880 1030 114940 1040
rect 112880 970 112890 1030
rect 112950 970 113110 1030
rect 113170 970 113330 1030
rect 113390 970 113550 1030
rect 113610 970 113770 1030
rect 113830 970 113990 1030
rect 114050 970 114210 1030
rect 114270 970 114430 1030
rect 114490 970 114650 1030
rect 114710 970 114870 1030
rect 114930 970 114940 1030
rect 112880 960 114940 970
rect 117220 980 117230 1040
rect 117290 980 117310 1040
rect 117370 980 117390 1040
rect 117450 980 117470 1040
rect 117530 980 117550 1040
rect 117610 980 117630 1040
rect 117690 980 117710 1040
rect 117770 980 117790 1040
rect 117850 980 117870 1040
rect 117930 980 117950 1040
rect 118010 980 118030 1040
rect 118090 980 118760 1040
rect 118820 980 119130 1040
rect 119190 980 119210 1040
rect 119270 980 119300 1040
rect 119360 980 119380 1040
rect 119440 980 119470 1040
rect 119530 980 119550 1040
rect 119610 980 119620 1040
rect 117220 960 119620 980
rect 107980 900 107990 960
rect 108050 900 108070 960
rect 108130 900 108160 960
rect 108220 900 108240 960
rect 108300 900 108330 960
rect 108390 900 108410 960
rect 108470 900 108780 960
rect 108840 900 109510 960
rect 109570 900 109590 960
rect 109650 900 109670 960
rect 109730 900 109750 960
rect 109810 900 109830 960
rect 109890 900 109910 960
rect 109970 900 109990 960
rect 110050 900 110070 960
rect 110130 900 110150 960
rect 110210 900 110230 960
rect 110290 900 110310 960
rect 110370 900 110380 960
rect 107980 880 110380 900
rect 107980 820 107990 880
rect 108050 820 108070 880
rect 108130 820 108160 880
rect 108220 820 108240 880
rect 108300 820 108330 880
rect 108390 820 108410 880
rect 108470 820 108780 880
rect 108840 820 109510 880
rect 109570 820 109590 880
rect 109650 820 109670 880
rect 109730 820 109750 880
rect 109810 820 109830 880
rect 109890 820 109910 880
rect 109970 820 109990 880
rect 110050 820 110070 880
rect 110130 820 110150 880
rect 110210 820 110230 880
rect 110290 820 110310 880
rect 110370 820 110380 880
rect 107980 810 110380 820
rect 117220 900 117230 960
rect 117290 900 117310 960
rect 117370 900 117390 960
rect 117450 900 117470 960
rect 117530 900 117550 960
rect 117610 900 117630 960
rect 117690 900 117710 960
rect 117770 900 117790 960
rect 117850 900 117870 960
rect 117930 900 117950 960
rect 118010 900 118030 960
rect 118090 900 118760 960
rect 118820 900 119130 960
rect 119190 900 119210 960
rect 119270 900 119300 960
rect 119360 900 119380 960
rect 119440 900 119470 960
rect 119530 900 119550 960
rect 119610 900 119620 960
rect 117220 880 119620 900
rect 117220 820 117230 880
rect 117290 820 117310 880
rect 117370 820 117390 880
rect 117450 820 117470 880
rect 117530 820 117550 880
rect 117610 820 117630 880
rect 117690 820 117710 880
rect 117770 820 117790 880
rect 117850 820 117870 880
rect 117930 820 117950 880
rect 118010 820 118030 880
rect 118090 820 118760 880
rect 118820 820 119130 880
rect 119190 820 119210 880
rect 119270 820 119300 880
rect 119360 820 119380 880
rect 119440 820 119470 880
rect 119530 820 119550 880
rect 119610 820 119620 880
rect 117220 810 119620 820
rect 108640 770 110280 780
rect 108640 710 108650 770
rect 108710 710 109610 770
rect 109670 710 109810 770
rect 109870 710 110010 770
rect 110070 710 110210 770
rect 110270 710 110280 770
rect 108640 700 110280 710
rect 117320 770 118960 780
rect 117320 710 117330 770
rect 117390 710 117530 770
rect 117590 710 117730 770
rect 117790 710 117930 770
rect 117990 710 118890 770
rect 118950 710 118960 770
rect 117320 700 118960 710
rect 108650 660 108720 670
rect 108650 580 108720 590
rect 108770 660 108840 670
rect 108770 580 108840 590
rect 118760 660 118830 670
rect 118760 580 118830 590
rect 118880 660 118950 670
rect 118880 580 118950 590
rect 112440 370 112520 380
rect 112440 310 112450 370
rect 112510 360 112520 370
rect 112550 370 112630 380
rect 112550 360 112560 370
rect 112510 320 112560 360
rect 112510 310 112520 320
rect 112440 300 112520 310
rect 112550 310 112560 320
rect 112620 360 112630 370
rect 112770 370 112850 380
rect 112770 360 112780 370
rect 112620 320 112780 360
rect 112620 310 112630 320
rect 112550 300 112630 310
rect 112770 310 112780 320
rect 112840 360 112850 370
rect 112990 370 113070 380
rect 112990 360 113000 370
rect 112840 320 113000 360
rect 112840 310 112850 320
rect 112770 300 112850 310
rect 112990 310 113000 320
rect 113060 360 113070 370
rect 113210 370 113290 380
rect 113210 360 113220 370
rect 113060 320 113220 360
rect 113060 310 113070 320
rect 112990 300 113070 310
rect 113210 310 113220 320
rect 113280 360 113290 370
rect 113430 370 113510 380
rect 113430 360 113440 370
rect 113280 320 113440 360
rect 113280 310 113290 320
rect 113210 300 113290 310
rect 113430 310 113440 320
rect 113500 360 113510 370
rect 113650 370 113730 380
rect 113650 360 113660 370
rect 113500 320 113660 360
rect 113500 310 113510 320
rect 113430 300 113510 310
rect 113650 310 113660 320
rect 113720 360 113730 370
rect 113870 370 113950 380
rect 113870 360 113880 370
rect 113720 320 113880 360
rect 113720 310 113730 320
rect 113650 300 113730 310
rect 113870 310 113880 320
rect 113940 360 113950 370
rect 114090 370 114170 380
rect 114090 360 114100 370
rect 113940 320 114100 360
rect 113940 310 113950 320
rect 113870 300 113950 310
rect 114090 310 114100 320
rect 114160 360 114170 370
rect 114310 370 114390 380
rect 114310 360 114320 370
rect 114160 320 114320 360
rect 114160 310 114170 320
rect 114090 300 114170 310
rect 114310 310 114320 320
rect 114380 360 114390 370
rect 114530 370 114610 380
rect 114530 360 114540 370
rect 114380 320 114540 360
rect 114380 310 114390 320
rect 114310 300 114390 310
rect 114530 310 114540 320
rect 114600 360 114610 370
rect 114750 370 114830 380
rect 114750 360 114760 370
rect 114600 320 114760 360
rect 114600 310 114610 320
rect 114530 300 114610 310
rect 114750 310 114760 320
rect 114820 360 114830 370
rect 114970 370 115050 380
rect 114970 360 114980 370
rect 114820 320 114980 360
rect 114820 310 114830 320
rect 114750 300 114830 310
rect 114970 310 114980 320
rect 115040 310 115050 370
rect 114970 300 115050 310
rect 112880 260 115660 270
rect 112880 200 112890 260
rect 112950 200 113110 260
rect 113170 200 113330 260
rect 113390 200 113550 260
rect 113610 200 113770 260
rect 113830 200 113990 260
rect 114050 200 114210 260
rect 114270 200 114430 260
rect 114490 200 114650 260
rect 114710 200 114870 260
rect 114930 200 115430 260
rect 115490 200 115510 260
rect 115570 200 115590 260
rect 115650 200 115660 260
rect 112880 180 115660 200
rect 112880 120 112890 180
rect 112950 120 113110 180
rect 113170 120 113330 180
rect 113390 120 113550 180
rect 113610 120 113770 180
rect 113830 120 113990 180
rect 114050 120 114210 180
rect 114270 120 114430 180
rect 114490 120 114650 180
rect 114710 120 114870 180
rect 114930 120 115430 180
rect 115490 120 115510 180
rect 115570 120 115590 180
rect 115650 120 115660 180
rect 112880 100 115660 120
rect 112880 40 112890 100
rect 112950 40 113110 100
rect 113170 40 113330 100
rect 113390 40 113550 100
rect 113610 40 113770 100
rect 113830 40 113990 100
rect 114050 40 114210 100
rect 114270 40 114430 100
rect 114490 40 114650 100
rect 114710 40 114870 100
rect 114930 40 115430 100
rect 115490 40 115510 100
rect 115570 40 115590 100
rect 115650 40 115660 100
rect 112880 30 115660 40
rect 114830 -10 114910 0
rect 114830 -70 114840 -10
rect 114900 -20 114910 -10
rect 115730 -10 115810 0
rect 115730 -20 115740 -10
rect 114900 -60 115740 -20
rect 114900 -70 114910 -60
rect 114830 -80 114910 -70
rect 115730 -70 115740 -60
rect 115800 -70 115810 -10
rect 115730 -80 115810 -70
rect 111340 -120 116260 -110
rect 111340 -180 111350 -120
rect 111410 -180 111430 -120
rect 111490 -180 111510 -120
rect 111570 -180 112670 -120
rect 112730 -180 116030 -120
rect 116090 -180 116110 -120
rect 116170 -180 116190 -120
rect 116250 -180 116260 -120
rect 111340 -200 116260 -180
rect 111340 -260 111350 -200
rect 111410 -260 111430 -200
rect 111490 -260 111510 -200
rect 111570 -260 112670 -200
rect 112730 -260 116030 -200
rect 116090 -260 116110 -200
rect 116170 -260 116190 -200
rect 116250 -260 116260 -200
rect 111340 -280 116260 -260
rect 111340 -340 111350 -280
rect 111410 -340 111430 -280
rect 111490 -340 111510 -280
rect 111570 -340 112670 -280
rect 112730 -340 116030 -280
rect 116090 -340 116110 -280
rect 116170 -340 116190 -280
rect 116250 -340 116260 -280
rect 111340 -350 116260 -340
rect 113080 -390 113160 -380
rect 113080 -450 113090 -390
rect 113150 -400 113160 -390
rect 113300 -390 113380 -380
rect 113300 -400 113310 -390
rect 113150 -440 113310 -400
rect 113150 -450 113160 -440
rect 113080 -460 113160 -450
rect 113300 -450 113310 -440
rect 113370 -400 113380 -390
rect 113740 -390 113820 -380
rect 113740 -400 113750 -390
rect 113370 -440 113750 -400
rect 113370 -450 113380 -440
rect 113300 -460 113380 -450
rect 113740 -450 113750 -440
rect 113810 -450 113820 -390
rect 113740 -460 113820 -450
rect 111690 -500 114160 -490
rect 111690 -560 111700 -500
rect 111760 -560 111780 -500
rect 111840 -560 112980 -500
rect 113040 -560 113200 -500
rect 113260 -560 113420 -500
rect 113480 -560 114090 -500
rect 114150 -560 114160 -500
rect 111690 -570 114160 -560
rect 109500 -730 110380 -720
rect 109500 -790 109510 -730
rect 109570 -790 109910 -730
rect 109970 -790 110310 -730
rect 110370 -790 110380 -730
rect 109500 -800 110380 -790
rect 111690 -930 112750 -570
rect 114430 -640 115660 -630
rect 114430 -650 115430 -640
rect 114490 -700 115430 -650
rect 115490 -700 115510 -640
rect 115570 -700 115590 -640
rect 115650 -700 115660 -640
rect 114490 -720 115660 -700
rect 114490 -780 115430 -720
rect 115490 -780 115510 -720
rect 115570 -780 115590 -720
rect 115650 -780 115660 -720
rect 114490 -800 115660 -780
rect 117220 -730 118100 -720
rect 117220 -790 117230 -730
rect 117290 -790 117630 -730
rect 117690 -790 118030 -730
rect 118090 -790 118100 -730
rect 117220 -800 118100 -790
rect 114490 -850 115430 -800
rect 114430 -860 115430 -850
rect 115490 -860 115510 -800
rect 115570 -860 115590 -800
rect 115650 -860 115660 -800
rect 114430 -870 115660 -860
rect 111690 -940 114160 -930
rect 111690 -1000 111700 -940
rect 111760 -1000 111780 -940
rect 111840 -1000 112980 -940
rect 113040 -1000 113200 -940
rect 113260 -1000 113420 -940
rect 113480 -1000 114090 -940
rect 114150 -1000 114160 -940
rect 111690 -1010 114160 -1000
rect 113080 -1050 113820 -1040
rect 113080 -1110 113090 -1050
rect 113150 -1110 113310 -1050
rect 113370 -1110 113750 -1050
rect 113810 -1110 113820 -1050
rect 113080 -1120 113820 -1110
rect 104580 -1160 123020 -1150
rect 104580 -1220 104590 -1160
rect 104650 -1220 104670 -1160
rect 104730 -1220 104750 -1160
rect 104810 -1220 105290 -1160
rect 105350 -1220 105370 -1160
rect 105430 -1220 105450 -1160
rect 105510 -1220 105990 -1160
rect 106050 -1220 106070 -1160
rect 106130 -1220 106150 -1160
rect 106210 -1220 106690 -1160
rect 106750 -1220 106770 -1160
rect 106830 -1220 106850 -1160
rect 106910 -1220 107390 -1160
rect 107450 -1220 107470 -1160
rect 107530 -1220 107550 -1160
rect 107610 -1220 107690 -1160
rect 107750 -1220 107770 -1160
rect 107830 -1220 107850 -1160
rect 107910 -1220 108090 -1160
rect 108150 -1220 108170 -1160
rect 108230 -1220 108250 -1160
rect 108310 -1220 108790 -1160
rect 108850 -1220 108870 -1160
rect 108930 -1220 108950 -1160
rect 109010 -1220 109310 -1160
rect 109370 -1220 109490 -1160
rect 109550 -1220 109570 -1160
rect 109630 -1220 109650 -1160
rect 109710 -1220 110190 -1160
rect 110250 -1220 110270 -1160
rect 110330 -1220 110350 -1160
rect 110410 -1220 110510 -1160
rect 110570 -1220 110890 -1160
rect 110950 -1220 110970 -1160
rect 111030 -1220 111050 -1160
rect 111110 -1220 111590 -1160
rect 111650 -1220 111670 -1160
rect 111730 -1220 111750 -1160
rect 111810 -1220 112290 -1160
rect 112350 -1220 112370 -1160
rect 112430 -1220 112450 -1160
rect 112510 -1220 112870 -1160
rect 112930 -1220 112990 -1160
rect 113050 -1220 113070 -1160
rect 113130 -1220 113150 -1160
rect 113210 -1220 113530 -1160
rect 113590 -1220 113690 -1160
rect 113750 -1220 113770 -1160
rect 113830 -1220 113850 -1160
rect 113910 -1220 114390 -1160
rect 114450 -1220 114470 -1160
rect 114530 -1220 114550 -1160
rect 114610 -1220 114980 -1160
rect 115040 -1220 115090 -1160
rect 115150 -1220 115170 -1160
rect 115230 -1220 115250 -1160
rect 115310 -1220 115790 -1160
rect 115850 -1220 115870 -1160
rect 115930 -1220 115950 -1160
rect 116010 -1220 116490 -1160
rect 116550 -1220 116570 -1160
rect 116630 -1220 116650 -1160
rect 116710 -1220 117030 -1160
rect 117090 -1220 117190 -1160
rect 117250 -1220 117270 -1160
rect 117330 -1220 117350 -1160
rect 117410 -1220 117890 -1160
rect 117950 -1220 117970 -1160
rect 118030 -1220 118050 -1160
rect 118110 -1220 118230 -1160
rect 118290 -1220 118750 -1160
rect 118810 -1220 118830 -1160
rect 118890 -1220 118910 -1160
rect 118970 -1220 119290 -1160
rect 119350 -1220 119370 -1160
rect 119430 -1220 119450 -1160
rect 119510 -1220 119690 -1160
rect 119750 -1220 119770 -1160
rect 119830 -1220 119850 -1160
rect 119910 -1220 119990 -1160
rect 120050 -1220 120070 -1160
rect 120130 -1220 120150 -1160
rect 120210 -1220 120690 -1160
rect 120750 -1220 120770 -1160
rect 120830 -1220 120850 -1160
rect 120910 -1220 121390 -1160
rect 121450 -1220 121470 -1160
rect 121530 -1220 121550 -1160
rect 121610 -1220 122090 -1160
rect 122150 -1220 122170 -1160
rect 122230 -1220 122250 -1160
rect 122310 -1220 122790 -1160
rect 122850 -1220 122870 -1160
rect 122930 -1220 122950 -1160
rect 123010 -1220 123020 -1160
rect 104580 -1240 123020 -1220
rect 104580 -1300 104590 -1240
rect 104650 -1300 104670 -1240
rect 104730 -1300 104750 -1240
rect 104810 -1300 105290 -1240
rect 105350 -1300 105370 -1240
rect 105430 -1300 105450 -1240
rect 105510 -1300 105990 -1240
rect 106050 -1300 106070 -1240
rect 106130 -1300 106150 -1240
rect 106210 -1300 106690 -1240
rect 106750 -1300 106770 -1240
rect 106830 -1300 106850 -1240
rect 106910 -1300 107390 -1240
rect 107450 -1300 107470 -1240
rect 107530 -1300 107550 -1240
rect 107610 -1300 107690 -1240
rect 107750 -1300 107770 -1240
rect 107830 -1300 107850 -1240
rect 107910 -1300 108090 -1240
rect 108150 -1300 108170 -1240
rect 108230 -1300 108250 -1240
rect 108310 -1300 108790 -1240
rect 108850 -1300 108870 -1240
rect 108930 -1300 108950 -1240
rect 109010 -1300 109310 -1240
rect 109370 -1300 109490 -1240
rect 109550 -1300 109570 -1240
rect 109630 -1300 109650 -1240
rect 109710 -1300 110190 -1240
rect 110250 -1300 110270 -1240
rect 110330 -1300 110350 -1240
rect 110410 -1300 110510 -1240
rect 110570 -1300 110890 -1240
rect 110950 -1300 110970 -1240
rect 111030 -1300 111050 -1240
rect 111110 -1300 111590 -1240
rect 111650 -1300 111670 -1240
rect 111730 -1300 111750 -1240
rect 111810 -1300 112290 -1240
rect 112350 -1300 112370 -1240
rect 112430 -1300 112450 -1240
rect 112510 -1300 112870 -1240
rect 112930 -1300 112990 -1240
rect 113050 -1300 113070 -1240
rect 113130 -1300 113150 -1240
rect 113210 -1300 113530 -1240
rect 113590 -1300 113690 -1240
rect 113750 -1300 113770 -1240
rect 113830 -1300 113850 -1240
rect 113910 -1300 114390 -1240
rect 114450 -1300 114470 -1240
rect 114530 -1300 114550 -1240
rect 114610 -1300 114980 -1240
rect 115040 -1300 115090 -1240
rect 115150 -1300 115170 -1240
rect 115230 -1300 115250 -1240
rect 115310 -1300 115790 -1240
rect 115850 -1300 115870 -1240
rect 115930 -1300 115950 -1240
rect 116010 -1300 116490 -1240
rect 116550 -1300 116570 -1240
rect 116630 -1300 116650 -1240
rect 116710 -1300 117030 -1240
rect 117090 -1300 117190 -1240
rect 117250 -1300 117270 -1240
rect 117330 -1300 117350 -1240
rect 117410 -1300 117890 -1240
rect 117950 -1300 117970 -1240
rect 118030 -1300 118050 -1240
rect 118110 -1300 118230 -1240
rect 118290 -1300 118750 -1240
rect 118810 -1300 118830 -1240
rect 118890 -1300 118910 -1240
rect 118970 -1300 119290 -1240
rect 119350 -1300 119370 -1240
rect 119430 -1300 119450 -1240
rect 119510 -1300 119690 -1240
rect 119750 -1300 119770 -1240
rect 119830 -1300 119850 -1240
rect 119910 -1300 119990 -1240
rect 120050 -1300 120070 -1240
rect 120130 -1300 120150 -1240
rect 120210 -1300 120690 -1240
rect 120750 -1300 120770 -1240
rect 120830 -1300 120850 -1240
rect 120910 -1300 121390 -1240
rect 121450 -1300 121470 -1240
rect 121530 -1300 121550 -1240
rect 121610 -1300 122090 -1240
rect 122150 -1300 122170 -1240
rect 122230 -1300 122250 -1240
rect 122310 -1300 122790 -1240
rect 122850 -1300 122870 -1240
rect 122930 -1300 122950 -1240
rect 123010 -1300 123020 -1240
rect 104580 -1320 123020 -1300
rect 104580 -1380 104590 -1320
rect 104650 -1380 104670 -1320
rect 104730 -1380 104750 -1320
rect 104810 -1380 105290 -1320
rect 105350 -1380 105370 -1320
rect 105430 -1380 105450 -1320
rect 105510 -1380 105990 -1320
rect 106050 -1380 106070 -1320
rect 106130 -1380 106150 -1320
rect 106210 -1380 106690 -1320
rect 106750 -1380 106770 -1320
rect 106830 -1380 106850 -1320
rect 106910 -1380 107390 -1320
rect 107450 -1380 107470 -1320
rect 107530 -1380 107550 -1320
rect 107610 -1380 107690 -1320
rect 107750 -1380 107770 -1320
rect 107830 -1380 107850 -1320
rect 107910 -1380 108090 -1320
rect 108150 -1380 108170 -1320
rect 108230 -1380 108250 -1320
rect 108310 -1380 108790 -1320
rect 108850 -1380 108870 -1320
rect 108930 -1380 108950 -1320
rect 109010 -1380 109310 -1320
rect 109370 -1380 109490 -1320
rect 109550 -1380 109570 -1320
rect 109630 -1380 109650 -1320
rect 109710 -1380 110190 -1320
rect 110250 -1380 110270 -1320
rect 110330 -1380 110350 -1320
rect 110410 -1380 110510 -1320
rect 110570 -1380 110890 -1320
rect 110950 -1380 110970 -1320
rect 111030 -1380 111050 -1320
rect 111110 -1380 111590 -1320
rect 111650 -1380 111670 -1320
rect 111730 -1380 111750 -1320
rect 111810 -1380 112290 -1320
rect 112350 -1380 112370 -1320
rect 112430 -1380 112450 -1320
rect 112510 -1380 112870 -1320
rect 112930 -1380 112990 -1320
rect 113050 -1380 113070 -1320
rect 113130 -1380 113150 -1320
rect 113210 -1380 113530 -1320
rect 113590 -1380 113690 -1320
rect 113750 -1380 113770 -1320
rect 113830 -1380 113850 -1320
rect 113910 -1380 114390 -1320
rect 114450 -1380 114470 -1320
rect 114530 -1380 114550 -1320
rect 114610 -1380 114980 -1320
rect 115040 -1380 115090 -1320
rect 115150 -1380 115170 -1320
rect 115230 -1380 115250 -1320
rect 115310 -1380 115790 -1320
rect 115850 -1380 115870 -1320
rect 115930 -1380 115950 -1320
rect 116010 -1380 116490 -1320
rect 116550 -1380 116570 -1320
rect 116630 -1380 116650 -1320
rect 116710 -1380 117030 -1320
rect 117090 -1380 117190 -1320
rect 117250 -1380 117270 -1320
rect 117330 -1380 117350 -1320
rect 117410 -1380 117890 -1320
rect 117950 -1380 117970 -1320
rect 118030 -1380 118050 -1320
rect 118110 -1380 118230 -1320
rect 118290 -1380 118750 -1320
rect 118810 -1380 118830 -1320
rect 118890 -1380 118910 -1320
rect 118970 -1380 119290 -1320
rect 119350 -1380 119370 -1320
rect 119430 -1380 119450 -1320
rect 119510 -1380 119690 -1320
rect 119750 -1380 119770 -1320
rect 119830 -1380 119850 -1320
rect 119910 -1380 119990 -1320
rect 120050 -1380 120070 -1320
rect 120130 -1380 120150 -1320
rect 120210 -1380 120690 -1320
rect 120750 -1380 120770 -1320
rect 120830 -1380 120850 -1320
rect 120910 -1380 121390 -1320
rect 121450 -1380 121470 -1320
rect 121530 -1380 121550 -1320
rect 121610 -1380 122090 -1320
rect 122150 -1380 122170 -1320
rect 122230 -1380 122250 -1320
rect 122310 -1380 122790 -1320
rect 122850 -1380 122870 -1320
rect 122930 -1380 122950 -1320
rect 123010 -1380 123020 -1320
rect 104580 -1390 123020 -1380
<< via2 >>
rect 108520 6690 108580 6750
rect 119020 6690 119080 6750
rect 108000 3360 108060 3420
rect 108100 3360 108160 3420
rect 108200 3360 108260 3420
rect 108300 3360 108360 3420
rect 108400 3360 108460 3420
rect 108000 3260 108060 3320
rect 108100 3260 108160 3320
rect 108200 3260 108260 3320
rect 108300 3260 108360 3320
rect 108400 3260 108460 3320
rect 119140 3360 119200 3420
rect 119240 3360 119300 3420
rect 119340 3360 119400 3420
rect 119440 3360 119500 3420
rect 119540 3360 119600 3420
rect 108000 3160 108060 3220
rect 108100 3160 108160 3220
rect 108200 3160 108260 3220
rect 108300 3160 108360 3220
rect 108400 3160 108460 3220
rect 119140 3260 119200 3320
rect 119240 3260 119300 3320
rect 119340 3260 119400 3320
rect 119440 3260 119500 3320
rect 119540 3260 119600 3320
rect 119140 3160 119200 3220
rect 119240 3160 119300 3220
rect 119340 3160 119400 3220
rect 119440 3160 119500 3220
rect 119540 3160 119600 3220
<< metal3 >>
rect 104120 11040 104580 11210
rect 104820 11040 105280 11210
rect 105520 11040 105980 11210
rect 106220 11040 106680 11210
rect 106920 11040 107380 11210
rect 107620 11040 108080 11210
rect 108320 11040 108780 11210
rect 109020 11040 109480 11210
rect 109720 11040 110180 11210
rect 110420 11040 110880 11210
rect 111120 11040 111580 11210
rect 111820 11040 112280 11210
rect 112520 11040 112980 11210
rect 113220 11040 113680 11210
rect 104120 10940 113680 11040
rect 104120 10750 104580 10940
rect 104820 10750 105280 10940
rect 105520 10750 105980 10940
rect 106220 10750 106680 10940
rect 106920 10750 107380 10940
rect 107620 10750 108080 10940
rect 108320 10750 108780 10940
rect 109020 10750 109480 10940
rect 109720 10750 110180 10940
rect 110420 10750 110880 10940
rect 111120 10750 111580 10940
rect 111820 10750 112280 10940
rect 112520 10750 112980 10940
rect 113220 10750 113680 10940
rect 113920 11040 114380 11210
rect 114620 11040 115080 11210
rect 115320 11040 115780 11210
rect 116020 11040 116480 11210
rect 116720 11040 117180 11210
rect 117420 11040 117880 11210
rect 118120 11040 118580 11210
rect 118820 11040 119280 11210
rect 119520 11040 119980 11210
rect 120220 11040 120680 11210
rect 120920 11040 121380 11210
rect 121620 11040 122080 11210
rect 122320 11040 122780 11210
rect 123020 11040 123480 11210
rect 113920 10940 123480 11040
rect 113920 10750 114380 10940
rect 114620 10750 115080 10940
rect 115320 10750 115780 10940
rect 116020 10750 116480 10940
rect 116720 10750 117180 10940
rect 117420 10750 117880 10940
rect 118120 10750 118580 10940
rect 118820 10750 119280 10940
rect 119520 10750 119980 10940
rect 120220 10750 120680 10940
rect 120920 10750 121380 10940
rect 121620 10750 122080 10940
rect 122320 10750 122780 10940
rect 123020 10750 123480 10940
rect 105700 10510 105800 10750
rect 107800 10510 107900 10750
rect 108500 10510 108600 10750
rect 109200 10510 109300 10750
rect 109900 10510 110000 10750
rect 110600 10510 110700 10750
rect 111300 10510 111400 10750
rect 116200 10510 116300 10750
rect 116900 10510 117000 10750
rect 117600 10510 117700 10750
rect 118300 10510 118400 10750
rect 119000 10510 119100 10750
rect 119700 10510 119800 10750
rect 121800 10510 121900 10750
rect 104120 10340 104580 10510
rect 104820 10340 105280 10510
rect 105520 10340 105980 10510
rect 106220 10340 106680 10510
rect 106920 10340 107380 10510
rect 104120 10240 107380 10340
rect 104120 10050 104580 10240
rect 104820 10050 105280 10240
rect 105520 10050 105980 10240
rect 106220 10050 106680 10240
rect 106920 10050 107380 10240
rect 107620 10050 108080 10510
rect 108320 10050 108780 10510
rect 109020 10050 109480 10510
rect 109720 10050 110180 10510
rect 110420 10050 110880 10510
rect 111120 10050 111580 10510
rect 116020 10050 116480 10510
rect 116720 10050 117180 10510
rect 117420 10050 117880 10510
rect 118120 10050 118580 10510
rect 118820 10050 119280 10510
rect 119520 10050 119980 10510
rect 120220 10340 120680 10510
rect 120920 10340 121380 10510
rect 121620 10340 122080 10510
rect 122320 10340 122780 10510
rect 123020 10340 123480 10510
rect 120220 10240 123480 10340
rect 120220 10050 120680 10240
rect 120920 10050 121380 10240
rect 121620 10050 122080 10240
rect 122320 10050 122780 10240
rect 123020 10050 123480 10240
rect 105700 9810 105800 10050
rect 107800 9810 107900 10050
rect 108500 9810 108600 10050
rect 109200 9810 109300 10050
rect 109900 9810 110000 10050
rect 110600 9810 110700 10050
rect 116900 9810 117000 10050
rect 117600 9810 117700 10050
rect 118300 9810 118400 10050
rect 119000 9810 119100 10050
rect 119700 9810 119800 10050
rect 121800 9810 121900 10050
rect 104120 9640 104580 9810
rect 104820 9640 105280 9810
rect 105520 9640 105980 9810
rect 106220 9640 106680 9810
rect 106920 9640 107380 9810
rect 104120 9540 107380 9640
rect 104120 9350 104580 9540
rect 104820 9350 105280 9540
rect 105520 9350 105980 9540
rect 106220 9350 106680 9540
rect 106920 9350 107380 9540
rect 107620 9350 108080 9810
rect 108320 9350 108780 9810
rect 109020 9350 109480 9810
rect 109720 9350 110180 9810
rect 110420 9350 110880 9810
rect 116720 9350 117180 9810
rect 117420 9350 117880 9810
rect 118120 9350 118580 9810
rect 118820 9350 119280 9810
rect 119520 9350 119980 9810
rect 120220 9640 120680 9810
rect 120920 9640 121380 9810
rect 121620 9640 122080 9810
rect 122320 9640 122780 9810
rect 123020 9640 123480 9810
rect 120220 9540 123480 9640
rect 120220 9350 120680 9540
rect 120920 9350 121380 9540
rect 121620 9350 122080 9540
rect 122320 9350 122780 9540
rect 123020 9350 123480 9540
rect 105700 9110 105800 9350
rect 104120 8940 104580 9110
rect 104820 8940 105280 9110
rect 105520 8940 105980 9110
rect 106220 8940 106680 9110
rect 106920 8940 107380 9110
rect 104120 8840 107380 8940
rect 104120 8650 104580 8840
rect 104820 8650 105280 8840
rect 105520 8650 105980 8840
rect 106220 8650 106680 8840
rect 106920 8650 107380 8840
rect 105700 8410 105800 8650
rect 104120 8240 104580 8410
rect 104820 8240 105280 8410
rect 105520 8240 105980 8410
rect 106220 8240 106680 8410
rect 106920 8240 107380 8410
rect 104120 8140 107380 8240
rect 104120 7950 104580 8140
rect 104820 7950 105280 8140
rect 105520 7950 105980 8140
rect 106220 7950 106680 8140
rect 106920 7950 107380 8140
rect 105700 7710 105800 7950
rect 104120 7540 104580 7710
rect 104820 7540 105280 7710
rect 105520 7540 105980 7710
rect 106220 7540 106680 7710
rect 106920 7540 107380 7710
rect 104120 7440 107380 7540
rect 104120 7250 104580 7440
rect 104820 7250 105280 7440
rect 105520 7250 105980 7440
rect 106220 7250 106680 7440
rect 106920 7250 107380 7440
rect 105700 7010 105800 7250
rect 104120 6840 104580 7010
rect 104820 6840 105280 7010
rect 105520 6840 105980 7010
rect 106220 6840 106680 7010
rect 106920 6840 107380 7010
rect 104120 6740 107380 6840
rect 104120 6550 104580 6740
rect 104820 6550 105280 6740
rect 105520 6550 105980 6740
rect 106220 6550 106680 6740
rect 106920 6550 107380 6740
rect 108510 6750 108590 9350
rect 108510 6690 108520 6750
rect 108580 6690 108590 6750
rect 108510 6680 108590 6690
rect 119010 6750 119090 9350
rect 121800 9110 121900 9350
rect 120220 8940 120680 9110
rect 120920 8940 121380 9110
rect 121620 8940 122080 9110
rect 122320 8940 122780 9110
rect 123020 8940 123480 9110
rect 120220 8840 123480 8940
rect 120220 8650 120680 8840
rect 120920 8650 121380 8840
rect 121620 8650 122080 8840
rect 122320 8650 122780 8840
rect 123020 8650 123480 8840
rect 121800 8410 121900 8650
rect 120220 8240 120680 8410
rect 120920 8240 121380 8410
rect 121620 8240 122080 8410
rect 122320 8240 122780 8410
rect 123020 8240 123480 8410
rect 120220 8140 123480 8240
rect 120220 7950 120680 8140
rect 120920 7950 121380 8140
rect 121620 7950 122080 8140
rect 122320 7950 122780 8140
rect 123020 7950 123480 8140
rect 121800 7710 121900 7950
rect 120220 7540 120680 7710
rect 120920 7540 121380 7710
rect 121620 7540 122080 7710
rect 122320 7540 122780 7710
rect 123020 7540 123480 7710
rect 120220 7440 123480 7540
rect 120220 7250 120680 7440
rect 120920 7250 121380 7440
rect 121620 7250 122080 7440
rect 122320 7250 122780 7440
rect 123020 7250 123480 7440
rect 121800 7010 121900 7250
rect 119010 6690 119020 6750
rect 119080 6690 119090 6750
rect 119010 6680 119090 6690
rect 120220 6840 120680 7010
rect 120920 6840 121380 7010
rect 121620 6840 122080 7010
rect 122320 6840 122780 7010
rect 123020 6840 123480 7010
rect 120220 6740 123480 6840
rect 120220 6550 120680 6740
rect 120920 6550 121380 6740
rect 121620 6550 122080 6740
rect 122320 6550 122780 6740
rect 123020 6550 123480 6740
rect 105700 6310 105800 6550
rect 121800 6310 121900 6550
rect 104120 6140 104580 6310
rect 104820 6140 105280 6310
rect 105520 6140 105980 6310
rect 106220 6140 106680 6310
rect 106920 6140 107380 6310
rect 104120 6040 107380 6140
rect 104120 5850 104580 6040
rect 104820 5850 105280 6040
rect 105520 5850 105980 6040
rect 106220 5850 106680 6040
rect 106920 5850 107380 6040
rect 120220 6140 120680 6310
rect 120920 6140 121380 6310
rect 121620 6140 122080 6310
rect 122320 6140 122780 6310
rect 123020 6140 123480 6310
rect 120220 6040 123480 6140
rect 120220 5850 120680 6040
rect 120920 5850 121380 6040
rect 121620 5850 122080 6040
rect 122320 5850 122780 6040
rect 123020 5850 123480 6040
rect 105700 5610 105800 5850
rect 121800 5610 121900 5850
rect 104120 5440 104580 5610
rect 104820 5440 105280 5610
rect 105520 5440 105980 5610
rect 106220 5440 106680 5610
rect 106920 5440 107380 5610
rect 104120 5340 107380 5440
rect 104120 5150 104580 5340
rect 104820 5150 105280 5340
rect 105520 5150 105980 5340
rect 106220 5150 106680 5340
rect 106920 5150 107380 5340
rect 120220 5440 120680 5610
rect 120920 5440 121380 5610
rect 121620 5440 122080 5610
rect 122320 5440 122780 5610
rect 123020 5440 123480 5610
rect 120220 5340 123480 5440
rect 120220 5150 120680 5340
rect 120920 5150 121380 5340
rect 121620 5150 122080 5340
rect 122320 5150 122780 5340
rect 123020 5150 123480 5340
rect 105700 4910 105800 5150
rect 121800 4910 121900 5150
rect 104120 4740 104580 4910
rect 104820 4740 105280 4910
rect 105520 4740 105980 4910
rect 106220 4740 106680 4910
rect 106920 4740 107380 4910
rect 104120 4640 107380 4740
rect 104120 4450 104580 4640
rect 104820 4450 105280 4640
rect 105520 4450 105980 4640
rect 106220 4450 106680 4640
rect 106920 4450 107380 4640
rect 120220 4740 120680 4910
rect 120920 4740 121380 4910
rect 121620 4740 122080 4910
rect 122320 4740 122780 4910
rect 123020 4740 123480 4910
rect 120220 4640 123480 4740
rect 120220 4450 120680 4640
rect 120920 4450 121380 4640
rect 121620 4450 122080 4640
rect 122320 4450 122780 4640
rect 123020 4450 123480 4640
rect 105700 4210 105800 4450
rect 121800 4210 121900 4450
rect 104120 4040 104580 4210
rect 104820 4040 105280 4210
rect 105520 4040 105980 4210
rect 106220 4040 106680 4210
rect 106920 4040 107380 4210
rect 104120 3940 107380 4040
rect 104120 3750 104580 3940
rect 104820 3750 105280 3940
rect 105520 3750 105980 3940
rect 106220 3750 106680 3940
rect 106920 3750 107380 3940
rect 120220 4040 120680 4210
rect 120920 4040 121380 4210
rect 121620 4040 122080 4210
rect 122320 4040 122780 4210
rect 123020 4040 123480 4210
rect 120220 3940 123480 4040
rect 120220 3750 120680 3940
rect 120920 3750 121380 3940
rect 121620 3750 122080 3940
rect 122320 3750 122780 3940
rect 123020 3750 123480 3940
rect 105700 3510 105800 3750
rect 121800 3510 121900 3750
rect 104120 3340 104580 3510
rect 104820 3340 105280 3510
rect 105520 3340 105980 3510
rect 106220 3340 106680 3510
rect 106920 3340 107380 3510
rect 104120 3240 107380 3340
rect 104120 3050 104580 3240
rect 104820 3050 105280 3240
rect 105520 3050 105980 3240
rect 106220 3050 106680 3240
rect 106920 3050 107380 3240
rect 107980 3430 108480 3440
rect 107980 3350 107990 3430
rect 108070 3350 108090 3430
rect 108170 3350 108190 3430
rect 108270 3350 108290 3430
rect 108370 3350 108390 3430
rect 108470 3350 108480 3430
rect 107980 3330 108480 3350
rect 107980 3250 107990 3330
rect 108070 3250 108090 3330
rect 108170 3250 108190 3330
rect 108270 3250 108290 3330
rect 108370 3250 108390 3330
rect 108470 3250 108480 3330
rect 107980 3230 108480 3250
rect 107980 3150 107990 3230
rect 108070 3150 108090 3230
rect 108170 3150 108190 3230
rect 108270 3150 108290 3230
rect 108370 3150 108390 3230
rect 108470 3150 108480 3230
rect 107980 3140 108480 3150
rect 119120 3430 119620 3440
rect 119120 3350 119130 3430
rect 119210 3350 119230 3430
rect 119310 3350 119330 3430
rect 119410 3350 119430 3430
rect 119510 3350 119530 3430
rect 119610 3350 119620 3430
rect 119120 3330 119620 3350
rect 119120 3250 119130 3330
rect 119210 3250 119230 3330
rect 119310 3250 119330 3330
rect 119410 3250 119430 3330
rect 119510 3250 119530 3330
rect 119610 3250 119620 3330
rect 119120 3230 119620 3250
rect 119120 3150 119130 3230
rect 119210 3150 119230 3230
rect 119310 3150 119330 3230
rect 119410 3150 119430 3230
rect 119510 3150 119530 3230
rect 119610 3150 119620 3230
rect 119120 3140 119620 3150
rect 120220 3340 120680 3510
rect 120920 3340 121380 3510
rect 121620 3340 122080 3510
rect 122320 3340 122780 3510
rect 123020 3340 123480 3510
rect 120220 3240 123480 3340
rect 120220 3050 120680 3240
rect 120920 3050 121380 3240
rect 121620 3050 122080 3240
rect 122320 3050 122780 3240
rect 123020 3050 123480 3240
rect 105700 2810 105800 3050
rect 121800 2810 121900 3050
rect 104120 2640 104580 2810
rect 104820 2640 105280 2810
rect 105520 2640 105980 2810
rect 106220 2640 106680 2810
rect 106920 2640 107380 2810
rect 104120 2540 107380 2640
rect 104120 2350 104580 2540
rect 104820 2350 105280 2540
rect 105520 2350 105980 2540
rect 106220 2350 106680 2540
rect 106920 2350 107380 2540
rect 120220 2640 120680 2810
rect 120920 2640 121380 2810
rect 121620 2640 122080 2810
rect 122320 2640 122780 2810
rect 123020 2640 123480 2810
rect 120220 2540 123480 2640
rect 120220 2350 120680 2540
rect 120920 2350 121380 2540
rect 121620 2350 122080 2540
rect 122320 2350 122780 2540
rect 123020 2350 123480 2540
rect 105700 2110 105800 2350
rect 121800 2110 121900 2350
rect 104120 1940 104580 2110
rect 104820 1940 105280 2110
rect 105520 1940 105980 2110
rect 106220 1940 106680 2110
rect 106920 1940 107380 2110
rect 104120 1840 107380 1940
rect 104120 1650 104580 1840
rect 104820 1650 105280 1840
rect 105520 1650 105980 1840
rect 106220 1650 106680 1840
rect 106920 1650 107380 1840
rect 120220 1940 120680 2110
rect 120920 1940 121380 2110
rect 121620 1940 122080 2110
rect 122320 1940 122780 2110
rect 123020 1940 123480 2110
rect 120220 1840 123480 1940
rect 120220 1650 120680 1840
rect 120920 1650 121380 1840
rect 121620 1650 122080 1840
rect 122320 1650 122780 1840
rect 123020 1650 123480 1840
rect 105700 1410 105800 1650
rect 121800 1410 121900 1650
rect 104120 1240 104580 1410
rect 104820 1240 105280 1410
rect 105520 1240 105980 1410
rect 106220 1240 106680 1410
rect 106920 1240 107380 1410
rect 104120 1140 107380 1240
rect 104120 950 104580 1140
rect 104820 950 105280 1140
rect 105520 950 105980 1140
rect 106220 950 106680 1140
rect 106920 950 107380 1140
rect 120220 1240 120680 1410
rect 120920 1240 121380 1410
rect 121620 1240 122080 1410
rect 122320 1240 122780 1410
rect 123020 1240 123480 1410
rect 120220 1140 123480 1240
rect 120220 950 120680 1140
rect 120920 950 121380 1140
rect 121620 950 122080 1140
rect 122320 950 122780 1140
rect 123020 950 123480 1140
rect 105700 710 105800 950
rect 121800 710 121900 950
rect 104120 540 104580 710
rect 104820 540 105280 710
rect 105520 540 105980 710
rect 106220 540 106680 710
rect 106920 540 107380 710
rect 104120 440 107380 540
rect 104120 250 104580 440
rect 104820 250 105280 440
rect 105520 250 105980 440
rect 106220 250 106680 440
rect 106920 250 107380 440
rect 120220 540 120680 710
rect 120920 540 121380 710
rect 121620 540 122080 710
rect 122320 540 122780 710
rect 123020 540 123480 710
rect 120220 440 123480 540
rect 120220 250 120680 440
rect 120920 250 121380 440
rect 121620 250 122080 440
rect 122320 250 122780 440
rect 123020 250 123480 440
rect 105700 10 105800 250
rect 121800 10 121900 250
rect 104120 -160 104580 10
rect 104820 -160 105280 10
rect 105520 -160 105980 10
rect 106220 -160 106680 10
rect 106920 -160 107380 10
rect 104120 -260 107380 -160
rect 104120 -450 104580 -260
rect 104820 -450 105280 -260
rect 105520 -450 105980 -260
rect 106220 -450 106680 -260
rect 106920 -450 107380 -260
rect 120220 -160 120680 10
rect 120920 -160 121380 10
rect 121620 -160 122080 10
rect 122320 -160 122780 10
rect 123020 -160 123480 10
rect 120220 -260 123480 -160
rect 120220 -450 120680 -260
rect 120920 -450 121380 -260
rect 121620 -450 122080 -260
rect 122320 -450 122780 -260
rect 123020 -450 123480 -260
rect 105700 -690 105800 -450
rect 121800 -690 121900 -450
rect 104120 -860 104580 -690
rect 104820 -860 105280 -690
rect 105520 -860 105980 -690
rect 106220 -860 106680 -690
rect 106920 -860 107380 -690
rect 104120 -960 107380 -860
rect 104120 -1150 104580 -960
rect 104820 -1150 105280 -960
rect 105520 -1150 105980 -960
rect 106220 -1150 106680 -960
rect 106920 -1150 107380 -960
rect 120220 -860 120680 -690
rect 120920 -860 121380 -690
rect 121620 -860 122080 -690
rect 122320 -860 122780 -690
rect 123020 -860 123480 -690
rect 120220 -960 123480 -860
rect 120220 -1150 120680 -960
rect 120920 -1150 121380 -960
rect 121620 -1150 122080 -960
rect 122320 -1150 122780 -960
rect 123020 -1150 123480 -960
rect 105700 -1390 105800 -1150
rect 121800 -1390 121900 -1150
rect 104120 -1560 104580 -1390
rect 104820 -1560 105280 -1390
rect 105520 -1560 105980 -1390
rect 106220 -1560 106680 -1390
rect 106920 -1560 107380 -1390
rect 107620 -1560 108080 -1390
rect 108320 -1560 108780 -1390
rect 109020 -1560 109480 -1390
rect 109720 -1560 110180 -1390
rect 110420 -1560 110880 -1390
rect 111120 -1560 111580 -1390
rect 111820 -1560 112280 -1390
rect 112520 -1560 112980 -1390
rect 113220 -1560 113680 -1390
rect 104120 -1660 113680 -1560
rect 104120 -1850 104580 -1660
rect 104820 -1850 105280 -1660
rect 105520 -1850 105980 -1660
rect 106220 -1850 106680 -1660
rect 106920 -1850 107380 -1660
rect 107620 -1850 108080 -1660
rect 108320 -1850 108780 -1660
rect 109020 -1850 109480 -1660
rect 109720 -1850 110180 -1660
rect 110420 -1850 110880 -1660
rect 111120 -1850 111580 -1660
rect 111820 -1850 112280 -1660
rect 112520 -1850 112980 -1660
rect 113220 -1850 113680 -1660
rect 113920 -1560 114380 -1390
rect 114620 -1560 115080 -1390
rect 115320 -1560 115780 -1390
rect 116020 -1560 116480 -1390
rect 116720 -1560 117180 -1390
rect 117420 -1560 117880 -1390
rect 118120 -1560 118580 -1390
rect 118820 -1560 119280 -1390
rect 119520 -1560 119980 -1390
rect 120220 -1560 120680 -1390
rect 120920 -1560 121380 -1390
rect 121620 -1560 122080 -1390
rect 122320 -1560 122780 -1390
rect 123020 -1560 123480 -1390
rect 113920 -1660 123480 -1560
rect 113920 -1850 114380 -1660
rect 114620 -1850 115080 -1660
rect 115320 -1850 115780 -1660
rect 116020 -1850 116480 -1660
rect 116720 -1850 117180 -1660
rect 117420 -1850 117880 -1660
rect 118120 -1850 118580 -1660
rect 118820 -1850 119280 -1660
rect 119520 -1850 119980 -1660
rect 120220 -1850 120680 -1660
rect 120920 -1850 121380 -1660
rect 121620 -1850 122080 -1660
rect 122320 -1850 122780 -1660
rect 123020 -1850 123480 -1660
rect 105700 -2090 105800 -1850
rect 106400 -2090 106500 -1850
rect 107100 -2090 107200 -1850
rect 107800 -2090 107900 -1850
rect 108500 -2090 108600 -1850
rect 109200 -2090 109300 -1850
rect 109900 -2090 110000 -1850
rect 110600 -2090 110700 -1850
rect 111300 -2090 111400 -1850
rect 112000 -2090 112100 -1850
rect 112700 -2090 112800 -1850
rect 113400 -2090 113500 -1850
rect 114100 -2090 114200 -1850
rect 114800 -2090 114900 -1850
rect 115500 -2090 115600 -1850
rect 116200 -2090 116300 -1850
rect 116900 -2090 117000 -1850
rect 117600 -2090 117700 -1850
rect 118300 -2090 118400 -1850
rect 119000 -2090 119100 -1850
rect 119700 -2090 119800 -1850
rect 120400 -2090 120500 -1850
rect 121100 -2090 121200 -1850
rect 121800 -2090 121900 -1850
rect 104120 -2260 104580 -2090
rect 104820 -2260 105280 -2090
rect 105520 -2260 105980 -2090
rect 104120 -2360 105980 -2260
rect 104120 -2550 104580 -2360
rect 104820 -2550 105280 -2360
rect 105520 -2550 105980 -2360
rect 106220 -2550 106680 -2090
rect 106920 -2550 107380 -2090
rect 107620 -2550 108080 -2090
rect 108320 -2550 108780 -2090
rect 109020 -2550 109480 -2090
rect 109720 -2550 110180 -2090
rect 110420 -2550 110880 -2090
rect 111120 -2550 111580 -2090
rect 111820 -2550 112280 -2090
rect 112520 -2550 112980 -2090
rect 113220 -2550 113680 -2090
rect 113920 -2550 114380 -2090
rect 114620 -2550 115080 -2090
rect 115320 -2550 115780 -2090
rect 116020 -2550 116480 -2090
rect 116720 -2550 117180 -2090
rect 117420 -2550 117880 -2090
rect 118120 -2550 118580 -2090
rect 118820 -2550 119280 -2090
rect 119520 -2550 119980 -2090
rect 120220 -2550 120680 -2090
rect 120920 -2550 121380 -2090
rect 121620 -2260 122080 -2090
rect 122320 -2260 122780 -2090
rect 123020 -2260 123480 -2090
rect 121620 -2360 123480 -2260
rect 121620 -2550 122080 -2360
rect 122320 -2550 122780 -2360
rect 123020 -2550 123480 -2360
<< via3 >>
rect 107990 3420 108070 3430
rect 107990 3360 108000 3420
rect 108000 3360 108060 3420
rect 108060 3360 108070 3420
rect 107990 3350 108070 3360
rect 108090 3420 108170 3430
rect 108090 3360 108100 3420
rect 108100 3360 108160 3420
rect 108160 3360 108170 3420
rect 108090 3350 108170 3360
rect 108190 3420 108270 3430
rect 108190 3360 108200 3420
rect 108200 3360 108260 3420
rect 108260 3360 108270 3420
rect 108190 3350 108270 3360
rect 108290 3420 108370 3430
rect 108290 3360 108300 3420
rect 108300 3360 108360 3420
rect 108360 3360 108370 3420
rect 108290 3350 108370 3360
rect 108390 3420 108470 3430
rect 108390 3360 108400 3420
rect 108400 3360 108460 3420
rect 108460 3360 108470 3420
rect 108390 3350 108470 3360
rect 107990 3320 108070 3330
rect 107990 3260 108000 3320
rect 108000 3260 108060 3320
rect 108060 3260 108070 3320
rect 107990 3250 108070 3260
rect 108090 3320 108170 3330
rect 108090 3260 108100 3320
rect 108100 3260 108160 3320
rect 108160 3260 108170 3320
rect 108090 3250 108170 3260
rect 108190 3320 108270 3330
rect 108190 3260 108200 3320
rect 108200 3260 108260 3320
rect 108260 3260 108270 3320
rect 108190 3250 108270 3260
rect 108290 3320 108370 3330
rect 108290 3260 108300 3320
rect 108300 3260 108360 3320
rect 108360 3260 108370 3320
rect 108290 3250 108370 3260
rect 108390 3320 108470 3330
rect 108390 3260 108400 3320
rect 108400 3260 108460 3320
rect 108460 3260 108470 3320
rect 108390 3250 108470 3260
rect 107990 3220 108070 3230
rect 107990 3160 108000 3220
rect 108000 3160 108060 3220
rect 108060 3160 108070 3220
rect 107990 3150 108070 3160
rect 108090 3220 108170 3230
rect 108090 3160 108100 3220
rect 108100 3160 108160 3220
rect 108160 3160 108170 3220
rect 108090 3150 108170 3160
rect 108190 3220 108270 3230
rect 108190 3160 108200 3220
rect 108200 3160 108260 3220
rect 108260 3160 108270 3220
rect 108190 3150 108270 3160
rect 108290 3220 108370 3230
rect 108290 3160 108300 3220
rect 108300 3160 108360 3220
rect 108360 3160 108370 3220
rect 108290 3150 108370 3160
rect 108390 3220 108470 3230
rect 108390 3160 108400 3220
rect 108400 3160 108460 3220
rect 108460 3160 108470 3220
rect 108390 3150 108470 3160
rect 119130 3420 119210 3430
rect 119130 3360 119140 3420
rect 119140 3360 119200 3420
rect 119200 3360 119210 3420
rect 119130 3350 119210 3360
rect 119230 3420 119310 3430
rect 119230 3360 119240 3420
rect 119240 3360 119300 3420
rect 119300 3360 119310 3420
rect 119230 3350 119310 3360
rect 119330 3420 119410 3430
rect 119330 3360 119340 3420
rect 119340 3360 119400 3420
rect 119400 3360 119410 3420
rect 119330 3350 119410 3360
rect 119430 3420 119510 3430
rect 119430 3360 119440 3420
rect 119440 3360 119500 3420
rect 119500 3360 119510 3420
rect 119430 3350 119510 3360
rect 119530 3420 119610 3430
rect 119530 3360 119540 3420
rect 119540 3360 119600 3420
rect 119600 3360 119610 3420
rect 119530 3350 119610 3360
rect 119130 3320 119210 3330
rect 119130 3260 119140 3320
rect 119140 3260 119200 3320
rect 119200 3260 119210 3320
rect 119130 3250 119210 3260
rect 119230 3320 119310 3330
rect 119230 3260 119240 3320
rect 119240 3260 119300 3320
rect 119300 3260 119310 3320
rect 119230 3250 119310 3260
rect 119330 3320 119410 3330
rect 119330 3260 119340 3320
rect 119340 3260 119400 3320
rect 119400 3260 119410 3320
rect 119330 3250 119410 3260
rect 119430 3320 119510 3330
rect 119430 3260 119440 3320
rect 119440 3260 119500 3320
rect 119500 3260 119510 3320
rect 119430 3250 119510 3260
rect 119530 3320 119610 3330
rect 119530 3260 119540 3320
rect 119540 3260 119600 3320
rect 119600 3260 119610 3320
rect 119530 3250 119610 3260
rect 119130 3220 119210 3230
rect 119130 3160 119140 3220
rect 119140 3160 119200 3220
rect 119200 3160 119210 3220
rect 119130 3150 119210 3160
rect 119230 3220 119310 3230
rect 119230 3160 119240 3220
rect 119240 3160 119300 3220
rect 119300 3160 119310 3220
rect 119230 3150 119310 3160
rect 119330 3220 119410 3230
rect 119330 3160 119340 3220
rect 119340 3160 119400 3220
rect 119400 3160 119410 3220
rect 119330 3150 119410 3160
rect 119430 3220 119510 3230
rect 119430 3160 119440 3220
rect 119440 3160 119500 3220
rect 119500 3160 119510 3220
rect 119430 3150 119510 3160
rect 119530 3220 119610 3230
rect 119530 3160 119540 3220
rect 119540 3160 119600 3220
rect 119600 3160 119610 3220
rect 119530 3150 119610 3160
<< mimcap >>
rect 104150 11030 104550 11180
rect 104150 10950 104310 11030
rect 104390 10950 104550 11030
rect 104150 10780 104550 10950
rect 104850 11030 105250 11180
rect 104850 10950 105010 11030
rect 105090 10950 105250 11030
rect 104850 10780 105250 10950
rect 105550 11030 105950 11180
rect 105550 10950 105710 11030
rect 105790 10950 105950 11030
rect 105550 10780 105950 10950
rect 106250 11030 106650 11180
rect 106250 10950 106410 11030
rect 106490 10950 106650 11030
rect 106250 10780 106650 10950
rect 106950 11030 107350 11180
rect 106950 10950 107110 11030
rect 107190 10950 107350 11030
rect 106950 10780 107350 10950
rect 107650 11030 108050 11180
rect 107650 10950 107810 11030
rect 107890 10950 108050 11030
rect 107650 10780 108050 10950
rect 108350 11030 108750 11180
rect 108350 10950 108510 11030
rect 108590 10950 108750 11030
rect 108350 10780 108750 10950
rect 109050 11030 109450 11180
rect 109050 10950 109210 11030
rect 109290 10950 109450 11030
rect 109050 10780 109450 10950
rect 109750 11030 110150 11180
rect 109750 10950 109910 11030
rect 109990 10950 110150 11030
rect 109750 10780 110150 10950
rect 110450 11030 110850 11180
rect 110450 10950 110610 11030
rect 110690 10950 110850 11030
rect 110450 10780 110850 10950
rect 111150 11030 111550 11180
rect 111150 10950 111310 11030
rect 111390 10950 111550 11030
rect 111150 10780 111550 10950
rect 111850 11030 112250 11180
rect 111850 10950 112010 11030
rect 112090 10950 112250 11030
rect 111850 10780 112250 10950
rect 112550 11030 112950 11180
rect 112550 10950 112710 11030
rect 112790 10950 112950 11030
rect 112550 10780 112950 10950
rect 113250 11030 113650 11180
rect 113250 10950 113410 11030
rect 113490 10950 113650 11030
rect 113250 10780 113650 10950
rect 113950 11030 114350 11180
rect 113950 10950 114110 11030
rect 114190 10950 114350 11030
rect 113950 10780 114350 10950
rect 114650 11030 115050 11180
rect 114650 10950 114810 11030
rect 114890 10950 115050 11030
rect 114650 10780 115050 10950
rect 115350 11030 115750 11180
rect 115350 10950 115510 11030
rect 115590 10950 115750 11030
rect 115350 10780 115750 10950
rect 116050 11030 116450 11180
rect 116050 10950 116210 11030
rect 116290 10950 116450 11030
rect 116050 10780 116450 10950
rect 116750 11030 117150 11180
rect 116750 10950 116910 11030
rect 116990 10950 117150 11030
rect 116750 10780 117150 10950
rect 117450 11030 117850 11180
rect 117450 10950 117610 11030
rect 117690 10950 117850 11030
rect 117450 10780 117850 10950
rect 118150 11030 118550 11180
rect 118150 10950 118310 11030
rect 118390 10950 118550 11030
rect 118150 10780 118550 10950
rect 118850 11030 119250 11180
rect 118850 10950 119010 11030
rect 119090 10950 119250 11030
rect 118850 10780 119250 10950
rect 119550 11030 119950 11180
rect 119550 10950 119710 11030
rect 119790 10950 119950 11030
rect 119550 10780 119950 10950
rect 120250 11030 120650 11180
rect 120250 10950 120410 11030
rect 120490 10950 120650 11030
rect 120250 10780 120650 10950
rect 120950 11030 121350 11180
rect 120950 10950 121110 11030
rect 121190 10950 121350 11030
rect 120950 10780 121350 10950
rect 121650 11030 122050 11180
rect 121650 10950 121810 11030
rect 121890 10950 122050 11030
rect 121650 10780 122050 10950
rect 122350 11030 122750 11180
rect 122350 10950 122510 11030
rect 122590 10950 122750 11030
rect 122350 10780 122750 10950
rect 123050 11030 123450 11180
rect 123050 10950 123210 11030
rect 123290 10950 123450 11030
rect 123050 10780 123450 10950
rect 104150 10330 104550 10480
rect 104150 10250 104310 10330
rect 104390 10250 104550 10330
rect 104150 10080 104550 10250
rect 104850 10330 105250 10480
rect 104850 10250 105010 10330
rect 105090 10250 105250 10330
rect 104850 10080 105250 10250
rect 105550 10330 105950 10480
rect 105550 10250 105710 10330
rect 105790 10250 105950 10330
rect 105550 10080 105950 10250
rect 106250 10330 106650 10480
rect 106250 10250 106410 10330
rect 106490 10250 106650 10330
rect 106250 10080 106650 10250
rect 106950 10330 107350 10480
rect 106950 10250 107110 10330
rect 107190 10250 107350 10330
rect 106950 10080 107350 10250
rect 107650 10330 108050 10480
rect 107650 10250 107810 10330
rect 107890 10250 108050 10330
rect 107650 10080 108050 10250
rect 108350 10330 108750 10480
rect 108350 10250 108510 10330
rect 108590 10250 108750 10330
rect 108350 10080 108750 10250
rect 109050 10330 109450 10480
rect 109050 10250 109210 10330
rect 109290 10250 109450 10330
rect 109050 10080 109450 10250
rect 109750 10330 110150 10480
rect 109750 10250 109910 10330
rect 109990 10250 110150 10330
rect 109750 10080 110150 10250
rect 110450 10310 110850 10480
rect 110450 10230 110610 10310
rect 110690 10230 110850 10310
rect 110450 10080 110850 10230
rect 111150 10310 111550 10480
rect 111150 10230 111310 10310
rect 111390 10230 111550 10310
rect 111150 10080 111550 10230
rect 116050 10310 116450 10480
rect 116050 10230 116210 10310
rect 116290 10230 116450 10310
rect 116050 10080 116450 10230
rect 116750 10310 117150 10480
rect 116750 10230 116910 10310
rect 116990 10230 117150 10310
rect 116750 10080 117150 10230
rect 117450 10330 117850 10480
rect 117450 10250 117610 10330
rect 117690 10250 117850 10330
rect 117450 10080 117850 10250
rect 118150 10330 118550 10480
rect 118150 10250 118310 10330
rect 118390 10250 118550 10330
rect 118150 10080 118550 10250
rect 118850 10330 119250 10480
rect 118850 10250 119010 10330
rect 119090 10250 119250 10330
rect 118850 10080 119250 10250
rect 119550 10330 119950 10480
rect 119550 10250 119710 10330
rect 119790 10250 119950 10330
rect 119550 10080 119950 10250
rect 120250 10330 120650 10480
rect 120250 10250 120410 10330
rect 120490 10250 120650 10330
rect 120250 10080 120650 10250
rect 120950 10330 121350 10480
rect 120950 10250 121110 10330
rect 121190 10250 121350 10330
rect 120950 10080 121350 10250
rect 121650 10330 122050 10480
rect 121650 10250 121810 10330
rect 121890 10250 122050 10330
rect 121650 10080 122050 10250
rect 122350 10330 122750 10480
rect 122350 10250 122510 10330
rect 122590 10250 122750 10330
rect 122350 10080 122750 10250
rect 123050 10330 123450 10480
rect 123050 10250 123210 10330
rect 123290 10250 123450 10330
rect 123050 10080 123450 10250
rect 104150 9630 104550 9780
rect 104150 9550 104310 9630
rect 104390 9550 104550 9630
rect 104150 9380 104550 9550
rect 104850 9630 105250 9780
rect 104850 9550 105010 9630
rect 105090 9550 105250 9630
rect 104850 9380 105250 9550
rect 105550 9630 105950 9780
rect 105550 9550 105710 9630
rect 105790 9550 105950 9630
rect 105550 9380 105950 9550
rect 106250 9630 106650 9780
rect 106250 9550 106410 9630
rect 106490 9550 106650 9630
rect 106250 9380 106650 9550
rect 106950 9630 107350 9780
rect 106950 9550 107110 9630
rect 107190 9550 107350 9630
rect 106950 9380 107350 9550
rect 107650 9630 108050 9780
rect 107650 9550 107810 9630
rect 107890 9550 108050 9630
rect 107650 9380 108050 9550
rect 108350 9630 108750 9780
rect 108350 9550 108510 9630
rect 108590 9550 108750 9630
rect 108350 9380 108750 9550
rect 109050 9630 109450 9780
rect 109050 9550 109210 9630
rect 109290 9550 109450 9630
rect 109050 9380 109450 9550
rect 109750 9630 110150 9780
rect 109750 9550 109910 9630
rect 109990 9550 110150 9630
rect 109750 9380 110150 9550
rect 110450 9610 110850 9780
rect 110450 9530 110610 9610
rect 110690 9530 110850 9610
rect 110450 9380 110850 9530
rect 116750 9610 117150 9780
rect 116750 9530 116910 9610
rect 116990 9530 117150 9610
rect 116750 9380 117150 9530
rect 117450 9630 117850 9780
rect 117450 9550 117610 9630
rect 117690 9550 117850 9630
rect 117450 9380 117850 9550
rect 118150 9630 118550 9780
rect 118150 9550 118310 9630
rect 118390 9550 118550 9630
rect 118150 9380 118550 9550
rect 118850 9630 119250 9780
rect 118850 9550 119010 9630
rect 119090 9550 119250 9630
rect 118850 9380 119250 9550
rect 119550 9630 119950 9780
rect 119550 9550 119710 9630
rect 119790 9550 119950 9630
rect 119550 9380 119950 9550
rect 120250 9630 120650 9780
rect 120250 9550 120410 9630
rect 120490 9550 120650 9630
rect 120250 9380 120650 9550
rect 120950 9630 121350 9780
rect 120950 9550 121110 9630
rect 121190 9550 121350 9630
rect 120950 9380 121350 9550
rect 121650 9630 122050 9780
rect 121650 9550 121810 9630
rect 121890 9550 122050 9630
rect 121650 9380 122050 9550
rect 122350 9630 122750 9780
rect 122350 9550 122510 9630
rect 122590 9550 122750 9630
rect 122350 9380 122750 9550
rect 123050 9630 123450 9780
rect 123050 9550 123210 9630
rect 123290 9550 123450 9630
rect 123050 9380 123450 9550
rect 104150 8930 104550 9080
rect 104150 8850 104310 8930
rect 104390 8850 104550 8930
rect 104150 8680 104550 8850
rect 104850 8930 105250 9080
rect 104850 8850 105010 8930
rect 105090 8850 105250 8930
rect 104850 8680 105250 8850
rect 105550 8930 105950 9080
rect 105550 8850 105710 8930
rect 105790 8850 105950 8930
rect 105550 8680 105950 8850
rect 106250 8930 106650 9080
rect 106250 8850 106410 8930
rect 106490 8850 106650 8930
rect 106250 8680 106650 8850
rect 106950 8930 107350 9080
rect 106950 8850 107110 8930
rect 107190 8850 107350 8930
rect 106950 8680 107350 8850
rect 120250 8930 120650 9080
rect 120250 8850 120410 8930
rect 120490 8850 120650 8930
rect 120250 8680 120650 8850
rect 120950 8930 121350 9080
rect 120950 8850 121110 8930
rect 121190 8850 121350 8930
rect 120950 8680 121350 8850
rect 121650 8930 122050 9080
rect 121650 8850 121810 8930
rect 121890 8850 122050 8930
rect 121650 8680 122050 8850
rect 122350 8930 122750 9080
rect 122350 8850 122510 8930
rect 122590 8850 122750 8930
rect 122350 8680 122750 8850
rect 123050 8930 123450 9080
rect 123050 8850 123210 8930
rect 123290 8850 123450 8930
rect 123050 8680 123450 8850
rect 104150 8230 104550 8380
rect 104150 8150 104310 8230
rect 104390 8150 104550 8230
rect 104150 7980 104550 8150
rect 104850 8230 105250 8380
rect 104850 8150 105010 8230
rect 105090 8150 105250 8230
rect 104850 7980 105250 8150
rect 105550 8230 105950 8380
rect 105550 8150 105710 8230
rect 105790 8150 105950 8230
rect 105550 7980 105950 8150
rect 106250 8230 106650 8380
rect 106250 8150 106410 8230
rect 106490 8150 106650 8230
rect 106250 7980 106650 8150
rect 106950 8230 107350 8380
rect 106950 8150 107110 8230
rect 107190 8150 107350 8230
rect 106950 7980 107350 8150
rect 120250 8230 120650 8380
rect 120250 8150 120410 8230
rect 120490 8150 120650 8230
rect 120250 7980 120650 8150
rect 120950 8230 121350 8380
rect 120950 8150 121110 8230
rect 121190 8150 121350 8230
rect 120950 7980 121350 8150
rect 121650 8230 122050 8380
rect 121650 8150 121810 8230
rect 121890 8150 122050 8230
rect 121650 7980 122050 8150
rect 122350 8230 122750 8380
rect 122350 8150 122510 8230
rect 122590 8150 122750 8230
rect 122350 7980 122750 8150
rect 123050 8230 123450 8380
rect 123050 8150 123210 8230
rect 123290 8150 123450 8230
rect 123050 7980 123450 8150
rect 104150 7530 104550 7680
rect 104150 7450 104310 7530
rect 104390 7450 104550 7530
rect 104150 7280 104550 7450
rect 104850 7530 105250 7680
rect 104850 7450 105010 7530
rect 105090 7450 105250 7530
rect 104850 7280 105250 7450
rect 105550 7530 105950 7680
rect 105550 7450 105710 7530
rect 105790 7450 105950 7530
rect 105550 7280 105950 7450
rect 106250 7530 106650 7680
rect 106250 7450 106410 7530
rect 106490 7450 106650 7530
rect 106250 7280 106650 7450
rect 106950 7530 107350 7680
rect 106950 7450 107110 7530
rect 107190 7450 107350 7530
rect 106950 7280 107350 7450
rect 120250 7530 120650 7680
rect 120250 7450 120410 7530
rect 120490 7450 120650 7530
rect 120250 7280 120650 7450
rect 120950 7530 121350 7680
rect 120950 7450 121110 7530
rect 121190 7450 121350 7530
rect 120950 7280 121350 7450
rect 121650 7530 122050 7680
rect 121650 7450 121810 7530
rect 121890 7450 122050 7530
rect 121650 7280 122050 7450
rect 122350 7530 122750 7680
rect 122350 7450 122510 7530
rect 122590 7450 122750 7530
rect 122350 7280 122750 7450
rect 123050 7530 123450 7680
rect 123050 7450 123210 7530
rect 123290 7450 123450 7530
rect 123050 7280 123450 7450
rect 104150 6830 104550 6980
rect 104150 6750 104310 6830
rect 104390 6750 104550 6830
rect 104150 6580 104550 6750
rect 104850 6830 105250 6980
rect 104850 6750 105010 6830
rect 105090 6750 105250 6830
rect 104850 6580 105250 6750
rect 105550 6830 105950 6980
rect 105550 6750 105710 6830
rect 105790 6750 105950 6830
rect 105550 6580 105950 6750
rect 106250 6830 106650 6980
rect 106250 6750 106410 6830
rect 106490 6750 106650 6830
rect 106250 6580 106650 6750
rect 106950 6830 107350 6980
rect 106950 6750 107110 6830
rect 107190 6750 107350 6830
rect 106950 6580 107350 6750
rect 120250 6830 120650 6980
rect 120250 6750 120410 6830
rect 120490 6750 120650 6830
rect 120250 6580 120650 6750
rect 120950 6830 121350 6980
rect 120950 6750 121110 6830
rect 121190 6750 121350 6830
rect 120950 6580 121350 6750
rect 121650 6830 122050 6980
rect 121650 6750 121810 6830
rect 121890 6750 122050 6830
rect 121650 6580 122050 6750
rect 122350 6830 122750 6980
rect 122350 6750 122510 6830
rect 122590 6750 122750 6830
rect 122350 6580 122750 6750
rect 123050 6830 123450 6980
rect 123050 6750 123210 6830
rect 123290 6750 123450 6830
rect 123050 6580 123450 6750
rect 104150 6130 104550 6280
rect 104150 6050 104310 6130
rect 104390 6050 104550 6130
rect 104150 5880 104550 6050
rect 104850 6130 105250 6280
rect 104850 6050 105010 6130
rect 105090 6050 105250 6130
rect 104850 5880 105250 6050
rect 105550 6130 105950 6280
rect 105550 6050 105710 6130
rect 105790 6050 105950 6130
rect 105550 5880 105950 6050
rect 106250 6130 106650 6280
rect 106250 6050 106410 6130
rect 106490 6050 106650 6130
rect 106250 5880 106650 6050
rect 106950 6130 107350 6280
rect 106950 6050 107110 6130
rect 107190 6050 107350 6130
rect 106950 5880 107350 6050
rect 120250 6130 120650 6280
rect 120250 6050 120410 6130
rect 120490 6050 120650 6130
rect 120250 5880 120650 6050
rect 120950 6130 121350 6280
rect 120950 6050 121110 6130
rect 121190 6050 121350 6130
rect 120950 5880 121350 6050
rect 121650 6130 122050 6280
rect 121650 6050 121810 6130
rect 121890 6050 122050 6130
rect 121650 5880 122050 6050
rect 122350 6130 122750 6280
rect 122350 6050 122510 6130
rect 122590 6050 122750 6130
rect 122350 5880 122750 6050
rect 123050 6130 123450 6280
rect 123050 6050 123210 6130
rect 123290 6050 123450 6130
rect 123050 5880 123450 6050
rect 104150 5430 104550 5580
rect 104150 5350 104310 5430
rect 104390 5350 104550 5430
rect 104150 5180 104550 5350
rect 104850 5430 105250 5580
rect 104850 5350 105010 5430
rect 105090 5350 105250 5430
rect 104850 5180 105250 5350
rect 105550 5430 105950 5580
rect 105550 5350 105710 5430
rect 105790 5350 105950 5430
rect 105550 5180 105950 5350
rect 106250 5430 106650 5580
rect 106250 5350 106410 5430
rect 106490 5350 106650 5430
rect 106250 5180 106650 5350
rect 106950 5430 107350 5580
rect 106950 5350 107110 5430
rect 107190 5350 107350 5430
rect 106950 5180 107350 5350
rect 120250 5430 120650 5580
rect 120250 5350 120410 5430
rect 120490 5350 120650 5430
rect 120250 5180 120650 5350
rect 120950 5430 121350 5580
rect 120950 5350 121110 5430
rect 121190 5350 121350 5430
rect 120950 5180 121350 5350
rect 121650 5430 122050 5580
rect 121650 5350 121810 5430
rect 121890 5350 122050 5430
rect 121650 5180 122050 5350
rect 122350 5430 122750 5580
rect 122350 5350 122510 5430
rect 122590 5350 122750 5430
rect 122350 5180 122750 5350
rect 123050 5430 123450 5580
rect 123050 5350 123210 5430
rect 123290 5350 123450 5430
rect 123050 5180 123450 5350
rect 104150 4730 104550 4880
rect 104150 4650 104310 4730
rect 104390 4650 104550 4730
rect 104150 4480 104550 4650
rect 104850 4730 105250 4880
rect 104850 4650 105010 4730
rect 105090 4650 105250 4730
rect 104850 4480 105250 4650
rect 105550 4730 105950 4880
rect 105550 4650 105710 4730
rect 105790 4650 105950 4730
rect 105550 4480 105950 4650
rect 106250 4730 106650 4880
rect 106250 4650 106410 4730
rect 106490 4650 106650 4730
rect 106250 4480 106650 4650
rect 106950 4730 107350 4880
rect 106950 4650 107110 4730
rect 107190 4650 107350 4730
rect 106950 4480 107350 4650
rect 120250 4730 120650 4880
rect 120250 4650 120410 4730
rect 120490 4650 120650 4730
rect 120250 4480 120650 4650
rect 120950 4730 121350 4880
rect 120950 4650 121110 4730
rect 121190 4650 121350 4730
rect 120950 4480 121350 4650
rect 121650 4730 122050 4880
rect 121650 4650 121810 4730
rect 121890 4650 122050 4730
rect 121650 4480 122050 4650
rect 122350 4730 122750 4880
rect 122350 4650 122510 4730
rect 122590 4650 122750 4730
rect 122350 4480 122750 4650
rect 123050 4730 123450 4880
rect 123050 4650 123210 4730
rect 123290 4650 123450 4730
rect 123050 4480 123450 4650
rect 104150 4030 104550 4180
rect 104150 3950 104310 4030
rect 104390 3950 104550 4030
rect 104150 3780 104550 3950
rect 104850 4030 105250 4180
rect 104850 3950 105010 4030
rect 105090 3950 105250 4030
rect 104850 3780 105250 3950
rect 105550 4030 105950 4180
rect 105550 3950 105710 4030
rect 105790 3950 105950 4030
rect 105550 3780 105950 3950
rect 106250 4030 106650 4180
rect 106250 3950 106410 4030
rect 106490 3950 106650 4030
rect 106250 3780 106650 3950
rect 106950 4030 107350 4180
rect 106950 3950 107110 4030
rect 107190 3950 107350 4030
rect 106950 3780 107350 3950
rect 120250 4030 120650 4180
rect 120250 3950 120410 4030
rect 120490 3950 120650 4030
rect 120250 3780 120650 3950
rect 120950 4030 121350 4180
rect 120950 3950 121110 4030
rect 121190 3950 121350 4030
rect 120950 3780 121350 3950
rect 121650 4030 122050 4180
rect 121650 3950 121810 4030
rect 121890 3950 122050 4030
rect 121650 3780 122050 3950
rect 122350 4030 122750 4180
rect 122350 3950 122510 4030
rect 122590 3950 122750 4030
rect 122350 3780 122750 3950
rect 123050 4030 123450 4180
rect 123050 3950 123210 4030
rect 123290 3950 123450 4030
rect 123050 3780 123450 3950
rect 104150 3330 104550 3480
rect 104150 3250 104310 3330
rect 104390 3250 104550 3330
rect 104150 3080 104550 3250
rect 104850 3330 105250 3480
rect 104850 3250 105010 3330
rect 105090 3250 105250 3330
rect 104850 3080 105250 3250
rect 105550 3330 105950 3480
rect 105550 3250 105710 3330
rect 105790 3250 105950 3330
rect 105550 3080 105950 3250
rect 106250 3330 106650 3480
rect 106250 3250 106410 3330
rect 106490 3250 106650 3330
rect 106250 3080 106650 3250
rect 106950 3330 107350 3480
rect 106950 3250 107110 3330
rect 107190 3250 107350 3330
rect 106950 3080 107350 3250
rect 120250 3330 120650 3480
rect 120250 3250 120410 3330
rect 120490 3250 120650 3330
rect 120250 3080 120650 3250
rect 120950 3330 121350 3480
rect 120950 3250 121110 3330
rect 121190 3250 121350 3330
rect 120950 3080 121350 3250
rect 121650 3330 122050 3480
rect 121650 3250 121810 3330
rect 121890 3250 122050 3330
rect 121650 3080 122050 3250
rect 122350 3330 122750 3480
rect 122350 3250 122510 3330
rect 122590 3250 122750 3330
rect 122350 3080 122750 3250
rect 123050 3330 123450 3480
rect 123050 3250 123210 3330
rect 123290 3250 123450 3330
rect 123050 3080 123450 3250
rect 104150 2630 104550 2780
rect 104150 2550 104310 2630
rect 104390 2550 104550 2630
rect 104150 2380 104550 2550
rect 104850 2630 105250 2780
rect 104850 2550 105010 2630
rect 105090 2550 105250 2630
rect 104850 2380 105250 2550
rect 105550 2630 105950 2780
rect 105550 2550 105710 2630
rect 105790 2550 105950 2630
rect 105550 2380 105950 2550
rect 106250 2630 106650 2780
rect 106250 2550 106410 2630
rect 106490 2550 106650 2630
rect 106250 2380 106650 2550
rect 106950 2630 107350 2780
rect 106950 2550 107110 2630
rect 107190 2550 107350 2630
rect 106950 2380 107350 2550
rect 120250 2630 120650 2780
rect 120250 2550 120410 2630
rect 120490 2550 120650 2630
rect 120250 2380 120650 2550
rect 120950 2630 121350 2780
rect 120950 2550 121110 2630
rect 121190 2550 121350 2630
rect 120950 2380 121350 2550
rect 121650 2630 122050 2780
rect 121650 2550 121810 2630
rect 121890 2550 122050 2630
rect 121650 2380 122050 2550
rect 122350 2630 122750 2780
rect 122350 2550 122510 2630
rect 122590 2550 122750 2630
rect 122350 2380 122750 2550
rect 123050 2630 123450 2780
rect 123050 2550 123210 2630
rect 123290 2550 123450 2630
rect 123050 2380 123450 2550
rect 104150 1930 104550 2080
rect 104150 1850 104310 1930
rect 104390 1850 104550 1930
rect 104150 1680 104550 1850
rect 104850 1930 105250 2080
rect 104850 1850 105010 1930
rect 105090 1850 105250 1930
rect 104850 1680 105250 1850
rect 105550 1930 105950 2080
rect 105550 1850 105710 1930
rect 105790 1850 105950 1930
rect 105550 1680 105950 1850
rect 106250 1930 106650 2080
rect 106250 1850 106410 1930
rect 106490 1850 106650 1930
rect 106250 1680 106650 1850
rect 106950 1930 107350 2080
rect 106950 1850 107110 1930
rect 107190 1850 107350 1930
rect 106950 1680 107350 1850
rect 120250 1930 120650 2080
rect 120250 1850 120410 1930
rect 120490 1850 120650 1930
rect 120250 1680 120650 1850
rect 120950 1930 121350 2080
rect 120950 1850 121110 1930
rect 121190 1850 121350 1930
rect 120950 1680 121350 1850
rect 121650 1930 122050 2080
rect 121650 1850 121810 1930
rect 121890 1850 122050 1930
rect 121650 1680 122050 1850
rect 122350 1930 122750 2080
rect 122350 1850 122510 1930
rect 122590 1850 122750 1930
rect 122350 1680 122750 1850
rect 123050 1930 123450 2080
rect 123050 1850 123210 1930
rect 123290 1850 123450 1930
rect 123050 1680 123450 1850
rect 104150 1230 104550 1380
rect 104150 1150 104310 1230
rect 104390 1150 104550 1230
rect 104150 980 104550 1150
rect 104850 1230 105250 1380
rect 104850 1150 105010 1230
rect 105090 1150 105250 1230
rect 104850 980 105250 1150
rect 105550 1230 105950 1380
rect 105550 1150 105710 1230
rect 105790 1150 105950 1230
rect 105550 980 105950 1150
rect 106250 1230 106650 1380
rect 106250 1150 106410 1230
rect 106490 1150 106650 1230
rect 106250 980 106650 1150
rect 106950 1230 107350 1380
rect 106950 1150 107110 1230
rect 107190 1150 107350 1230
rect 106950 980 107350 1150
rect 120250 1230 120650 1380
rect 120250 1150 120410 1230
rect 120490 1150 120650 1230
rect 120250 980 120650 1150
rect 120950 1230 121350 1380
rect 120950 1150 121110 1230
rect 121190 1150 121350 1230
rect 120950 980 121350 1150
rect 121650 1230 122050 1380
rect 121650 1150 121810 1230
rect 121890 1150 122050 1230
rect 121650 980 122050 1150
rect 122350 1230 122750 1380
rect 122350 1150 122510 1230
rect 122590 1150 122750 1230
rect 122350 980 122750 1150
rect 123050 1230 123450 1380
rect 123050 1150 123210 1230
rect 123290 1150 123450 1230
rect 123050 980 123450 1150
rect 104150 530 104550 680
rect 104150 450 104310 530
rect 104390 450 104550 530
rect 104150 280 104550 450
rect 104850 530 105250 680
rect 104850 450 105010 530
rect 105090 450 105250 530
rect 104850 280 105250 450
rect 105550 530 105950 680
rect 105550 450 105710 530
rect 105790 450 105950 530
rect 105550 280 105950 450
rect 106250 530 106650 680
rect 106250 450 106410 530
rect 106490 450 106650 530
rect 106250 280 106650 450
rect 106950 530 107350 680
rect 106950 450 107110 530
rect 107190 450 107350 530
rect 106950 280 107350 450
rect 120250 530 120650 680
rect 120250 450 120410 530
rect 120490 450 120650 530
rect 120250 280 120650 450
rect 120950 530 121350 680
rect 120950 450 121110 530
rect 121190 450 121350 530
rect 120950 280 121350 450
rect 121650 530 122050 680
rect 121650 450 121810 530
rect 121890 450 122050 530
rect 121650 280 122050 450
rect 122350 530 122750 680
rect 122350 450 122510 530
rect 122590 450 122750 530
rect 122350 280 122750 450
rect 123050 530 123450 680
rect 123050 450 123210 530
rect 123290 450 123450 530
rect 123050 280 123450 450
rect 104150 -170 104550 -20
rect 104150 -250 104310 -170
rect 104390 -250 104550 -170
rect 104150 -420 104550 -250
rect 104850 -170 105250 -20
rect 104850 -250 105010 -170
rect 105090 -250 105250 -170
rect 104850 -420 105250 -250
rect 105550 -170 105950 -20
rect 105550 -250 105710 -170
rect 105790 -250 105950 -170
rect 105550 -420 105950 -250
rect 106250 -170 106650 -20
rect 106250 -250 106410 -170
rect 106490 -250 106650 -170
rect 106250 -420 106650 -250
rect 106950 -170 107350 -20
rect 106950 -250 107110 -170
rect 107190 -250 107350 -170
rect 106950 -420 107350 -250
rect 120250 -170 120650 -20
rect 120250 -250 120410 -170
rect 120490 -250 120650 -170
rect 120250 -420 120650 -250
rect 120950 -170 121350 -20
rect 120950 -250 121110 -170
rect 121190 -250 121350 -170
rect 120950 -420 121350 -250
rect 121650 -170 122050 -20
rect 121650 -250 121810 -170
rect 121890 -250 122050 -170
rect 121650 -420 122050 -250
rect 122350 -170 122750 -20
rect 122350 -250 122510 -170
rect 122590 -250 122750 -170
rect 122350 -420 122750 -250
rect 123050 -170 123450 -20
rect 123050 -250 123210 -170
rect 123290 -250 123450 -170
rect 123050 -420 123450 -250
rect 104150 -870 104550 -720
rect 104150 -950 104310 -870
rect 104390 -950 104550 -870
rect 104150 -1120 104550 -950
rect 104850 -870 105250 -720
rect 104850 -950 105010 -870
rect 105090 -950 105250 -870
rect 104850 -1120 105250 -950
rect 105550 -870 105950 -720
rect 105550 -950 105710 -870
rect 105790 -950 105950 -870
rect 105550 -1120 105950 -950
rect 106250 -870 106650 -720
rect 106250 -950 106410 -870
rect 106490 -950 106650 -870
rect 106250 -1120 106650 -950
rect 106950 -870 107350 -720
rect 106950 -950 107110 -870
rect 107190 -950 107350 -870
rect 106950 -1120 107350 -950
rect 120250 -870 120650 -720
rect 120250 -950 120410 -870
rect 120490 -950 120650 -870
rect 120250 -1120 120650 -950
rect 120950 -870 121350 -720
rect 120950 -950 121110 -870
rect 121190 -950 121350 -870
rect 120950 -1120 121350 -950
rect 121650 -870 122050 -720
rect 121650 -950 121810 -870
rect 121890 -950 122050 -870
rect 121650 -1120 122050 -950
rect 122350 -870 122750 -720
rect 122350 -950 122510 -870
rect 122590 -950 122750 -870
rect 122350 -1120 122750 -950
rect 123050 -870 123450 -720
rect 123050 -950 123210 -870
rect 123290 -950 123450 -870
rect 123050 -1120 123450 -950
rect 104150 -1570 104550 -1420
rect 104150 -1650 104310 -1570
rect 104390 -1650 104550 -1570
rect 104150 -1820 104550 -1650
rect 104850 -1570 105250 -1420
rect 104850 -1650 105010 -1570
rect 105090 -1650 105250 -1570
rect 104850 -1820 105250 -1650
rect 105550 -1570 105950 -1420
rect 105550 -1650 105710 -1570
rect 105790 -1650 105950 -1570
rect 105550 -1820 105950 -1650
rect 106250 -1570 106650 -1420
rect 106250 -1650 106410 -1570
rect 106490 -1650 106650 -1570
rect 106250 -1820 106650 -1650
rect 106950 -1570 107350 -1420
rect 106950 -1650 107110 -1570
rect 107190 -1650 107350 -1570
rect 106950 -1820 107350 -1650
rect 107650 -1570 108050 -1420
rect 107650 -1650 107810 -1570
rect 107890 -1650 108050 -1570
rect 107650 -1820 108050 -1650
rect 108350 -1570 108750 -1420
rect 108350 -1650 108510 -1570
rect 108590 -1650 108750 -1570
rect 108350 -1820 108750 -1650
rect 109050 -1570 109450 -1420
rect 109050 -1650 109210 -1570
rect 109290 -1650 109450 -1570
rect 109050 -1820 109450 -1650
rect 109750 -1570 110150 -1420
rect 109750 -1650 109910 -1570
rect 109990 -1650 110150 -1570
rect 109750 -1820 110150 -1650
rect 110450 -1570 110850 -1420
rect 110450 -1650 110610 -1570
rect 110690 -1650 110850 -1570
rect 110450 -1820 110850 -1650
rect 111150 -1570 111550 -1420
rect 111150 -1650 111310 -1570
rect 111390 -1650 111550 -1570
rect 111150 -1820 111550 -1650
rect 111850 -1570 112250 -1420
rect 111850 -1650 112010 -1570
rect 112090 -1650 112250 -1570
rect 111850 -1820 112250 -1650
rect 112550 -1570 112950 -1420
rect 112550 -1650 112710 -1570
rect 112790 -1650 112950 -1570
rect 112550 -1820 112950 -1650
rect 113250 -1570 113650 -1420
rect 113250 -1650 113410 -1570
rect 113490 -1650 113650 -1570
rect 113250 -1820 113650 -1650
rect 113950 -1570 114350 -1420
rect 113950 -1650 114110 -1570
rect 114190 -1650 114350 -1570
rect 113950 -1820 114350 -1650
rect 114650 -1570 115050 -1420
rect 114650 -1650 114810 -1570
rect 114890 -1650 115050 -1570
rect 114650 -1820 115050 -1650
rect 115350 -1570 115750 -1420
rect 115350 -1650 115510 -1570
rect 115590 -1650 115750 -1570
rect 115350 -1820 115750 -1650
rect 116050 -1570 116450 -1420
rect 116050 -1650 116210 -1570
rect 116290 -1650 116450 -1570
rect 116050 -1820 116450 -1650
rect 116750 -1570 117150 -1420
rect 116750 -1650 116910 -1570
rect 116990 -1650 117150 -1570
rect 116750 -1820 117150 -1650
rect 117450 -1570 117850 -1420
rect 117450 -1650 117610 -1570
rect 117690 -1650 117850 -1570
rect 117450 -1820 117850 -1650
rect 118150 -1570 118550 -1420
rect 118150 -1650 118310 -1570
rect 118390 -1650 118550 -1570
rect 118150 -1820 118550 -1650
rect 118850 -1570 119250 -1420
rect 118850 -1650 119010 -1570
rect 119090 -1650 119250 -1570
rect 118850 -1820 119250 -1650
rect 119550 -1570 119950 -1420
rect 119550 -1650 119710 -1570
rect 119790 -1650 119950 -1570
rect 119550 -1820 119950 -1650
rect 120250 -1570 120650 -1420
rect 120250 -1650 120410 -1570
rect 120490 -1650 120650 -1570
rect 120250 -1820 120650 -1650
rect 120950 -1570 121350 -1420
rect 120950 -1650 121110 -1570
rect 121190 -1650 121350 -1570
rect 120950 -1820 121350 -1650
rect 121650 -1570 122050 -1420
rect 121650 -1650 121810 -1570
rect 121890 -1650 122050 -1570
rect 121650 -1820 122050 -1650
rect 122350 -1570 122750 -1420
rect 122350 -1650 122510 -1570
rect 122590 -1650 122750 -1570
rect 122350 -1820 122750 -1650
rect 123050 -1570 123450 -1420
rect 123050 -1650 123210 -1570
rect 123290 -1650 123450 -1570
rect 123050 -1820 123450 -1650
rect 104150 -2270 104550 -2120
rect 104150 -2350 104310 -2270
rect 104390 -2350 104550 -2270
rect 104150 -2520 104550 -2350
rect 104850 -2270 105250 -2120
rect 104850 -2350 105010 -2270
rect 105090 -2350 105250 -2270
rect 104850 -2520 105250 -2350
rect 105550 -2270 105950 -2120
rect 105550 -2350 105710 -2270
rect 105790 -2350 105950 -2270
rect 105550 -2520 105950 -2350
rect 106250 -2270 106650 -2120
rect 106250 -2350 106410 -2270
rect 106490 -2350 106650 -2270
rect 106250 -2520 106650 -2350
rect 106950 -2270 107350 -2120
rect 106950 -2350 107110 -2270
rect 107190 -2350 107350 -2270
rect 106950 -2520 107350 -2350
rect 107650 -2270 108050 -2120
rect 107650 -2350 107810 -2270
rect 107890 -2350 108050 -2270
rect 107650 -2520 108050 -2350
rect 108350 -2270 108750 -2120
rect 108350 -2350 108510 -2270
rect 108590 -2350 108750 -2270
rect 108350 -2520 108750 -2350
rect 109050 -2270 109450 -2120
rect 109050 -2350 109210 -2270
rect 109290 -2350 109450 -2270
rect 109050 -2520 109450 -2350
rect 109750 -2270 110150 -2120
rect 109750 -2350 109910 -2270
rect 109990 -2350 110150 -2270
rect 109750 -2520 110150 -2350
rect 110450 -2270 110850 -2120
rect 110450 -2350 110610 -2270
rect 110690 -2350 110850 -2270
rect 110450 -2520 110850 -2350
rect 111150 -2270 111550 -2120
rect 111150 -2350 111310 -2270
rect 111390 -2350 111550 -2270
rect 111150 -2520 111550 -2350
rect 111850 -2270 112250 -2120
rect 111850 -2350 112010 -2270
rect 112090 -2350 112250 -2270
rect 111850 -2520 112250 -2350
rect 112550 -2270 112950 -2120
rect 112550 -2350 112710 -2270
rect 112790 -2350 112950 -2270
rect 112550 -2520 112950 -2350
rect 113250 -2270 113650 -2120
rect 113250 -2350 113410 -2270
rect 113490 -2350 113650 -2270
rect 113250 -2520 113650 -2350
rect 113950 -2270 114350 -2120
rect 113950 -2350 114110 -2270
rect 114190 -2350 114350 -2270
rect 113950 -2520 114350 -2350
rect 114650 -2270 115050 -2120
rect 114650 -2350 114810 -2270
rect 114890 -2350 115050 -2270
rect 114650 -2520 115050 -2350
rect 115350 -2270 115750 -2120
rect 115350 -2350 115510 -2270
rect 115590 -2350 115750 -2270
rect 115350 -2520 115750 -2350
rect 116050 -2270 116450 -2120
rect 116050 -2350 116210 -2270
rect 116290 -2350 116450 -2270
rect 116050 -2520 116450 -2350
rect 116750 -2270 117150 -2120
rect 116750 -2350 116910 -2270
rect 116990 -2350 117150 -2270
rect 116750 -2520 117150 -2350
rect 117450 -2270 117850 -2120
rect 117450 -2350 117610 -2270
rect 117690 -2350 117850 -2270
rect 117450 -2520 117850 -2350
rect 118150 -2270 118550 -2120
rect 118150 -2350 118310 -2270
rect 118390 -2350 118550 -2270
rect 118150 -2520 118550 -2350
rect 118850 -2270 119250 -2120
rect 118850 -2350 119010 -2270
rect 119090 -2350 119250 -2270
rect 118850 -2520 119250 -2350
rect 119550 -2270 119950 -2120
rect 119550 -2350 119710 -2270
rect 119790 -2350 119950 -2270
rect 119550 -2520 119950 -2350
rect 120250 -2270 120650 -2120
rect 120250 -2350 120410 -2270
rect 120490 -2350 120650 -2270
rect 120250 -2520 120650 -2350
rect 120950 -2270 121350 -2120
rect 120950 -2350 121110 -2270
rect 121190 -2350 121350 -2270
rect 120950 -2520 121350 -2350
rect 121650 -2270 122050 -2120
rect 121650 -2350 121810 -2270
rect 121890 -2350 122050 -2270
rect 121650 -2520 122050 -2350
rect 122350 -2270 122750 -2120
rect 122350 -2350 122510 -2270
rect 122590 -2350 122750 -2270
rect 122350 -2520 122750 -2350
rect 123050 -2270 123450 -2120
rect 123050 -2350 123210 -2270
rect 123290 -2350 123450 -2270
rect 123050 -2520 123450 -2350
<< mimcapcontact >>
rect 104310 10950 104390 11030
rect 105010 10950 105090 11030
rect 105710 10950 105790 11030
rect 106410 10950 106490 11030
rect 107110 10950 107190 11030
rect 107810 10950 107890 11030
rect 108510 10950 108590 11030
rect 109210 10950 109290 11030
rect 109910 10950 109990 11030
rect 110610 10950 110690 11030
rect 111310 10950 111390 11030
rect 112010 10950 112090 11030
rect 112710 10950 112790 11030
rect 113410 10950 113490 11030
rect 114110 10950 114190 11030
rect 114810 10950 114890 11030
rect 115510 10950 115590 11030
rect 116210 10950 116290 11030
rect 116910 10950 116990 11030
rect 117610 10950 117690 11030
rect 118310 10950 118390 11030
rect 119010 10950 119090 11030
rect 119710 10950 119790 11030
rect 120410 10950 120490 11030
rect 121110 10950 121190 11030
rect 121810 10950 121890 11030
rect 122510 10950 122590 11030
rect 123210 10950 123290 11030
rect 104310 10250 104390 10330
rect 105010 10250 105090 10330
rect 105710 10250 105790 10330
rect 106410 10250 106490 10330
rect 107110 10250 107190 10330
rect 107810 10250 107890 10330
rect 108510 10250 108590 10330
rect 109210 10250 109290 10330
rect 109910 10250 109990 10330
rect 110610 10230 110690 10310
rect 111310 10230 111390 10310
rect 116210 10230 116290 10310
rect 116910 10230 116990 10310
rect 117610 10250 117690 10330
rect 118310 10250 118390 10330
rect 119010 10250 119090 10330
rect 119710 10250 119790 10330
rect 120410 10250 120490 10330
rect 121110 10250 121190 10330
rect 121810 10250 121890 10330
rect 122510 10250 122590 10330
rect 123210 10250 123290 10330
rect 104310 9550 104390 9630
rect 105010 9550 105090 9630
rect 105710 9550 105790 9630
rect 106410 9550 106490 9630
rect 107110 9550 107190 9630
rect 107810 9550 107890 9630
rect 108510 9550 108590 9630
rect 109210 9550 109290 9630
rect 109910 9550 109990 9630
rect 110610 9530 110690 9610
rect 116910 9530 116990 9610
rect 117610 9550 117690 9630
rect 118310 9550 118390 9630
rect 119010 9550 119090 9630
rect 119710 9550 119790 9630
rect 120410 9550 120490 9630
rect 121110 9550 121190 9630
rect 121810 9550 121890 9630
rect 122510 9550 122590 9630
rect 123210 9550 123290 9630
rect 104310 8850 104390 8930
rect 105010 8850 105090 8930
rect 105710 8850 105790 8930
rect 106410 8850 106490 8930
rect 107110 8850 107190 8930
rect 120410 8850 120490 8930
rect 121110 8850 121190 8930
rect 121810 8850 121890 8930
rect 122510 8850 122590 8930
rect 123210 8850 123290 8930
rect 104310 8150 104390 8230
rect 105010 8150 105090 8230
rect 105710 8150 105790 8230
rect 106410 8150 106490 8230
rect 107110 8150 107190 8230
rect 120410 8150 120490 8230
rect 121110 8150 121190 8230
rect 121810 8150 121890 8230
rect 122510 8150 122590 8230
rect 123210 8150 123290 8230
rect 104310 7450 104390 7530
rect 105010 7450 105090 7530
rect 105710 7450 105790 7530
rect 106410 7450 106490 7530
rect 107110 7450 107190 7530
rect 120410 7450 120490 7530
rect 121110 7450 121190 7530
rect 121810 7450 121890 7530
rect 122510 7450 122590 7530
rect 123210 7450 123290 7530
rect 104310 6750 104390 6830
rect 105010 6750 105090 6830
rect 105710 6750 105790 6830
rect 106410 6750 106490 6830
rect 107110 6750 107190 6830
rect 120410 6750 120490 6830
rect 121110 6750 121190 6830
rect 121810 6750 121890 6830
rect 122510 6750 122590 6830
rect 123210 6750 123290 6830
rect 104310 6050 104390 6130
rect 105010 6050 105090 6130
rect 105710 6050 105790 6130
rect 106410 6050 106490 6130
rect 107110 6050 107190 6130
rect 120410 6050 120490 6130
rect 121110 6050 121190 6130
rect 121810 6050 121890 6130
rect 122510 6050 122590 6130
rect 123210 6050 123290 6130
rect 104310 5350 104390 5430
rect 105010 5350 105090 5430
rect 105710 5350 105790 5430
rect 106410 5350 106490 5430
rect 107110 5350 107190 5430
rect 120410 5350 120490 5430
rect 121110 5350 121190 5430
rect 121810 5350 121890 5430
rect 122510 5350 122590 5430
rect 123210 5350 123290 5430
rect 104310 4650 104390 4730
rect 105010 4650 105090 4730
rect 105710 4650 105790 4730
rect 106410 4650 106490 4730
rect 107110 4650 107190 4730
rect 120410 4650 120490 4730
rect 121110 4650 121190 4730
rect 121810 4650 121890 4730
rect 122510 4650 122590 4730
rect 123210 4650 123290 4730
rect 104310 3950 104390 4030
rect 105010 3950 105090 4030
rect 105710 3950 105790 4030
rect 106410 3950 106490 4030
rect 107110 3950 107190 4030
rect 120410 3950 120490 4030
rect 121110 3950 121190 4030
rect 121810 3950 121890 4030
rect 122510 3950 122590 4030
rect 123210 3950 123290 4030
rect 104310 3250 104390 3330
rect 105010 3250 105090 3330
rect 105710 3250 105790 3330
rect 106410 3250 106490 3330
rect 107110 3250 107190 3330
rect 120410 3250 120490 3330
rect 121110 3250 121190 3330
rect 121810 3250 121890 3330
rect 122510 3250 122590 3330
rect 123210 3250 123290 3330
rect 104310 2550 104390 2630
rect 105010 2550 105090 2630
rect 105710 2550 105790 2630
rect 106410 2550 106490 2630
rect 107110 2550 107190 2630
rect 120410 2550 120490 2630
rect 121110 2550 121190 2630
rect 121810 2550 121890 2630
rect 122510 2550 122590 2630
rect 123210 2550 123290 2630
rect 104310 1850 104390 1930
rect 105010 1850 105090 1930
rect 105710 1850 105790 1930
rect 106410 1850 106490 1930
rect 107110 1850 107190 1930
rect 120410 1850 120490 1930
rect 121110 1850 121190 1930
rect 121810 1850 121890 1930
rect 122510 1850 122590 1930
rect 123210 1850 123290 1930
rect 104310 1150 104390 1230
rect 105010 1150 105090 1230
rect 105710 1150 105790 1230
rect 106410 1150 106490 1230
rect 107110 1150 107190 1230
rect 120410 1150 120490 1230
rect 121110 1150 121190 1230
rect 121810 1150 121890 1230
rect 122510 1150 122590 1230
rect 123210 1150 123290 1230
rect 104310 450 104390 530
rect 105010 450 105090 530
rect 105710 450 105790 530
rect 106410 450 106490 530
rect 107110 450 107190 530
rect 120410 450 120490 530
rect 121110 450 121190 530
rect 121810 450 121890 530
rect 122510 450 122590 530
rect 123210 450 123290 530
rect 104310 -250 104390 -170
rect 105010 -250 105090 -170
rect 105710 -250 105790 -170
rect 106410 -250 106490 -170
rect 107110 -250 107190 -170
rect 120410 -250 120490 -170
rect 121110 -250 121190 -170
rect 121810 -250 121890 -170
rect 122510 -250 122590 -170
rect 123210 -250 123290 -170
rect 104310 -950 104390 -870
rect 105010 -950 105090 -870
rect 105710 -950 105790 -870
rect 106410 -950 106490 -870
rect 107110 -950 107190 -870
rect 120410 -950 120490 -870
rect 121110 -950 121190 -870
rect 121810 -950 121890 -870
rect 122510 -950 122590 -870
rect 123210 -950 123290 -870
rect 104310 -1650 104390 -1570
rect 105010 -1650 105090 -1570
rect 105710 -1650 105790 -1570
rect 106410 -1650 106490 -1570
rect 107110 -1650 107190 -1570
rect 107810 -1650 107890 -1570
rect 108510 -1650 108590 -1570
rect 109210 -1650 109290 -1570
rect 109910 -1650 109990 -1570
rect 110610 -1650 110690 -1570
rect 111310 -1650 111390 -1570
rect 112010 -1650 112090 -1570
rect 112710 -1650 112790 -1570
rect 113410 -1650 113490 -1570
rect 114110 -1650 114190 -1570
rect 114810 -1650 114890 -1570
rect 115510 -1650 115590 -1570
rect 116210 -1650 116290 -1570
rect 116910 -1650 116990 -1570
rect 117610 -1650 117690 -1570
rect 118310 -1650 118390 -1570
rect 119010 -1650 119090 -1570
rect 119710 -1650 119790 -1570
rect 120410 -1650 120490 -1570
rect 121110 -1650 121190 -1570
rect 121810 -1650 121890 -1570
rect 122510 -1650 122590 -1570
rect 123210 -1650 123290 -1570
rect 104310 -2350 104390 -2270
rect 105010 -2350 105090 -2270
rect 105710 -2350 105790 -2270
rect 106410 -2350 106490 -2270
rect 107110 -2350 107190 -2270
rect 107810 -2350 107890 -2270
rect 108510 -2350 108590 -2270
rect 109210 -2350 109290 -2270
rect 109910 -2350 109990 -2270
rect 110610 -2350 110690 -2270
rect 111310 -2350 111390 -2270
rect 112010 -2350 112090 -2270
rect 112710 -2350 112790 -2270
rect 113410 -2350 113490 -2270
rect 114110 -2350 114190 -2270
rect 114810 -2350 114890 -2270
rect 115510 -2350 115590 -2270
rect 116210 -2350 116290 -2270
rect 116910 -2350 116990 -2270
rect 117610 -2350 117690 -2270
rect 118310 -2350 118390 -2270
rect 119010 -2350 119090 -2270
rect 119710 -2350 119790 -2270
rect 120410 -2350 120490 -2270
rect 121110 -2350 121190 -2270
rect 121810 -2350 121890 -2270
rect 122510 -2350 122590 -2270
rect 123210 -2350 123290 -2270
<< metal4 >>
rect 104300 11030 113500 11040
rect 104300 10950 104310 11030
rect 104390 10950 105010 11030
rect 105090 10950 105710 11030
rect 105790 10950 106410 11030
rect 106490 10950 107110 11030
rect 107190 10950 107810 11030
rect 107890 10950 108510 11030
rect 108590 10950 109210 11030
rect 109290 10950 109910 11030
rect 109990 10950 110610 11030
rect 110690 10950 111310 11030
rect 111390 10950 112010 11030
rect 112090 10950 112710 11030
rect 112790 10950 113410 11030
rect 113490 10950 113500 11030
rect 104300 10940 113500 10950
rect 114100 11030 123300 11040
rect 114100 10950 114110 11030
rect 114190 10950 114810 11030
rect 114890 10950 115510 11030
rect 115590 10950 116210 11030
rect 116290 10950 116910 11030
rect 116990 10950 117610 11030
rect 117690 10950 118310 11030
rect 118390 10950 119010 11030
rect 119090 10950 119710 11030
rect 119790 10950 120410 11030
rect 120490 10950 121110 11030
rect 121190 10950 121810 11030
rect 121890 10950 122510 11030
rect 122590 10950 123210 11030
rect 123290 10950 123300 11030
rect 114100 10940 123300 10950
rect 105700 10340 105800 10940
rect 104300 10330 107200 10340
rect 104300 10250 104310 10330
rect 104390 10250 105010 10330
rect 105090 10250 105710 10330
rect 105790 10250 106410 10330
rect 106490 10250 107110 10330
rect 107190 10250 107200 10330
rect 104300 10240 107200 10250
rect 107800 10330 107900 10940
rect 107800 10250 107810 10330
rect 107890 10250 107900 10330
rect 105700 9640 105800 10240
rect 104300 9630 107200 9640
rect 104300 9550 104310 9630
rect 104390 9550 105010 9630
rect 105090 9550 105710 9630
rect 105790 9550 106410 9630
rect 106490 9550 107110 9630
rect 107190 9550 107200 9630
rect 104300 9540 107200 9550
rect 107800 9630 107900 10250
rect 107800 9550 107810 9630
rect 107890 9550 107900 9630
rect 107800 9540 107900 9550
rect 108500 10330 108600 10940
rect 108500 10250 108510 10330
rect 108590 10250 108600 10330
rect 108500 9630 108600 10250
rect 108500 9550 108510 9630
rect 108590 9550 108600 9630
rect 108500 9540 108600 9550
rect 109200 10330 109300 10940
rect 109200 10250 109210 10330
rect 109290 10250 109300 10330
rect 109200 9630 109300 10250
rect 109200 9550 109210 9630
rect 109290 9550 109300 9630
rect 109200 9540 109300 9550
rect 109900 10330 110000 10940
rect 109900 10250 109910 10330
rect 109990 10250 110000 10330
rect 109900 9630 110000 10250
rect 109900 9550 109910 9630
rect 109990 9550 110000 9630
rect 109900 9540 110000 9550
rect 110600 10310 110700 10940
rect 110600 10230 110610 10310
rect 110690 10230 110700 10310
rect 110600 9610 110700 10230
rect 111300 10310 111400 10940
rect 111300 10230 111310 10310
rect 111390 10230 111400 10310
rect 111300 10220 111400 10230
rect 116200 10310 116300 10940
rect 116200 10230 116210 10310
rect 116290 10230 116300 10310
rect 116200 10220 116300 10230
rect 116900 10310 117000 10940
rect 116900 10230 116910 10310
rect 116990 10230 117000 10310
rect 105700 8940 105800 9540
rect 110600 9530 110610 9610
rect 110690 9530 110700 9610
rect 110600 9520 110700 9530
rect 116900 9610 117000 10230
rect 116900 9530 116910 9610
rect 116990 9530 117000 9610
rect 117600 10330 117700 10940
rect 117600 10250 117610 10330
rect 117690 10250 117700 10330
rect 117600 9630 117700 10250
rect 117600 9550 117610 9630
rect 117690 9550 117700 9630
rect 117600 9540 117700 9550
rect 118300 10330 118400 10940
rect 118300 10250 118310 10330
rect 118390 10250 118400 10330
rect 118300 9630 118400 10250
rect 118300 9550 118310 9630
rect 118390 9550 118400 9630
rect 118300 9540 118400 9550
rect 119000 10330 119100 10940
rect 119000 10250 119010 10330
rect 119090 10250 119100 10330
rect 119000 9630 119100 10250
rect 119000 9550 119010 9630
rect 119090 9550 119100 9630
rect 119000 9540 119100 9550
rect 119700 10330 119800 10940
rect 121800 10340 121900 10940
rect 119700 10250 119710 10330
rect 119790 10250 119800 10330
rect 119700 9630 119800 10250
rect 120400 10330 123300 10340
rect 120400 10250 120410 10330
rect 120490 10250 121110 10330
rect 121190 10250 121810 10330
rect 121890 10250 122510 10330
rect 122590 10250 123210 10330
rect 123290 10250 123300 10330
rect 120400 10240 123300 10250
rect 121800 9640 121900 10240
rect 119700 9550 119710 9630
rect 119790 9550 119800 9630
rect 119700 9540 119800 9550
rect 120400 9630 123300 9640
rect 120400 9550 120410 9630
rect 120490 9550 121110 9630
rect 121190 9550 121810 9630
rect 121890 9550 122510 9630
rect 122590 9550 123210 9630
rect 123290 9550 123300 9630
rect 120400 9540 123300 9550
rect 116900 9520 117000 9530
rect 121800 8940 121900 9540
rect 104300 8930 107200 8940
rect 104300 8850 104310 8930
rect 104390 8850 105010 8930
rect 105090 8850 105710 8930
rect 105790 8850 106410 8930
rect 106490 8850 107110 8930
rect 107190 8850 107200 8930
rect 104300 8840 107200 8850
rect 120400 8930 123300 8940
rect 120400 8850 120410 8930
rect 120490 8850 121110 8930
rect 121190 8850 121810 8930
rect 121890 8850 122510 8930
rect 122590 8850 123210 8930
rect 123290 8850 123300 8930
rect 120400 8840 123300 8850
rect 105700 8240 105800 8840
rect 121800 8240 121900 8840
rect 104300 8230 107200 8240
rect 104300 8150 104310 8230
rect 104390 8150 105010 8230
rect 105090 8150 105710 8230
rect 105790 8150 106410 8230
rect 106490 8150 107110 8230
rect 107190 8150 107200 8230
rect 104300 8140 107200 8150
rect 120400 8230 123300 8240
rect 120400 8150 120410 8230
rect 120490 8150 121110 8230
rect 121190 8150 121810 8230
rect 121890 8150 122510 8230
rect 122590 8150 123210 8230
rect 123290 8150 123300 8230
rect 120400 8140 123300 8150
rect 105700 7540 105800 8140
rect 121800 7540 121900 8140
rect 104300 7530 107200 7540
rect 104300 7450 104310 7530
rect 104390 7450 105010 7530
rect 105090 7450 105710 7530
rect 105790 7450 106410 7530
rect 106490 7450 107110 7530
rect 107190 7450 107200 7530
rect 104300 7440 107200 7450
rect 120400 7530 123300 7540
rect 120400 7450 120410 7530
rect 120490 7450 121110 7530
rect 121190 7450 121810 7530
rect 121890 7450 122510 7530
rect 122590 7450 123210 7530
rect 123290 7450 123300 7530
rect 120400 7440 123300 7450
rect 105700 6840 105800 7440
rect 121800 6840 121900 7440
rect 104300 6830 107200 6840
rect 104300 6750 104310 6830
rect 104390 6750 105010 6830
rect 105090 6750 105710 6830
rect 105790 6750 106410 6830
rect 106490 6750 107110 6830
rect 107190 6750 107200 6830
rect 104300 6740 107200 6750
rect 120400 6830 123300 6840
rect 120400 6750 120410 6830
rect 120490 6750 121110 6830
rect 121190 6750 121810 6830
rect 121890 6750 122510 6830
rect 122590 6750 123210 6830
rect 123290 6750 123300 6830
rect 120400 6740 123300 6750
rect 105700 6140 105800 6740
rect 121800 6140 121900 6740
rect 104300 6130 107200 6140
rect 104300 6050 104310 6130
rect 104390 6050 105010 6130
rect 105090 6050 105710 6130
rect 105790 6050 106410 6130
rect 106490 6050 107110 6130
rect 107190 6050 107200 6130
rect 104300 6040 107200 6050
rect 120400 6130 123300 6140
rect 120400 6050 120410 6130
rect 120490 6050 121110 6130
rect 121190 6050 121810 6130
rect 121890 6050 122510 6130
rect 122590 6050 123210 6130
rect 123290 6050 123300 6130
rect 120400 6040 123300 6050
rect 105700 5440 105800 6040
rect 121800 5440 121900 6040
rect 104300 5430 107200 5440
rect 104300 5350 104310 5430
rect 104390 5350 105010 5430
rect 105090 5350 105710 5430
rect 105790 5350 106410 5430
rect 106490 5350 107110 5430
rect 107190 5350 107200 5430
rect 104300 5340 107200 5350
rect 120400 5430 123300 5440
rect 120400 5350 120410 5430
rect 120490 5350 121110 5430
rect 121190 5350 121810 5430
rect 121890 5350 122510 5430
rect 122590 5350 123210 5430
rect 123290 5350 123300 5430
rect 120400 5340 123300 5350
rect 105700 4740 105800 5340
rect 121800 4740 121900 5340
rect 104300 4730 107200 4740
rect 104300 4650 104310 4730
rect 104390 4650 105010 4730
rect 105090 4650 105710 4730
rect 105790 4650 106410 4730
rect 106490 4650 107110 4730
rect 107190 4650 107200 4730
rect 104300 4640 107200 4650
rect 120400 4730 123300 4740
rect 120400 4650 120410 4730
rect 120490 4650 121110 4730
rect 121190 4650 121810 4730
rect 121890 4650 122510 4730
rect 122590 4650 123210 4730
rect 123290 4650 123300 4730
rect 120400 4640 123300 4650
rect 105700 4040 105800 4640
rect 121800 4040 121900 4640
rect 104300 4030 107200 4040
rect 104300 3950 104310 4030
rect 104390 3950 105010 4030
rect 105090 3950 105710 4030
rect 105790 3950 106410 4030
rect 106490 3950 107110 4030
rect 107190 3950 107200 4030
rect 104300 3940 107200 3950
rect 120400 4030 123300 4040
rect 120400 3950 120410 4030
rect 120490 3950 121110 4030
rect 121190 3950 121810 4030
rect 121890 3950 122510 4030
rect 122590 3950 123210 4030
rect 123290 3950 123300 4030
rect 120400 3940 123300 3950
rect 105700 3340 105800 3940
rect 107100 3430 108480 3440
rect 107100 3350 107990 3430
rect 108070 3350 108090 3430
rect 108170 3350 108190 3430
rect 108270 3350 108290 3430
rect 108370 3350 108390 3430
rect 108470 3350 108480 3430
rect 107100 3340 108480 3350
rect 104300 3330 108480 3340
rect 104300 3250 104310 3330
rect 104390 3250 105010 3330
rect 105090 3250 105710 3330
rect 105790 3250 106410 3330
rect 106490 3250 107110 3330
rect 107190 3250 107990 3330
rect 108070 3250 108090 3330
rect 108170 3250 108190 3330
rect 108270 3250 108290 3330
rect 108370 3250 108390 3330
rect 108470 3250 108480 3330
rect 104300 3240 108480 3250
rect 105700 2640 105800 3240
rect 107100 3230 108480 3240
rect 107100 3150 107990 3230
rect 108070 3150 108090 3230
rect 108170 3150 108190 3230
rect 108270 3150 108290 3230
rect 108370 3150 108390 3230
rect 108470 3150 108480 3230
rect 107100 3140 108480 3150
rect 119120 3430 120510 3440
rect 119120 3350 119130 3430
rect 119210 3350 119230 3430
rect 119310 3350 119330 3430
rect 119410 3350 119430 3430
rect 119510 3350 119530 3430
rect 119610 3350 120510 3430
rect 119120 3340 120510 3350
rect 121800 3340 121900 3940
rect 119120 3330 123300 3340
rect 119120 3250 119130 3330
rect 119210 3250 119230 3330
rect 119310 3250 119330 3330
rect 119410 3250 119430 3330
rect 119510 3250 119530 3330
rect 119610 3250 120410 3330
rect 120490 3250 121110 3330
rect 121190 3250 121810 3330
rect 121890 3250 122510 3330
rect 122590 3250 123210 3330
rect 123290 3250 123300 3330
rect 119120 3240 123300 3250
rect 119120 3230 120510 3240
rect 119120 3150 119130 3230
rect 119210 3150 119230 3230
rect 119310 3150 119330 3230
rect 119410 3150 119430 3230
rect 119510 3150 119530 3230
rect 119610 3150 120510 3230
rect 119120 3140 120510 3150
rect 121800 2640 121900 3240
rect 104300 2630 107200 2640
rect 104300 2550 104310 2630
rect 104390 2550 105010 2630
rect 105090 2550 105710 2630
rect 105790 2550 106410 2630
rect 106490 2550 107110 2630
rect 107190 2550 107200 2630
rect 104300 2540 107200 2550
rect 120400 2630 123300 2640
rect 120400 2550 120410 2630
rect 120490 2550 121110 2630
rect 121190 2550 121810 2630
rect 121890 2550 122510 2630
rect 122590 2550 123210 2630
rect 123290 2550 123300 2630
rect 120400 2540 123300 2550
rect 105700 1940 105800 2540
rect 121800 1940 121900 2540
rect 104300 1930 107200 1940
rect 104300 1850 104310 1930
rect 104390 1850 105010 1930
rect 105090 1850 105710 1930
rect 105790 1850 106410 1930
rect 106490 1850 107110 1930
rect 107190 1850 107200 1930
rect 104300 1840 107200 1850
rect 120400 1930 123300 1940
rect 120400 1850 120410 1930
rect 120490 1850 121110 1930
rect 121190 1850 121810 1930
rect 121890 1850 122510 1930
rect 122590 1850 123210 1930
rect 123290 1850 123300 1930
rect 120400 1840 123300 1850
rect 105700 1240 105800 1840
rect 121800 1240 121900 1840
rect 104300 1230 107200 1240
rect 104300 1150 104310 1230
rect 104390 1150 105010 1230
rect 105090 1150 105710 1230
rect 105790 1150 106410 1230
rect 106490 1150 107110 1230
rect 107190 1150 107200 1230
rect 104300 1140 107200 1150
rect 120400 1230 123300 1240
rect 120400 1150 120410 1230
rect 120490 1150 121110 1230
rect 121190 1150 121810 1230
rect 121890 1150 122510 1230
rect 122590 1150 123210 1230
rect 123290 1150 123300 1230
rect 120400 1140 123300 1150
rect 105700 540 105800 1140
rect 121800 540 121900 1140
rect 104300 530 107200 540
rect 104300 450 104310 530
rect 104390 450 105010 530
rect 105090 450 105710 530
rect 105790 450 106410 530
rect 106490 450 107110 530
rect 107190 450 107200 530
rect 104300 440 107200 450
rect 120400 530 123300 540
rect 120400 450 120410 530
rect 120490 450 121110 530
rect 121190 450 121810 530
rect 121890 450 122510 530
rect 122590 450 123210 530
rect 123290 450 123300 530
rect 120400 440 123300 450
rect 105700 -160 105800 440
rect 121800 -160 121900 440
rect 104300 -170 107200 -160
rect 104300 -250 104310 -170
rect 104390 -250 105010 -170
rect 105090 -250 105710 -170
rect 105790 -250 106410 -170
rect 106490 -250 107110 -170
rect 107190 -250 107200 -170
rect 104300 -260 107200 -250
rect 120400 -170 123300 -160
rect 120400 -250 120410 -170
rect 120490 -250 121110 -170
rect 121190 -250 121810 -170
rect 121890 -250 122510 -170
rect 122590 -250 123210 -170
rect 123290 -250 123300 -170
rect 120400 -260 123300 -250
rect 105700 -860 105800 -260
rect 121800 -860 121900 -260
rect 104300 -870 107200 -860
rect 104300 -950 104310 -870
rect 104390 -950 105010 -870
rect 105090 -950 105710 -870
rect 105790 -950 106410 -870
rect 106490 -950 107110 -870
rect 107190 -950 107200 -870
rect 104300 -960 107200 -950
rect 120400 -870 123300 -860
rect 120400 -950 120410 -870
rect 120490 -950 121110 -870
rect 121190 -950 121810 -870
rect 121890 -950 122510 -870
rect 122590 -950 123210 -870
rect 123290 -950 123300 -870
rect 120400 -960 123300 -950
rect 105700 -1560 105800 -960
rect 121800 -1560 121900 -960
rect 104300 -1570 113500 -1560
rect 104300 -1650 104310 -1570
rect 104390 -1650 105010 -1570
rect 105090 -1650 105710 -1570
rect 105790 -1650 106410 -1570
rect 106490 -1650 107110 -1570
rect 107190 -1650 107810 -1570
rect 107890 -1650 108510 -1570
rect 108590 -1650 109210 -1570
rect 109290 -1650 109910 -1570
rect 109990 -1650 110610 -1570
rect 110690 -1650 111310 -1570
rect 111390 -1650 112010 -1570
rect 112090 -1650 112710 -1570
rect 112790 -1650 113410 -1570
rect 113490 -1650 113500 -1570
rect 104300 -1660 113500 -1650
rect 105700 -2260 105800 -1660
rect 104300 -2270 105800 -2260
rect 104300 -2350 104310 -2270
rect 104390 -2350 105010 -2270
rect 105090 -2350 105710 -2270
rect 105790 -2350 105800 -2270
rect 104300 -2360 105800 -2350
rect 106400 -2270 106500 -1660
rect 106400 -2350 106410 -2270
rect 106490 -2350 106500 -2270
rect 106400 -2360 106500 -2350
rect 107100 -2270 107200 -1660
rect 107100 -2350 107110 -2270
rect 107190 -2350 107200 -2270
rect 107100 -2360 107200 -2350
rect 107800 -2270 107900 -1660
rect 107800 -2350 107810 -2270
rect 107890 -2350 107900 -2270
rect 107800 -2360 107900 -2350
rect 108500 -2270 108600 -1660
rect 108500 -2350 108510 -2270
rect 108590 -2350 108600 -2270
rect 108500 -2360 108600 -2350
rect 109200 -2270 109300 -1660
rect 109200 -2350 109210 -2270
rect 109290 -2350 109300 -2270
rect 109200 -2360 109300 -2350
rect 109900 -2270 110000 -1660
rect 109900 -2350 109910 -2270
rect 109990 -2350 110000 -2270
rect 109900 -2360 110000 -2350
rect 110600 -2270 110700 -1660
rect 110600 -2350 110610 -2270
rect 110690 -2350 110700 -2270
rect 110600 -2360 110700 -2350
rect 111300 -2270 111400 -1660
rect 111300 -2350 111310 -2270
rect 111390 -2350 111400 -2270
rect 111300 -2360 111400 -2350
rect 112000 -2270 112100 -1660
rect 112000 -2350 112010 -2270
rect 112090 -2350 112100 -2270
rect 112000 -2360 112100 -2350
rect 112700 -2270 112800 -1660
rect 112700 -2350 112710 -2270
rect 112790 -2350 112800 -2270
rect 112700 -2360 112800 -2350
rect 113400 -2270 113500 -1660
rect 113400 -2350 113410 -2270
rect 113490 -2350 113500 -2270
rect 113400 -2360 113500 -2350
rect 114100 -1570 123300 -1560
rect 114100 -1650 114110 -1570
rect 114190 -1650 114810 -1570
rect 114890 -1650 115510 -1570
rect 115590 -1650 116210 -1570
rect 116290 -1650 116910 -1570
rect 116990 -1650 117610 -1570
rect 117690 -1650 118310 -1570
rect 118390 -1650 119010 -1570
rect 119090 -1650 119710 -1570
rect 119790 -1650 120410 -1570
rect 120490 -1650 121110 -1570
rect 121190 -1650 121810 -1570
rect 121890 -1650 122510 -1570
rect 122590 -1650 123210 -1570
rect 123290 -1650 123300 -1570
rect 114100 -1660 123300 -1650
rect 114100 -2270 114200 -1660
rect 114100 -2350 114110 -2270
rect 114190 -2350 114200 -2270
rect 114100 -2360 114200 -2350
rect 114800 -2270 114900 -1660
rect 114800 -2350 114810 -2270
rect 114890 -2350 114900 -2270
rect 114800 -2360 114900 -2350
rect 115500 -2270 115600 -1660
rect 115500 -2350 115510 -2270
rect 115590 -2350 115600 -2270
rect 115500 -2360 115600 -2350
rect 116200 -2270 116300 -1660
rect 116200 -2350 116210 -2270
rect 116290 -2350 116300 -2270
rect 116200 -2360 116300 -2350
rect 116900 -2270 117000 -1660
rect 116900 -2350 116910 -2270
rect 116990 -2350 117000 -2270
rect 116900 -2360 117000 -2350
rect 117600 -2270 117700 -1660
rect 117600 -2350 117610 -2270
rect 117690 -2350 117700 -2270
rect 117600 -2360 117700 -2350
rect 118300 -2270 118400 -1660
rect 118300 -2350 118310 -2270
rect 118390 -2350 118400 -2270
rect 118300 -2360 118400 -2350
rect 119000 -2270 119100 -1660
rect 119000 -2350 119010 -2270
rect 119090 -2350 119100 -2270
rect 119000 -2360 119100 -2350
rect 119700 -2270 119800 -1660
rect 119700 -2350 119710 -2270
rect 119790 -2350 119800 -2270
rect 119700 -2360 119800 -2350
rect 120400 -2270 120500 -1660
rect 120400 -2350 120410 -2270
rect 120490 -2350 120500 -2270
rect 120400 -2360 120500 -2350
rect 121100 -2270 121200 -1660
rect 121100 -2350 121110 -2270
rect 121190 -2350 121200 -2270
rect 121100 -2360 121200 -2350
rect 121800 -2260 121900 -1660
rect 121800 -2270 123300 -2260
rect 121800 -2350 121810 -2270
rect 121890 -2350 122510 -2270
rect 122590 -2350 123210 -2270
rect 123290 -2350 123300 -2270
rect 121800 -2360 123300 -2350
<< labels >>
flabel metal1 113890 1310 113890 1310 7 FreeSans 480 0 -160 0 V_tail_gate
port 11 w
flabel metal2 115540 2560 115540 2560 3 FreeSans 480 0 160 0 VIN-
flabel metal2 112060 2560 112060 2560 7 FreeSans 480 0 -160 0 VIN+
flabel metal1 114860 2650 114860 2650 3 FreeSans 480 0 160 0 VD1
flabel metal1 112740 2650 112740 2650 7 FreeSans 480 0 -160 0 VD2
flabel metal2 114910 4930 114910 4930 7 FreeSans 480 0 -160 0 X
flabel metal2 115050 5330 115050 5330 1 FreeSans 480 0 0 160 err_amp_out
flabel metal2 114000 5420 114000 5420 3 FreeSans 480 0 160 0 err_amp_mir
flabel metal2 112730 5630 112730 5630 7 FreeSans 480 0 -160 0 V_err_amp_ref
port 12 w
flabel metal2 115160 5550 115160 5550 1 FreeSans 480 0 0 320 V_tot
flabel metal1 112690 4910 112690 4910 3 FreeSans 480 0 160 0 Y
flabel metal2 114360 6410 114360 6410 3 FreeSans 480 0 160 0 V_err_p
flabel metal1 113240 6410 113240 6410 7 FreeSans 480 0 -160 0 V_err_mir_p
flabel metal2 114250 5770 114250 5770 3 FreeSans 480 0 160 0 V_err_gate
port 13 e
flabel metal2 113600 -400 113600 -400 1 FreeSans 480 0 0 160 Vb1_2
flabel metal2 112920 -110 112920 -110 1 FreeSans 480 0 0 160 V_p_mir
flabel metal2 109010 3330 109010 3330 1 FreeSans 480 0 0 160 V_CMFB_S3
port 3 n
flabel metal2 109100 2960 109100 2960 1 FreeSans 480 0 0 160 V_CMFB_S4
port 8 n
flabel metal1 118500 2960 118500 2960 1 FreeSans 480 0 0 160 V_CMFB_S2
port 7 n
flabel metal1 118590 3330 118590 3330 1 FreeSans 480 0 0 160 V_CMFB_S1
port 2 n
flabel metal3 108510 6870 108510 6870 7 FreeSans 480 0 -160 0 cap_res_Y
flabel metal3 119080 6870 119080 6870 3 FreeSans 480 0 160 0 cap_res_X
flabel metal1 114440 1250 114440 1250 3 FreeSans 480 0 160 0 V_source
flabel metal1 119410 810 119410 810 5 FreeSans 480 0 0 -160 VOUT-
port 9 s
flabel metal2 115440 1100 115440 1100 5 FreeSans 400 0 0 -160 V_b_2nd_stage
flabel metal2 108190 810 108190 810 5 FreeSans 480 0 0 -160 VOUT+
port 10 s
flabel metal2 113800 3870 113800 3870 5 FreeSans 480 0 0 -160 Vb1
flabel metal1 113710 6870 113710 6870 5 FreeSans 400 0 0 -160 Vb2
port 5 s
flabel metal2 114000 6770 114000 6770 5 FreeSans 400 0 0 -160 Vb3
port 4 s
flabel metal2 111560 7900 111560 7900 5 FreeSans 480 0 0 -160 VD4
flabel metal2 116080 7900 116080 7900 5 FreeSans 480 0 0 -160 VD3
flabel metal2 112910 10120 112910 10120 1 FreeSans 480 0 0 160 Vb2_2
flabel metal2 114730 10120 114730 10120 1 FreeSans 480 0 0 160 Vb2_Vb3
<< end >>
