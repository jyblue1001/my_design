* PEX produced on Wed Jul  9 09:39:59 AM CEST 2025 using /foss/tools/osic-multitool/iic-pex.sh with m=3 and s=1
* NGSPICE file created from two_stage_opamp_dummy_magic.ext - technology: sky130A

.subckt two_stage_opamp_dummy_magic VDDA V_CMFB_S1 V_CMFB_S3 Vb3 Vb2 Vb1 V_CMFB_S2
+ V_CMFB_S4 VOUT- VOUT+ V_tail_gate V_err_amp_ref V_err_gate VIN+ VIN- GNDA
X0 VD4.t36 Vb2.t3 Y.t13 VD4.t35 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X1 VD1.t21 VIN-.t0 V_source.t27 GNDA.t8 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X2 VDDA.t124 Vb3.t2 VD3.t9 VDDA.t123 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X3 VOUT-.t16 X.t25 VDDA.t11 VDDA.t10 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X4 VOUT-.t19 cap_res_X.t138 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5 VOUT+.t19 cap_res_Y.t138 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6 VOUT-.t20 cap_res_X.t137 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7 VOUT+.t20 cap_res_Y.t137 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8 VOUT-.t21 cap_res_X.t136 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9 VOUT+.t21 cap_res_Y.t136 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X10 V_source.t14 V_tail_gate.t4 GNDA.t29 GNDA.t3 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X11 err_amp_out.t7 GNDA.t114 GNDA.t116 GNDA.t115 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X12 VDDA.t122 Vb3.t3 VD3.t7 VDDA.t121 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X13 VDDA.t54 X.t26 V_CMFB_S2.t10 GNDA.t0 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X14 VOUT+.t14 a_109990_5430# VDDA.t221 VDDA.t220 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=2.4 ps=12.8 w=6 l=0.15
X15 VDDA.t219 Y.t25 V_CMFB_S4.t10 GNDA.t0 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X16 VDDA.t43 V_err_gate.t12 V_err_p.t20 VDDA.t42 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X17 VDDA.t218 Y.t26 V_CMFB_S4.t9 GNDA.t0 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X18 Vb2_Vb3.t6 Vb2_Vb3.t3 Vb2_Vb3.t5 Vb2_Vb3.t4 sky130_fd_pr__pfet_01v8 ad=1.44 pd=8 as=0 ps=0 w=3.6 l=0.2
X19 VOUT+.t22 cap_res_Y.t135 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X20 VD1.t0 Vb1.t2 X.t0 GNDA.t1 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X21 VOUT-.t22 cap_res_X.t135 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X22 VOUT+.t23 cap_res_Y.t134 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X23 err_amp_mir.t16 V_tot.t4 V_err_p.t3 VDDA.t51 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X24 GNDA.t122 X.t27 V_CMFB_S1.t10 VDDA.t240 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X25 V_source.t34 VIN-.t1 VD1.t20 GNDA.t8 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X26 VOUT+.t24 cap_res_Y.t133 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X27 GNDA.t125 err_amp_mir.t17 err_amp_out.t8 GNDA.t124 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X28 GNDA.t113 GNDA.t112 VOUT+.t16 GNDA.t9 sky130_fd_pr__nfet_01v8 ad=2.8 pd=14.8 as=1.4 ps=7.4 w=7 l=0.6
X29 VD2.t21 Vb1.t3 Y.t24 GNDA.t1 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X30 VD4.t34 Vb2.t4 Y.t19 VD4.t33 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X31 VDDA.t120 Vb3.t4 VD3.t4 VDDA.t119 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X32 VOUT+.t25 cap_res_Y.t132 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X33 VOUT-.t23 cap_res_X.t134 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X34 VOUT-.t24 cap_res_X.t133 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X35 VOUT+.t26 cap_res_Y.t131 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X36 VOUT+.t27 cap_res_Y.t130 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X37 VOUT+.t28 cap_res_Y.t129 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X38 VOUT-.t25 cap_res_X.t132 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X39 VOUT-.t26 cap_res_X.t131 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X40 V_CMFB_S3.t10 Y.t27 GNDA.t67 VDDA.t217 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X41 VD3.t31 Vb2.t5 X.t20 VD3.t30 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X42 VOUT-.t15 X.t28 VDDA.t39 VDDA.t38 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X43 VDDA.t179 VDDA.t177 GNDA.t15 VDDA.t178 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X44 V_err_gate.t3 V_err_amp_ref.t0 V_err_mir_p.t4 VDDA.t27 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X45 VOUT+.t29 cap_res_Y.t128 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X46 Vb2_Vb3.t2 Vb2_Vb3.t0 Vb3.t1 Vb2_Vb3.t1 sky130_fd_pr__pfet_01v8 ad=1.44 pd=8 as=0.72 ps=4 w=3.6 l=0.2
X47 V_source.t37 V_tail_gate.t5 GNDA.t120 GNDA.t3 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X48 VOUT+.t30 cap_res_Y.t127 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X49 V_source.t11 V_tail_gate.t6 GNDA.t27 GNDA.t3 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X50 VDDA.t118 Vb3.t5 VD4.t4 VDDA.t117 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X51 VOUT+.t31 cap_res_Y.t126 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X52 VOUT+.t32 cap_res_Y.t125 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X53 VOUT+.t33 cap_res_Y.t124 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X54 VOUT+.t34 cap_res_Y.t123 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X55 VOUT-.t2 V_b_2nd_stage.t2 GNDA.t38 GNDA.t9 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X56 VDDA.t29 X.t29 V_CMFB_S2.t9 GNDA.t0 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X57 VDDA.t47 V_err_gate.t13 V_err_mir_p.t14 VDDA.t46 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X58 VOUT+.t35 cap_res_Y.t122 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X59 VOUT-.t27 cap_res_X.t130 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X60 VD3.t2 Vb3.t6 VDDA.t116 VDDA.t115 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X61 VDDA.t239 V_err_gate.t14 V_err_mir_p.t13 VDDA.t238 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X62 VD1.t4 Vb1.t4 X.t4 GNDA.t1 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X63 VOUT+.t36 cap_res_Y.t121 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X64 err_amp_mir.t15 V_tot.t5 V_err_p.t8 VDDA.t72 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X65 VOUT+.t37 cap_res_Y.t120 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X66 VDDA.t216 Y.t28 VOUT+.t13 VDDA.t215 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X67 VDDA.t82 a_111200_5430# VOUT+.t3 VDDA.t81 sky130_fd_pr__pfet_01v8 ad=2.4 pd=12.8 as=1.2 ps=6.4 w=6 l=0.15
X68 GNDA.t55 X.t30 V_CMFB_S1.t9 VDDA.t68 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X69 VDDA.t176 VDDA.t174 VDDA.t176 VDDA.t175 sky130_fd_pr__pfet_01v8 ad=0.71 pd=3.95 as=0 ps=0 w=3.55 l=0.2
X70 VOUT-.t28 cap_res_X.t129 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X71 V_source.t23 VIN+.t0 VD2.t9 GNDA.t8 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X72 VOUT+.t38 cap_res_Y.t119 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X73 VOUT+.t39 cap_res_Y.t118 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X74 VOUT+.t40 cap_res_Y.t117 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X75 GNDA.t111 GNDA.t110 V_source.t6 GNDA.t3 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=0.5 ps=2.9 w=2.5 l=0.15
X76 VDDA.t227 GNDA.t108 GNDA.t109 GNDA.t0 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=1.2 ps=6.8 w=3 l=0.15
X77 GNDA.t34 err_amp_mir.t8 err_amp_mir.t9 GNDA.t33 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X78 VOUT+.t41 cap_res_Y.t116 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X79 VDDA.t114 Vb3.t7 VD4.t10 VDDA.t113 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X80 GNDA.t107 GNDA.t105 err_amp_mir.t11 GNDA.t106 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X81 VOUT+.t42 cap_res_Y.t115 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X82 VOUT-.t29 cap_res_X.t128 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X83 VOUT-.t30 cap_res_X.t127 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X84 VOUT+.t43 cap_res_Y.t114 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X85 VOUT-.t31 cap_res_X.t126 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X86 VOUT+.t44 cap_res_Y.t113 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X87 VOUT+.t15 GNDA.t103 GNDA.t104 GNDA.t9 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=2.8 ps=14.8 w=7 l=0.6
X88 V_err_p.t19 V_err_gate.t15 VDDA.t18 VDDA.t17 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X89 VOUT+.t45 cap_res_Y.t112 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X90 VOUT-.t32 cap_res_X.t125 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X91 V_CMFB_S3.t9 Y.t29 GNDA.t69 VDDA.t214 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X92 GNDA.t102 GNDA.t101 V_tail_gate.t3 GNDA.t8 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X93 VD1.t19 VIN-.t2 V_source.t26 GNDA.t8 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X94 VOUT-.t14 X.t31 VDDA.t9 VDDA.t8 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X95 VOUT+.t46 cap_res_Y.t111 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X96 V_err_gate.t0 V_err_amp_ref.t1 V_err_mir_p.t3 VDDA.t19 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X97 VOUT+.t47 cap_res_Y.t110 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X98 VOUT-.t33 cap_res_X.t124 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X99 VOUT+.t0 V_b_2nd_stage.t3 GNDA.t10 GNDA.t9 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X100 VOUT+.t48 cap_res_Y.t109 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X101 VD3.t3 Vb3.t8 VDDA.t112 VDDA.t111 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X102 V_source.t25 V_tail_gate.t7 GNDA.t58 GNDA.t3 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X103 VOUT-.t34 cap_res_X.t123 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X104 VOUT+.t49 cap_res_Y.t108 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X105 VOUT+.t50 cap_res_Y.t107 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X106 VOUT-.t35 cap_res_X.t122 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X107 Vb3.t0 Vb2.t6 Vb2_Vb3.t10 Vb2_Vb3.t9 sky130_fd_pr__pfet_01v8 ad=0.72 pd=4 as=0.72 ps=4 w=3.6 l=0.2
X108 VOUT-.t36 cap_res_X.t121 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X109 VDDA.t14 X.t32 V_CMFB_S2.t8 GNDA.t0 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X110 VDDA.t26 V_err_gate.t16 V_err_mir_p.t12 VDDA.t25 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X111 VDDA.t23 V_err_gate.t17 V_err_p.t18 VDDA.t22 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X112 VOUT+.t18 V_b_2nd_stage.t4 GNDA.t132 GNDA.t9 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X113 err_amp_out.t4 V_err_amp_ref.t2 V_err_p.t5 VDDA.t61 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X114 VOUT-.t37 cap_res_X.t120 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X115 VOUT+.t51 cap_res_Y.t106 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X116 VDDA.t173 VDDA.t171 VD4.t37 VDDA.t172 sky130_fd_pr__pfet_01v8 ad=1.575 pd=7.9 as=0.7 ps=3.9 w=3.5 l=0.2
X117 VDDA.t213 Y.t30 VOUT+.t12 VDDA.t212 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X118 VOUT+.t52 cap_res_Y.t105 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X119 VOUT-.t38 cap_res_X.t119 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X120 GNDA.t14 X.t33 V_CMFB_S1.t8 VDDA.t12 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X121 VOUT-.t39 cap_res_X.t118 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X122 VOUT+.t53 cap_res_Y.t104 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X123 VOUT+.t54 cap_res_Y.t103 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X124 VOUT-.t40 cap_res_X.t117 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X125 VD3.t8 Vb3.t9 VDDA.t110 VDDA.t109 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X126 VOUT-.t41 cap_res_X.t116 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X127 VOUT+.t55 cap_res_Y.t102 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X128 GNDA.t53 V_tail_gate.t8 V_source.t21 GNDA.t3 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X129 X.t22 VD3.t35 VD3.t37 VD3.t36 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X130 GNDA.t129 err_amp_mir.t18 err_amp_out.t10 GNDA.t128 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X131 VOUT-.t42 cap_res_X.t115 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X132 VOUT+.t56 cap_res_Y.t101 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X133 VOUT+.t57 cap_res_Y.t100 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X134 GNDA.t30 V_b_2nd_stage.t5 VOUT-.t1 GNDA.t9 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X135 VOUT+.t58 cap_res_Y.t99 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X136 V_CMFB_S4.t8 Y.t31 VDDA.t211 GNDA.t0 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X137 GNDA.t100 GNDA.t99 VDDA.t226 GNDA.t0 sky130_fd_pr__nfet_01v8 ad=1.2 pd=6.8 as=0.6 ps=3.4 w=3 l=0.15
X138 V_err_mir_p.t11 V_err_gate.t18 VDDA.t70 VDDA.t69 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X139 VOUT+.t59 cap_res_Y.t98 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X140 VOUT-.t43 cap_res_X.t114 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X141 VOUT+.t60 cap_res_Y.t97 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X142 V_err_p.t0 V_err_amp_ref.t3 err_amp_out.t0 VDDA.t1 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X143 VOUT+.t61 cap_res_Y.t96 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X144 V_CMFB_S3.t8 Y.t32 GNDA.t68 VDDA.t210 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X145 VOUT-.t44 cap_res_X.t113 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X146 VOUT-.t45 cap_res_X.t112 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X147 VOUT+.t62 cap_res_Y.t95 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X148 VOUT-.t13 X.t34 VDDA.t76 VDDA.t75 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X149 V_p_mir.t3 VIN-.t3 V_tail_gate.t1 GNDA.t8 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X150 VD2.t8 VIN+.t1 V_source.t22 GNDA.t8 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X151 VOUT-.t46 cap_res_X.t111 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X152 V_err_gate.t9 V_tot.t6 V_err_mir_p.t19 VDDA.t80 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X153 VOUT-.t47 cap_res_X.t110 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X154 GNDA.t45 V_b_2nd_stage.t6 VOUT-.t3 GNDA.t9 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X155 VD4.t9 Vb3.t10 VDDA.t108 VDDA.t107 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X156 V_source.t10 V_tail_gate.t9 GNDA.t23 GNDA.t3 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X157 Y.t10 Vb1.t5 VD2.t20 GNDA.t1 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X158 VOUT+.t63 cap_res_Y.t94 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X159 VOUT-.t48 cap_res_X.t109 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X160 VDDA.t170 VDDA.t167 VDDA.t169 VDDA.t168 sky130_fd_pr__pfet_01v8 ad=0.252 pd=2.06 as=0 ps=0 w=0.63 l=0.2
X161 VOUT+.t64 cap_res_Y.t93 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X162 VDDA.t0 X.t35 V_CMFB_S2.t7 GNDA.t0 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X163 VDDA.t64 V_err_gate.t19 V_err_p.t17 VDDA.t63 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X164 VOUT-.t49 cap_res_X.t108 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X165 VOUT-.t50 cap_res_X.t107 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X166 VOUT+.t65 cap_res_Y.t92 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X167 VOUT-.t51 cap_res_X.t106 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X168 VOUT-.t52 cap_res_X.t105 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X169 VOUT-.t53 cap_res_X.t104 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X170 err_amp_mir.t10 VDDA.t164 VDDA.t166 VDDA.t165 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X171 VDDA.t209 Y.t33 VOUT+.t11 VDDA.t208 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X172 GNDA.t54 VDDA.t161 VDDA.t163 VDDA.t162 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X173 VOUT-.t54 cap_res_X.t103 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X174 VD4.t0 Vb3.t11 VDDA.t104 VDDA.t103 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X175 VOUT-.t55 cap_res_X.t102 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X176 GNDA.t48 V_tail_gate.t10 V_source.t17 GNDA.t3 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X177 VOUT+.t66 cap_res_Y.t91 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X178 V_CMFB_S4.t7 Y.t34 VDDA.t207 GNDA.t0 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X179 VOUT-.t56 cap_res_X.t101 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X180 VOUT-.t57 cap_res_X.t100 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X181 VOUT-.t58 cap_res_X.t99 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X182 VOUT-.t59 cap_res_X.t98 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X183 VOUT+.t67 cap_res_Y.t90 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X184 VD4.t6 Vb3.t12 VDDA.t106 VDDA.t105 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X185 VOUT-.t60 cap_res_X.t97 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X186 VOUT+.t68 cap_res_Y.t89 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X187 V_err_p.t7 V_tot.t7 err_amp_mir.t14 VDDA.t65 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X188 X.t7 Vb1.t6 VD1.t7 GNDA.t1 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X189 X.t19 Vb2.t7 VD3.t29 VD3.t28 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X190 VD2.t4 VIN+.t2 V_source.t5 GNDA.t8 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X191 V_CMFB_S1.t7 X.t36 GNDA.t117 VDDA.t230 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X192 VOUT-.t4 a_116370_5430# VDDA.t67 VDDA.t66 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=2.4 ps=12.8 w=6 l=0.15
X193 V_CMFB_S3.t7 Y.t35 GNDA.t66 VDDA.t206 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X194 VOUT-.t61 cap_res_X.t96 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X195 VD1.t18 VIN-.t4 V_source.t31 GNDA.t8 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X196 VDDA.t102 Vb3.t13 VD3.t5 VDDA.t101 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X197 V_err_gate.t7 V_err_amp_ref.t4 V_err_mir_p.t2 VDDA.t73 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X198 VOUT+.t69 cap_res_Y.t88 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X199 VDDA.t160 VDDA.t158 Vb2.t0 VDDA.t159 sky130_fd_pr__pfet_01v8 ad=0.252 pd=2.06 as=0.126 ps=1.03 w=0.63 l=0.2
X200 Y.t0 Vb1.t7 VD2.t19 GNDA.t1 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X201 VOUT-.t62 cap_res_X.t95 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X202 V_p_mir.t2 V_tail_gate.t11 GNDA.t4 GNDA.t3 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X203 Y.t1 Vb1.t8 VD2.t18 GNDA.t1 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X204 VOUT+.t70 cap_res_Y.t87 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X205 VOUT+.t71 cap_res_Y.t86 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X206 VOUT-.t63 cap_res_X.t94 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X207 VOUT-.t64 cap_res_X.t93 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X208 VOUT+.t72 cap_res_Y.t85 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X209 VOUT-.t65 cap_res_X.t92 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X210 VOUT+.t73 cap_res_Y.t84 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X211 VD4.t32 Vb2.t8 Y.t16 VD4.t31 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X212 VDDA.t231 X.t37 V_CMFB_S2.t6 GNDA.t0 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X213 VOUT-.t66 cap_res_X.t91 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X214 VOUT-.t67 cap_res_X.t90 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X215 cap_res_X.t0 X.t9 GNDA.t52 sky130_fd_pr__res_high_po_1p41 l=1.41
X216 VDDA.t229 X.t38 VOUT-.t12 VDDA.t228 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X217 VDDA.t205 Y.t36 VOUT+.t10 VDDA.t204 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X218 VOUT-.t68 cap_res_X.t89 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X219 VDDA.t157 VDDA.t155 VD3.t0 VDDA.t156 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X220 VD3.t27 Vb2.t9 X.t18 VD3.t26 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X221 VOUT+.t74 cap_res_Y.t83 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X222 VOUT-.t69 cap_res_X.t88 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X223 VOUT+.t75 cap_res_Y.t82 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X224 VOUT-.t70 cap_res_X.t87 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X225 VOUT-.t71 cap_res_X.t86 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X226 V_CMFB_S4.t6 Y.t37 VDDA.t203 GNDA.t0 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X227 V_err_p.t16 V_err_gate.t20 VDDA.t250 VDDA.t249 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X228 VOUT+.t76 cap_res_Y.t81 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X229 X.t5 Vb1.t9 VD1.t5 GNDA.t1 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X230 X.t2 Vb1.t10 VD1.t2 GNDA.t1 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X231 V_b_2nd_stage.t0 a_109420_966.t0 GNDA.t11 sky130_fd_pr__res_xhigh_po_0p35 l=2.63
X232 VDDA.t154 VDDA.t152 err_amp_out.t6 VDDA.t153 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X233 VD1.t17 VIN-.t5 V_source.t32 GNDA.t8 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X234 V_CMFB_S1.t6 X.t39 GNDA.t118 VDDA.t232 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X235 VDDA.t151 VDDA.t149 GNDA.t126 VDDA.t150 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X236 VDDA.t100 Vb3.t14 VD4.t2 VDDA.t99 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X237 V_CMFB_S3.t6 Y.t38 GNDA.t65 VDDA.t202 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X238 VOUT-.t72 cap_res_X.t85 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X239 VOUT+.t77 cap_res_Y.t80 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X240 VD1.t16 VIN-.t6 V_source.t35 GNDA.t8 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X241 VOUT+.t78 cap_res_Y.t79 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X242 VOUT+.t79 cap_res_Y.t78 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X243 VD2.t7 VIN+.t3 V_source.t19 GNDA.t8 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X244 V_err_gate.t11 VDDA.t146 VDDA.t148 VDDA.t147 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X245 V_err_gate.t6 V_tot.t8 V_err_mir_p.t18 VDDA.t71 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X246 VOUT+.t80 cap_res_Y.t77 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X247 VOUT+.t81 cap_res_Y.t76 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X248 VOUT+.t82 cap_res_Y.t75 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X249 a_109020_3958.t1 V_tot.t0 GNDA.t7 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X250 Y.t23 Vb1.t11 VD2.t17 GNDA.t1 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X251 V_source.t39 V_tail_gate.t12 GNDA.t127 GNDA.t3 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X252 Vb2.t2 Vb2.t1 VDDA.t223 VDDA.t222 sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.03 as=0.126 ps=1.03 w=0.63 l=0.2
X253 VOUT+.t83 cap_res_Y.t74 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X254 VOUT-.t73 cap_res_X.t84 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X255 VDDA.t225 GNDA.t97 GNDA.t98 GNDA.t0 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=1.2 ps=6.8 w=3 l=0.15
X256 VD3.t25 Vb2.t10 X.t17 VD3.t24 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X257 VDDA.t242 V_err_gate.t21 V_err_p.t15 VDDA.t241 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X258 Y.t3 VD4.t14 VD4.t16 VD4.t15 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X259 V_source.t33 VIN-.t7 VD1.t15 GNDA.t8 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X260 VDDA.t234 X.t40 VOUT-.t11 VDDA.t233 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X261 VOUT-.t74 cap_res_X.t83 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X262 VDDA.t78 a_117580_5430# VOUT-.t5 VDDA.t77 sky130_fd_pr__pfet_01v8 ad=2.4 pd=12.8 as=1.2 ps=6.4 w=6 l=0.15
X263 VOUT+.t84 cap_res_Y.t73 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X264 VOUT-.t75 cap_res_X.t82 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X265 VOUT+.t85 cap_res_Y.t72 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X266 VDDA.t201 Y.t39 VOUT+.t9 VDDA.t200 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X267 VOUT-.t6 a_117950_966.t1 GNDA.t39 sky130_fd_pr__res_xhigh_po_0p35 l=2.63
X268 VOUT+.t86 cap_res_Y.t71 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X269 VOUT-.t76 cap_res_X.t81 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X270 VOUT+.t87 cap_res_Y.t70 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X271 GNDA.t28 V_tail_gate.t13 V_source.t13 GNDA.t3 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X272 GNDA.t135 err_amp_mir.t19 err_amp_out.t11 GNDA.t134 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X273 VOUT+.t88 cap_res_Y.t69 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X274 VOUT-.t77 cap_res_X.t80 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X275 V_source.t20 Vb1.t0 Vb1.t1 GNDA.t50 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=2.9
X276 VOUT+.t89 cap_res_Y.t68 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X277 V_CMFB_S2.t5 X.t41 VDDA.t235 GNDA.t0 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X278 VOUT+.t90 cap_res_Y.t67 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X279 VDDA.t98 Vb3.t15 VD4.t7 VDDA.t97 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X280 VOUT+.t91 cap_res_Y.t66 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X281 V_CMFB_S4.t5 Y.t40 VDDA.t197 GNDA.t0 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X282 V_err_mir_p.t10 V_err_gate.t22 VDDA.t246 VDDA.t245 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X283 VD3.t23 Vb2.t11 X.t16 VD3.t22 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X284 VOUT+.t92 cap_res_Y.t65 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X285 VOUT+.t93 cap_res_Y.t64 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X286 VOUT-.t78 cap_res_X.t79 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X287 VOUT+.t94 cap_res_Y.t63 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X288 X.t1 Vb1.t12 VD1.t1 GNDA.t1 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X289 VOUT+.t95 cap_res_Y.t62 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X290 V_err_p.t2 V_tot.t9 err_amp_mir.t13 VDDA.t13 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X291 VOUT+.t96 cap_res_Y.t61 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X292 VD3.t6 Vb3.t16 VDDA.t96 VDDA.t95 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X293 VD2.t11 GNDA.t95 GNDA.t96 GNDA.t8 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X294 V_CMFB_S1.t5 X.t42 GNDA.t35 VDDA.t30 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X295 VOUT+.t97 cap_res_Y.t60 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X296 VD2.t1 VIN+.t4 V_source.t2 GNDA.t8 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X297 VOUT-.t79 cap_res_X.t78 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X298 err_amp_mir.t7 err_amp_mir.t6 GNDA.t44 GNDA.t43 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X299 VOUT+.t98 cap_res_Y.t59 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X300 VOUT-.t80 cap_res_X.t77 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X301 Y.t20 Vb2.t12 VD4.t30 VD4.t29 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X302 Y.t5 Vb1.t13 VD2.t16 GNDA.t1 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X303 VOUT+.t99 cap_res_Y.t58 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X304 V_source.t15 V_tail_gate.t14 GNDA.t37 GNDA.t3 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X305 a_118270_3958.t0 V_CMFB_S2.t0 GNDA.t20 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X306 VOUT-.t81 cap_res_X.t76 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X307 VOUT+.t100 cap_res_Y.t57 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X308 VOUT-.t82 cap_res_X.t75 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X309 VOUT-.t83 cap_res_X.t74 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X310 X.t15 Vb2.t13 VD3.t21 VD3.t20 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X311 VDDA.t32 X.t43 VOUT-.t10 VDDA.t31 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X312 VOUT-.t84 cap_res_X.t73 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X313 VOUT-.t85 cap_res_X.t72 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X314 VDDA.t145 VDDA.t143 V_err_gate.t10 VDDA.t144 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X315 VOUT+.t101 cap_res_Y.t56 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X316 VOUT-.t86 cap_res_X.t71 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X317 GNDA.t40 V_tail_gate.t15 V_source.t16 GNDA.t3 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X318 Y.t17 Vb2.t14 VD4.t28 VD4.t27 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X319 VOUT-.t87 cap_res_X.t70 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X320 VOUT+.t102 cap_res_Y.t55 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X321 VOUT+.t103 cap_res_Y.t54 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X322 VOUT+.t104 cap_res_Y.t53 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X323 VOUT+.t105 cap_res_Y.t52 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X324 GNDA.t94 GNDA.t93 VDDA.t224 GNDA.t0 sky130_fd_pr__nfet_01v8 ad=1.2 pd=6.8 as=0.6 ps=3.4 w=3 l=0.15
X325 V_CMFB_S2.t4 X.t44 VDDA.t33 GNDA.t0 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X326 VOUT+.t106 cap_res_Y.t51 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X327 VOUT-.t88 cap_res_X.t69 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X328 VOUT+.t107 cap_res_Y.t50 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X329 VOUT+.t1 a_109420_966.t1 GNDA.t32 sky130_fd_pr__res_xhigh_po_0p35 l=2.63
X330 V_CMFB_S4.t4 Y.t41 VDDA.t199 GNDA.t0 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X331 V_err_p.t14 V_err_gate.t23 VDDA.t248 VDDA.t247 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X332 V_err_p.t13 V_err_gate.t24 VDDA.t41 VDDA.t40 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X333 VOUT-.t89 cap_res_X.t68 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X334 VOUT-.t90 cap_res_X.t67 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X335 X.t8 Vb1.t14 VD1.t8 GNDA.t1 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X336 a_118390_3958.t0 V_tot.t1 GNDA.t20 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X337 V_CMFB_S1.t4 X.t45 GNDA.t36 VDDA.t34 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X338 VD1.t14 VIN-.t8 V_source.t29 GNDA.t8 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X339 a_109020_3958.t0 V_CMFB_S3.t0 GNDA.t2 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X340 err_amp_out.t2 err_amp_mir.t20 GNDA.t42 GNDA.t41 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X341 VOUT+.t108 cap_res_Y.t49 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X342 VOUT+.t109 cap_res_Y.t48 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X343 Y.t4 GNDA.t91 GNDA.t92 GNDA.t1 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X344 VOUT-.t91 cap_res_X.t66 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X345 VOUT-.t92 cap_res_X.t65 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X346 VOUT-.t93 cap_res_X.t64 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X347 VOUT+.t110 cap_res_Y.t47 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X348 VOUT-.t94 cap_res_X.t63 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X349 X.t14 Vb2.t15 VD3.t19 VD3.t18 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X350 VOUT+.t111 cap_res_Y.t46 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X351 VDDA.t142 VDDA.t140 V_err_p.t10 VDDA.t141 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X352 VOUT-.t95 cap_res_X.t62 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X353 VOUT+.t112 cap_res_Y.t45 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X354 VOUT-.t96 cap_res_X.t61 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X355 VOUT-.t97 cap_res_X.t60 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X356 VD1.t9 Vb1.t15 X.t10 GNDA.t1 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X357 VOUT-.t98 cap_res_X.t59 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X358 GNDA.t63 Y.t42 V_CMFB_S3.t5 VDDA.t198 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X359 GNDA.t84 GNDA.t83 VOUT-.t18 GNDA.t9 sky130_fd_pr__nfet_01v8 ad=2.8 pd=14.8 as=1.4 ps=7.4 w=7 l=0.6
X360 GNDA.t90 GNDA.t89 VD1.t10 GNDA.t8 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X361 VDDA.t59 X.t46 VOUT-.t9 VDDA.t58 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X362 VOUT-.t99 cap_res_X.t58 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X363 VOUT-.t100 cap_res_X.t57 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X364 V_err_mir_p.t1 V_err_amp_ref.t5 V_err_gate.t8 VDDA.t74 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X365 V_err_mir_p.t17 V_tot.t10 V_err_gate.t2 VDDA.t21 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X366 VOUT-.t101 cap_res_X.t56 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X367 VOUT-.t102 cap_res_X.t55 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X368 GNDA.t119 V_tail_gate.t16 V_source.t36 GNDA.t3 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X369 GNDA.t16 V_tail_gate.t17 V_source.t7 GNDA.t3 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X370 VD4.t5 Vb3.t17 VDDA.t94 VDDA.t93 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X371 VOUT-.t103 cap_res_X.t54 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X372 VOUT-.t104 cap_res_X.t53 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X373 VOUT-.t105 cap_res_X.t52 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X374 X.t13 Vb2.t16 VD3.t17 VD3.t16 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X375 VOUT-.t106 cap_res_X.t51 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X376 VOUT-.t107 cap_res_X.t50 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X377 VOUT-.t108 cap_res_X.t49 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X378 VD4.t3 VDDA.t137 VDDA.t139 VDDA.t138 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X379 VOUT-.t109 cap_res_X.t48 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X380 V_CMFB_S2.t3 X.t47 VDDA.t60 GNDA.t0 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X381 V_err_mir_p.t9 V_err_gate.t25 VDDA.t45 VDDA.t44 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X382 VOUT-.t110 cap_res_X.t47 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X383 V_err_p.t6 V_err_amp_ref.t6 err_amp_out.t5 VDDA.t62 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X384 X.t24 GNDA.t87 GNDA.t88 GNDA.t1 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X385 VOUT+.t113 cap_res_Y.t44 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X386 GNDA.t121 V_b_2nd_stage.t7 VOUT+.t17 GNDA.t9 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X387 VOUT+.t8 Y.t43 VDDA.t196 VDDA.t195 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X388 VOUT+.t114 cap_res_Y.t43 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X389 VOUT-.t111 cap_res_X.t46 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X390 VD2.t10 GNDA.t85 GNDA.t86 GNDA.t8 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X391 VD4.t26 Vb2.t17 Y.t15 VD4.t25 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X392 a_118390_3958.t1 V_CMFB_S1.t0 GNDA.t20 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X393 VOUT+.t115 cap_res_Y.t42 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X394 VOUT-.t112 cap_res_X.t45 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X395 err_amp_mir.t5 err_amp_mir.t4 GNDA.t131 GNDA.t130 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X396 V_source.t0 err_amp_out.t12 GNDA.t5 GNDA.t3 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X397 err_amp_mir.t3 err_amp_mir.t2 GNDA.t19 GNDA.t18 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X398 VOUT-.t113 cap_res_X.t44 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X399 VOUT-.t114 cap_res_X.t43 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X400 VOUT+.t116 cap_res_Y.t41 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X401 VOUT+.t117 cap_res_Y.t40 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X402 GNDA.t51 V_b_2nd_stage.t8 VOUT+.t2 GNDA.t9 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X403 VDDA.t237 V_err_gate.t26 V_err_mir_p.t8 VDDA.t236 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X404 VOUT+.t118 cap_res_Y.t39 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X405 VOUT-.t115 cap_res_X.t42 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X406 VOUT-.t116 cap_res_X.t41 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X407 GNDA.t61 Y.t44 V_CMFB_S3.t4 VDDA.t194 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X408 VOUT+.t119 cap_res_Y.t38 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X409 V_tail_gate.t0 VIN+.t5 V_p_mir.t0 GNDA.t8 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X410 V_source.t4 VIN+.t6 VD2.t3 GNDA.t8 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X411 V_err_mir_p.t16 V_tot.t11 V_err_gate.t4 VDDA.t28 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X412 VOUT+.t120 cap_res_Y.t37 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X413 VOUT-.t17 GNDA.t81 GNDA.t82 GNDA.t9 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=2.8 ps=14.8 w=7 l=0.6
X414 VD4.t24 Vb2.t18 Y.t14 VD4.t23 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X415 VOUT-.t117 cap_res_X.t40 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X416 GNDA.t22 V_tail_gate.t18 V_source.t9 GNDA.t3 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X417 GNDA.t80 GNDA.t79 Y.t12 GNDA.t1 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X418 GNDA.t17 V_tail_gate.t19 V_source.t8 GNDA.t3 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X419 VOUT-.t118 cap_res_X.t39 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X420 V_err_mir_p.t7 V_err_gate.t27 VDDA.t3 VDDA.t2 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X421 V_CMFB_S2.t2 X.t48 VDDA.t35 GNDA.t0 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X422 VOUT-.t119 cap_res_X.t38 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X423 VOUT+.t121 cap_res_Y.t36 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X424 VOUT+.t122 cap_res_Y.t35 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X425 VOUT-.t120 cap_res_X.t37 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X426 VOUT+.t123 cap_res_Y.t34 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X427 VOUT-.t0 V_b_2nd_stage.t9 GNDA.t26 GNDA.t9 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X428 a_118270_3958.t1 V_tot.t3 GNDA.t20 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X429 VOUT+.t7 Y.t45 VDDA.t193 VDDA.t192 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X430 V_err_p.t1 V_tot.t12 err_amp_mir.t12 VDDA.t6 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X431 VOUT+.t124 cap_res_Y.t33 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X432 a_108900_3958.t1 V_CMFB_S4.t0 GNDA.t47 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X433 V_CMFB_S1.t3 X.t49 GNDA.t21 VDDA.t24 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X434 VOUT+.t125 cap_res_Y.t32 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X435 VOUT+.t126 cap_res_Y.t31 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X436 V_source.t24 V_tail_gate.t20 GNDA.t57 GNDA.t3 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X437 VD3.t15 Vb2.t19 X.t12 VD3.t14 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X438 err_amp_out.t1 err_amp_mir.t21 GNDA.t13 GNDA.t12 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X439 VOUT+.t127 cap_res_Y.t30 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X440 VDDA.t187 Y.t46 V_CMFB_S4.t3 GNDA.t0 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X441 VOUT+.t128 cap_res_Y.t29 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X442 VDDA.t5 V_err_gate.t28 V_err_p.t12 VDDA.t4 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X443 VOUT+.t129 cap_res_Y.t28 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X444 VDDA.t92 Vb3.t18 VD4.t8 VDDA.t91 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X445 VD4.t13 VD4.t11 Y.t9 VD4.t12 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X446 err_amp_out.t3 V_err_amp_ref.t7 V_err_p.t4 VDDA.t57 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X447 GNDA.t78 GNDA.t77 X.t23 GNDA.t1 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X448 VOUT+.t130 cap_res_Y.t27 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X449 VOUT+.t131 cap_res_Y.t26 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X450 V_source.t18 VIN+.t7 VD2.t6 GNDA.t8 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X451 VDDA.t53 X.t50 VOUT-.t8 VDDA.t52 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X452 GNDA.t60 Y.t47 V_CMFB_S3.t3 VDDA.t191 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X453 VOUT-.t121 cap_res_X.t36 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X454 V_tail_gate.t2 GNDA.t75 GNDA.t76 GNDA.t8 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X455 VOUT+.t132 cap_res_Y.t25 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X456 cap_res_Y.t0 Y.t8 GNDA.t46 sky130_fd_pr__res_high_po_1p41 l=1.41
X457 GNDA.t74 GNDA.t73 VD1.t11 GNDA.t8 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X458 VD3.t1 VDDA.t134 VDDA.t136 VDDA.t135 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X459 V_err_mir_p.t0 V_err_amp_ref.t8 V_err_gate.t5 VDDA.t48 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X460 VD3.t34 VD3.t32 X.t21 VD3.t33 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X461 GNDA.t49 V_tail_gate.t21 V_p_mir.t1 GNDA.t3 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X462 VD2.t15 Vb1.t16 Y.t7 GNDA.t1 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X463 VOUT-.t122 cap_res_X.t35 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X464 Vb2_Vb3.t8 VDDA.t131 VDDA.t133 VDDA.t132 sky130_fd_pr__pfet_01v8 ad=0.71 pd=3.95 as=1.42 ps=7.9 w=3.55 l=0.2
X465 VOUT+.t133 cap_res_Y.t24 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X466 VOUT+.t134 cap_res_Y.t23 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X467 V_err_p.t9 VDDA.t128 VDDA.t130 VDDA.t129 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X468 VOUT+.t135 cap_res_Y.t22 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X469 VOUT+.t136 cap_res_Y.t21 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X470 VOUT-.t123 cap_res_X.t34 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X471 VOUT+.t137 cap_res_Y.t20 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X472 VOUT-.t124 cap_res_X.t33 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X473 VOUT-.t125 cap_res_X.t32 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X474 VOUT-.t126 cap_res_X.t31 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X475 VOUT-.t127 cap_res_X.t30 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X476 VOUT+.t6 Y.t48 VDDA.t181 VDDA.t180 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X477 Y.t21 Vb2.t20 VD4.t22 VD4.t21 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X478 VOUT+.t138 cap_res_Y.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X479 VOUT+.t139 cap_res_Y.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X480 VOUT+.t140 cap_res_Y.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X481 VOUT-.t128 cap_res_X.t29 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X482 VOUT+.t141 cap_res_Y.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X483 VOUT+.t142 cap_res_Y.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X484 VOUT+.t143 cap_res_Y.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X485 VDDA.t188 Y.t49 V_CMFB_S4.t2 GNDA.t0 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X486 VOUT-.t129 cap_res_X.t28 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X487 VOUT-.t130 cap_res_X.t27 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X488 VOUT-.t131 cap_res_X.t26 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X489 VOUT+.t144 cap_res_Y.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X490 VOUT+.t145 cap_res_Y.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X491 VD1.t3 Vb1.t17 X.t3 GNDA.t1 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X492 GNDA.t6 X.t51 V_CMFB_S1.t2 VDDA.t7 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X493 V_source.t28 VIN-.t9 VD1.t13 GNDA.t8 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X494 Y.t18 Vb2.t21 VD4.t20 VD4.t19 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X495 GNDA.t62 Y.t50 V_CMFB_S3.t2 VDDA.t190 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X496 GNDA.t64 Y.t51 V_CMFB_S3.t1 VDDA.t189 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X497 VOUT-.t132 cap_res_X.t25 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X498 V_source.t30 VIN-.t10 VD1.t12 GNDA.t8 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X499 V_source.t1 VIN+.t8 VD2.t0 GNDA.t8 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X500 V_err_mir_p.t15 V_tot.t13 V_err_gate.t1 VDDA.t20 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X501 VOUT+.t146 cap_res_Y.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X502 VOUT+.t147 cap_res_Y.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X503 VOUT-.t133 cap_res_X.t24 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X504 GNDA.t72 GNDA.t70 GNDA.t71 GNDA.t3 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=0 ps=0 w=2.5 l=0.15
X505 VD2.t14 Vb1.t18 Y.t2 GNDA.t1 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X506 VD2.t13 Vb1.t19 Y.t6 GNDA.t1 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X507 VOUT-.t134 cap_res_X.t23 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X508 VOUT-.t135 cap_res_X.t22 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X509 VOUT-.t136 cap_res_X.t21 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X510 VOUT+.t148 cap_res_Y.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X511 Y.t22 Vb2.t22 VD4.t18 VD4.t17 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X512 VOUT-.t137 cap_res_X.t20 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X513 V_CMFB_S2.t1 X.t52 VDDA.t244 GNDA.t0 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X514 VOUT-.t138 cap_res_X.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X515 VD3.t10 Vb3.t19 VDDA.t90 VDDA.t89 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X516 V_err_mir_p.t6 V_err_gate.t29 VDDA.t16 VDDA.t15 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X517 VOUT-.t139 cap_res_X.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X518 VOUT-.t7 X.t53 VDDA.t37 VDDA.t36 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X519 VOUT+.t5 Y.t52 VDDA.t186 VDDA.t185 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X520 VOUT+.t4 Y.t53 VDDA.t184 VDDA.t183 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X521 VOUT+.t149 cap_res_Y.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X522 VOUT-.t140 cap_res_X.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X523 X.t11 Vb2.t23 VD3.t13 VD3.t12 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X524 VOUT-.t141 cap_res_X.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X525 VOUT-.t142 cap_res_X.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X526 V_source.t40 V_tail_gate.t22 GNDA.t133 GNDA.t3 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X527 a_108900_3958.t0 V_tot.t2 GNDA.t31 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X528 VOUT-.t143 cap_res_X.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X529 VOUT+.t150 cap_res_Y.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X530 VOUT-.t144 cap_res_X.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X531 VOUT+.t151 cap_res_Y.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X532 VD4.t1 Vb3.t20 VDDA.t88 VDDA.t87 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X533 VOUT-.t145 cap_res_X.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X534 VDDA.t182 Y.t54 V_CMFB_S4.t1 GNDA.t0 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X535 VDDA.t56 V_err_gate.t30 V_err_mir_p.t5 VDDA.t55 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X536 VD1.t6 Vb1.t20 X.t6 GNDA.t1 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X537 err_amp_out.t9 V_err_amp_ref.t9 V_err_p.t21 VDDA.t243 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X538 VOUT-.t146 cap_res_X.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X539 VDDA.t86 Vb3.t21 VD3.t11 VDDA.t85 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X540 VOUT+.t152 cap_res_Y.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X541 VOUT-.t147 cap_res_X.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X542 V_b_2nd_stage.t1 a_117950_966.t0 GNDA.t39 sky130_fd_pr__res_xhigh_po_0p35 l=2.63
X543 V_source.t12 VIN+.t9 VD2.t5 GNDA.t8 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X544 GNDA.t59 X.t54 V_CMFB_S1.t1 VDDA.t79 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X545 V_source.t3 VIN+.t10 VD2.t2 GNDA.t8 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X546 VOUT-.t148 cap_res_X.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X547 VOUT-.t149 cap_res_X.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X548 VOUT+.t153 cap_res_Y.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X549 GNDA.t25 err_amp_mir.t0 err_amp_mir.t1 GNDA.t24 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X550 VOUT-.t150 cap_res_X.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X551 VDDA.t84 Vb3.t22 Vb2_Vb3.t7 VDDA.t83 sky130_fd_pr__pfet_01v8 ad=0.71 pd=3.95 as=0.71 ps=3.95 w=3.55 l=0.2
X552 VOUT-.t151 cap_res_X.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X553 VD2.t12 Vb1.t21 Y.t11 GNDA.t1 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X554 VOUT-.t152 cap_res_X.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X555 GNDA.t123 V_tail_gate.t23 V_source.t38 GNDA.t3 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X556 VOUT-.t153 cap_res_X.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X557 VOUT+.t154 cap_res_Y.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X558 GNDA.t56 VDDA.t125 VDDA.t127 VDDA.t126 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X559 V_err_p.t11 V_err_gate.t31 VDDA.t50 VDDA.t49 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X560 VOUT-.t154 cap_res_X.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X561 VOUT-.t155 cap_res_X.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X562 VOUT+.t155 cap_res_Y.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X563 VOUT+.t156 cap_res_Y.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X564 VOUT-.t156 cap_res_X.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
R0 Vb2.n2 Vb2.t6 677.534
R1 Vb2.n1 Vb2.n0 620.841
R2 Vb2.n16 Vb2.t8 611.739
R3 Vb2.n12 Vb2.t21 611.739
R4 Vb2.n7 Vb2.t9 611.739
R5 Vb2.n3 Vb2.t16 611.739
R6 Vb2.n16 Vb2.t12 421.75
R7 Vb2.n17 Vb2.t17 421.75
R8 Vb2.n18 Vb2.t20 421.75
R9 Vb2.n19 Vb2.t3 421.75
R10 Vb2.n12 Vb2.t18 421.75
R11 Vb2.n13 Vb2.t14 421.75
R12 Vb2.n14 Vb2.t4 421.75
R13 Vb2.n15 Vb2.t22 421.75
R14 Vb2.n7 Vb2.t13 421.75
R15 Vb2.n8 Vb2.t10 421.75
R16 Vb2.n9 Vb2.t15 421.75
R17 Vb2.n10 Vb2.t19 421.75
R18 Vb2.n3 Vb2.t11 421.75
R19 Vb2.n4 Vb2.t7 421.75
R20 Vb2.n5 Vb2.t5 421.75
R21 Vb2.n6 Vb2.t23 421.75
R22 Vb2.n1 Vb2.t1 288.166
R23 Vb2.n21 Vb2.n11 169.405
R24 Vb2.n21 Vb2.n20 168.843
R25 Vb2.n17 Vb2.n16 167.094
R26 Vb2.n18 Vb2.n17 167.094
R27 Vb2.n19 Vb2.n18 167.094
R28 Vb2.n13 Vb2.n12 167.094
R29 Vb2.n14 Vb2.n13 167.094
R30 Vb2.n15 Vb2.n14 167.094
R31 Vb2.n8 Vb2.n7 167.094
R32 Vb2.n9 Vb2.n8 167.094
R33 Vb2.n10 Vb2.n9 167.094
R34 Vb2.n4 Vb2.n3 167.094
R35 Vb2.n5 Vb2.n4 167.094
R36 Vb2.n6 Vb2.n5 167.094
R37 Vb2.n0 Vb2.t0 62.5402
R38 Vb2.n0 Vb2.t2 62.5402
R39 Vb2.n20 Vb2.n19 47.1294
R40 Vb2.n20 Vb2.n15 47.1294
R41 Vb2.n11 Vb2.n10 47.1294
R42 Vb2.n11 Vb2.n6 47.1294
R43 Vb2.n2 Vb2.n1 17.8942
R44 Vb2.n22 Vb2.n2 8.59425
R45 Vb2.n22 Vb2.n21 4.5005
R46 Vb2 Vb2.n22 0.063
R47 Y.n49 Y.t39 1172.87
R48 Y.n43 Y.t53 1172.87
R49 Y.n50 Y.t36 996.134
R50 Y.n49 Y.t52 996.134
R51 Y.n43 Y.t28 996.134
R52 Y.n44 Y.t43 996.134
R53 Y.n45 Y.t30 996.134
R54 Y.n46 Y.t45 996.134
R55 Y.n47 Y.t33 996.134
R56 Y.n48 Y.t48 996.134
R57 Y.n32 Y.t41 690.867
R58 Y.n31 Y.t26 690.867
R59 Y.n23 Y.t38 530.201
R60 Y.n22 Y.t51 530.201
R61 Y.n32 Y.t25 514.134
R62 Y.n33 Y.t40 514.134
R63 Y.n34 Y.t54 514.134
R64 Y.n35 Y.t37 514.134
R65 Y.n36 Y.t49 514.134
R66 Y.n37 Y.t34 514.134
R67 Y.n38 Y.t46 514.134
R68 Y.n31 Y.t31 514.134
R69 Y.n29 Y.t42 353.467
R70 Y.n28 Y.t29 353.467
R71 Y.n27 Y.t44 353.467
R72 Y.n26 Y.t32 353.467
R73 Y.n25 Y.t47 353.467
R74 Y.n24 Y.t35 353.467
R75 Y.n23 Y.t50 353.467
R76 Y.n22 Y.t27 353.467
R77 Y.n50 Y.n49 176.733
R78 Y.n44 Y.n43 176.733
R79 Y.n45 Y.n44 176.733
R80 Y.n46 Y.n45 176.733
R81 Y.n47 Y.n46 176.733
R82 Y.n48 Y.n47 176.733
R83 Y.n29 Y.n28 176.733
R84 Y.n28 Y.n27 176.733
R85 Y.n27 Y.n26 176.733
R86 Y.n26 Y.n25 176.733
R87 Y.n25 Y.n24 176.733
R88 Y.n24 Y.n23 176.733
R89 Y.n38 Y.n37 176.733
R90 Y.n37 Y.n36 176.733
R91 Y.n36 Y.n35 176.733
R92 Y.n35 Y.n34 176.733
R93 Y.n34 Y.n33 176.733
R94 Y.n33 Y.n32 176.733
R95 Y.n52 Y.n51 166.436
R96 Y.n40 Y.n30 161.843
R97 Y.n40 Y.n39 161.718
R98 Y.n13 Y.n11 160.427
R99 Y.n19 Y.n18 159.802
R100 Y.n17 Y.n16 159.802
R101 Y.n15 Y.n14 159.802
R102 Y.n13 Y.n12 159.802
R103 Y.n21 Y.n20 155.302
R104 Y.n9 Y.n8 114.689
R105 Y.n3 Y.n1 114.689
R106 Y.n7 Y.n6 114.126
R107 Y.n5 Y.n4 114.126
R108 Y.n3 Y.n2 114.126
R109 Y.n10 Y.n0 109.626
R110 Y.n51 Y.n50 51.9494
R111 Y.n51 Y.n48 51.9494
R112 Y.n30 Y.n29 51.9494
R113 Y.n30 Y.n22 51.9494
R114 Y.n39 Y.n38 51.9494
R115 Y.n39 Y.n31 51.9494
R116 Y.t8 Y.n52 49.4594
R117 Y.n41 Y.n21 17.438
R118 Y.n8 Y.t24 16.0005
R119 Y.n8 Y.t4 16.0005
R120 Y.n6 Y.t2 16.0005
R121 Y.n6 Y.t23 16.0005
R122 Y.n4 Y.t6 16.0005
R123 Y.n4 Y.t0 16.0005
R124 Y.n2 Y.t7 16.0005
R125 Y.n2 Y.t1 16.0005
R126 Y.n1 Y.t12 16.0005
R127 Y.n1 Y.t10 16.0005
R128 Y.n0 Y.t11 16.0005
R129 Y.n0 Y.t5 16.0005
R130 Y.n41 Y.n40 13.938
R131 Y.n20 Y.t16 11.2576
R132 Y.n20 Y.t3 11.2576
R133 Y.n18 Y.t15 11.2576
R134 Y.n18 Y.t20 11.2576
R135 Y.n16 Y.t13 11.2576
R136 Y.n16 Y.t21 11.2576
R137 Y.n14 Y.t19 11.2576
R138 Y.n14 Y.t22 11.2576
R139 Y.n12 Y.t14 11.2576
R140 Y.n12 Y.t17 11.2576
R141 Y.n11 Y.t9 11.2576
R142 Y.n11 Y.t18 11.2576
R143 Y.n42 Y.n10 9.313
R144 Y.n21 Y.n19 5.1255
R145 Y.n10 Y.n9 4.5005
R146 Y.n42 Y.n41 4.5005
R147 Y.n52 Y.n42 3.3755
R148 Y.n15 Y.n13 0.6255
R149 Y.n17 Y.n15 0.6255
R150 Y.n19 Y.n17 0.6255
R151 Y.n5 Y.n3 0.563
R152 Y.n7 Y.n5 0.563
R153 Y.n9 Y.n7 0.563
R154 VD4.n38 VD4.t14 680.832
R155 VD4.n28 VD4.t11 680.832
R156 VD4.n50 VD4.n2 585
R157 VD4.n31 VD4.n30 585
R158 VD4.n37 VD4.n2 290.233
R159 VD4.n44 VD4.n2 290.233
R160 VD4.n39 VD4.n2 290.233
R161 VD4.n30 VD4.n18 290.233
R162 VD4.n30 VD4.n23 290.233
R163 VD4.n30 VD4.n29 290.233
R164 VD4.n50 VD4.n49 238.367
R165 VD4.n38 VD4.n35 238.367
R166 VD4.n28 VD4.n7 238.367
R167 VD4.n4 VD4.n3 185
R168 VD4.n47 VD4.n46 185
R169 VD4.n48 VD4.n47 185
R170 VD4.n45 VD4.n36 185
R171 VD4.n43 VD4.n42 185
R172 VD4.n41 VD4.n40 185
R173 VD4.n32 VD4.n31 185
R174 VD4.n33 VD4.n32 185
R175 VD4.n17 VD4.n8 185
R176 VD4.n20 VD4.n19 185
R177 VD4.n22 VD4.n21 185
R178 VD4.n25 VD4.n24 185
R179 VD4.n27 VD4.n26 185
R180 VD4.t12 VD4.n33 170.513
R181 VD4.n48 VD4.t15 170.513
R182 VD4.n54 VD4.n52 160.427
R183 VD4.n12 VD4.n11 159.804
R184 VD4.n14 VD4.n13 159.803
R185 VD4.n16 VD4.n15 159.803
R186 VD4.n1 VD4.n0 159.803
R187 VD4.n10 VD4.n9 159.803
R188 VD4.n62 VD4.n61 159.802
R189 VD4.n60 VD4.n59 159.802
R190 VD4.n58 VD4.n57 159.802
R191 VD4.n56 VD4.n55 159.802
R192 VD4.n54 VD4.n53 159.802
R193 VD4.n47 VD4.n4 150
R194 VD4.n47 VD4.n36 150
R195 VD4.n42 VD4.n41 150
R196 VD4.n32 VD4.n8 150
R197 VD4.n21 VD4.n20 150
R198 VD4.n26 VD4.n25 150
R199 VD4.t19 VD4.t12 146.155
R200 VD4.t23 VD4.t19 146.155
R201 VD4.t27 VD4.t23 146.155
R202 VD4.t33 VD4.t27 146.155
R203 VD4.t17 VD4.t33 146.155
R204 VD4.t35 VD4.t17 146.155
R205 VD4.t21 VD4.t35 146.155
R206 VD4.t25 VD4.t21 146.155
R207 VD4.t29 VD4.t25 146.155
R208 VD4.t31 VD4.t29 146.155
R209 VD4.t15 VD4.t31 146.155
R210 VD4.n49 VD4.n48 65.8183
R211 VD4.n48 VD4.n34 65.8183
R212 VD4.n48 VD4.n35 65.8183
R213 VD4.n33 VD4.n5 65.8183
R214 VD4.n33 VD4.n6 65.8183
R215 VD4.n33 VD4.n7 65.8183
R216 VD4.n36 VD4.n34 53.3664
R217 VD4.n41 VD4.n35 53.3664
R218 VD4.n49 VD4.n4 53.3664
R219 VD4.n42 VD4.n34 53.3664
R220 VD4.n8 VD4.n5 53.3664
R221 VD4.n21 VD4.n6 53.3664
R222 VD4.n26 VD4.n7 53.3664
R223 VD4.n20 VD4.n5 53.3664
R224 VD4.n25 VD4.n6 53.3664
R225 VD4.n31 VD4.n16 37.2826
R226 VD4.n51 VD4.n50 36.6576
R227 VD4.n13 VD4.t28 11.2576
R228 VD4.n13 VD4.t34 11.2576
R229 VD4.n15 VD4.t20 11.2576
R230 VD4.n15 VD4.t24 11.2576
R231 VD4.n30 VD4.t13 11.2576
R232 VD4.n2 VD4.t16 11.2576
R233 VD4.n61 VD4.t37 11.2576
R234 VD4.n61 VD4.t0 11.2576
R235 VD4.n59 VD4.t10 11.2576
R236 VD4.n59 VD4.t5 11.2576
R237 VD4.n57 VD4.t7 11.2576
R238 VD4.n57 VD4.t6 11.2576
R239 VD4.n55 VD4.t2 11.2576
R240 VD4.n55 VD4.t9 11.2576
R241 VD4.n53 VD4.t4 11.2576
R242 VD4.n53 VD4.t1 11.2576
R243 VD4.n52 VD4.t8 11.2576
R244 VD4.n52 VD4.t3 11.2576
R245 VD4.n0 VD4.t30 11.2576
R246 VD4.n0 VD4.t32 11.2576
R247 VD4.n9 VD4.t22 11.2576
R248 VD4.n9 VD4.t26 11.2576
R249 VD4.n11 VD4.t18 11.2576
R250 VD4.n11 VD4.t36 11.2576
R251 VD4.n50 VD4.n3 9.14336
R252 VD4.n46 VD4.n45 9.14336
R253 VD4.n43 VD4.n40 9.14336
R254 VD4.n31 VD4.n17 9.14336
R255 VD4.n22 VD4.n19 9.14336
R256 VD4.n27 VD4.n24 9.14336
R257 VD4 VD4.n62 8.5005
R258 VD4 VD4.n51 5.188
R259 VD4.n37 VD4.n3 4.53698
R260 VD4.n45 VD4.n44 4.53698
R261 VD4.n40 VD4.n39 4.53698
R262 VD4.n46 VD4.n37 4.53698
R263 VD4.n44 VD4.n43 4.53698
R264 VD4.n39 VD4.n38 4.53698
R265 VD4.n18 VD4.n17 4.53698
R266 VD4.n23 VD4.n22 4.53698
R267 VD4.n29 VD4.n27 4.53698
R268 VD4.n19 VD4.n18 4.53698
R269 VD4.n24 VD4.n23 4.53698
R270 VD4.n29 VD4.n28 4.53698
R271 VD4.n56 VD4.n54 0.6255
R272 VD4.n58 VD4.n56 0.6255
R273 VD4.n60 VD4.n58 0.6255
R274 VD4.n62 VD4.n60 0.6255
R275 VD4.n12 VD4.n10 0.6255
R276 VD4.n10 VD4.n1 0.6255
R277 VD4.n51 VD4.n1 0.6255
R278 VD4.n16 VD4.n14 0.6255
R279 VD4.n14 VD4.n12 0.6255
R280 VIN-.n4 VIN-.t3 485.021
R281 VIN-.n1 VIN-.t4 484.159
R282 VIN-.n5 VIN-.t2 483.358
R283 VIN-.n8 VIN-.t5 431.536
R284 VIN-.n2 VIN-.t8 431.536
R285 VIN-.n6 VIN-.t0 431.257
R286 VIN-.n0 VIN-.t6 431.257
R287 VIN-.n6 VIN-.t7 289.908
R288 VIN-.n0 VIN-.t10 289.908
R289 VIN-.n8 VIN-.t9 279.183
R290 VIN-.n2 VIN-.t1 279.183
R291 VIN-.n7 VIN-.n6 233.374
R292 VIN-.n1 VIN-.n0 233.374
R293 VIN-.n9 VIN-.n8 188.989
R294 VIN-.n3 VIN-.n2 188.989
R295 VIN-.n4 VIN-.n3 2.463
R296 VIN- VIN-.n9 1.78175
R297 VIN-.n5 VIN-.n4 1.563
R298 VIN-.n3 VIN-.n1 1.2755
R299 VIN-.n9 VIN-.n7 1.2755
R300 VIN-.n7 VIN-.n5 0.8005
R301 V_source.n7 V_source.t20 205.97
R302 V_source.n25 V_source.n23 118.168
R303 V_source.n19 V_source.n17 117.831
R304 V_source.n31 V_source.n30 117.269
R305 V_source.n29 V_source.n28 117.269
R306 V_source.n27 V_source.n26 117.269
R307 V_source.n25 V_source.n24 117.269
R308 V_source.n0 V_source.n22 117.269
R309 V_source.n21 V_source.n20 117.269
R310 V_source.n19 V_source.n18 117.269
R311 V_source.n32 V_source.n16 113.136
R312 V_source.n37 V_source.n36 99.7419
R313 V_source.n3 V_source.n1 99.647
R314 V_source.n36 V_source.n35 99.0845
R315 V_source.n14 V_source.n13 99.0845
R316 V_source.n12 V_source.n11 99.0845
R317 V_source.n10 V_source.n9 99.0845
R318 V_source.n5 V_source.n4 99.0845
R319 V_source.n3 V_source.n2 99.0845
R320 V_source.n33 V_source.n15 94.5845
R321 V_source.n7 V_source.n6 94.5845
R322 V_source.n30 V_source.t26 16.0005
R323 V_source.n30 V_source.t4 16.0005
R324 V_source.n28 V_source.t22 16.0005
R325 V_source.n28 V_source.t33 16.0005
R326 V_source.n26 V_source.t27 16.0005
R327 V_source.n26 V_source.t18 16.0005
R328 V_source.n24 V_source.t5 16.0005
R329 V_source.n24 V_source.t28 16.0005
R330 V_source.n23 V_source.t32 16.0005
R331 V_source.n23 V_source.t12 16.0005
R332 V_source.n22 V_source.t2 16.0005
R333 V_source.n22 V_source.t34 16.0005
R334 V_source.n20 V_source.t35 16.0005
R335 V_source.n20 V_source.t3 16.0005
R336 V_source.n18 V_source.t19 16.0005
R337 V_source.n18 V_source.t30 16.0005
R338 V_source.n17 V_source.t31 16.0005
R339 V_source.n17 V_source.t1 16.0005
R340 V_source.n16 V_source.t29 16.0005
R341 V_source.n16 V_source.t23 16.0005
R342 V_source.n35 V_source.t21 9.6005
R343 V_source.n35 V_source.t24 9.6005
R344 V_source.n15 V_source.t17 9.6005
R345 V_source.n15 V_source.t11 9.6005
R346 V_source.n13 V_source.t7 9.6005
R347 V_source.n13 V_source.t25 9.6005
R348 V_source.n11 V_source.t8 9.6005
R349 V_source.n11 V_source.t40 9.6005
R350 V_source.n9 V_source.t13 9.6005
R351 V_source.n9 V_source.t14 9.6005
R352 V_source.n6 V_source.t16 9.6005
R353 V_source.n6 V_source.t37 9.6005
R354 V_source.n4 V_source.t36 9.6005
R355 V_source.n4 V_source.t39 9.6005
R356 V_source.n2 V_source.t38 9.6005
R357 V_source.n2 V_source.t15 9.6005
R358 V_source.n1 V_source.t9 9.6005
R359 V_source.n1 V_source.t10 9.6005
R360 V_source.n37 V_source.t6 9.6005
R361 V_source.t0 V_source.n37 9.6005
R362 V_source.n32 V_source.n0 4.5005
R363 V_source.n8 V_source.n7 4.5005
R364 V_source.n34 V_source.n33 4.5005
R365 V_source.n0 V_source.n31 3.65675
R366 V_source.n33 V_source.n32 1.34425
R367 V_source.n0 V_source.n21 1.09425
R368 V_source.n27 V_source.n25 0.563
R369 V_source.n29 V_source.n27 0.563
R370 V_source.n31 V_source.n29 0.563
R371 V_source.n21 V_source.n19 0.563
R372 V_source.n5 V_source.n3 0.563
R373 V_source.n8 V_source.n5 0.563
R374 V_source.n10 V_source.n8 0.563
R375 V_source.n12 V_source.n10 0.563
R376 V_source.n14 V_source.n12 0.563
R377 V_source.n34 V_source.n14 0.563
R378 V_source.n36 V_source.n34 0.563
R379 VD1.n10 VD1.n9 114.719
R380 VD1.n6 VD1.n4 114.719
R381 VD1.n8 VD1.n7 114.156
R382 VD1.n6 VD1.n5 114.156
R383 VD1.n2 VD1.n0 113.081
R384 VD1.n16 VD1.n15 111.769
R385 VD1.n18 VD1.n17 111.769
R386 VD1 VD1.n19 111.769
R387 VD1.n2 VD1.n1 111.769
R388 VD1.n11 VD1.n3 109.656
R389 VD1.n13 VD1.n12 107.267
R390 VD1.n15 VD1.t10 16.0005
R391 VD1.n15 VD1.t19 16.0005
R392 VD1.n17 VD1.t15 16.0005
R393 VD1.n17 VD1.t21 16.0005
R394 VD1.n19 VD1.t13 16.0005
R395 VD1.n19 VD1.t17 16.0005
R396 VD1.n1 VD1.t12 16.0005
R397 VD1.n1 VD1.t16 16.0005
R398 VD1.n0 VD1.t11 16.0005
R399 VD1.n0 VD1.t18 16.0005
R400 VD1.n9 VD1.t8 16.0005
R401 VD1.n9 VD1.t4 16.0005
R402 VD1.n7 VD1.t5 16.0005
R403 VD1.n7 VD1.t6 16.0005
R404 VD1.n5 VD1.t2 16.0005
R405 VD1.n5 VD1.t9 16.0005
R406 VD1.n4 VD1.t7 16.0005
R407 VD1.n4 VD1.t3 16.0005
R408 VD1.n3 VD1.t1 16.0005
R409 VD1.n3 VD1.t0 16.0005
R410 VD1.n12 VD1.t20 16.0005
R411 VD1.n12 VD1.t14 16.0005
R412 VD1.n11 VD1.n10 4.5005
R413 VD1.n14 VD1.n13 4.5005
R414 VD1.n16 VD1.n14 3.563
R415 VD1.n18 VD1.n16 1.313
R416 VD1.n14 VD1.n2 1.2505
R417 VD1 VD1.n18 1.2505
R418 VD1.n8 VD1.n6 0.563
R419 VD1.n10 VD1.n8 0.563
R420 VD1.n13 VD1.n11 0.21925
R421 GNDA.n243 GNDA.n237 12249
R422 GNDA.n252 GNDA.n251 12249
R423 GNDA.n245 GNDA.n221 12151.5
R424 GNDA.n248 GNDA.n247 11440
R425 GNDA.n245 GNDA.n219 11275
R426 GNDA.n218 GNDA.n217 10236.5
R427 GNDA.n247 GNDA.n245 9418.75
R428 GNDA.n247 GNDA.n246 9418.75
R429 GNDA.n244 GNDA.n222 8257.53
R430 GNDA.n222 GNDA.n215 8257.53
R431 GNDA.n249 GNDA.n216 7745.63
R432 GNDA.n221 GNDA.n218 6534.33
R433 GNDA.n248 GNDA.n218 5447.23
R434 GNDA.n250 GNDA.n249 5404.35
R435 GNDA.n246 GNDA.n216 5183.79
R436 GNDA.n245 GNDA.n244 3806
R437 GNDA.n246 GNDA.n215 3806
R438 GNDA.n249 GNDA.n248 3714.29
R439 GNDA.n221 GNDA.n220 3488.99
R440 GNDA.n244 GNDA.n243 2971.52
R441 GNDA.n252 GNDA.n215 2971.52
R442 GNDA.n220 GNDA.n219 2695.83
R443 GNDA.n236 GNDA.n222 2640
R444 GNDA.n220 GNDA.n217 2510.03
R445 GNDA.n251 GNDA.n216 1388.09
R446 GNDA.n243 GNDA.n242 1309.92
R447 GNDA.n253 GNDA.n252 1309.92
R448 GNDA.t1 GNDA.n208 1272.11
R449 GNDA.t1 GNDA.n207 1272.11
R450 GNDA.n250 GNDA.n217 924.639
R451 GNDA.t52 GNDA.n219 845.833
R452 GNDA.n251 GNDA.n250 813.446
R453 GNDA.n237 GNDA.t52 754.168
R454 GNDA.n192 GNDA.t93 734.418
R455 GNDA.n269 GNDA.t97 734.418
R456 GNDA.n296 GNDA.t99 734.418
R457 GNDA.n294 GNDA.t108 734.418
R458 GNDA.n99 GNDA.t70 682.201
R459 GNDA.n237 GNDA.n236 666.668
R460 GNDA.n136 GNDA.t110 666.134
R461 GNDA.n279 GNDA.n278 590.789
R462 GNDA.n282 GNDA.n175 590.789
R463 GNDA.n281 GNDA.n280 590.789
R464 GNDA.n285 GNDA.n284 590.789
R465 GNDA.n76 GNDA.n75 585
R466 GNDA.n384 GNDA.n76 585
R467 GNDA.n392 GNDA.n391 585
R468 GNDA.n391 GNDA.n390 585
R469 GNDA.n74 GNDA.n73 585
R470 GNDA.n377 GNDA.n73 585
R471 GNDA.n397 GNDA.n396 585
R472 GNDA.n398 GNDA.n397 585
R473 GNDA.n60 GNDA.n59 585
R474 GNDA.n371 GNDA.n60 585
R475 GNDA.n409 GNDA.n408 585
R476 GNDA.n408 GNDA.n407 585
R477 GNDA.n57 GNDA.n56 585
R478 GNDA.n64 GNDA.n56 585
R479 GNDA.n414 GNDA.n413 585
R480 GNDA.n415 GNDA.n414 585
R481 GNDA.n45 GNDA.n44 585
R482 GNDA.n46 GNDA.n45 585
R483 GNDA.n430 GNDA.n429 585
R484 GNDA.n429 GNDA.n428 585
R485 GNDA.n42 GNDA.n41 585
R486 GNDA.n41 GNDA.n38 585
R487 GNDA.n436 GNDA.n435 585
R488 GNDA.n437 GNDA.n436 585
R489 GNDA.n434 GNDA.n31 585
R490 GNDA.n31 GNDA.n28 585
R491 GNDA.n449 GNDA.n448 585
R492 GNDA.n450 GNDA.n449 585
R493 GNDA.n128 GNDA.n127 585
R494 GNDA.n127 GNDA.n77 585
R495 GNDA.n126 GNDA.n125 585
R496 GNDA.n126 GNDA.n80 585
R497 GNDA.n131 GNDA.n124 585
R498 GNDA.n124 GNDA.t3 585
R499 GNDA.n133 GNDA.n132 585
R500 GNDA.n133 GNDA.n72 585
R501 GNDA.n135 GNDA.n134 585
R502 GNDA.n134 GNDA.n61 585
R503 GNDA.n91 GNDA.n90 585
R504 GNDA.n90 GNDA.n77 585
R505 GNDA.n89 GNDA.n88 585
R506 GNDA.n89 GNDA.n80 585
R507 GNDA.n94 GNDA.n87 585
R508 GNDA.n87 GNDA.t3 585
R509 GNDA.n96 GNDA.n95 585
R510 GNDA.n96 GNDA.n72 585
R511 GNDA.n98 GNDA.n97 585
R512 GNDA.n97 GNDA.n61 585
R513 GNDA.n328 GNDA.n323 585
R514 GNDA.n384 GNDA.n323 585
R515 GNDA.n327 GNDA.n78 585
R516 GNDA.n390 GNDA.n78 585
R517 GNDA.n376 GNDA.n375 585
R518 GNDA.n377 GNDA.n376 585
R519 GNDA.n374 GNDA.n70 585
R520 GNDA.n398 GNDA.n70 585
R521 GNDA.n373 GNDA.n372 585
R522 GNDA.n372 GNDA.n371 585
R523 GNDA.n344 GNDA.n62 585
R524 GNDA.n407 GNDA.n62 585
R525 GNDA.n343 GNDA.n342 585
R526 GNDA.n342 GNDA.n64 585
R527 GNDA.n341 GNDA.n54 585
R528 GNDA.n415 GNDA.n54 585
R529 GNDA.n340 GNDA.n339 585
R530 GNDA.n339 GNDA.n46 585
R531 GNDA.n338 GNDA.n47 585
R532 GNDA.n428 GNDA.n47 585
R533 GNDA.n36 GNDA.n35 585
R534 GNDA.n38 GNDA.n36 585
R535 GNDA.n439 GNDA.n438 585
R536 GNDA.n438 GNDA.n437 585
R537 GNDA.n37 GNDA.n33 585
R538 GNDA.n37 GNDA.n28 585
R539 GNDA.n442 GNDA.n29 585
R540 GNDA.n450 GNDA.n29 585
R541 GNDA.n386 GNDA.n385 585
R542 GNDA.n385 GNDA.n384 585
R543 GNDA.n389 GNDA.n388 585
R544 GNDA.n390 GNDA.n389 585
R545 GNDA.n69 GNDA.n68 585
R546 GNDA.n377 GNDA.n69 585
R547 GNDA.n400 GNDA.n399 585
R548 GNDA.n399 GNDA.n398 585
R549 GNDA.n66 GNDA.n65 585
R550 GNDA.n371 GNDA.n65 585
R551 GNDA.n406 GNDA.n405 585
R552 GNDA.n407 GNDA.n406 585
R553 GNDA.n53 GNDA.n52 585
R554 GNDA.n64 GNDA.n53 585
R555 GNDA.n417 GNDA.n416 585
R556 GNDA.n416 GNDA.n415 585
R557 GNDA.n51 GNDA.n49 585
R558 GNDA.n49 GNDA.n46 585
R559 GNDA.n427 GNDA.n426 585
R560 GNDA.n428 GNDA.n427 585
R561 GNDA.n425 GNDA.n50 585
R562 GNDA.n50 GNDA.n38 585
R563 GNDA.n424 GNDA.n40 585
R564 GNDA.n437 GNDA.n40 585
R565 GNDA.n423 GNDA.n27 585
R566 GNDA.n28 GNDA.n27 585
R567 GNDA.n452 GNDA.n451 585
R568 GNDA.n451 GNDA.n450 585
R569 GNDA.n383 GNDA.n382 585
R570 GNDA.n384 GNDA.n383 585
R571 GNDA.n324 GNDA.n79 585
R572 GNDA.n390 GNDA.n79 585
R573 GNDA.n379 GNDA.n378 585
R574 GNDA.n378 GNDA.n377 585
R575 GNDA.n326 GNDA.n71 585
R576 GNDA.n398 GNDA.n71 585
R577 GNDA.n370 GNDA.n369 585
R578 GNDA.n371 GNDA.n370 585
R579 GNDA.n368 GNDA.n63 585
R580 GNDA.n407 GNDA.n63 585
R581 GNDA.n367 GNDA.n366 585
R582 GNDA.n366 GNDA.n64 585
R583 GNDA.n365 GNDA.n55 585
R584 GNDA.n415 GNDA.n55 585
R585 GNDA.n364 GNDA.n363 585
R586 GNDA.n363 GNDA.n46 585
R587 GNDA.n362 GNDA.n48 585
R588 GNDA.n428 GNDA.n48 585
R589 GNDA.n361 GNDA.n360 585
R590 GNDA.n360 GNDA.n38 585
R591 GNDA.n359 GNDA.n39 585
R592 GNDA.n437 GNDA.n39 585
R593 GNDA.n358 GNDA.n357 585
R594 GNDA.n357 GNDA.n28 585
R595 GNDA.n355 GNDA.n30 585
R596 GNDA.n450 GNDA.n30 585
R597 GNDA.n283 GNDA.n282 585
R598 GNDA.n177 GNDA.n176 585
R599 GNDA.n178 GNDA.n177 585
R600 GNDA.n306 GNDA.n305 585
R601 GNDA.n305 GNDA.n304 585
R602 GNDA.n173 GNDA.n171 585
R603 GNDA.n171 GNDA.n146 585
R604 GNDA.n311 GNDA.n310 585
R605 GNDA.n312 GNDA.n311 585
R606 GNDA.n174 GNDA.n172 585
R607 GNDA.n172 GNDA.t8 585
R608 GNDA.n170 GNDA.n169 585
R609 GNDA.n312 GNDA.n170 585
R610 GNDA.n168 GNDA.n84 585
R611 GNDA.n84 GNDA.t8 585
R612 GNDA.n321 GNDA.n320 585
R613 GNDA.n322 GNDA.n321 585
R614 GNDA.n314 GNDA.n313 585
R615 GNDA.n313 GNDA.n312 585
R616 GNDA.n145 GNDA.n142 585
R617 GNDA.n145 GNDA.t8 585
R618 GNDA.n317 GNDA.n81 585
R619 GNDA.n322 GNDA.n81 585
R620 GNDA.n166 GNDA.n165 585
R621 GNDA.n312 GNDA.n166 585
R622 GNDA.n160 GNDA.n157 585
R623 GNDA.n157 GNDA.t8 585
R624 GNDA.n162 GNDA.n83 585
R625 GNDA.n322 GNDA.n83 585
R626 GNDA.n154 GNDA.n153 585
R627 GNDA.n312 GNDA.n154 585
R628 GNDA.n152 GNDA.n148 585
R629 GNDA.n148 GNDA.t8 585
R630 GNDA.n150 GNDA.n82 585
R631 GNDA.n322 GNDA.n82 585
R632 GNDA.n283 GNDA.n279 585
R633 GNDA.n190 GNDA.n189 585
R634 GNDA.n189 GNDA.n178 585
R635 GNDA.n276 GNDA.n179 585
R636 GNDA.n304 GNDA.n179 585
R637 GNDA.n275 GNDA.n274 585
R638 GNDA.n274 GNDA.n146 585
R639 GNDA.n273 GNDA.n147 585
R640 GNDA.n312 GNDA.n147 585
R641 GNDA.n271 GNDA.n270 585
R642 GNDA.n270 GNDA.t8 585
R643 GNDA.n283 GNDA.n281 585
R644 GNDA.n183 GNDA.n181 585
R645 GNDA.n181 GNDA.n178 585
R646 GNDA.n303 GNDA.n302 585
R647 GNDA.n304 GNDA.n303 585
R648 GNDA.n301 GNDA.n182 585
R649 GNDA.n182 GNDA.n146 585
R650 GNDA.n300 GNDA.n156 585
R651 GNDA.n312 GNDA.n156 585
R652 GNDA.n298 GNDA.n297 585
R653 GNDA.n297 GNDA.t8 585
R654 GNDA.n284 GNDA.n283 585
R655 GNDA.n188 GNDA.n187 585
R656 GNDA.n188 GNDA.n178 585
R657 GNDA.n287 GNDA.n180 585
R658 GNDA.n304 GNDA.n180 585
R659 GNDA.n289 GNDA.n288 585
R660 GNDA.n288 GNDA.n146 585
R661 GNDA.n186 GNDA.n155 585
R662 GNDA.n312 GNDA.n155 585
R663 GNDA.n293 GNDA.n292 585
R664 GNDA.n292 GNDA.t8 585
R665 GNDA.n239 GNDA.n196 585
R666 GNDA.t1 GNDA.n196 585
R667 GNDA.n264 GNDA.n263 585
R668 GNDA.n263 GNDA.n262 585
R669 GNDA.n232 GNDA.n228 585
R670 GNDA.n228 GNDA.t1 585
R671 GNDA.n230 GNDA.n209 585
R672 GNDA.n262 GNDA.n209 585
R673 GNDA.n224 GNDA.n211 585
R674 GNDA.n211 GNDA.t1 585
R675 GNDA.n261 GNDA.n260 585
R676 GNDA.n262 GNDA.n261 585
R677 GNDA.n214 GNDA.n213 585
R678 GNDA.n214 GNDA.t1 585
R679 GNDA.n258 GNDA.n210 585
R680 GNDA.n262 GNDA.n210 585
R681 GNDA.n241 GNDA.n240 585
R682 GNDA.n242 GNDA.n241 585
R683 GNDA.n234 GNDA.n233 585
R684 GNDA.n235 GNDA.n234 585
R685 GNDA.n226 GNDA.n225 585
R686 GNDA.n227 GNDA.n226 585
R687 GNDA.n255 GNDA.n254 585
R688 GNDA.n254 GNDA.n253 585
R689 GNDA.n386 GNDA.t112 555.914
R690 GNDA.n382 GNDA.t103 555.914
R691 GNDA.n75 GNDA.t83 555.914
R692 GNDA.n328 GNDA.t81 555.914
R693 GNDA.n240 GNDA.t77 514.141
R694 GNDA.n233 GNDA.t87 514.141
R695 GNDA.n225 GNDA.t79 514.141
R696 GNDA.n255 GNDA.t91 514.141
R697 GNDA.n169 GNDA.t73 514.141
R698 GNDA.n153 GNDA.t95 514.141
R699 GNDA.n143 GNDA.t101 510.483
R700 GNDA.n143 GNDA.t85 510.483
R701 GNDA.n158 GNDA.t89 510.483
R702 GNDA.n158 GNDA.t75 510.483
R703 GNDA.n242 GNDA.t1 453.435
R704 GNDA.n253 GNDA.t1 453.435
R705 GNDA.t43 GNDA.t24 369.466
R706 GNDA.t124 GNDA.t41 369.466
R707 GNDA.n207 GNDA.t114 349.817
R708 GNDA.n208 GNDA.t105 349.817
R709 GNDA.n307 GNDA.n175 267.125
R710 GNDA.n309 GNDA.n308 267.125
R711 GNDA.n278 GNDA.n277 267.125
R712 GNDA.n272 GNDA.n191 267.125
R713 GNDA.n280 GNDA.n184 267.125
R714 GNDA.n299 GNDA.n185 267.125
R715 GNDA.n286 GNDA.n285 267.125
R716 GNDA.n291 GNDA.n290 267.125
R717 GNDA.n387 GNDA.n67 267.125
R718 GNDA.n422 GNDA.n26 267.125
R719 GNDA.n381 GNDA.n380 267.125
R720 GNDA.n356 GNDA.n352 267.125
R721 GNDA.n394 GNDA.n393 267.125
R722 GNDA.n433 GNDA.n32 267.125
R723 GNDA.n330 GNDA.n329 267.125
R724 GNDA.n441 GNDA.n440 267.125
R725 GNDA.n384 GNDA.n322 258.046
R726 GNDA.n254 GNDA.n214 246.25
R727 GNDA.n214 GNDA.n210 246.25
R728 GNDA.n226 GNDA.n211 246.25
R729 GNDA.n261 GNDA.n211 246.25
R730 GNDA.n234 GNDA.n228 246.25
R731 GNDA.n228 GNDA.n209 246.25
R732 GNDA.n241 GNDA.n196 246.25
R733 GNDA.n263 GNDA.n196 246.25
R734 GNDA.n284 GNDA.n188 246.25
R735 GNDA.n188 GNDA.n180 246.25
R736 GNDA.n288 GNDA.n180 246.25
R737 GNDA.n288 GNDA.n155 246.25
R738 GNDA.n292 GNDA.n155 246.25
R739 GNDA.n281 GNDA.n181 246.25
R740 GNDA.n303 GNDA.n181 246.25
R741 GNDA.n303 GNDA.n182 246.25
R742 GNDA.n182 GNDA.n156 246.25
R743 GNDA.n297 GNDA.n156 246.25
R744 GNDA.n279 GNDA.n189 246.25
R745 GNDA.n189 GNDA.n179 246.25
R746 GNDA.n274 GNDA.n179 246.25
R747 GNDA.n274 GNDA.n147 246.25
R748 GNDA.n270 GNDA.n147 246.25
R749 GNDA.n154 GNDA.n148 246.25
R750 GNDA.n148 GNDA.n82 246.25
R751 GNDA.n166 GNDA.n157 246.25
R752 GNDA.n157 GNDA.n83 246.25
R753 GNDA.n313 GNDA.n145 246.25
R754 GNDA.n145 GNDA.n81 246.25
R755 GNDA.n170 GNDA.n84 246.25
R756 GNDA.n321 GNDA.n84 246.25
R757 GNDA.n282 GNDA.n177 246.25
R758 GNDA.n305 GNDA.n177 246.25
R759 GNDA.n305 GNDA.n171 246.25
R760 GNDA.n311 GNDA.n171 246.25
R761 GNDA.n311 GNDA.n172 246.25
R762 GNDA.n383 GNDA.n79 246.25
R763 GNDA.n378 GNDA.n79 246.25
R764 GNDA.n378 GNDA.n71 246.25
R765 GNDA.n370 GNDA.n71 246.25
R766 GNDA.n370 GNDA.n63 246.25
R767 GNDA.n366 GNDA.n63 246.25
R768 GNDA.n366 GNDA.n55 246.25
R769 GNDA.n363 GNDA.n55 246.25
R770 GNDA.n363 GNDA.n48 246.25
R771 GNDA.n360 GNDA.n48 246.25
R772 GNDA.n360 GNDA.n39 246.25
R773 GNDA.n357 GNDA.n39 246.25
R774 GNDA.n357 GNDA.n30 246.25
R775 GNDA.n389 GNDA.n385 246.25
R776 GNDA.n389 GNDA.n69 246.25
R777 GNDA.n399 GNDA.n69 246.25
R778 GNDA.n399 GNDA.n65 246.25
R779 GNDA.n406 GNDA.n65 246.25
R780 GNDA.n406 GNDA.n53 246.25
R781 GNDA.n416 GNDA.n53 246.25
R782 GNDA.n416 GNDA.n49 246.25
R783 GNDA.n427 GNDA.n49 246.25
R784 GNDA.n427 GNDA.n50 246.25
R785 GNDA.n50 GNDA.n40 246.25
R786 GNDA.n40 GNDA.n27 246.25
R787 GNDA.n451 GNDA.n27 246.25
R788 GNDA.n323 GNDA.n78 246.25
R789 GNDA.n376 GNDA.n78 246.25
R790 GNDA.n376 GNDA.n70 246.25
R791 GNDA.n372 GNDA.n70 246.25
R792 GNDA.n372 GNDA.n62 246.25
R793 GNDA.n342 GNDA.n62 246.25
R794 GNDA.n342 GNDA.n54 246.25
R795 GNDA.n339 GNDA.n54 246.25
R796 GNDA.n339 GNDA.n47 246.25
R797 GNDA.n47 GNDA.n36 246.25
R798 GNDA.n438 GNDA.n36 246.25
R799 GNDA.n438 GNDA.n37 246.25
R800 GNDA.n37 GNDA.n29 246.25
R801 GNDA.n90 GNDA.n89 246.25
R802 GNDA.n89 GNDA.n87 246.25
R803 GNDA.n96 GNDA.n87 246.25
R804 GNDA.n97 GNDA.n96 246.25
R805 GNDA.n127 GNDA.n126 246.25
R806 GNDA.n126 GNDA.n124 246.25
R807 GNDA.n133 GNDA.n124 246.25
R808 GNDA.n134 GNDA.n133 246.25
R809 GNDA.n391 GNDA.n76 246.25
R810 GNDA.n391 GNDA.n73 246.25
R811 GNDA.n397 GNDA.n73 246.25
R812 GNDA.n397 GNDA.n60 246.25
R813 GNDA.n408 GNDA.n60 246.25
R814 GNDA.n408 GNDA.n56 246.25
R815 GNDA.n414 GNDA.n56 246.25
R816 GNDA.n414 GNDA.n45 246.25
R817 GNDA.n429 GNDA.n45 246.25
R818 GNDA.n429 GNDA.n41 246.25
R819 GNDA.n436 GNDA.n41 246.25
R820 GNDA.n436 GNDA.n31 246.25
R821 GNDA.n449 GNDA.n31 246.25
R822 GNDA.t12 GNDA.t1 235.115
R823 GNDA.t33 GNDA.t1 235.115
R824 GNDA.n208 GNDA.t107 233
R825 GNDA.n207 GNDA.t116 233
R826 GNDA.n198 GNDA.n197 226.534
R827 GNDA.n200 GNDA.n199 226.534
R828 GNDA.n202 GNDA.n201 226.534
R829 GNDA.n204 GNDA.n203 226.534
R830 GNDA.n206 GNDA.n205 226.534
R831 GNDA.n235 GNDA.t12 218.321
R832 GNDA.n227 GNDA.t33 218.321
R833 GNDA.n14 GNDA.n12 206.052
R834 GNDA.n3 GNDA.n1 206.052
R835 GNDA.n22 GNDA.n21 205.488
R836 GNDA.n20 GNDA.n19 205.488
R837 GNDA.n18 GNDA.n17 205.488
R838 GNDA.n16 GNDA.n15 205.488
R839 GNDA.n14 GNDA.n13 205.488
R840 GNDA.n11 GNDA.n10 205.488
R841 GNDA.n9 GNDA.n8 205.488
R842 GNDA.n7 GNDA.n6 205.488
R843 GNDA.n5 GNDA.n4 205.488
R844 GNDA.n3 GNDA.n2 205.488
R845 GNDA.n233 GNDA.n229 185
R846 GNDA.n225 GNDA.n223 185
R847 GNDA.n256 GNDA.n255 185
R848 GNDA.n240 GNDA.n238 185
R849 GNDA.n315 GNDA.n314 185
R850 GNDA.n317 GNDA.n141 185
R851 GNDA.n165 GNDA.n164 185
R852 GNDA.n162 GNDA.n161 185
R853 GNDA.n153 GNDA.n149 185
R854 GNDA.n169 GNDA.n167 185
R855 GNDA.n277 GNDA.n276 185
R856 GNDA.n275 GNDA.n191 185
R857 GNDA.n307 GNDA.n306 185
R858 GNDA.n308 GNDA.n173 185
R859 GNDA.n92 GNDA.n91 185
R860 GNDA.n302 GNDA.n184 185
R861 GNDA.n301 GNDA.n185 185
R862 GNDA.n287 GNDA.n286 185
R863 GNDA.n290 GNDA.n289 185
R864 GNDA.n68 GNDA.n67 185
R865 GNDA.n401 GNDA.n400 185
R866 GNDA.n402 GNDA.n66 185
R867 GNDA.n405 GNDA.n404 185
R868 GNDA.n403 GNDA.n52 185
R869 GNDA.n418 GNDA.n417 185
R870 GNDA.n419 GNDA.n51 185
R871 GNDA.n426 GNDA.n420 185
R872 GNDA.n425 GNDA.n421 185
R873 GNDA.n424 GNDA.n422 185
R874 GNDA.n380 GNDA.n379 185
R875 GNDA.n326 GNDA.n325 185
R876 GNDA.n369 GNDA.n345 185
R877 GNDA.n368 GNDA.n346 185
R878 GNDA.n367 GNDA.n347 185
R879 GNDA.n365 GNDA.n348 185
R880 GNDA.n364 GNDA.n349 185
R881 GNDA.n362 GNDA.n350 185
R882 GNDA.n361 GNDA.n351 185
R883 GNDA.n359 GNDA.n352 185
R884 GNDA.n129 GNDA.n128 185
R885 GNDA.n375 GNDA.n330 185
R886 GNDA.n374 GNDA.n331 185
R887 GNDA.n373 GNDA.n332 185
R888 GNDA.n344 GNDA.n333 185
R889 GNDA.n343 GNDA.n334 185
R890 GNDA.n341 GNDA.n335 185
R891 GNDA.n340 GNDA.n336 185
R892 GNDA.n338 GNDA.n337 185
R893 GNDA.n35 GNDA.n34 185
R894 GNDA.n440 GNDA.n439 185
R895 GNDA.n394 GNDA.n74 185
R896 GNDA.n396 GNDA.n395 185
R897 GNDA.n59 GNDA.n58 185
R898 GNDA.n410 GNDA.n409 185
R899 GNDA.n411 GNDA.n57 185
R900 GNDA.n413 GNDA.n412 185
R901 GNDA.n44 GNDA.n43 185
R902 GNDA.n431 GNDA.n430 185
R903 GNDA.n432 GNDA.n42 185
R904 GNDA.n435 GNDA.n433 185
R905 GNDA.n236 GNDA.t43 184.733
R906 GNDA.n236 GNDA.t124 184.733
R907 GNDA.t24 GNDA.n235 151.145
R908 GNDA.t41 GNDA.n227 151.145
R909 GNDA.n401 GNDA.n67 150
R910 GNDA.n402 GNDA.n401 150
R911 GNDA.n404 GNDA.n402 150
R912 GNDA.n404 GNDA.n403 150
R913 GNDA.n419 GNDA.n418 150
R914 GNDA.n420 GNDA.n419 150
R915 GNDA.n421 GNDA.n420 150
R916 GNDA.n422 GNDA.n421 150
R917 GNDA.n380 GNDA.n325 150
R918 GNDA.n345 GNDA.n325 150
R919 GNDA.n346 GNDA.n345 150
R920 GNDA.n347 GNDA.n346 150
R921 GNDA.n349 GNDA.n348 150
R922 GNDA.n350 GNDA.n349 150
R923 GNDA.n351 GNDA.n350 150
R924 GNDA.n352 GNDA.n351 150
R925 GNDA.n395 GNDA.n394 150
R926 GNDA.n395 GNDA.n58 150
R927 GNDA.n410 GNDA.n58 150
R928 GNDA.n411 GNDA.n410 150
R929 GNDA.n412 GNDA.n43 150
R930 GNDA.n431 GNDA.n43 150
R931 GNDA.n432 GNDA.n431 150
R932 GNDA.n433 GNDA.n432 150
R933 GNDA.n331 GNDA.n330 150
R934 GNDA.n332 GNDA.n331 150
R935 GNDA.n333 GNDA.n332 150
R936 GNDA.n334 GNDA.n333 150
R937 GNDA.n336 GNDA.n335 150
R938 GNDA.n337 GNDA.n336 150
R939 GNDA.n337 GNDA.n34 150
R940 GNDA.n440 GNDA.n34 150
R941 GNDA.n262 GNDA.t20 102.888
R942 GNDA.n122 GNDA.n121 99.0842
R943 GNDA.n120 GNDA.n119 99.0842
R944 GNDA.n118 GNDA.n117 99.0842
R945 GNDA.n116 GNDA.n115 99.0842
R946 GNDA.n114 GNDA.n113 99.0842
R947 GNDA.n112 GNDA.n111 99.0842
R948 GNDA.n110 GNDA.n109 99.0842
R949 GNDA.n108 GNDA.n107 99.0842
R950 GNDA.n106 GNDA.n105 99.0842
R951 GNDA.n104 GNDA.n103 99.0842
R952 GNDA.n102 GNDA.n101 99.0842
R953 GNDA.n25 GNDA.n24 94.601
R954 GNDA.n354 GNDA.n353 94.601
R955 GNDA.n447 GNDA.n446 94.601
R956 GNDA.n445 GNDA.n444 94.601
R957 GNDA.n316 GNDA.n315 91.069
R958 GNDA.n144 GNDA.n141 91.069
R959 GNDA.n164 GNDA.n163 91.069
R960 GNDA.n161 GNDA.n159 91.069
R961 GNDA.n231 GNDA.n229 90.2704
R962 GNDA.n223 GNDA.n212 90.2704
R963 GNDA.n257 GNDA.n256 90.2704
R964 GNDA.n238 GNDA.n195 90.2704
R965 GNDA.n151 GNDA.n149 90.2704
R966 GNDA.n167 GNDA.n85 90.2704
R967 GNDA.n93 GNDA.n92 90.2704
R968 GNDA.n92 GNDA.n86 90.2704
R969 GNDA.n130 GNDA.n129 90.2704
R970 GNDA.n129 GNDA.n123 90.2704
R971 GNDA.t1 GNDA.t106 85.4967
R972 GNDA.t1 GNDA.t18 85.4967
R973 GNDA.t1 GNDA.t128 85.4967
R974 GNDA.t1 GNDA.t130 85.4967
R975 GNDA.t1 GNDA.t134 85.4967
R976 GNDA.t1 GNDA.t115 85.4967
R977 GNDA.t94 GNDA.n307 75.0005
R978 GNDA.n308 GNDA.t94 75.0005
R979 GNDA.n277 GNDA.t98 75.0005
R980 GNDA.n191 GNDA.t98 75.0005
R981 GNDA.t100 GNDA.n184 75.0005
R982 GNDA.n185 GNDA.t100 75.0005
R983 GNDA.n286 GNDA.t109 75.0005
R984 GNDA.n290 GNDA.t109 75.0005
R985 GNDA.n403 GNDA.t113 75.0005
R986 GNDA.n418 GNDA.t113 75.0005
R987 GNDA.t104 GNDA.n347 75.0005
R988 GNDA.n348 GNDA.t104 75.0005
R989 GNDA.t84 GNDA.n411 75.0005
R990 GNDA.n412 GNDA.t84 75.0005
R991 GNDA.t82 GNDA.n334 75.0005
R992 GNDA.n335 GNDA.t82 75.0005
R993 GNDA.n251 GNDA.t32 70.0746
R994 GNDA.t11 GNDA.t47 52.1486
R995 GNDA.n197 GNDA.t19 48.0005
R996 GNDA.n197 GNDA.t129 48.0005
R997 GNDA.n199 GNDA.t13 48.0005
R998 GNDA.n199 GNDA.t25 48.0005
R999 GNDA.n201 GNDA.t44 48.0005
R1000 GNDA.n201 GNDA.t125 48.0005
R1001 GNDA.n203 GNDA.t42 48.0005
R1002 GNDA.n203 GNDA.t34 48.0005
R1003 GNDA.n205 GNDA.t131 48.0005
R1004 GNDA.n205 GNDA.t135 48.0005
R1005 GNDA.n150 GNDA.n140 41.7462
R1006 GNDA.n259 GNDA.n258 40.6576
R1007 GNDA.t32 GNDA.t11 39.1116
R1008 GNDA.t2 GNDA.t7 39.1116
R1009 GNDA.t7 GNDA.t31 39.1116
R1010 GNDA.n355 GNDA.n354 37.7826
R1011 GNDA.n448 GNDA.n447 37.7826
R1012 GNDA.n320 GNDA.n319 37.4545
R1013 GNDA.n230 GNDA.n194 36.6576
R1014 GNDA.n260 GNDA.n259 36.6576
R1015 GNDA.n265 GNDA.n264 36.6576
R1016 GNDA.n453 GNDA.n452 36.6576
R1017 GNDA.n443 GNDA.n442 36.6576
R1018 GNDA.n318 GNDA.n317 36.1246
R1019 GNDA.n162 GNDA.n140 36.1246
R1020 GNDA.n456 GNDA.n11 35.938
R1021 GNDA.n455 GNDA.n22 35.688
R1022 GNDA.n207 GNDA.n206 33.563
R1023 GNDA.n262 GNDA.t1 33.0832
R1024 GNDA.n283 GNDA.n178 33.0832
R1025 GNDA.n304 GNDA.n178 33.0832
R1026 GNDA.n312 GNDA.n146 33.0832
R1027 GNDA.n312 GNDA.t8 33.0832
R1028 GNDA.n322 GNDA.t8 33.0832
R1029 GNDA.n407 GNDA.n64 33.0832
R1030 GNDA.n428 GNDA.n46 33.0832
R1031 GNDA.n428 GNDA.n38 33.0832
R1032 GNDA.n437 GNDA.n38 33.0832
R1033 GNDA.n450 GNDA.n28 33.0832
R1034 GNDA.n208 GNDA.n193 33.0005
R1035 GNDA.n236 GNDA.t1 29.7749
R1036 GNDA.t46 GNDA.t2 24.119
R1037 GNDA.t50 GNDA.n28 23.1584
R1038 GNDA.n99 GNDA.n98 22.8576
R1039 GNDA.n136 GNDA.n135 22.8576
R1040 GNDA GNDA.n457 22.617
R1041 GNDA.n271 GNDA.n269 20.7243
R1042 GNDA.n192 GNDA.n174 20.7243
R1043 GNDA.n298 GNDA.n296 20.7243
R1044 GNDA.n294 GNDA.n293 20.7243
R1045 GNDA.n21 GNDA.t65 19.7005
R1046 GNDA.n21 GNDA.t56 19.7005
R1047 GNDA.n19 GNDA.t66 19.7005
R1048 GNDA.n19 GNDA.t62 19.7005
R1049 GNDA.n17 GNDA.t68 19.7005
R1050 GNDA.n17 GNDA.t60 19.7005
R1051 GNDA.n15 GNDA.t69 19.7005
R1052 GNDA.n15 GNDA.t61 19.7005
R1053 GNDA.n13 GNDA.t67 19.7005
R1054 GNDA.n13 GNDA.t63 19.7005
R1055 GNDA.n12 GNDA.t15 19.7005
R1056 GNDA.n12 GNDA.t64 19.7005
R1057 GNDA.n10 GNDA.t126 19.7005
R1058 GNDA.n10 GNDA.t59 19.7005
R1059 GNDA.n8 GNDA.t35 19.7005
R1060 GNDA.n8 GNDA.t122 19.7005
R1061 GNDA.n6 GNDA.t36 19.7005
R1062 GNDA.n6 GNDA.t55 19.7005
R1063 GNDA.n4 GNDA.t117 19.7005
R1064 GNDA.n4 GNDA.t6 19.7005
R1065 GNDA.n2 GNDA.t118 19.7005
R1066 GNDA.n2 GNDA.t14 19.7005
R1067 GNDA.n1 GNDA.t21 19.7005
R1068 GNDA.n1 GNDA.t54 19.7005
R1069 GNDA.n251 GNDA.t39 19.1885
R1070 GNDA.n268 GNDA.n192 18.0765
R1071 GNDA.n295 GNDA.n294 18.0765
R1072 GNDA.n304 GNDA.t0 16.5419
R1073 GNDA.t0 GNDA.n146 16.5419
R1074 GNDA.n384 GNDA.n77 16.5419
R1075 GNDA.n390 GNDA.n77 16.5419
R1076 GNDA.n390 GNDA.n80 16.5419
R1077 GNDA.n377 GNDA.n80 16.5419
R1078 GNDA.n377 GNDA.t3 16.5419
R1079 GNDA.n398 GNDA.t3 16.5419
R1080 GNDA.n398 GNDA.n72 16.5419
R1081 GNDA.n371 GNDA.n72 16.5419
R1082 GNDA.n371 GNDA.n61 16.5419
R1083 GNDA.n407 GNDA.n61 16.5419
R1084 GNDA.n64 GNDA.t9 16.5419
R1085 GNDA.n415 GNDA.t9 16.5419
R1086 GNDA.n238 GNDA.t78 16.0005
R1087 GNDA.n229 GNDA.t88 16.0005
R1088 GNDA.n223 GNDA.t80 16.0005
R1089 GNDA.n256 GNDA.t92 16.0005
R1090 GNDA.n167 GNDA.t74 16.0005
R1091 GNDA.n141 GNDA.t102 16.0005
R1092 GNDA.n315 GNDA.t86 16.0005
R1093 GNDA.n161 GNDA.t90 16.0005
R1094 GNDA.n164 GNDA.t76 16.0005
R1095 GNDA.n149 GNDA.t96 16.0005
R1096 GNDA.t47 GNDA.t46 14.9931
R1097 GNDA.n269 GNDA.n268 14.0401
R1098 GNDA.n296 GNDA.n295 14.0401
R1099 GNDA.n100 GNDA.n99 13.8005
R1100 GNDA.n137 GNDA.n136 13.8005
R1101 GNDA.n456 GNDA.n455 13.313
R1102 GNDA.n415 GNDA.t39 12.2411
R1103 GNDA.n266 GNDA.n193 11.1567
R1104 GNDA.n437 GNDA.t50 9.92531
R1105 GNDA.n129 GNDA.t111 9.6005
R1106 GNDA.n121 GNDA.t5 9.6005
R1107 GNDA.n121 GNDA.t53 9.6005
R1108 GNDA.n119 GNDA.t57 9.6005
R1109 GNDA.n119 GNDA.t48 9.6005
R1110 GNDA.n117 GNDA.t27 9.6005
R1111 GNDA.n117 GNDA.t16 9.6005
R1112 GNDA.n115 GNDA.t58 9.6005
R1113 GNDA.n115 GNDA.t17 9.6005
R1114 GNDA.n113 GNDA.t133 9.6005
R1115 GNDA.n113 GNDA.t28 9.6005
R1116 GNDA.n111 GNDA.t29 9.6005
R1117 GNDA.n111 GNDA.t40 9.6005
R1118 GNDA.n109 GNDA.t120 9.6005
R1119 GNDA.n109 GNDA.t119 9.6005
R1120 GNDA.n107 GNDA.t127 9.6005
R1121 GNDA.n107 GNDA.t123 9.6005
R1122 GNDA.n105 GNDA.t37 9.6005
R1123 GNDA.n105 GNDA.t22 9.6005
R1124 GNDA.n103 GNDA.t23 9.6005
R1125 GNDA.n103 GNDA.t49 9.6005
R1126 GNDA.n101 GNDA.t4 9.6005
R1127 GNDA.n101 GNDA.t71 9.6005
R1128 GNDA.n92 GNDA.t72 9.6005
R1129 GNDA.n283 GNDA.t20 9.59449
R1130 GNDA.n233 GNDA.n232 9.14336
R1131 GNDA.n225 GNDA.n224 9.14336
R1132 GNDA.n255 GNDA.n213 9.14336
R1133 GNDA.n240 GNDA.n239 9.14336
R1134 GNDA.n153 GNDA.n152 9.14336
R1135 GNDA.n169 GNDA.n168 9.14336
R1136 GNDA.n276 GNDA.n190 9.14336
R1137 GNDA.n276 GNDA.n275 9.14336
R1138 GNDA.n275 GNDA.n273 9.14336
R1139 GNDA.n306 GNDA.n176 9.14336
R1140 GNDA.n306 GNDA.n173 9.14336
R1141 GNDA.n310 GNDA.n173 9.14336
R1142 GNDA.n91 GNDA.n88 9.14336
R1143 GNDA.n95 GNDA.n94 9.14336
R1144 GNDA.n302 GNDA.n183 9.14336
R1145 GNDA.n302 GNDA.n301 9.14336
R1146 GNDA.n301 GNDA.n300 9.14336
R1147 GNDA.n287 GNDA.n187 9.14336
R1148 GNDA.n289 GNDA.n287 9.14336
R1149 GNDA.n289 GNDA.n186 9.14336
R1150 GNDA.n388 GNDA.n68 9.14336
R1151 GNDA.n400 GNDA.n68 9.14336
R1152 GNDA.n400 GNDA.n66 9.14336
R1153 GNDA.n405 GNDA.n66 9.14336
R1154 GNDA.n405 GNDA.n52 9.14336
R1155 GNDA.n417 GNDA.n52 9.14336
R1156 GNDA.n417 GNDA.n51 9.14336
R1157 GNDA.n426 GNDA.n51 9.14336
R1158 GNDA.n426 GNDA.n425 9.14336
R1159 GNDA.n425 GNDA.n424 9.14336
R1160 GNDA.n424 GNDA.n423 9.14336
R1161 GNDA.n379 GNDA.n324 9.14336
R1162 GNDA.n379 GNDA.n326 9.14336
R1163 GNDA.n369 GNDA.n326 9.14336
R1164 GNDA.n369 GNDA.n368 9.14336
R1165 GNDA.n368 GNDA.n367 9.14336
R1166 GNDA.n367 GNDA.n365 9.14336
R1167 GNDA.n365 GNDA.n364 9.14336
R1168 GNDA.n364 GNDA.n362 9.14336
R1169 GNDA.n362 GNDA.n361 9.14336
R1170 GNDA.n361 GNDA.n359 9.14336
R1171 GNDA.n359 GNDA.n358 9.14336
R1172 GNDA.n128 GNDA.n125 9.14336
R1173 GNDA.n132 GNDA.n131 9.14336
R1174 GNDA.n375 GNDA.n327 9.14336
R1175 GNDA.n375 GNDA.n374 9.14336
R1176 GNDA.n374 GNDA.n373 9.14336
R1177 GNDA.n373 GNDA.n344 9.14336
R1178 GNDA.n344 GNDA.n343 9.14336
R1179 GNDA.n343 GNDA.n341 9.14336
R1180 GNDA.n341 GNDA.n340 9.14336
R1181 GNDA.n340 GNDA.n338 9.14336
R1182 GNDA.n338 GNDA.n35 9.14336
R1183 GNDA.n439 GNDA.n35 9.14336
R1184 GNDA.n439 GNDA.n33 9.14336
R1185 GNDA.n392 GNDA.n74 9.14336
R1186 GNDA.n396 GNDA.n74 9.14336
R1187 GNDA.n396 GNDA.n59 9.14336
R1188 GNDA.n409 GNDA.n59 9.14336
R1189 GNDA.n409 GNDA.n57 9.14336
R1190 GNDA.n413 GNDA.n57 9.14336
R1191 GNDA.n413 GNDA.n44 9.14336
R1192 GNDA.n430 GNDA.n44 9.14336
R1193 GNDA.n430 GNDA.n42 9.14336
R1194 GNDA.n435 GNDA.n42 9.14336
R1195 GNDA.n435 GNDA.n434 9.14336
R1196 GNDA.n295 GNDA.n23 9.1255
R1197 GNDA.n138 GNDA.n137 7.15675
R1198 GNDA.n100 GNDA.n23 7.03175
R1199 GNDA.n266 GNDA.n265 5.938
R1200 GNDA.n272 GNDA.n271 5.78934
R1201 GNDA.n309 GNDA.n174 5.78934
R1202 GNDA.n299 GNDA.n298 5.78934
R1203 GNDA.n293 GNDA.n291 5.78934
R1204 GNDA.n387 GNDA.n386 5.78934
R1205 GNDA.n452 GNDA.n26 5.78934
R1206 GNDA.n382 GNDA.n381 5.78934
R1207 GNDA.n356 GNDA.n355 5.78934
R1208 GNDA.n329 GNDA.n328 5.78934
R1209 GNDA.n442 GNDA.n441 5.78934
R1210 GNDA.n393 GNDA.n75 5.78934
R1211 GNDA.n448 GNDA.n32 5.78934
R1212 GNDA.n268 GNDA.n267 5.688
R1213 GNDA.n319 GNDA.n139 5.67758
R1214 GNDA.n443 GNDA.n0 5.563
R1215 GNDA.n454 GNDA.n453 5.313
R1216 GNDA.n455 GNDA.n454 5.03175
R1217 GNDA.n457 GNDA.n456 4.5005
R1218 GNDA.n232 GNDA.n231 4.46219
R1219 GNDA.n231 GNDA.n230 4.46219
R1220 GNDA.n224 GNDA.n212 4.46219
R1221 GNDA.n260 GNDA.n212 4.46219
R1222 GNDA.n257 GNDA.n213 4.46219
R1223 GNDA.n258 GNDA.n257 4.46219
R1224 GNDA.n239 GNDA.n195 4.46219
R1225 GNDA.n264 GNDA.n195 4.46219
R1226 GNDA.n152 GNDA.n151 4.46219
R1227 GNDA.n151 GNDA.n150 4.46219
R1228 GNDA.n168 GNDA.n85 4.46219
R1229 GNDA.n320 GNDA.n85 4.46219
R1230 GNDA.n93 GNDA.n88 4.46219
R1231 GNDA.n95 GNDA.n86 4.46219
R1232 GNDA.n94 GNDA.n93 4.46219
R1233 GNDA.n98 GNDA.n86 4.46219
R1234 GNDA.n130 GNDA.n125 4.46219
R1235 GNDA.n132 GNDA.n123 4.46219
R1236 GNDA.n131 GNDA.n130 4.46219
R1237 GNDA.n135 GNDA.n123 4.46219
R1238 GNDA.n319 GNDA.n318 4.29217
R1239 GNDA.n265 GNDA.n194 4.0005
R1240 GNDA.n24 GNDA.t132 3.42907
R1241 GNDA.n24 GNDA.t51 3.42907
R1242 GNDA.n353 GNDA.t10 3.42907
R1243 GNDA.n353 GNDA.t121 3.42907
R1244 GNDA.n446 GNDA.t38 3.42907
R1245 GNDA.n446 GNDA.t45 3.42907
R1246 GNDA.n444 GNDA.t26 3.42907
R1247 GNDA.n444 GNDA.t30 3.42907
R1248 GNDA.n278 GNDA.n190 3.19754
R1249 GNDA.n273 GNDA.n272 3.19754
R1250 GNDA.n176 GNDA.n175 3.19754
R1251 GNDA.n310 GNDA.n309 3.19754
R1252 GNDA.n280 GNDA.n183 3.19754
R1253 GNDA.n300 GNDA.n299 3.19754
R1254 GNDA.n285 GNDA.n187 3.19754
R1255 GNDA.n291 GNDA.n186 3.19754
R1256 GNDA.n388 GNDA.n387 3.19754
R1257 GNDA.n423 GNDA.n26 3.19754
R1258 GNDA.n381 GNDA.n324 3.19754
R1259 GNDA.n358 GNDA.n356 3.19754
R1260 GNDA.n329 GNDA.n327 3.19754
R1261 GNDA.n441 GNDA.n33 3.19754
R1262 GNDA.n393 GNDA.n392 3.19754
R1263 GNDA.n434 GNDA.n32 3.19754
R1264 GNDA.n144 GNDA.n142 2.86505
R1265 GNDA.n316 GNDA.n142 2.86505
R1266 GNDA.n317 GNDA.n316 2.86505
R1267 GNDA.n314 GNDA.n144 2.86505
R1268 GNDA.n160 GNDA.n159 2.86505
R1269 GNDA.n163 GNDA.n160 2.86505
R1270 GNDA.n163 GNDA.n162 2.86505
R1271 GNDA.n165 GNDA.n159 2.86505
R1272 GNDA.n267 GNDA.n266 2.84425
R1273 GNDA.n139 GNDA.n138 2.813
R1274 GNDA.n454 GNDA.n23 2.53175
R1275 GNDA.n138 GNDA.n0 2.46925
R1276 GNDA.n314 GNDA.n143 2.32777
R1277 GNDA.n165 GNDA.n158 2.32777
R1278 GNDA.n318 GNDA.n140 1.79217
R1279 GNDA.n259 GNDA.n194 1.688
R1280 GNDA.n251 GNDA.n46 1.65464
R1281 GNDA.n354 GNDA.n25 1.1255
R1282 GNDA.n453 GNDA.n25 1.1255
R1283 GNDA.n445 GNDA.n443 1.1255
R1284 GNDA.n447 GNDA.n445 1.1255
R1285 GNDA.n267 GNDA.n139 0.813
R1286 GNDA.n137 GNDA.n122 0.59425
R1287 GNDA.n16 GNDA.n14 0.563
R1288 GNDA.n18 GNDA.n16 0.563
R1289 GNDA.n20 GNDA.n18 0.563
R1290 GNDA.n22 GNDA.n20 0.563
R1291 GNDA.n5 GNDA.n3 0.563
R1292 GNDA.n7 GNDA.n5 0.563
R1293 GNDA.n9 GNDA.n7 0.563
R1294 GNDA.n11 GNDA.n9 0.563
R1295 GNDA.n104 GNDA.n102 0.563
R1296 GNDA.n106 GNDA.n104 0.563
R1297 GNDA.n108 GNDA.n106 0.563
R1298 GNDA.n110 GNDA.n108 0.563
R1299 GNDA.n112 GNDA.n110 0.563
R1300 GNDA.n114 GNDA.n112 0.563
R1301 GNDA.n116 GNDA.n114 0.563
R1302 GNDA.n118 GNDA.n116 0.563
R1303 GNDA.n120 GNDA.n118 0.563
R1304 GNDA.n122 GNDA.n120 0.563
R1305 GNDA.n206 GNDA.n204 0.563
R1306 GNDA.n204 GNDA.n202 0.563
R1307 GNDA.n202 GNDA.n200 0.563
R1308 GNDA.n200 GNDA.n198 0.563
R1309 GNDA.n198 GNDA.n193 0.563
R1310 GNDA.n457 GNDA.n0 0.53175
R1311 GNDA.n102 GNDA.n100 0.28175
R1312 Vb3.n19 Vb3.t22 661.375
R1313 Vb3.n13 Vb3.t18 611.739
R1314 Vb3.n9 Vb3.t11 611.739
R1315 Vb3.n4 Vb3.t21 611.739
R1316 Vb3.n0 Vb3.t9 611.739
R1317 Vb3.n13 Vb3.t20 421.75
R1318 Vb3.n14 Vb3.t5 421.75
R1319 Vb3.n15 Vb3.t10 421.75
R1320 Vb3.n16 Vb3.t14 421.75
R1321 Vb3.n9 Vb3.t7 421.75
R1322 Vb3.n10 Vb3.t17 421.75
R1323 Vb3.n11 Vb3.t15 421.75
R1324 Vb3.n12 Vb3.t12 421.75
R1325 Vb3.n4 Vb3.t6 421.75
R1326 Vb3.n5 Vb3.t3 421.75
R1327 Vb3.n6 Vb3.t8 421.75
R1328 Vb3.n7 Vb3.t13 421.75
R1329 Vb3.n0 Vb3.t4 421.75
R1330 Vb3.n1 Vb3.t19 421.75
R1331 Vb3.n2 Vb3.t2 421.75
R1332 Vb3.n3 Vb3.t16 421.75
R1333 Vb3.n19 Vb3.n18 181.37
R1334 Vb3.n20 Vb3.n17 176.25
R1335 Vb3 Vb3.n8 175.415
R1336 Vb3.n14 Vb3.n13 167.094
R1337 Vb3.n15 Vb3.n14 167.094
R1338 Vb3.n16 Vb3.n15 167.094
R1339 Vb3.n10 Vb3.n9 167.094
R1340 Vb3.n11 Vb3.n10 167.094
R1341 Vb3.n12 Vb3.n11 167.094
R1342 Vb3.n5 Vb3.n4 167.094
R1343 Vb3.n6 Vb3.n5 167.094
R1344 Vb3.n7 Vb3.n6 167.094
R1345 Vb3.n1 Vb3.n0 167.094
R1346 Vb3.n2 Vb3.n1 167.094
R1347 Vb3.n3 Vb3.n2 167.094
R1348 Vb3.n17 Vb3.n16 47.1294
R1349 Vb3.n17 Vb3.n12 47.1294
R1350 Vb3.n8 Vb3.n7 47.1294
R1351 Vb3.n8 Vb3.n3 47.1294
R1352 Vb3.n18 Vb3.t1 10.9449
R1353 Vb3.n18 Vb3.t0 10.9449
R1354 Vb3.n20 Vb3.n19 9.5005
R1355 Vb3 Vb3.n20 0.28175
R1356 VD3.n35 VD3.t32 680.832
R1357 VD3.n1 VD3.t35 680.832
R1358 VD3.n38 VD3.n37 585
R1359 VD3.n63 VD3.n1 585
R1360 VD3.n37 VD3.n20 290.233
R1361 VD3.n37 VD3.n21 290.233
R1362 VD3.n37 VD3.n36 290.233
R1363 VD3.n63 VD3.n0 290.233
R1364 VD3.n63 VD3.n62 290.233
R1365 VD3.n63 VD3.n2 290.233
R1366 VD3.n35 VD3.n34 238.367
R1367 VD3.n51 VD3.n50 238.367
R1368 VD3.n38 VD3.n18 185
R1369 VD3.n33 VD3.n18 185
R1370 VD3.n24 VD3.n19 185
R1371 VD3.n27 VD3.n26 185
R1372 VD3.n29 VD3.n28 185
R1373 VD3.n31 VD3.n30 185
R1374 VD3.n23 VD3.n22 185
R1375 VD3.n5 VD3.n4 185
R1376 VD3.n61 VD3.n60 185
R1377 VD3.n6 VD3.n3 185
R1378 VD3.n56 VD3.n55 185
R1379 VD3.n54 VD3.n53 185
R1380 VD3.n52 VD3.n1 185
R1381 VD3.n58 VD3.n52 185
R1382 VD3.n33 VD3.t33 170.513
R1383 VD3.n58 VD3.t36 170.513
R1384 VD3.n9 VD3.n7 160.427
R1385 VD3.n49 VD3.n48 159.803
R1386 VD3.n47 VD3.n46 159.803
R1387 VD3.n45 VD3.n44 159.803
R1388 VD3.n43 VD3.n42 159.803
R1389 VD3.n41 VD3.n40 159.803
R1390 VD3.n17 VD3.n16 159.802
R1391 VD3.n15 VD3.n14 159.802
R1392 VD3.n13 VD3.n12 159.802
R1393 VD3.n11 VD3.n10 159.802
R1394 VD3.n9 VD3.n8 159.802
R1395 VD3.n60 VD3.n5 150
R1396 VD3.n56 VD3.n6 150
R1397 VD3.n54 VD3.n52 150
R1398 VD3.n24 VD3.n18 150
R1399 VD3.n29 VD3.n26 150
R1400 VD3.n31 VD3.n23 150
R1401 VD3.t33 VD3.t16 146.155
R1402 VD3.t16 VD3.t22 146.155
R1403 VD3.t22 VD3.t28 146.155
R1404 VD3.t28 VD3.t30 146.155
R1405 VD3.t30 VD3.t12 146.155
R1406 VD3.t12 VD3.t14 146.155
R1407 VD3.t14 VD3.t18 146.155
R1408 VD3.t18 VD3.t24 146.155
R1409 VD3.t24 VD3.t20 146.155
R1410 VD3.t20 VD3.t26 146.155
R1411 VD3.t26 VD3.t36 146.155
R1412 VD3.n33 VD3.n25 65.8183
R1413 VD3.n33 VD3.n32 65.8183
R1414 VD3.n34 VD3.n33 65.8183
R1415 VD3.n58 VD3.n51 65.8183
R1416 VD3.n59 VD3.n58 65.8183
R1417 VD3.n58 VD3.n57 65.8183
R1418 VD3.n51 VD3.n5 53.3664
R1419 VD3.n60 VD3.n59 53.3664
R1420 VD3.n57 VD3.n56 53.3664
R1421 VD3.n25 VD3.n24 53.3664
R1422 VD3.n32 VD3.n29 53.3664
R1423 VD3.n34 VD3.n23 53.3664
R1424 VD3.n26 VD3.n25 53.3664
R1425 VD3.n32 VD3.n31 53.3664
R1426 VD3.n59 VD3.n6 53.3664
R1427 VD3.n57 VD3.n54 53.3664
R1428 VD3.n50 VD3.n49 37.2826
R1429 VD3.n39 VD3.n38 36.6576
R1430 VD3.n39 VD3.n17 13.688
R1431 VD3.n48 VD3.t21 11.2576
R1432 VD3.n48 VD3.t27 11.2576
R1433 VD3.n46 VD3.t19 11.2576
R1434 VD3.n46 VD3.t25 11.2576
R1435 VD3.n44 VD3.t13 11.2576
R1436 VD3.n44 VD3.t15 11.2576
R1437 VD3.n42 VD3.t29 11.2576
R1438 VD3.n42 VD3.t31 11.2576
R1439 VD3.n40 VD3.t17 11.2576
R1440 VD3.n40 VD3.t23 11.2576
R1441 VD3.n37 VD3.t34 11.2576
R1442 VD3.n16 VD3.t11 11.2576
R1443 VD3.n16 VD3.t1 11.2576
R1444 VD3.n14 VD3.t7 11.2576
R1445 VD3.n14 VD3.t2 11.2576
R1446 VD3.n12 VD3.t5 11.2576
R1447 VD3.n12 VD3.t3 11.2576
R1448 VD3.n10 VD3.t9 11.2576
R1449 VD3.n10 VD3.t6 11.2576
R1450 VD3.n8 VD3.t4 11.2576
R1451 VD3.n8 VD3.t10 11.2576
R1452 VD3.n7 VD3.t0 11.2576
R1453 VD3.n7 VD3.t8 11.2576
R1454 VD3.t37 VD3.n63 11.2576
R1455 VD3.n38 VD3.n19 9.14336
R1456 VD3.n28 VD3.n27 9.14336
R1457 VD3.n30 VD3.n22 9.14336
R1458 VD3.n61 VD3.n4 9.14336
R1459 VD3.n55 VD3.n3 9.14336
R1460 VD3.n53 VD3.n1 9.14336
R1461 VD3.n20 VD3.n19 4.53698
R1462 VD3.n28 VD3.n21 4.53698
R1463 VD3.n36 VD3.n22 4.53698
R1464 VD3.n27 VD3.n20 4.53698
R1465 VD3.n30 VD3.n21 4.53698
R1466 VD3.n36 VD3.n35 4.53698
R1467 VD3.n4 VD3.n0 4.53698
R1468 VD3.n62 VD3.n61 4.53698
R1469 VD3.n55 VD3.n2 4.53698
R1470 VD3.n62 VD3.n3 4.53698
R1471 VD3.n53 VD3.n2 4.53698
R1472 VD3.n50 VD3.n0 4.53698
R1473 VD3.n11 VD3.n9 0.6255
R1474 VD3.n13 VD3.n11 0.6255
R1475 VD3.n15 VD3.n13 0.6255
R1476 VD3.n17 VD3.n15 0.6255
R1477 VD3.n41 VD3.n39 0.6255
R1478 VD3.n43 VD3.n41 0.6255
R1479 VD3.n45 VD3.n43 0.6255
R1480 VD3.n47 VD3.n45 0.6255
R1481 VD3.n49 VD3.n47 0.6255
R1482 VDDA.n326 VDDA.t141 1095.3
R1483 VDDA.t129 VDDA.n325 1095.3
R1484 VDDA.t165 VDDA.n213 1095.3
R1485 VDDA.t144 VDDA.n35 1095.3
R1486 VDDA.n215 VDDA.t153 1082.5
R1487 VDDA.n36 VDDA.t147 1082.5
R1488 VDDA.t159 VDDA.n393 1003.33
R1489 VDDA.n394 VDDA.t168 1003.33
R1490 VDDA.n390 VDDA.t131 713.83
R1491 VDDA.n389 VDDA.t174 713.83
R1492 VDDA.n363 VDDA.t137 680.832
R1493 VDDA.n159 VDDA.t134 680.832
R1494 VDDA.n149 VDDA.t155 680.832
R1495 VDDA.n353 VDDA.t171 680.588
R1496 VDDA.n326 VDDA.t142 663.801
R1497 VDDA.n325 VDDA.t130 663.801
R1498 VDDA.n214 VDDA.t154 663.801
R1499 VDDA.n213 VDDA.t166 663.801
R1500 VDDA.n35 VDDA.t145 663.801
R1501 VDDA.n34 VDDA.t148 663.801
R1502 VDDA.n393 VDDA.t160 647.54
R1503 VDDA.n394 VDDA.t170 647.54
R1504 VDDA.n386 VDDA.n385 633.573
R1505 VDDA.n306 VDDA.n305 626.534
R1506 VDDA.n308 VDDA.n307 626.534
R1507 VDDA.n310 VDDA.n309 626.534
R1508 VDDA.n312 VDDA.n311 626.534
R1509 VDDA.n314 VDDA.n313 626.534
R1510 VDDA.n316 VDDA.n315 626.534
R1511 VDDA.n318 VDDA.n317 626.534
R1512 VDDA.n320 VDDA.n319 626.534
R1513 VDDA.n322 VDDA.n321 626.534
R1514 VDDA.n324 VDDA.n323 626.534
R1515 VDDA.n195 VDDA.t149 594.475
R1516 VDDA.n17 VDDA.t125 594.475
R1517 VDDA.n264 VDDA.n236 587.407
R1518 VDDA.n249 VDDA.n245 587.407
R1519 VDDA.n275 VDDA.n219 587.407
R1520 VDDA.n283 VDDA.n282 587.407
R1521 VDDA.n96 VDDA.n40 587.407
R1522 VDDA.n104 VDDA.n103 587.407
R1523 VDDA.n90 VDDA.n89 587.407
R1524 VDDA.n70 VDDA.n69 587.407
R1525 VDDA.n375 VDDA.n333 585
R1526 VDDA.n356 VDDA.n355 585
R1527 VDDA.n299 VDDA.n275 585
R1528 VDDA.n298 VDDA.n276 585
R1529 VDDA.n297 VDDA.n277 585
R1530 VDDA.n294 VDDA.n278 585
R1531 VDDA.n293 VDDA.n279 585
R1532 VDDA.n290 VDDA.n280 585
R1533 VDDA.n289 VDDA.n281 585
R1534 VDDA.n286 VDDA.n282 585
R1535 VDDA.n262 VDDA.n236 585
R1536 VDDA.n261 VDDA.n260 585
R1537 VDDA.n259 VDDA.n239 585
R1538 VDDA.n258 VDDA.n257 585
R1539 VDDA.n256 VDDA.n255 585
R1540 VDDA.n254 VDDA.n244 585
R1541 VDDA.n253 VDDA.n252 585
R1542 VDDA.n251 VDDA.n245 585
R1543 VDDA.n171 VDDA.n129 585
R1544 VDDA.n152 VDDA.n151 585
R1545 VDDA.n120 VDDA.n96 585
R1546 VDDA.n119 VDDA.n97 585
R1547 VDDA.n118 VDDA.n98 585
R1548 VDDA.n115 VDDA.n99 585
R1549 VDDA.n114 VDDA.n100 585
R1550 VDDA.n111 VDDA.n101 585
R1551 VDDA.n110 VDDA.n102 585
R1552 VDDA.n107 VDDA.n103 585
R1553 VDDA.n89 VDDA.n88 585
R1554 VDDA.n85 VDDA.n63 585
R1555 VDDA.n84 VDDA.n64 585
R1556 VDDA.n81 VDDA.n65 585
R1557 VDDA.n80 VDDA.n66 585
R1558 VDDA.n77 VDDA.n67 585
R1559 VDDA.n76 VDDA.n68 585
R1560 VDDA.n73 VDDA.n69 585
R1561 VDDA.t141 VDDA.t17 580.557
R1562 VDDA.t17 VDDA.t236 580.557
R1563 VDDA.t236 VDDA.t69 580.557
R1564 VDDA.t69 VDDA.t4 580.557
R1565 VDDA.t4 VDDA.t40 580.557
R1566 VDDA.t40 VDDA.t238 580.557
R1567 VDDA.t238 VDDA.t44 580.557
R1568 VDDA.t44 VDDA.t22 580.557
R1569 VDDA.t22 VDDA.t249 580.557
R1570 VDDA.t249 VDDA.t55 580.557
R1571 VDDA.t55 VDDA.t245 580.557
R1572 VDDA.t245 VDDA.t42 580.557
R1573 VDDA.t42 VDDA.t247 580.557
R1574 VDDA.t247 VDDA.t46 580.557
R1575 VDDA.t46 VDDA.t15 580.557
R1576 VDDA.t15 VDDA.t241 580.557
R1577 VDDA.t241 VDDA.t49 580.557
R1578 VDDA.t49 VDDA.t25 580.557
R1579 VDDA.t25 VDDA.t2 580.557
R1580 VDDA.t2 VDDA.t63 580.557
R1581 VDDA.t63 VDDA.t129 580.557
R1582 VDDA.t153 VDDA.t243 580.557
R1583 VDDA.t243 VDDA.t13 580.557
R1584 VDDA.t13 VDDA.t51 580.557
R1585 VDDA.t51 VDDA.t1 580.557
R1586 VDDA.t1 VDDA.t57 580.557
R1587 VDDA.t57 VDDA.t65 580.557
R1588 VDDA.t65 VDDA.t72 580.557
R1589 VDDA.t72 VDDA.t62 580.557
R1590 VDDA.t62 VDDA.t61 580.557
R1591 VDDA.t61 VDDA.t6 580.557
R1592 VDDA.t6 VDDA.t165 580.557
R1593 VDDA.t27 VDDA.t144 580.557
R1594 VDDA.t21 VDDA.t27 580.557
R1595 VDDA.t71 VDDA.t21 580.557
R1596 VDDA.t74 VDDA.t71 580.557
R1597 VDDA.t19 VDDA.t74 580.557
R1598 VDDA.t28 VDDA.t19 580.557
R1599 VDDA.t80 VDDA.t28 580.557
R1600 VDDA.t48 VDDA.t80 580.557
R1601 VDDA.t73 VDDA.t48 580.557
R1602 VDDA.t20 VDDA.t73 580.557
R1603 VDDA.t147 VDDA.t20 580.557
R1604 VDDA.n211 VDDA.t161 573.75
R1605 VDDA.n32 VDDA.t177 573.75
R1606 VDDA.t222 VDDA.t159 542.857
R1607 VDDA.t168 VDDA.t222 542.857
R1608 VDDA.n199 VDDA.t151 464.281
R1609 VDDA.t151 VDDA.n198 464.281
R1610 VDDA.n206 VDDA.t163 464.281
R1611 VDDA.t163 VDDA.n190 464.281
R1612 VDDA.n27 VDDA.t179 464.281
R1613 VDDA.t179 VDDA.n11 464.281
R1614 VDDA.n21 VDDA.t127 464.281
R1615 VDDA.t127 VDDA.n20 464.281
R1616 VDDA.n325 VDDA.t128 349.817
R1617 VDDA.n326 VDDA.t140 349.817
R1618 VDDA.n214 VDDA.t152 349.817
R1619 VDDA.n213 VDDA.t164 349.817
R1620 VDDA.n35 VDDA.t143 349.817
R1621 VDDA.n34 VDDA.t146 349.817
R1622 VDDA.n394 VDDA.t167 335.729
R1623 VDDA.n393 VDDA.t158 335.729
R1624 VDDA.n355 VDDA.n343 290.384
R1625 VDDA.n355 VDDA.n348 290.384
R1626 VDDA.n355 VDDA.n354 290.384
R1627 VDDA.n362 VDDA.n333 290.233
R1628 VDDA.n369 VDDA.n333 290.233
R1629 VDDA.n364 VDDA.n333 290.233
R1630 VDDA.n158 VDDA.n129 290.233
R1631 VDDA.n165 VDDA.n129 290.233
R1632 VDDA.n160 VDDA.n129 290.233
R1633 VDDA.n151 VDDA.n139 290.233
R1634 VDDA.n151 VDDA.n144 290.233
R1635 VDDA.n151 VDDA.n150 290.233
R1636 VDDA.t150 VDDA.n201 267.188
R1637 VDDA.n208 VDDA.t162 267.188
R1638 VDDA.n29 VDDA.t178 267.188
R1639 VDDA.t126 VDDA.n23 267.188
R1640 VDDA.n260 VDDA.n236 246.25
R1641 VDDA.n260 VDDA.n259 246.25
R1642 VDDA.n259 VDDA.n258 246.25
R1643 VDDA.n255 VDDA.n254 246.25
R1644 VDDA.n254 VDDA.n253 246.25
R1645 VDDA.n253 VDDA.n245 246.25
R1646 VDDA.n276 VDDA.n275 246.25
R1647 VDDA.n277 VDDA.n276 246.25
R1648 VDDA.n278 VDDA.n277 246.25
R1649 VDDA.n280 VDDA.n279 246.25
R1650 VDDA.n281 VDDA.n280 246.25
R1651 VDDA.n282 VDDA.n281 246.25
R1652 VDDA.n97 VDDA.n96 246.25
R1653 VDDA.n98 VDDA.n97 246.25
R1654 VDDA.n99 VDDA.n98 246.25
R1655 VDDA.n101 VDDA.n100 246.25
R1656 VDDA.n102 VDDA.n101 246.25
R1657 VDDA.n103 VDDA.n102 246.25
R1658 VDDA.n89 VDDA.n63 246.25
R1659 VDDA.n64 VDDA.n63 246.25
R1660 VDDA.n65 VDDA.n64 246.25
R1661 VDDA.n67 VDDA.n66 246.25
R1662 VDDA.n68 VDDA.n67 246.25
R1663 VDDA.n69 VDDA.n68 246.25
R1664 VDDA.n200 VDDA.n199 243.698
R1665 VDDA.n22 VDDA.n21 243.698
R1666 VDDA.n375 VDDA.n374 238.367
R1667 VDDA.n363 VDDA.n360 238.367
R1668 VDDA.n353 VDDA.n338 238.367
R1669 VDDA.n303 VDDA.n302 238.367
R1670 VDDA.n195 VDDA.n192 238.367
R1671 VDDA.n171 VDDA.n170 238.367
R1672 VDDA.n159 VDDA.n156 238.367
R1673 VDDA.n149 VDDA.n134 238.367
R1674 VDDA.n124 VDDA.n123 238.367
R1675 VDDA.n17 VDDA.n14 238.367
R1676 VDDA.t79 VDDA.t150 217.708
R1677 VDDA.t30 VDDA.t79 217.708
R1678 VDDA.t240 VDDA.t30 217.708
R1679 VDDA.t34 VDDA.t240 217.708
R1680 VDDA.t68 VDDA.t34 217.708
R1681 VDDA.t230 VDDA.t68 217.708
R1682 VDDA.t7 VDDA.t230 217.708
R1683 VDDA.t232 VDDA.t7 217.708
R1684 VDDA.t12 VDDA.t232 217.708
R1685 VDDA.t24 VDDA.t12 217.708
R1686 VDDA.t162 VDDA.t24 217.708
R1687 VDDA.t178 VDDA.t189 217.708
R1688 VDDA.t189 VDDA.t217 217.708
R1689 VDDA.t217 VDDA.t198 217.708
R1690 VDDA.t198 VDDA.t214 217.708
R1691 VDDA.t214 VDDA.t194 217.708
R1692 VDDA.t194 VDDA.t210 217.708
R1693 VDDA.t210 VDDA.t191 217.708
R1694 VDDA.t191 VDDA.t206 217.708
R1695 VDDA.t206 VDDA.t190 217.708
R1696 VDDA.t190 VDDA.t202 217.708
R1697 VDDA.t202 VDDA.t126 217.708
R1698 VDDA.n283 VDDA.n272 190.333
R1699 VDDA.n249 VDDA.n226 190.333
R1700 VDDA.n207 VDDA.n206 190.333
R1701 VDDA.n104 VDDA.n46 190.333
R1702 VDDA.n70 VDDA.n52 190.333
R1703 VDDA.n28 VDDA.n27 190.333
R1704 VDDA.t175 VDDA.n389 188.889
R1705 VDDA.n390 VDDA.t132 188.889
R1706 VDDA.n335 VDDA.n334 185
R1707 VDDA.n372 VDDA.n371 185
R1708 VDDA.n373 VDDA.n372 185
R1709 VDDA.n370 VDDA.n361 185
R1710 VDDA.n368 VDDA.n367 185
R1711 VDDA.n366 VDDA.n365 185
R1712 VDDA.n357 VDDA.n356 185
R1713 VDDA.n358 VDDA.n357 185
R1714 VDDA.n342 VDDA.n339 185
R1715 VDDA.n345 VDDA.n344 185
R1716 VDDA.n347 VDDA.n346 185
R1717 VDDA.n350 VDDA.n349 185
R1718 VDDA.n352 VDDA.n351 185
R1719 VDDA.n274 VDDA.n220 185
R1720 VDDA.n300 VDDA.n299 185
R1721 VDDA.n301 VDDA.n300 185
R1722 VDDA.n298 VDDA.n273 185
R1723 VDDA.n297 VDDA.n296 185
R1724 VDDA.n295 VDDA.n294 185
R1725 VDDA.n293 VDDA.n292 185
R1726 VDDA.n291 VDDA.n290 185
R1727 VDDA.n289 VDDA.n288 185
R1728 VDDA.n287 VDDA.n286 185
R1729 VDDA.n285 VDDA.n284 185
R1730 VDDA.n301 VDDA.n272 185
R1731 VDDA.n266 VDDA.n265 185
R1732 VDDA.n267 VDDA.n266 185
R1733 VDDA.n263 VDDA.n227 185
R1734 VDDA.n262 VDDA.n237 185
R1735 VDDA.n261 VDDA.n238 185
R1736 VDDA.n240 VDDA.n239 185
R1737 VDDA.n257 VDDA.n241 185
R1738 VDDA.n256 VDDA.n242 185
R1739 VDDA.n244 VDDA.n243 185
R1740 VDDA.n252 VDDA.n246 185
R1741 VDDA.n251 VDDA.n247 185
R1742 VDDA.n250 VDDA.n248 185
R1743 VDDA.n267 VDDA.n226 185
R1744 VDDA.n194 VDDA.n193 185
R1745 VDDA.n197 VDDA.n196 185
R1746 VDDA.n208 VDDA.n207 185
R1747 VDDA.n205 VDDA.n203 185
R1748 VDDA.n204 VDDA.n191 185
R1749 VDDA.n210 VDDA.n209 185
R1750 VDDA.n209 VDDA.n208 185
R1751 VDDA.n131 VDDA.n130 185
R1752 VDDA.n168 VDDA.n167 185
R1753 VDDA.n169 VDDA.n168 185
R1754 VDDA.n166 VDDA.n157 185
R1755 VDDA.n164 VDDA.n163 185
R1756 VDDA.n162 VDDA.n161 185
R1757 VDDA.n153 VDDA.n152 185
R1758 VDDA.n154 VDDA.n153 185
R1759 VDDA.n138 VDDA.n135 185
R1760 VDDA.n141 VDDA.n140 185
R1761 VDDA.n143 VDDA.n142 185
R1762 VDDA.n146 VDDA.n145 185
R1763 VDDA.n148 VDDA.n147 185
R1764 VDDA.n95 VDDA.n41 185
R1765 VDDA.n121 VDDA.n120 185
R1766 VDDA.n122 VDDA.n121 185
R1767 VDDA.n119 VDDA.n94 185
R1768 VDDA.n118 VDDA.n117 185
R1769 VDDA.n116 VDDA.n115 185
R1770 VDDA.n114 VDDA.n113 185
R1771 VDDA.n112 VDDA.n111 185
R1772 VDDA.n110 VDDA.n109 185
R1773 VDDA.n108 VDDA.n107 185
R1774 VDDA.n106 VDDA.n105 185
R1775 VDDA.n122 VDDA.n46 185
R1776 VDDA.n92 VDDA.n91 185
R1777 VDDA.n93 VDDA.n92 185
R1778 VDDA.n62 VDDA.n53 185
R1779 VDDA.n88 VDDA.n87 185
R1780 VDDA.n86 VDDA.n85 185
R1781 VDDA.n84 VDDA.n83 185
R1782 VDDA.n82 VDDA.n81 185
R1783 VDDA.n80 VDDA.n79 185
R1784 VDDA.n78 VDDA.n77 185
R1785 VDDA.n76 VDDA.n75 185
R1786 VDDA.n74 VDDA.n73 185
R1787 VDDA.n72 VDDA.n71 185
R1788 VDDA.n93 VDDA.n52 185
R1789 VDDA.n16 VDDA.n15 185
R1790 VDDA.n19 VDDA.n18 185
R1791 VDDA.n29 VDDA.n28 185
R1792 VDDA.n26 VDDA.n24 185
R1793 VDDA.n25 VDDA.n12 185
R1794 VDDA.n31 VDDA.n30 185
R1795 VDDA.n30 VDDA.n29 185
R1796 VDDA.t172 VDDA.n358 182.692
R1797 VDDA.n388 VDDA.n387 173.733
R1798 VDDA.n373 VDDA.t138 170.513
R1799 VDDA.t156 VDDA.n154 170.513
R1800 VDDA.n169 VDDA.t135 170.513
R1801 VDDA.n332 VDDA.n331 159.803
R1802 VDDA.n341 VDDA.n340 159.803
R1803 VDDA.n377 VDDA.n376 159.803
R1804 VDDA.n379 VDDA.n378 159.803
R1805 VDDA.n128 VDDA.n127 159.803
R1806 VDDA.n137 VDDA.n136 159.803
R1807 VDDA.n173 VDDA.n172 159.803
R1808 VDDA.n175 VDDA.n174 159.803
R1809 VDDA.n382 VDDA.n381 155.303
R1810 VDDA.n178 VDDA.n177 155.303
R1811 VDDA.n372 VDDA.n335 150
R1812 VDDA.n372 VDDA.n361 150
R1813 VDDA.n367 VDDA.n366 150
R1814 VDDA.n357 VDDA.n339 150
R1815 VDDA.n346 VDDA.n345 150
R1816 VDDA.n351 VDDA.n350 150
R1817 VDDA.n300 VDDA.n220 150
R1818 VDDA.n300 VDDA.n273 150
R1819 VDDA.n296 VDDA.n295 150
R1820 VDDA.n292 VDDA.n291 150
R1821 VDDA.n288 VDDA.n287 150
R1822 VDDA.n284 VDDA.n272 150
R1823 VDDA.n266 VDDA.n227 150
R1824 VDDA.n238 VDDA.n237 150
R1825 VDDA.n241 VDDA.n240 150
R1826 VDDA.n243 VDDA.n242 150
R1827 VDDA.n247 VDDA.n246 150
R1828 VDDA.n248 VDDA.n226 150
R1829 VDDA.n196 VDDA.n193 150
R1830 VDDA.n207 VDDA.n203 150
R1831 VDDA.n209 VDDA.n191 150
R1832 VDDA.n168 VDDA.n131 150
R1833 VDDA.n168 VDDA.n157 150
R1834 VDDA.n163 VDDA.n162 150
R1835 VDDA.n153 VDDA.n135 150
R1836 VDDA.n142 VDDA.n141 150
R1837 VDDA.n147 VDDA.n146 150
R1838 VDDA.n121 VDDA.n41 150
R1839 VDDA.n121 VDDA.n94 150
R1840 VDDA.n117 VDDA.n116 150
R1841 VDDA.n113 VDDA.n112 150
R1842 VDDA.n109 VDDA.n108 150
R1843 VDDA.n105 VDDA.n46 150
R1844 VDDA.n92 VDDA.n53 150
R1845 VDDA.n87 VDDA.n86 150
R1846 VDDA.n83 VDDA.n82 150
R1847 VDDA.n79 VDDA.n78 150
R1848 VDDA.n75 VDDA.n74 150
R1849 VDDA.n71 VDDA.n52 150
R1850 VDDA.n18 VDDA.n15 150
R1851 VDDA.n28 VDDA.n24 150
R1852 VDDA.n30 VDDA.n12 150
R1853 VDDA.t103 VDDA.t172 146.155
R1854 VDDA.t113 VDDA.t103 146.155
R1855 VDDA.t93 VDDA.t113 146.155
R1856 VDDA.t97 VDDA.t93 146.155
R1857 VDDA.t105 VDDA.t97 146.155
R1858 VDDA.t99 VDDA.t105 146.155
R1859 VDDA.t107 VDDA.t99 146.155
R1860 VDDA.t117 VDDA.t107 146.155
R1861 VDDA.t87 VDDA.t117 146.155
R1862 VDDA.t91 VDDA.t87 146.155
R1863 VDDA.t138 VDDA.t91 146.155
R1864 VDDA.t109 VDDA.t156 146.155
R1865 VDDA.t119 VDDA.t109 146.155
R1866 VDDA.t89 VDDA.t119 146.155
R1867 VDDA.t123 VDDA.t89 146.155
R1868 VDDA.t95 VDDA.t123 146.155
R1869 VDDA.t101 VDDA.t95 146.155
R1870 VDDA.t111 VDDA.t101 146.155
R1871 VDDA.t121 VDDA.t111 146.155
R1872 VDDA.t115 VDDA.t121 146.155
R1873 VDDA.t85 VDDA.t115 146.155
R1874 VDDA.t135 VDDA.t85 146.155
R1875 VDDA.n218 VDDA.n217 145.429
R1876 VDDA.n229 VDDA.n228 145.429
R1877 VDDA.n231 VDDA.n230 145.429
R1878 VDDA.n233 VDDA.n232 145.429
R1879 VDDA.n235 VDDA.n234 145.429
R1880 VDDA.n39 VDDA.n38 145.429
R1881 VDDA.n55 VDDA.n54 145.429
R1882 VDDA.n57 VDDA.n56 145.429
R1883 VDDA.n59 VDDA.n58 145.429
R1884 VDDA.n61 VDDA.n60 145.429
R1885 VDDA.t83 VDDA.t175 126.668
R1886 VDDA.t132 VDDA.t83 126.668
R1887 VDDA.n258 VDDA.t78 123.126
R1888 VDDA.n255 VDDA.t78 123.126
R1889 VDDA.t67 VDDA.n278 123.126
R1890 VDDA.n279 VDDA.t67 123.126
R1891 VDDA.t82 VDDA.n99 123.126
R1892 VDDA.n100 VDDA.t82 123.126
R1893 VDDA.t221 VDDA.n65 123.126
R1894 VDDA.n66 VDDA.t221 123.126
R1895 VDDA.t77 VDDA.n267 100.195
R1896 VDDA.n301 VDDA.t66 100.195
R1897 VDDA.n122 VDDA.t81 100.195
R1898 VDDA.t220 VDDA.n93 100.195
R1899 VDDA.n181 VDDA.n179 97.4034
R1900 VDDA.n2 VDDA.n0 97.4034
R1901 VDDA.n189 VDDA.n188 96.8409
R1902 VDDA.n187 VDDA.n186 96.8409
R1903 VDDA.n185 VDDA.n184 96.8409
R1904 VDDA.n183 VDDA.n182 96.8409
R1905 VDDA.n181 VDDA.n180 96.8409
R1906 VDDA.n10 VDDA.n9 96.8409
R1907 VDDA.n8 VDDA.n7 96.8409
R1908 VDDA.n6 VDDA.n5 96.8409
R1909 VDDA.n4 VDDA.n3 96.8409
R1910 VDDA.n2 VDDA.n1 96.8409
R1911 VDDA.t10 VDDA.t77 81.6411
R1912 VDDA.t31 VDDA.t10 81.6411
R1913 VDDA.t38 VDDA.t31 81.6411
R1914 VDDA.t58 VDDA.t38 81.6411
R1915 VDDA.t8 VDDA.t58 81.6411
R1916 VDDA.t228 VDDA.t8 81.6411
R1917 VDDA.t36 VDDA.t228 81.6411
R1918 VDDA.t233 VDDA.t36 81.6411
R1919 VDDA.t75 VDDA.t233 81.6411
R1920 VDDA.t52 VDDA.t75 81.6411
R1921 VDDA.t66 VDDA.t52 81.6411
R1922 VDDA.t81 VDDA.t183 81.6411
R1923 VDDA.t183 VDDA.t215 81.6411
R1924 VDDA.t215 VDDA.t195 81.6411
R1925 VDDA.t195 VDDA.t212 81.6411
R1926 VDDA.t212 VDDA.t192 81.6411
R1927 VDDA.t192 VDDA.t208 81.6411
R1928 VDDA.t208 VDDA.t180 81.6411
R1929 VDDA.t180 VDDA.t204 81.6411
R1930 VDDA.t204 VDDA.t185 81.6411
R1931 VDDA.t185 VDDA.t200 81.6411
R1932 VDDA.t200 VDDA.t220 81.6411
R1933 VDDA.n305 VDDA.t18 78.8005
R1934 VDDA.n305 VDDA.t237 78.8005
R1935 VDDA.n307 VDDA.t70 78.8005
R1936 VDDA.n307 VDDA.t5 78.8005
R1937 VDDA.n309 VDDA.t41 78.8005
R1938 VDDA.n309 VDDA.t239 78.8005
R1939 VDDA.n311 VDDA.t45 78.8005
R1940 VDDA.n311 VDDA.t23 78.8005
R1941 VDDA.n313 VDDA.t250 78.8005
R1942 VDDA.n313 VDDA.t56 78.8005
R1943 VDDA.n315 VDDA.t246 78.8005
R1944 VDDA.n315 VDDA.t43 78.8005
R1945 VDDA.n317 VDDA.t248 78.8005
R1946 VDDA.n317 VDDA.t47 78.8005
R1947 VDDA.n319 VDDA.t16 78.8005
R1948 VDDA.n319 VDDA.t242 78.8005
R1949 VDDA.n321 VDDA.t50 78.8005
R1950 VDDA.n321 VDDA.t26 78.8005
R1951 VDDA.n323 VDDA.t3 78.8005
R1952 VDDA.n323 VDDA.t64 78.8005
R1953 VDDA.n389 VDDA.t176 76.0991
R1954 VDDA.n390 VDDA.t133 76.0991
R1955 VDDA.n374 VDDA.n373 65.8183
R1956 VDDA.n373 VDDA.n359 65.8183
R1957 VDDA.n373 VDDA.n360 65.8183
R1958 VDDA.n358 VDDA.n336 65.8183
R1959 VDDA.n358 VDDA.n337 65.8183
R1960 VDDA.n358 VDDA.n338 65.8183
R1961 VDDA.n302 VDDA.n301 65.8183
R1962 VDDA.n301 VDDA.n268 65.8183
R1963 VDDA.n301 VDDA.n269 65.8183
R1964 VDDA.n301 VDDA.n270 65.8183
R1965 VDDA.n301 VDDA.n271 65.8183
R1966 VDDA.n267 VDDA.n221 65.8183
R1967 VDDA.n267 VDDA.n222 65.8183
R1968 VDDA.n267 VDDA.n223 65.8183
R1969 VDDA.n267 VDDA.n224 65.8183
R1970 VDDA.n267 VDDA.n225 65.8183
R1971 VDDA.n201 VDDA.n200 65.8183
R1972 VDDA.n201 VDDA.n192 65.8183
R1973 VDDA.n208 VDDA.n202 65.8183
R1974 VDDA.n170 VDDA.n169 65.8183
R1975 VDDA.n169 VDDA.n155 65.8183
R1976 VDDA.n169 VDDA.n156 65.8183
R1977 VDDA.n154 VDDA.n132 65.8183
R1978 VDDA.n154 VDDA.n133 65.8183
R1979 VDDA.n154 VDDA.n134 65.8183
R1980 VDDA.n123 VDDA.n122 65.8183
R1981 VDDA.n122 VDDA.n42 65.8183
R1982 VDDA.n122 VDDA.n43 65.8183
R1983 VDDA.n122 VDDA.n44 65.8183
R1984 VDDA.n122 VDDA.n45 65.8183
R1985 VDDA.n93 VDDA.n47 65.8183
R1986 VDDA.n93 VDDA.n48 65.8183
R1987 VDDA.n93 VDDA.n49 65.8183
R1988 VDDA.n93 VDDA.n50 65.8183
R1989 VDDA.n93 VDDA.n51 65.8183
R1990 VDDA.n23 VDDA.n22 65.8183
R1991 VDDA.n23 VDDA.n14 65.8183
R1992 VDDA.n29 VDDA.n13 65.8183
R1993 VDDA.n389 VDDA.n387 65.7076
R1994 VDDA.n391 VDDA.n390 65.4576
R1995 VDDA.n385 VDDA.t223 62.5402
R1996 VDDA.n385 VDDA.t169 62.5402
R1997 VDDA.n361 VDDA.n359 53.3664
R1998 VDDA.n366 VDDA.n360 53.3664
R1999 VDDA.n374 VDDA.n335 53.3664
R2000 VDDA.n367 VDDA.n359 53.3664
R2001 VDDA.n339 VDDA.n336 53.3664
R2002 VDDA.n346 VDDA.n337 53.3664
R2003 VDDA.n351 VDDA.n338 53.3664
R2004 VDDA.n345 VDDA.n336 53.3664
R2005 VDDA.n350 VDDA.n337 53.3664
R2006 VDDA.n273 VDDA.n268 53.3664
R2007 VDDA.n295 VDDA.n269 53.3664
R2008 VDDA.n291 VDDA.n270 53.3664
R2009 VDDA.n287 VDDA.n271 53.3664
R2010 VDDA.n302 VDDA.n220 53.3664
R2011 VDDA.n296 VDDA.n268 53.3664
R2012 VDDA.n292 VDDA.n269 53.3664
R2013 VDDA.n288 VDDA.n270 53.3664
R2014 VDDA.n284 VDDA.n271 53.3664
R2015 VDDA.n227 VDDA.n221 53.3664
R2016 VDDA.n238 VDDA.n222 53.3664
R2017 VDDA.n241 VDDA.n223 53.3664
R2018 VDDA.n243 VDDA.n224 53.3664
R2019 VDDA.n247 VDDA.n225 53.3664
R2020 VDDA.n237 VDDA.n221 53.3664
R2021 VDDA.n240 VDDA.n222 53.3664
R2022 VDDA.n242 VDDA.n223 53.3664
R2023 VDDA.n246 VDDA.n224 53.3664
R2024 VDDA.n248 VDDA.n225 53.3664
R2025 VDDA.n200 VDDA.n193 53.3664
R2026 VDDA.n196 VDDA.n192 53.3664
R2027 VDDA.n203 VDDA.n202 53.3664
R2028 VDDA.n202 VDDA.n191 53.3664
R2029 VDDA.n157 VDDA.n155 53.3664
R2030 VDDA.n162 VDDA.n156 53.3664
R2031 VDDA.n170 VDDA.n131 53.3664
R2032 VDDA.n163 VDDA.n155 53.3664
R2033 VDDA.n135 VDDA.n132 53.3664
R2034 VDDA.n142 VDDA.n133 53.3664
R2035 VDDA.n147 VDDA.n134 53.3664
R2036 VDDA.n141 VDDA.n132 53.3664
R2037 VDDA.n146 VDDA.n133 53.3664
R2038 VDDA.n94 VDDA.n42 53.3664
R2039 VDDA.n116 VDDA.n43 53.3664
R2040 VDDA.n112 VDDA.n44 53.3664
R2041 VDDA.n108 VDDA.n45 53.3664
R2042 VDDA.n123 VDDA.n41 53.3664
R2043 VDDA.n117 VDDA.n42 53.3664
R2044 VDDA.n113 VDDA.n43 53.3664
R2045 VDDA.n109 VDDA.n44 53.3664
R2046 VDDA.n105 VDDA.n45 53.3664
R2047 VDDA.n53 VDDA.n47 53.3664
R2048 VDDA.n86 VDDA.n48 53.3664
R2049 VDDA.n82 VDDA.n49 53.3664
R2050 VDDA.n78 VDDA.n50 53.3664
R2051 VDDA.n74 VDDA.n51 53.3664
R2052 VDDA.n87 VDDA.n47 53.3664
R2053 VDDA.n83 VDDA.n48 53.3664
R2054 VDDA.n79 VDDA.n49 53.3664
R2055 VDDA.n75 VDDA.n50 53.3664
R2056 VDDA.n71 VDDA.n51 53.3664
R2057 VDDA.n22 VDDA.n15 53.3664
R2058 VDDA.n18 VDDA.n14 53.3664
R2059 VDDA.n24 VDDA.n13 53.3664
R2060 VDDA.n13 VDDA.n12 53.3664
R2061 VDDA.n395 VDDA.n394 41.5034
R2062 VDDA.n377 VDDA.n375 37.2826
R2063 VDDA.n173 VDDA.n171 37.2826
R2064 VDDA.n152 VDDA.n137 37.2826
R2065 VDDA.n265 VDDA.n235 37.2201
R2066 VDDA.n91 VDDA.n61 37.2201
R2067 VDDA.n356 VDDA.n341 37.0388
R2068 VDDA.n393 VDDA.n392 37.0034
R2069 VDDA.n304 VDDA.n303 36.6576
R2070 VDDA.n125 VDDA.n124 36.6576
R2071 VDDA.n325 VDDA.n324 33.563
R2072 VDDA.n327 VDDA.n326 33.0005
R2073 VDDA VDDA.n396 25.2335
R2074 VDDA.n211 VDDA.n210 20.7243
R2075 VDDA.n216 VDDA.n215 19.7067
R2076 VDDA.n37 VDDA.n36 19.6755
R2077 VDDA.n33 VDDA.n32 19.238
R2078 VDDA.n212 VDDA.n211 19.2067
R2079 VDDA.n32 VDDA.n31 18.591
R2080 VDDA.n383 VDDA.n330 13.5943
R2081 VDDA.n215 VDDA.n214 12.8005
R2082 VDDA.n36 VDDA.n34 12.8005
R2083 VDDA.n381 VDDA.t106 11.2576
R2084 VDDA.n381 VDDA.t100 11.2576
R2085 VDDA.n331 VDDA.t94 11.2576
R2086 VDDA.n331 VDDA.t98 11.2576
R2087 VDDA.n340 VDDA.t104 11.2576
R2088 VDDA.n340 VDDA.t114 11.2576
R2089 VDDA.n355 VDDA.t173 11.2576
R2090 VDDA.n333 VDDA.t139 11.2576
R2091 VDDA.n376 VDDA.t88 11.2576
R2092 VDDA.n376 VDDA.t92 11.2576
R2093 VDDA.n378 VDDA.t108 11.2576
R2094 VDDA.n378 VDDA.t118 11.2576
R2095 VDDA.n177 VDDA.t96 11.2576
R2096 VDDA.n177 VDDA.t102 11.2576
R2097 VDDA.n127 VDDA.t90 11.2576
R2098 VDDA.n127 VDDA.t124 11.2576
R2099 VDDA.n136 VDDA.t110 11.2576
R2100 VDDA.n136 VDDA.t120 11.2576
R2101 VDDA.n151 VDDA.t157 11.2576
R2102 VDDA.n129 VDDA.t136 11.2576
R2103 VDDA.n172 VDDA.t116 11.2576
R2104 VDDA.n172 VDDA.t86 11.2576
R2105 VDDA.n174 VDDA.t112 11.2576
R2106 VDDA.n174 VDDA.t122 11.2576
R2107 VDDA.t176 VDDA.n388 11.0991
R2108 VDDA.n388 VDDA.t84 11.0991
R2109 VDDA.n330 VDDA.n329 9.5005
R2110 VDDA.n392 VDDA.n391 9.23175
R2111 VDDA.n33 VDDA.n10 9.15675
R2112 VDDA.n375 VDDA.n334 9.14336
R2113 VDDA.n371 VDDA.n370 9.14336
R2114 VDDA.n368 VDDA.n365 9.14336
R2115 VDDA.n299 VDDA.n274 9.14336
R2116 VDDA.n299 VDDA.n298 9.14336
R2117 VDDA.n298 VDDA.n297 9.14336
R2118 VDDA.n297 VDDA.n294 9.14336
R2119 VDDA.n294 VDDA.n293 9.14336
R2120 VDDA.n293 VDDA.n290 9.14336
R2121 VDDA.n290 VDDA.n289 9.14336
R2122 VDDA.n289 VDDA.n286 9.14336
R2123 VDDA.n286 VDDA.n285 9.14336
R2124 VDDA.n263 VDDA.n262 9.14336
R2125 VDDA.n262 VDDA.n261 9.14336
R2126 VDDA.n261 VDDA.n239 9.14336
R2127 VDDA.n257 VDDA.n239 9.14336
R2128 VDDA.n257 VDDA.n256 9.14336
R2129 VDDA.n256 VDDA.n244 9.14336
R2130 VDDA.n252 VDDA.n244 9.14336
R2131 VDDA.n252 VDDA.n251 9.14336
R2132 VDDA.n251 VDDA.n250 9.14336
R2133 VDDA.n197 VDDA.n194 9.14336
R2134 VDDA.n205 VDDA.n204 9.14336
R2135 VDDA.n171 VDDA.n130 9.14336
R2136 VDDA.n167 VDDA.n166 9.14336
R2137 VDDA.n164 VDDA.n161 9.14336
R2138 VDDA.n152 VDDA.n138 9.14336
R2139 VDDA.n143 VDDA.n140 9.14336
R2140 VDDA.n148 VDDA.n145 9.14336
R2141 VDDA.n120 VDDA.n95 9.14336
R2142 VDDA.n120 VDDA.n119 9.14336
R2143 VDDA.n119 VDDA.n118 9.14336
R2144 VDDA.n118 VDDA.n115 9.14336
R2145 VDDA.n115 VDDA.n114 9.14336
R2146 VDDA.n114 VDDA.n111 9.14336
R2147 VDDA.n111 VDDA.n110 9.14336
R2148 VDDA.n110 VDDA.n107 9.14336
R2149 VDDA.n107 VDDA.n106 9.14336
R2150 VDDA.n88 VDDA.n62 9.14336
R2151 VDDA.n88 VDDA.n85 9.14336
R2152 VDDA.n85 VDDA.n84 9.14336
R2153 VDDA.n84 VDDA.n81 9.14336
R2154 VDDA.n81 VDDA.n80 9.14336
R2155 VDDA.n80 VDDA.n77 9.14336
R2156 VDDA.n77 VDDA.n76 9.14336
R2157 VDDA.n76 VDDA.n73 9.14336
R2158 VDDA.n73 VDDA.n72 9.14336
R2159 VDDA.n19 VDDA.n16 9.14336
R2160 VDDA.n26 VDDA.n25 9.14336
R2161 VDDA.n212 VDDA.n189 9.1255
R2162 VDDA.n356 VDDA.n342 8.53383
R2163 VDDA.n347 VDDA.n344 8.53383
R2164 VDDA.n352 VDDA.n349 8.53383
R2165 VDDA.n188 VDDA.t244 8.0005
R2166 VDDA.n188 VDDA.t225 8.0005
R2167 VDDA.n186 VDDA.t33 8.0005
R2168 VDDA.n186 VDDA.t231 8.0005
R2169 VDDA.n184 VDDA.t235 8.0005
R2170 VDDA.n184 VDDA.t54 8.0005
R2171 VDDA.n182 VDDA.t35 8.0005
R2172 VDDA.n182 VDDA.t0 8.0005
R2173 VDDA.n180 VDDA.t60 8.0005
R2174 VDDA.n180 VDDA.t14 8.0005
R2175 VDDA.n179 VDDA.t224 8.0005
R2176 VDDA.n179 VDDA.t29 8.0005
R2177 VDDA.n9 VDDA.t226 8.0005
R2178 VDDA.n9 VDDA.t218 8.0005
R2179 VDDA.n7 VDDA.t211 8.0005
R2180 VDDA.n7 VDDA.t187 8.0005
R2181 VDDA.n5 VDDA.t207 8.0005
R2182 VDDA.n5 VDDA.t188 8.0005
R2183 VDDA.n3 VDDA.t203 8.0005
R2184 VDDA.n3 VDDA.t182 8.0005
R2185 VDDA.n1 VDDA.t197 8.0005
R2186 VDDA.n1 VDDA.t219 8.0005
R2187 VDDA.n0 VDDA.t199 8.0005
R2188 VDDA.n0 VDDA.t227 8.0005
R2189 VDDA.n383 VDDA.n382 7.8755
R2190 VDDA.n330 VDDA.n178 7.84425
R2191 VDDA.n396 VDDA.n395 6.6255
R2192 VDDA.n217 VDDA.t76 6.56717
R2193 VDDA.n217 VDDA.t53 6.56717
R2194 VDDA.n228 VDDA.t37 6.56717
R2195 VDDA.n228 VDDA.t234 6.56717
R2196 VDDA.n230 VDDA.t9 6.56717
R2197 VDDA.n230 VDDA.t229 6.56717
R2198 VDDA.n232 VDDA.t39 6.56717
R2199 VDDA.n232 VDDA.t59 6.56717
R2200 VDDA.n234 VDDA.t11 6.56717
R2201 VDDA.n234 VDDA.t32 6.56717
R2202 VDDA.n38 VDDA.t184 6.56717
R2203 VDDA.n38 VDDA.t216 6.56717
R2204 VDDA.n54 VDDA.t196 6.56717
R2205 VDDA.n54 VDDA.t213 6.56717
R2206 VDDA.n56 VDDA.t193 6.56717
R2207 VDDA.n56 VDDA.t209 6.56717
R2208 VDDA.n58 VDDA.t181 6.56717
R2209 VDDA.n58 VDDA.t205 6.56717
R2210 VDDA.n60 VDDA.t186 6.56717
R2211 VDDA.n60 VDDA.t201 6.56717
R2212 VDDA.n126 VDDA.n125 5.438
R2213 VDDA.n265 VDDA.n264 5.33286
R2214 VDDA.n303 VDDA.n219 5.33286
R2215 VDDA.n198 VDDA.n195 5.33286
R2216 VDDA.n210 VDDA.n190 5.33286
R2217 VDDA.n124 VDDA.n40 5.33286
R2218 VDDA.n91 VDDA.n90 5.33286
R2219 VDDA.n20 VDDA.n17 5.33286
R2220 VDDA.n31 VDDA.n11 5.33286
R2221 VDDA.n392 VDDA.n386 5.1255
R2222 VDDA.n384 VDDA.n126 5.0005
R2223 VDDA.n362 VDDA.n334 4.53698
R2224 VDDA.n370 VDDA.n369 4.53698
R2225 VDDA.n365 VDDA.n364 4.53698
R2226 VDDA.n371 VDDA.n362 4.53698
R2227 VDDA.n369 VDDA.n368 4.53698
R2228 VDDA.n364 VDDA.n363 4.53698
R2229 VDDA.n158 VDDA.n130 4.53698
R2230 VDDA.n166 VDDA.n165 4.53698
R2231 VDDA.n161 VDDA.n160 4.53698
R2232 VDDA.n167 VDDA.n158 4.53698
R2233 VDDA.n165 VDDA.n164 4.53698
R2234 VDDA.n160 VDDA.n159 4.53698
R2235 VDDA.n139 VDDA.n138 4.53698
R2236 VDDA.n144 VDDA.n143 4.53698
R2237 VDDA.n150 VDDA.n148 4.53698
R2238 VDDA.n140 VDDA.n139 4.53698
R2239 VDDA.n145 VDDA.n144 4.53698
R2240 VDDA.n150 VDDA.n149 4.53698
R2241 VDDA.n382 VDDA.n380 4.5005
R2242 VDDA.n329 VDDA.n328 4.5005
R2243 VDDA.n178 VDDA.n176 4.5005
R2244 VDDA.n384 VDDA.n383 4.5005
R2245 VDDA.n216 VDDA.n212 4.34425
R2246 VDDA.n37 VDDA.n33 4.34425
R2247 VDDA.n343 VDDA.n342 4.23677
R2248 VDDA.n348 VDDA.n347 4.23677
R2249 VDDA.n354 VDDA.n352 4.23677
R2250 VDDA.n344 VDDA.n343 4.23677
R2251 VDDA.n349 VDDA.n348 4.23677
R2252 VDDA.n354 VDDA.n353 4.23677
R2253 VDDA.n274 VDDA.n219 3.75335
R2254 VDDA.n285 VDDA.n283 3.75335
R2255 VDDA.n264 VDDA.n263 3.75335
R2256 VDDA.n250 VDDA.n249 3.75335
R2257 VDDA.n199 VDDA.n194 3.75335
R2258 VDDA.n198 VDDA.n197 3.75335
R2259 VDDA.n206 VDDA.n205 3.75335
R2260 VDDA.n204 VDDA.n190 3.75335
R2261 VDDA.n95 VDDA.n40 3.75335
R2262 VDDA.n106 VDDA.n104 3.75335
R2263 VDDA.n90 VDDA.n62 3.75335
R2264 VDDA.n72 VDDA.n70 3.75335
R2265 VDDA.n21 VDDA.n16 3.75335
R2266 VDDA.n20 VDDA.n19 3.75335
R2267 VDDA.n27 VDDA.n26 3.75335
R2268 VDDA.n25 VDDA.n11 3.75335
R2269 VDDA.n329 VDDA.n216 3.09425
R2270 VDDA.n126 VDDA.n37 3.09425
R2271 VDDA.n328 VDDA.n327 2.96925
R2272 VDDA.n396 VDDA.n384 1.95675
R2273 VDDA.n328 VDDA.n304 0.90675
R2274 VDDA.n391 VDDA.n387 0.6255
R2275 VDDA.n380 VDDA.n379 0.6255
R2276 VDDA.n379 VDDA.n377 0.6255
R2277 VDDA.n341 VDDA.n332 0.6255
R2278 VDDA.n380 VDDA.n332 0.6255
R2279 VDDA.n176 VDDA.n175 0.6255
R2280 VDDA.n175 VDDA.n173 0.6255
R2281 VDDA.n137 VDDA.n128 0.6255
R2282 VDDA.n176 VDDA.n128 0.6255
R2283 VDDA.n324 VDDA.n322 0.563
R2284 VDDA.n322 VDDA.n320 0.563
R2285 VDDA.n320 VDDA.n318 0.563
R2286 VDDA.n318 VDDA.n316 0.563
R2287 VDDA.n316 VDDA.n314 0.563
R2288 VDDA.n314 VDDA.n312 0.563
R2289 VDDA.n312 VDDA.n310 0.563
R2290 VDDA.n310 VDDA.n308 0.563
R2291 VDDA.n308 VDDA.n306 0.563
R2292 VDDA.n327 VDDA.n306 0.563
R2293 VDDA.n235 VDDA.n233 0.563
R2294 VDDA.n233 VDDA.n231 0.563
R2295 VDDA.n231 VDDA.n229 0.563
R2296 VDDA.n229 VDDA.n218 0.563
R2297 VDDA.n304 VDDA.n218 0.563
R2298 VDDA.n183 VDDA.n181 0.563
R2299 VDDA.n185 VDDA.n183 0.563
R2300 VDDA.n187 VDDA.n185 0.563
R2301 VDDA.n189 VDDA.n187 0.563
R2302 VDDA.n61 VDDA.n59 0.563
R2303 VDDA.n59 VDDA.n57 0.563
R2304 VDDA.n57 VDDA.n55 0.563
R2305 VDDA.n55 VDDA.n39 0.563
R2306 VDDA.n125 VDDA.n39 0.563
R2307 VDDA.n4 VDDA.n2 0.563
R2308 VDDA.n6 VDDA.n4 0.563
R2309 VDDA.n8 VDDA.n6 0.563
R2310 VDDA.n10 VDDA.n8 0.563
R2311 VDDA.n395 VDDA.n386 0.2505
R2312 X.n13 X.t50 1172.87
R2313 X.n11 X.t25 1172.87
R2314 X.n18 X.t46 996.134
R2315 X.n17 X.t31 996.134
R2316 X.n16 X.t38 996.134
R2317 X.n15 X.t53 996.134
R2318 X.n14 X.t40 996.134
R2319 X.n13 X.t34 996.134
R2320 X.n11 X.t43 996.134
R2321 X.n12 X.t28 996.134
R2322 X.n48 X.t52 690.867
R2323 X.n41 X.t29 690.867
R2324 X.n39 X.t49 530.201
R2325 X.n32 X.t54 530.201
R2326 X.n48 X.t37 514.134
R2327 X.n47 X.t44 514.134
R2328 X.n46 X.t26 514.134
R2329 X.n45 X.t41 514.134
R2330 X.n44 X.t35 514.134
R2331 X.n43 X.t48 514.134
R2332 X.n42 X.t32 514.134
R2333 X.n41 X.t47 514.134
R2334 X.n39 X.t33 353.467
R2335 X.n32 X.t42 353.467
R2336 X.n33 X.t27 353.467
R2337 X.n34 X.t45 353.467
R2338 X.n35 X.t30 353.467
R2339 X.n36 X.t36 353.467
R2340 X.n37 X.t51 353.467
R2341 X.n38 X.t39 353.467
R2342 X.n18 X.n17 176.733
R2343 X.n17 X.n16 176.733
R2344 X.n16 X.n15 176.733
R2345 X.n15 X.n14 176.733
R2346 X.n14 X.n13 176.733
R2347 X.n12 X.n11 176.733
R2348 X.n33 X.n32 176.733
R2349 X.n34 X.n33 176.733
R2350 X.n35 X.n34 176.733
R2351 X.n36 X.n35 176.733
R2352 X.n37 X.n36 176.733
R2353 X.n38 X.n37 176.733
R2354 X.n42 X.n41 176.733
R2355 X.n43 X.n42 176.733
R2356 X.n44 X.n43 176.733
R2357 X.n45 X.n44 176.733
R2358 X.n46 X.n45 176.733
R2359 X.n47 X.n46 176.733
R2360 X.n20 X.n19 166.436
R2361 X.n50 X.n40 161.843
R2362 X.n50 X.n49 161.718
R2363 X.n23 X.n21 160.427
R2364 X.n29 X.n28 159.802
R2365 X.n27 X.n26 159.802
R2366 X.n25 X.n24 159.802
R2367 X.n23 X.n22 159.802
R2368 X.n31 X.n30 155.302
R2369 X.n4 X.n2 114.689
R2370 X.n9 X.n1 114.689
R2371 X.n8 X.n7 114.126
R2372 X.n6 X.n5 114.126
R2373 X.n4 X.n3 114.126
R2374 X.n10 X.n0 109.626
R2375 X.n19 X.n18 51.9494
R2376 X.n19 X.n12 51.9494
R2377 X.n40 X.n39 51.9494
R2378 X.n40 X.n38 51.9494
R2379 X.n49 X.n48 51.9494
R2380 X.n49 X.n47 51.9494
R2381 X.n20 X.t9 49.4585
R2382 X.n51 X.n31 17.438
R2383 X.n7 X.t10 16.0005
R2384 X.n7 X.t5 16.0005
R2385 X.n5 X.t6 16.0005
R2386 X.n5 X.t1 16.0005
R2387 X.n3 X.t0 16.0005
R2388 X.n3 X.t8 16.0005
R2389 X.n2 X.t4 16.0005
R2390 X.n2 X.t24 16.0005
R2391 X.n1 X.t23 16.0005
R2392 X.n1 X.t7 16.0005
R2393 X.n0 X.t3 16.0005
R2394 X.n0 X.t2 16.0005
R2395 X.n51 X.n50 13.938
R2396 X.n30 X.t21 11.2576
R2397 X.n30 X.t13 11.2576
R2398 X.n28 X.t16 11.2576
R2399 X.n28 X.t19 11.2576
R2400 X.n26 X.t20 11.2576
R2401 X.n26 X.t11 11.2576
R2402 X.n24 X.t12 11.2576
R2403 X.n24 X.t14 11.2576
R2404 X.n22 X.t17 11.2576
R2405 X.n22 X.t15 11.2576
R2406 X.n21 X.t18 11.2576
R2407 X.n21 X.t22 11.2576
R2408 X.n53 X.n52 7.53175
R2409 X.n31 X.n29 5.1255
R2410 X.n10 X.n9 4.5005
R2411 X.n52 X.n51 4.5005
R2412 X.n52 X.n20 3.3755
R2413 X.n53 X.n10 1.71925
R2414 X.n25 X.n23 0.6255
R2415 X.n27 X.n25 0.6255
R2416 X.n29 X.n27 0.6255
R2417 X.n6 X.n4 0.563
R2418 X.n8 X.n6 0.563
R2419 X.n9 X.n8 0.563
R2420 X X.n53 0.063
R2421 VOUT-.n2 VOUT-.n0 145.989
R2422 VOUT-.n8 VOUT-.n7 145.989
R2423 VOUT-.n6 VOUT-.n5 145.427
R2424 VOUT-.n4 VOUT-.n3 145.427
R2425 VOUT-.n2 VOUT-.n1 145.427
R2426 VOUT-.n10 VOUT-.n9 140.927
R2427 VOUT-.n96 VOUT-.t6 113.192
R2428 VOUT-.n93 VOUT-.n91 95.7303
R2429 VOUT-.n95 VOUT-.n94 94.6053
R2430 VOUT-.n93 VOUT-.n92 94.6053
R2431 VOUT-.n90 VOUT-.n10 20.813
R2432 VOUT-.n90 VOUT-.n89 11.6871
R2433 VOUT-.n97 VOUT-.n96 7.46925
R2434 VOUT-.n9 VOUT-.t11 6.56717
R2435 VOUT-.n9 VOUT-.t13 6.56717
R2436 VOUT-.n7 VOUT-.t8 6.56717
R2437 VOUT-.n7 VOUT-.t4 6.56717
R2438 VOUT-.n5 VOUT-.t12 6.56717
R2439 VOUT-.n5 VOUT-.t7 6.56717
R2440 VOUT-.n3 VOUT-.t9 6.56717
R2441 VOUT-.n3 VOUT-.t14 6.56717
R2442 VOUT-.n1 VOUT-.t10 6.56717
R2443 VOUT-.n1 VOUT-.t15 6.56717
R2444 VOUT-.n0 VOUT-.t5 6.56717
R2445 VOUT-.n0 VOUT-.t16 6.56717
R2446 VOUT-.n37 VOUT-.t36 4.8295
R2447 VOUT-.n46 VOUT-.t74 4.8295
R2448 VOUT-.n44 VOUT-.t116 4.8295
R2449 VOUT-.n42 VOUT-.t147 4.8295
R2450 VOUT-.n40 VOUT-.t59 4.8295
R2451 VOUT-.n39 VOUT-.t139 4.8295
R2452 VOUT-.n59 VOUT-.t31 4.8295
R2453 VOUT-.n60 VOUT-.t94 4.8295
R2454 VOUT-.n62 VOUT-.t71 4.8295
R2455 VOUT-.n63 VOUT-.t128 4.8295
R2456 VOUT-.n65 VOUT-.t27 4.8295
R2457 VOUT-.n66 VOUT-.t88 4.8295
R2458 VOUT-.n68 VOUT-.t126 4.8295
R2459 VOUT-.n69 VOUT-.t51 4.8295
R2460 VOUT-.n71 VOUT-.t26 4.8295
R2461 VOUT-.n72 VOUT-.t82 4.8295
R2462 VOUT-.n74 VOUT-.t121 4.8295
R2463 VOUT-.n75 VOUT-.t44 4.8295
R2464 VOUT-.n77 VOUT-.t79 4.8295
R2465 VOUT-.n78 VOUT-.t148 4.8295
R2466 VOUT-.n80 VOUT-.t41 4.8295
R2467 VOUT-.n81 VOUT-.t112 4.8295
R2468 VOUT-.n83 VOUT-.t76 4.8295
R2469 VOUT-.n84 VOUT-.t141 4.8295
R2470 VOUT-.n11 VOUT-.t77 4.8295
R2471 VOUT-.n13 VOUT-.t49 4.8295
R2472 VOUT-.n25 VOUT-.t125 4.8295
R2473 VOUT-.n26 VOUT-.t118 4.8295
R2474 VOUT-.n28 VOUT-.t131 4.8295
R2475 VOUT-.n29 VOUT-.t57 4.8295
R2476 VOUT-.n31 VOUT-.t30 4.8295
R2477 VOUT-.n32 VOUT-.t91 4.8295
R2478 VOUT-.n34 VOUT-.t137 4.8295
R2479 VOUT-.n35 VOUT-.t64 4.8295
R2480 VOUT-.n86 VOUT-.t34 4.8295
R2481 VOUT-.n48 VOUT-.t68 4.8154
R2482 VOUT-.n49 VOUT-.t99 4.8154
R2483 VOUT-.n50 VOUT-.t132 4.8154
R2484 VOUT-.n51 VOUT-.t28 4.8154
R2485 VOUT-.n48 VOUT-.t101 4.806
R2486 VOUT-.n49 VOUT-.t138 4.806
R2487 VOUT-.n50 VOUT-.t33 4.806
R2488 VOUT-.n51 VOUT-.t73 4.806
R2489 VOUT-.n52 VOUT-.t53 4.806
R2490 VOUT-.n53 VOUT-.t87 4.806
R2491 VOUT-.n54 VOUT-.t127 4.806
R2492 VOUT-.n55 VOUT-.t111 4.806
R2493 VOUT-.n56 VOUT-.t145 4.806
R2494 VOUT-.n57 VOUT-.t122 4.806
R2495 VOUT-.n14 VOUT-.t115 4.806
R2496 VOUT-.n15 VOUT-.t146 4.806
R2497 VOUT-.n16 VOUT-.t38 4.806
R2498 VOUT-.n17 VOUT-.t75 4.806
R2499 VOUT-.n18 VOUT-.t123 4.806
R2500 VOUT-.n19 VOUT-.t24 4.806
R2501 VOUT-.n20 VOUT-.t58 4.806
R2502 VOUT-.n21 VOUT-.t114 4.806
R2503 VOUT-.n22 VOUT-.t144 4.806
R2504 VOUT-.n23 VOUT-.t97 4.806
R2505 VOUT-.n37 VOUT-.t140 4.5005
R2506 VOUT-.n38 VOUT-.t109 4.5005
R2507 VOUT-.n46 VOUT-.t119 4.5005
R2508 VOUT-.n47 VOUT-.t78 4.5005
R2509 VOUT-.n44 VOUT-.t155 4.5005
R2510 VOUT-.n45 VOUT-.t120 4.5005
R2511 VOUT-.n42 VOUT-.t43 4.5005
R2512 VOUT-.n43 VOUT-.t156 4.5005
R2513 VOUT-.n40 VOUT-.t93 4.5005
R2514 VOUT-.n41 VOUT-.t63 4.5005
R2515 VOUT-.n39 VOUT-.t102 4.5005
R2516 VOUT-.n58 VOUT-.t67 4.5005
R2517 VOUT-.n57 VOUT-.t81 4.5005
R2518 VOUT-.n56 VOUT-.t110 4.5005
R2519 VOUT-.n55 VOUT-.t69 4.5005
R2520 VOUT-.n54 VOUT-.t85 4.5005
R2521 VOUT-.n53 VOUT-.t48 4.5005
R2522 VOUT-.n52 VOUT-.t20 4.5005
R2523 VOUT-.n51 VOUT-.t32 4.5005
R2524 VOUT-.n50 VOUT-.t133 4.5005
R2525 VOUT-.n49 VOUT-.t98 4.5005
R2526 VOUT-.n48 VOUT-.t62 4.5005
R2527 VOUT-.n59 VOUT-.t136 4.5005
R2528 VOUT-.n61 VOUT-.t108 4.5005
R2529 VOUT-.n60 VOUT-.t52 4.5005
R2530 VOUT-.n62 VOUT-.t29 4.5005
R2531 VOUT-.n64 VOUT-.t134 4.5005
R2532 VOUT-.n63 VOUT-.t83 4.5005
R2533 VOUT-.n65 VOUT-.t130 4.5005
R2534 VOUT-.n67 VOUT-.t95 4.5005
R2535 VOUT-.n66 VOUT-.t45 4.5005
R2536 VOUT-.n68 VOUT-.t90 4.5005
R2537 VOUT-.n70 VOUT-.t60 4.5005
R2538 VOUT-.n69 VOUT-.t149 4.5005
R2539 VOUT-.n71 VOUT-.t124 4.5005
R2540 VOUT-.n73 VOUT-.t89 4.5005
R2541 VOUT-.n72 VOUT-.t39 4.5005
R2542 VOUT-.n74 VOUT-.t84 4.5005
R2543 VOUT-.n76 VOUT-.t54 4.5005
R2544 VOUT-.n75 VOUT-.t142 4.5005
R2545 VOUT-.n77 VOUT-.t47 4.5005
R2546 VOUT-.n79 VOUT-.t21 4.5005
R2547 VOUT-.n78 VOUT-.t104 4.5005
R2548 VOUT-.n80 VOUT-.t151 4.5005
R2549 VOUT-.n82 VOUT-.t117 4.5005
R2550 VOUT-.n81 VOUT-.t65 4.5005
R2551 VOUT-.n83 VOUT-.t40 4.5005
R2552 VOUT-.n85 VOUT-.t150 4.5005
R2553 VOUT-.n84 VOUT-.t92 4.5005
R2554 VOUT-.n11 VOUT-.t42 4.5005
R2555 VOUT-.n12 VOUT-.t153 4.5005
R2556 VOUT-.n13 VOUT-.t100 4.5005
R2557 VOUT-.n24 VOUT-.t152 4.5005
R2558 VOUT-.n23 VOUT-.t23 4.5005
R2559 VOUT-.n22 VOUT-.t25 4.5005
R2560 VOUT-.n21 VOUT-.t72 4.5005
R2561 VOUT-.n20 VOUT-.t80 4.5005
R2562 VOUT-.n19 VOUT-.t129 4.5005
R2563 VOUT-.n18 VOUT-.t37 4.5005
R2564 VOUT-.n17 VOUT-.t55 4.5005
R2565 VOUT-.n16 VOUT-.t105 4.5005
R2566 VOUT-.n15 VOUT-.t154 4.5005
R2567 VOUT-.n14 VOUT-.t61 4.5005
R2568 VOUT-.n25 VOUT-.t35 4.5005
R2569 VOUT-.n27 VOUT-.t86 4.5005
R2570 VOUT-.n26 VOUT-.t46 4.5005
R2571 VOUT-.n28 VOUT-.t96 4.5005
R2572 VOUT-.n30 VOUT-.t66 4.5005
R2573 VOUT-.n29 VOUT-.t19 4.5005
R2574 VOUT-.n31 VOUT-.t135 4.5005
R2575 VOUT-.n33 VOUT-.t107 4.5005
R2576 VOUT-.n32 VOUT-.t50 4.5005
R2577 VOUT-.n34 VOUT-.t106 4.5005
R2578 VOUT-.n36 VOUT-.t70 4.5005
R2579 VOUT-.n35 VOUT-.t22 4.5005
R2580 VOUT-.n86 VOUT-.t143 4.5005
R2581 VOUT-.n87 VOUT-.t113 4.5005
R2582 VOUT-.n88 VOUT-.t56 4.5005
R2583 VOUT-.n89 VOUT-.t103 4.5005
R2584 VOUT-.n10 VOUT-.n8 4.5005
R2585 VOUT-.n97 VOUT-.n90 3.84425
R2586 VOUT-.n94 VOUT-.t18 3.42907
R2587 VOUT-.n94 VOUT-.t2 3.42907
R2588 VOUT-.n92 VOUT-.t3 3.42907
R2589 VOUT-.n92 VOUT-.t0 3.42907
R2590 VOUT-.n91 VOUT-.t1 3.42907
R2591 VOUT-.n91 VOUT-.t17 3.42907
R2592 VOUT-.n96 VOUT-.n95 2.03175
R2593 VOUT-.n95 VOUT-.n93 1.1255
R2594 VOUT-.n4 VOUT-.n2 0.563
R2595 VOUT-.n6 VOUT-.n4 0.563
R2596 VOUT-.n8 VOUT-.n6 0.563
R2597 VOUT-.n38 VOUT-.n37 0.3295
R2598 VOUT-.n47 VOUT-.n46 0.3295
R2599 VOUT-.n45 VOUT-.n44 0.3295
R2600 VOUT-.n43 VOUT-.n42 0.3295
R2601 VOUT-.n41 VOUT-.n40 0.3295
R2602 VOUT-.n58 VOUT-.n39 0.3295
R2603 VOUT-.n58 VOUT-.n57 0.3295
R2604 VOUT-.n57 VOUT-.n56 0.3295
R2605 VOUT-.n56 VOUT-.n55 0.3295
R2606 VOUT-.n55 VOUT-.n54 0.3295
R2607 VOUT-.n54 VOUT-.n53 0.3295
R2608 VOUT-.n53 VOUT-.n52 0.3295
R2609 VOUT-.n52 VOUT-.n51 0.3295
R2610 VOUT-.n51 VOUT-.n50 0.3295
R2611 VOUT-.n50 VOUT-.n49 0.3295
R2612 VOUT-.n49 VOUT-.n48 0.3295
R2613 VOUT-.n61 VOUT-.n59 0.3295
R2614 VOUT-.n61 VOUT-.n60 0.3295
R2615 VOUT-.n64 VOUT-.n62 0.3295
R2616 VOUT-.n64 VOUT-.n63 0.3295
R2617 VOUT-.n67 VOUT-.n65 0.3295
R2618 VOUT-.n67 VOUT-.n66 0.3295
R2619 VOUT-.n70 VOUT-.n68 0.3295
R2620 VOUT-.n70 VOUT-.n69 0.3295
R2621 VOUT-.n73 VOUT-.n71 0.3295
R2622 VOUT-.n73 VOUT-.n72 0.3295
R2623 VOUT-.n76 VOUT-.n74 0.3295
R2624 VOUT-.n76 VOUT-.n75 0.3295
R2625 VOUT-.n79 VOUT-.n77 0.3295
R2626 VOUT-.n79 VOUT-.n78 0.3295
R2627 VOUT-.n82 VOUT-.n80 0.3295
R2628 VOUT-.n82 VOUT-.n81 0.3295
R2629 VOUT-.n85 VOUT-.n83 0.3295
R2630 VOUT-.n85 VOUT-.n84 0.3295
R2631 VOUT-.n12 VOUT-.n11 0.3295
R2632 VOUT-.n24 VOUT-.n13 0.3295
R2633 VOUT-.n24 VOUT-.n23 0.3295
R2634 VOUT-.n23 VOUT-.n22 0.3295
R2635 VOUT-.n22 VOUT-.n21 0.3295
R2636 VOUT-.n21 VOUT-.n20 0.3295
R2637 VOUT-.n20 VOUT-.n19 0.3295
R2638 VOUT-.n19 VOUT-.n18 0.3295
R2639 VOUT-.n18 VOUT-.n17 0.3295
R2640 VOUT-.n17 VOUT-.n16 0.3295
R2641 VOUT-.n16 VOUT-.n15 0.3295
R2642 VOUT-.n15 VOUT-.n14 0.3295
R2643 VOUT-.n27 VOUT-.n25 0.3295
R2644 VOUT-.n27 VOUT-.n26 0.3295
R2645 VOUT-.n30 VOUT-.n28 0.3295
R2646 VOUT-.n30 VOUT-.n29 0.3295
R2647 VOUT-.n33 VOUT-.n31 0.3295
R2648 VOUT-.n33 VOUT-.n32 0.3295
R2649 VOUT-.n36 VOUT-.n34 0.3295
R2650 VOUT-.n36 VOUT-.n35 0.3295
R2651 VOUT-.n87 VOUT-.n86 0.3295
R2652 VOUT-.n88 VOUT-.n87 0.3295
R2653 VOUT-.n89 VOUT-.n88 0.3295
R2654 VOUT-.n52 VOUT-.n47 0.306
R2655 VOUT-.n53 VOUT-.n45 0.306
R2656 VOUT-.n54 VOUT-.n43 0.306
R2657 VOUT-.n55 VOUT-.n41 0.306
R2658 VOUT-.n58 VOUT-.n38 0.2825
R2659 VOUT-.n61 VOUT-.n58 0.2825
R2660 VOUT-.n64 VOUT-.n61 0.2825
R2661 VOUT-.n67 VOUT-.n64 0.2825
R2662 VOUT-.n70 VOUT-.n67 0.2825
R2663 VOUT-.n73 VOUT-.n70 0.2825
R2664 VOUT-.n76 VOUT-.n73 0.2825
R2665 VOUT-.n79 VOUT-.n76 0.2825
R2666 VOUT-.n82 VOUT-.n79 0.2825
R2667 VOUT-.n85 VOUT-.n82 0.2825
R2668 VOUT-.n24 VOUT-.n12 0.2825
R2669 VOUT-.n27 VOUT-.n24 0.2825
R2670 VOUT-.n30 VOUT-.n27 0.2825
R2671 VOUT-.n33 VOUT-.n30 0.2825
R2672 VOUT-.n36 VOUT-.n33 0.2825
R2673 VOUT-.n87 VOUT-.n36 0.2825
R2674 VOUT-.n87 VOUT-.n85 0.2825
R2675 VOUT- VOUT-.n97 0.063
R2676 cap_res_X.t0 cap_res_X.t10 50.1603
R2677 cap_res_X.t95 cap_res_X.t89 0.1603
R2678 cap_res_X.t59 cap_res_X.t58 0.1603
R2679 cap_res_X.t24 cap_res_X.t25 0.1603
R2680 cap_res_X.t125 cap_res_X.t129 0.1603
R2681 cap_res_X.t38 cap_res_X.t83 0.1603
R2682 cap_res_X.t79 cap_res_X.t38 0.1603
R2683 cap_res_X.t137 cap_res_X.t79 0.1603
R2684 cap_res_X.t2 cap_res_X.t41 0.1603
R2685 cap_res_X.t37 cap_res_X.t2 0.1603
R2686 cap_res_X.t109 cap_res_X.t37 0.1603
R2687 cap_res_X.t55 cap_res_X.t18 0.1603
R2688 cap_res_X.t17 cap_res_X.t121 0.1603
R2689 cap_res_X.t105 cap_res_X.t63 0.1603
R2690 cap_res_X.t21 cap_res_X.t126 0.1603
R2691 cap_res_X.t74 cap_res_X.t29 0.1603
R2692 cap_res_X.t128 cap_res_X.t86 0.1603
R2693 cap_res_X.t112 cap_res_X.t69 0.1603
R2694 cap_res_X.t27 cap_res_X.t130 0.1603
R2695 cap_res_X.t8 cap_res_X.t106 0.1603
R2696 cap_res_X.t67 cap_res_X.t31 0.1603
R2697 cap_res_X.t118 cap_res_X.t75 0.1603
R2698 cap_res_X.t33 cap_res_X.t131 0.1603
R2699 cap_res_X.t15 cap_res_X.t113 0.1603
R2700 cap_res_X.t73 cap_res_X.t36 0.1603
R2701 cap_res_X.t53 cap_res_X.t9 0.1603
R2702 cap_res_X.t110 cap_res_X.t78 0.1603
R2703 cap_res_X.t92 cap_res_X.t45 0.1603
R2704 cap_res_X.t6 cap_res_X.t116 0.1603
R2705 cap_res_X.t65 cap_res_X.t16 0.1603
R2706 cap_res_X.t117 cap_res_X.t81 0.1603
R2707 cap_res_X.t101 cap_res_X.t54 0.1603
R2708 cap_res_X.t14 cap_res_X.t123 0.1603
R2709 cap_res_X.t135 cap_res_X.t93 0.1603
R2710 cap_res_X.t51 cap_res_X.t20 0.1603
R2711 cap_res_X.t107 cap_res_X.t66 0.1603
R2712 cap_res_X.t22 cap_res_X.t127 0.1603
R2713 cap_res_X.t138 cap_res_X.t100 0.1603
R2714 cap_res_X.t61 cap_res_X.t26 0.1603
R2715 cap_res_X.t111 cap_res_X.t39 0.1603
R2716 cap_res_X.t122 cap_res_X.t32 0.1603
R2717 cap_res_X.t96 cap_res_X.t42 0.1603
R2718 cap_res_X.t3 cap_res_X.t11 0.1603
R2719 cap_res_X.t52 cap_res_X.t119 0.1603
R2720 cap_res_X.t102 cap_res_X.t82 0.1603
R2721 cap_res_X.t120 cap_res_X.t34 0.1603
R2722 cap_res_X.t28 cap_res_X.t133 0.1603
R2723 cap_res_X.t77 cap_res_X.t99 0.1603
R2724 cap_res_X.t85 cap_res_X.t43 0.1603
R2725 cap_res_X.t132 cap_res_X.t13 0.1603
R2726 cap_res_X.t134 cap_res_X.t60 0.1603
R2727 cap_res_X.t57 cap_res_X.t108 0.1603
R2728 cap_res_X.t115 cap_res_X.t80 0.1603
R2729 cap_res_X.t64 cap_res_X.t98 0.1603
R2730 cap_res_X.t94 cap_res_X.t64 0.1603
R2731 cap_res_X.t88 cap_res_X.t94 0.1603
R2732 cap_res_X.t1 cap_res_X.t72 0.1603
R2733 cap_res_X.t114 cap_res_X.t1 0.1603
R2734 cap_res_X.t10 cap_res_X.t114 0.1603
R2735 cap_res_X.n29 cap_res_X.t56 0.159278
R2736 cap_res_X.n30 cap_res_X.t19 0.159278
R2737 cap_res_X.n31 cap_res_X.t124 0.159278
R2738 cap_res_X.n32 cap_res_X.t84 0.159278
R2739 cap_res_X.n33 cap_res_X.t104 0.159278
R2740 cap_res_X.n34 cap_res_X.t70 0.159278
R2741 cap_res_X.n25 cap_res_X.t48 0.159278
R2742 cap_res_X.t5 cap_res_X.n9 0.159278
R2743 cap_res_X.t71 cap_res_X.n10 0.159278
R2744 cap_res_X.t91 cap_res_X.n11 0.159278
R2745 cap_res_X.t50 cap_res_X.n12 0.159278
R2746 cap_res_X.t87 cap_res_X.n13 0.159278
R2747 cap_res_X.t44 cap_res_X.n14 0.159278
R2748 cap_res_X.t7 cap_res_X.n15 0.159278
R2749 cap_res_X.t40 cap_res_X.n16 0.159278
R2750 cap_res_X.t136 cap_res_X.n17 0.159278
R2751 cap_res_X.t103 cap_res_X.n18 0.159278
R2752 cap_res_X.t68 cap_res_X.n19 0.159278
R2753 cap_res_X.t97 cap_res_X.n20 0.159278
R2754 cap_res_X.t62 cap_res_X.n21 0.159278
R2755 cap_res_X.t23 cap_res_X.n22 0.159278
R2756 cap_res_X.t49 cap_res_X.n23 0.159278
R2757 cap_res_X.t90 cap_res_X.n24 0.159278
R2758 cap_res_X.n26 cap_res_X.t35 0.159278
R2759 cap_res_X.n27 cap_res_X.t12 0.159278
R2760 cap_res_X.n28 cap_res_X.t46 0.159278
R2761 cap_res_X.n35 cap_res_X.t30 0.159278
R2762 cap_res_X.t48 cap_res_X.t17 0.137822
R2763 cap_res_X.n25 cap_res_X.t55 0.1368
R2764 cap_res_X.n24 cap_res_X.t105 0.1368
R2765 cap_res_X.n24 cap_res_X.t21 0.1368
R2766 cap_res_X.n23 cap_res_X.t74 0.1368
R2767 cap_res_X.n23 cap_res_X.t128 0.1368
R2768 cap_res_X.n22 cap_res_X.t112 0.1368
R2769 cap_res_X.n22 cap_res_X.t27 0.1368
R2770 cap_res_X.n21 cap_res_X.t8 0.1368
R2771 cap_res_X.n21 cap_res_X.t67 0.1368
R2772 cap_res_X.n20 cap_res_X.t118 0.1368
R2773 cap_res_X.n20 cap_res_X.t33 0.1368
R2774 cap_res_X.n19 cap_res_X.t15 0.1368
R2775 cap_res_X.n19 cap_res_X.t73 0.1368
R2776 cap_res_X.n18 cap_res_X.t53 0.1368
R2777 cap_res_X.n18 cap_res_X.t110 0.1368
R2778 cap_res_X.n17 cap_res_X.t92 0.1368
R2779 cap_res_X.n17 cap_res_X.t6 0.1368
R2780 cap_res_X.n16 cap_res_X.t65 0.1368
R2781 cap_res_X.n16 cap_res_X.t117 0.1368
R2782 cap_res_X.n15 cap_res_X.t101 0.1368
R2783 cap_res_X.n15 cap_res_X.t14 0.1368
R2784 cap_res_X.n14 cap_res_X.t135 0.1368
R2785 cap_res_X.n14 cap_res_X.t51 0.1368
R2786 cap_res_X.n13 cap_res_X.t107 0.1368
R2787 cap_res_X.n13 cap_res_X.t22 0.1368
R2788 cap_res_X.n12 cap_res_X.t138 0.1368
R2789 cap_res_X.n12 cap_res_X.t61 0.1368
R2790 cap_res_X.n11 cap_res_X.t111 0.1368
R2791 cap_res_X.n11 cap_res_X.t122 0.1368
R2792 cap_res_X.n10 cap_res_X.t57 0.1368
R2793 cap_res_X.n9 cap_res_X.t115 0.1368
R2794 cap_res_X.n0 cap_res_X.t96 0.114322
R2795 cap_res_X.n30 cap_res_X.n29 0.1133
R2796 cap_res_X.n31 cap_res_X.n30 0.1133
R2797 cap_res_X.n32 cap_res_X.n31 0.1133
R2798 cap_res_X.n33 cap_res_X.n32 0.1133
R2799 cap_res_X.n34 cap_res_X.n33 0.1133
R2800 cap_res_X.n1 cap_res_X.n0 0.1133
R2801 cap_res_X.n2 cap_res_X.n1 0.1133
R2802 cap_res_X.n3 cap_res_X.n2 0.1133
R2803 cap_res_X.n4 cap_res_X.n3 0.1133
R2804 cap_res_X.n5 cap_res_X.n4 0.1133
R2805 cap_res_X.n6 cap_res_X.n5 0.1133
R2806 cap_res_X.n7 cap_res_X.n6 0.1133
R2807 cap_res_X.n8 cap_res_X.n7 0.1133
R2808 cap_res_X.n10 cap_res_X.n8 0.1133
R2809 cap_res_X.n26 cap_res_X.n25 0.1133
R2810 cap_res_X.n27 cap_res_X.n26 0.1133
R2811 cap_res_X.n28 cap_res_X.n27 0.1133
R2812 cap_res_X.n35 cap_res_X.n28 0.1133
R2813 cap_res_X.n35 cap_res_X.n34 0.1133
R2814 cap_res_X.n29 cap_res_X.t95 0.00152174
R2815 cap_res_X.n30 cap_res_X.t59 0.00152174
R2816 cap_res_X.n31 cap_res_X.t24 0.00152174
R2817 cap_res_X.n32 cap_res_X.t125 0.00152174
R2818 cap_res_X.n33 cap_res_X.t137 0.00152174
R2819 cap_res_X.n34 cap_res_X.t109 0.00152174
R2820 cap_res_X.n0 cap_res_X.t3 0.00152174
R2821 cap_res_X.n1 cap_res_X.t52 0.00152174
R2822 cap_res_X.n2 cap_res_X.t102 0.00152174
R2823 cap_res_X.n3 cap_res_X.t120 0.00152174
R2824 cap_res_X.n4 cap_res_X.t28 0.00152174
R2825 cap_res_X.n5 cap_res_X.t77 0.00152174
R2826 cap_res_X.n6 cap_res_X.t85 0.00152174
R2827 cap_res_X.n7 cap_res_X.t132 0.00152174
R2828 cap_res_X.n8 cap_res_X.t134 0.00152174
R2829 cap_res_X.n9 cap_res_X.t4 0.00152174
R2830 cap_res_X.n10 cap_res_X.t5 0.00152174
R2831 cap_res_X.n11 cap_res_X.t71 0.00152174
R2832 cap_res_X.n12 cap_res_X.t91 0.00152174
R2833 cap_res_X.n13 cap_res_X.t50 0.00152174
R2834 cap_res_X.n14 cap_res_X.t87 0.00152174
R2835 cap_res_X.n15 cap_res_X.t44 0.00152174
R2836 cap_res_X.n16 cap_res_X.t7 0.00152174
R2837 cap_res_X.n17 cap_res_X.t40 0.00152174
R2838 cap_res_X.n18 cap_res_X.t136 0.00152174
R2839 cap_res_X.n19 cap_res_X.t103 0.00152174
R2840 cap_res_X.n20 cap_res_X.t68 0.00152174
R2841 cap_res_X.n21 cap_res_X.t97 0.00152174
R2842 cap_res_X.n22 cap_res_X.t62 0.00152174
R2843 cap_res_X.n23 cap_res_X.t23 0.00152174
R2844 cap_res_X.n24 cap_res_X.t49 0.00152174
R2845 cap_res_X.n25 cap_res_X.t90 0.00152174
R2846 cap_res_X.n26 cap_res_X.t76 0.00152174
R2847 cap_res_X.n27 cap_res_X.t47 0.00152174
R2848 cap_res_X.n28 cap_res_X.t88 0.00152174
R2849 cap_res_X.t72 cap_res_X.n35 0.00152174
R2850 VOUT+.n8 VOUT+.n0 145.989
R2851 VOUT+.n3 VOUT+.n1 145.989
R2852 VOUT+.n7 VOUT+.n6 145.427
R2853 VOUT+.n5 VOUT+.n4 145.427
R2854 VOUT+.n3 VOUT+.n2 145.427
R2855 VOUT+.n10 VOUT+.n9 140.927
R2856 VOUT+.n96 VOUT+.t1 113.192
R2857 VOUT+.n93 VOUT+.n91 95.7303
R2858 VOUT+.n95 VOUT+.n94 94.6053
R2859 VOUT+.n93 VOUT+.n92 94.6053
R2860 VOUT+.n90 VOUT+.n10 20.813
R2861 VOUT+.n90 VOUT+.n89 11.6871
R2862 VOUT+.n97 VOUT+.n96 7.34425
R2863 VOUT+.n9 VOUT+.t13 6.56717
R2864 VOUT+.n9 VOUT+.t8 6.56717
R2865 VOUT+.n6 VOUT+.t12 6.56717
R2866 VOUT+.n6 VOUT+.t7 6.56717
R2867 VOUT+.n4 VOUT+.t11 6.56717
R2868 VOUT+.n4 VOUT+.t6 6.56717
R2869 VOUT+.n2 VOUT+.t10 6.56717
R2870 VOUT+.n2 VOUT+.t5 6.56717
R2871 VOUT+.n1 VOUT+.t9 6.56717
R2872 VOUT+.n1 VOUT+.t14 6.56717
R2873 VOUT+.n0 VOUT+.t3 6.56717
R2874 VOUT+.n0 VOUT+.t4 6.56717
R2875 VOUT+.n37 VOUT+.t56 4.8295
R2876 VOUT+.n39 VOUT+.t107 4.8295
R2877 VOUT+.n41 VOUT+.t137 4.8295
R2878 VOUT+.n43 VOUT+.t50 4.8295
R2879 VOUT+.n45 VOUT+.t144 4.8295
R2880 VOUT+.n57 VOUT+.t151 4.8295
R2881 VOUT+.n59 VOUT+.t73 4.8295
R2882 VOUT+.n60 VOUT+.t60 4.8295
R2883 VOUT+.n62 VOUT+.t110 4.8295
R2884 VOUT+.n63 VOUT+.t92 4.8295
R2885 VOUT+.n65 VOUT+.t67 4.8295
R2886 VOUT+.n66 VOUT+.t51 4.8295
R2887 VOUT+.n68 VOUT+.t23 4.8295
R2888 VOUT+.n69 VOUT+.t149 4.8295
R2889 VOUT+.n71 VOUT+.t65 4.8295
R2890 VOUT+.n72 VOUT+.t46 4.8295
R2891 VOUT+.n74 VOUT+.t19 4.8295
R2892 VOUT+.n75 VOUT+.t147 4.8295
R2893 VOUT+.n77 VOUT+.t120 4.8295
R2894 VOUT+.n78 VOUT+.t109 4.8295
R2895 VOUT+.n80 VOUT+.t82 4.8295
R2896 VOUT+.n81 VOUT+.t66 4.8295
R2897 VOUT+.n83 VOUT+.t115 4.8295
R2898 VOUT+.n84 VOUT+.t103 4.8295
R2899 VOUT+.n11 VOUT+.t106 4.8295
R2900 VOUT+.n23 VOUT+.t90 4.8295
R2901 VOUT+.n25 VOUT+.t117 4.8295
R2902 VOUT+.n26 VOUT+.t88 4.8295
R2903 VOUT+.n28 VOUT+.t27 4.8295
R2904 VOUT+.n29 VOUT+.t152 4.8295
R2905 VOUT+.n31 VOUT+.t72 4.8295
R2906 VOUT+.n32 VOUT+.t59 4.8295
R2907 VOUT+.n34 VOUT+.t33 4.8295
R2908 VOUT+.n35 VOUT+.t155 4.8295
R2909 VOUT+.n86 VOUT+.t64 4.8295
R2910 VOUT+.n50 VOUT+.t44 4.8154
R2911 VOUT+.n49 VOUT+.t98 4.8154
R2912 VOUT+.n48 VOUT+.t126 4.8154
R2913 VOUT+.n47 VOUT+.t21 4.8154
R2914 VOUT+.n56 VOUT+.t112 4.806
R2915 VOUT+.n55 VOUT+.t146 4.806
R2916 VOUT+.n54 VOUT+.t45 4.806
R2917 VOUT+.n53 VOUT+.t79 4.806
R2918 VOUT+.n52 VOUT+.t63 4.806
R2919 VOUT+.n51 VOUT+.t38 4.806
R2920 VOUT+.n50 VOUT+.t76 4.806
R2921 VOUT+.n49 VOUT+.t62 4.806
R2922 VOUT+.n48 VOUT+.t99 4.806
R2923 VOUT+.n47 VOUT+.t131 4.806
R2924 VOUT+.n22 VOUT+.t83 4.806
R2925 VOUT+.n21 VOUT+.t116 4.806
R2926 VOUT+.n20 VOUT+.t150 4.806
R2927 VOUT+.n19 VOUT+.t49 4.806
R2928 VOUT+.n18 VOUT+.t101 4.806
R2929 VOUT+.n17 VOUT+.t57 4.806
R2930 VOUT+.n16 VOUT+.t89 4.806
R2931 VOUT+.n15 VOUT+.t138 4.806
R2932 VOUT+.n14 VOUT+.t29 4.806
R2933 VOUT+.n13 VOUT+.t69 4.806
R2934 VOUT+.n38 VOUT+.t127 4.5005
R2935 VOUT+.n37 VOUT+.t96 4.5005
R2936 VOUT+.n39 VOUT+.t141 4.5005
R2937 VOUT+.n40 VOUT+.t111 4.5005
R2938 VOUT+.n41 VOUT+.t34 4.5005
R2939 VOUT+.n42 VOUT+.t143 4.5005
R2940 VOUT+.n43 VOUT+.t87 4.5005
R2941 VOUT+.n44 VOUT+.t55 4.5005
R2942 VOUT+.n45 VOUT+.t43 4.5005
R2943 VOUT+.n46 VOUT+.t148 4.5005
R2944 VOUT+.n47 VOUT+.t97 4.5005
R2945 VOUT+.n48 VOUT+.t58 4.5005
R2946 VOUT+.n49 VOUT+.t153 4.5005
R2947 VOUT+.n50 VOUT+.t36 4.5005
R2948 VOUT+.n51 VOUT+.t139 4.5005
R2949 VOUT+.n52 VOUT+.t154 4.5005
R2950 VOUT+.n53 VOUT+.t41 4.5005
R2951 VOUT+.n54 VOUT+.t145 4.5005
R2952 VOUT+.n55 VOUT+.t108 4.5005
R2953 VOUT+.n56 VOUT+.t68 4.5005
R2954 VOUT+.n58 VOUT+.t91 4.5005
R2955 VOUT+.n57 VOUT+.t53 4.5005
R2956 VOUT+.n59 VOUT+.t32 4.5005
R2957 VOUT+.n61 VOUT+.t123 4.5005
R2958 VOUT+.n60 VOUT+.t94 4.5005
R2959 VOUT+.n62 VOUT+.t71 4.5005
R2960 VOUT+.n64 VOUT+.t156 4.5005
R2961 VOUT+.n63 VOUT+.t122 4.5005
R2962 VOUT+.n65 VOUT+.t26 4.5005
R2963 VOUT+.n67 VOUT+.t119 4.5005
R2964 VOUT+.n66 VOUT+.t85 4.5005
R2965 VOUT+.n68 VOUT+.t130 4.5005
R2966 VOUT+.n70 VOUT+.t78 4.5005
R2967 VOUT+.n69 VOUT+.t47 4.5005
R2968 VOUT+.n71 VOUT+.t22 4.5005
R2969 VOUT+.n73 VOUT+.t114 4.5005
R2970 VOUT+.n72 VOUT+.t77 4.5005
R2971 VOUT+.n74 VOUT+.t124 4.5005
R2972 VOUT+.n76 VOUT+.t74 4.5005
R2973 VOUT+.n75 VOUT+.t39 4.5005
R2974 VOUT+.n77 VOUT+.t86 4.5005
R2975 VOUT+.n79 VOUT+.t30 4.5005
R2976 VOUT+.n78 VOUT+.t140 4.5005
R2977 VOUT+.n80 VOUT+.t48 4.5005
R2978 VOUT+.n82 VOUT+.t134 4.5005
R2979 VOUT+.n81 VOUT+.t104 4.5005
R2980 VOUT+.n83 VOUT+.t80 4.5005
R2981 VOUT+.n85 VOUT+.t25 4.5005
R2982 VOUT+.n84 VOUT+.t133 4.5005
R2983 VOUT+.n12 VOUT+.t28 4.5005
R2984 VOUT+.n11 VOUT+.t136 4.5005
R2985 VOUT+.n13 VOUT+.t81 4.5005
R2986 VOUT+.n14 VOUT+.t128 4.5005
R2987 VOUT+.n15 VOUT+.t37 4.5005
R2988 VOUT+.n16 VOUT+.t54 4.5005
R2989 VOUT+.n17 VOUT+.t102 4.5005
R2990 VOUT+.n18 VOUT+.t105 4.5005
R2991 VOUT+.n19 VOUT+.t113 4.5005
R2992 VOUT+.n20 VOUT+.t20 4.5005
R2993 VOUT+.n21 VOUT+.t70 4.5005
R2994 VOUT+.n22 VOUT+.t118 4.5005
R2995 VOUT+.n24 VOUT+.t132 4.5005
R2996 VOUT+.n23 VOUT+.t40 4.5005
R2997 VOUT+.n25 VOUT+.t24 4.5005
R2998 VOUT+.n27 VOUT+.t125 4.5005
R2999 VOUT+.n26 VOUT+.t35 4.5005
R3000 VOUT+.n28 VOUT+.t135 4.5005
R3001 VOUT+.n30 VOUT+.t84 4.5005
R3002 VOUT+.n29 VOUT+.t52 4.5005
R3003 VOUT+.n31 VOUT+.t31 4.5005
R3004 VOUT+.n33 VOUT+.t121 4.5005
R3005 VOUT+.n32 VOUT+.t93 4.5005
R3006 VOUT+.n34 VOUT+.t142 4.5005
R3007 VOUT+.n36 VOUT+.t95 4.5005
R3008 VOUT+.n35 VOUT+.t61 4.5005
R3009 VOUT+.n89 VOUT+.t75 4.5005
R3010 VOUT+.n88 VOUT+.t42 4.5005
R3011 VOUT+.n87 VOUT+.t129 4.5005
R3012 VOUT+.n86 VOUT+.t100 4.5005
R3013 VOUT+.n10 VOUT+.n8 4.5005
R3014 VOUT+.n97 VOUT+.n90 3.84425
R3015 VOUT+.n94 VOUT+.t17 3.42907
R3016 VOUT+.n94 VOUT+.t15 3.42907
R3017 VOUT+.n92 VOUT+.t2 3.42907
R3018 VOUT+.n92 VOUT+.t0 3.42907
R3019 VOUT+.n91 VOUT+.t16 3.42907
R3020 VOUT+.n91 VOUT+.t18 3.42907
R3021 VOUT+.n96 VOUT+.n95 2.15675
R3022 VOUT+.n95 VOUT+.n93 1.1255
R3023 VOUT+.n5 VOUT+.n3 0.563
R3024 VOUT+.n7 VOUT+.n5 0.563
R3025 VOUT+.n8 VOUT+.n7 0.563
R3026 VOUT+.n38 VOUT+.n37 0.3295
R3027 VOUT+.n40 VOUT+.n39 0.3295
R3028 VOUT+.n42 VOUT+.n41 0.3295
R3029 VOUT+.n44 VOUT+.n43 0.3295
R3030 VOUT+.n46 VOUT+.n45 0.3295
R3031 VOUT+.n48 VOUT+.n47 0.3295
R3032 VOUT+.n49 VOUT+.n48 0.3295
R3033 VOUT+.n50 VOUT+.n49 0.3295
R3034 VOUT+.n51 VOUT+.n50 0.3295
R3035 VOUT+.n52 VOUT+.n51 0.3295
R3036 VOUT+.n53 VOUT+.n52 0.3295
R3037 VOUT+.n54 VOUT+.n53 0.3295
R3038 VOUT+.n55 VOUT+.n54 0.3295
R3039 VOUT+.n56 VOUT+.n55 0.3295
R3040 VOUT+.n58 VOUT+.n56 0.3295
R3041 VOUT+.n58 VOUT+.n57 0.3295
R3042 VOUT+.n61 VOUT+.n59 0.3295
R3043 VOUT+.n61 VOUT+.n60 0.3295
R3044 VOUT+.n64 VOUT+.n62 0.3295
R3045 VOUT+.n64 VOUT+.n63 0.3295
R3046 VOUT+.n67 VOUT+.n65 0.3295
R3047 VOUT+.n67 VOUT+.n66 0.3295
R3048 VOUT+.n70 VOUT+.n68 0.3295
R3049 VOUT+.n70 VOUT+.n69 0.3295
R3050 VOUT+.n73 VOUT+.n71 0.3295
R3051 VOUT+.n73 VOUT+.n72 0.3295
R3052 VOUT+.n76 VOUT+.n74 0.3295
R3053 VOUT+.n76 VOUT+.n75 0.3295
R3054 VOUT+.n79 VOUT+.n77 0.3295
R3055 VOUT+.n79 VOUT+.n78 0.3295
R3056 VOUT+.n82 VOUT+.n80 0.3295
R3057 VOUT+.n82 VOUT+.n81 0.3295
R3058 VOUT+.n85 VOUT+.n83 0.3295
R3059 VOUT+.n85 VOUT+.n84 0.3295
R3060 VOUT+.n12 VOUT+.n11 0.3295
R3061 VOUT+.n14 VOUT+.n13 0.3295
R3062 VOUT+.n15 VOUT+.n14 0.3295
R3063 VOUT+.n16 VOUT+.n15 0.3295
R3064 VOUT+.n17 VOUT+.n16 0.3295
R3065 VOUT+.n18 VOUT+.n17 0.3295
R3066 VOUT+.n19 VOUT+.n18 0.3295
R3067 VOUT+.n20 VOUT+.n19 0.3295
R3068 VOUT+.n21 VOUT+.n20 0.3295
R3069 VOUT+.n22 VOUT+.n21 0.3295
R3070 VOUT+.n24 VOUT+.n22 0.3295
R3071 VOUT+.n24 VOUT+.n23 0.3295
R3072 VOUT+.n27 VOUT+.n25 0.3295
R3073 VOUT+.n27 VOUT+.n26 0.3295
R3074 VOUT+.n30 VOUT+.n28 0.3295
R3075 VOUT+.n30 VOUT+.n29 0.3295
R3076 VOUT+.n33 VOUT+.n31 0.3295
R3077 VOUT+.n33 VOUT+.n32 0.3295
R3078 VOUT+.n36 VOUT+.n34 0.3295
R3079 VOUT+.n36 VOUT+.n35 0.3295
R3080 VOUT+.n89 VOUT+.n88 0.3295
R3081 VOUT+.n88 VOUT+.n87 0.3295
R3082 VOUT+.n87 VOUT+.n86 0.3295
R3083 VOUT+.n54 VOUT+.n40 0.306
R3084 VOUT+.n53 VOUT+.n42 0.306
R3085 VOUT+.n52 VOUT+.n44 0.306
R3086 VOUT+.n51 VOUT+.n46 0.306
R3087 VOUT+.n58 VOUT+.n38 0.2825
R3088 VOUT+.n61 VOUT+.n58 0.2825
R3089 VOUT+.n64 VOUT+.n61 0.2825
R3090 VOUT+.n67 VOUT+.n64 0.2825
R3091 VOUT+.n70 VOUT+.n67 0.2825
R3092 VOUT+.n73 VOUT+.n70 0.2825
R3093 VOUT+.n76 VOUT+.n73 0.2825
R3094 VOUT+.n79 VOUT+.n76 0.2825
R3095 VOUT+.n82 VOUT+.n79 0.2825
R3096 VOUT+.n85 VOUT+.n82 0.2825
R3097 VOUT+.n24 VOUT+.n12 0.2825
R3098 VOUT+.n27 VOUT+.n24 0.2825
R3099 VOUT+.n30 VOUT+.n27 0.2825
R3100 VOUT+.n33 VOUT+.n30 0.2825
R3101 VOUT+.n36 VOUT+.n33 0.2825
R3102 VOUT+.n87 VOUT+.n36 0.2825
R3103 VOUT+.n87 VOUT+.n85 0.2825
R3104 VOUT+ VOUT+.n97 0.063
R3105 cap_res_Y cap_res_Y.t0 49.2388
R3106 cap_res_Y cap_res_Y.t20 0.922875
R3107 cap_res_Y.t104 cap_res_Y.t6 0.1603
R3108 cap_res_Y.t61 cap_res_Y.t101 0.1603
R3109 cap_res_Y.t63 cap_res_Y.t97 0.1603
R3110 cap_res_Y.t125 cap_res_Y.t84 0.1603
R3111 cap_res_Y.t35 cap_res_Y.t65 0.1603
R3112 cap_res_Y.t86 cap_res_Y.t47 0.1603
R3113 cap_res_Y.t72 cap_res_Y.t106 0.1603
R3114 cap_res_Y.t131 cap_res_Y.t90 0.1603
R3115 cap_res_Y.t110 cap_res_Y.t8 0.1603
R3116 cap_res_Y.t27 cap_res_Y.t134 0.1603
R3117 cap_res_Y.t80 cap_res_Y.t111 0.1603
R3118 cap_res_Y.t135 cap_res_Y.t92 0.1603
R3119 cap_res_Y.t118 cap_res_Y.t10 0.1603
R3120 cap_res_Y.t33 cap_res_Y.t138 0.1603
R3121 cap_res_Y.t17 cap_res_Y.t48 0.1603
R3122 cap_res_Y.t71 cap_res_Y.t37 0.1603
R3123 cap_res_Y.t53 cap_res_Y.t91 0.1603
R3124 cap_res_Y.t109 cap_res_Y.t75 0.1603
R3125 cap_res_Y.t24 cap_res_Y.t54 0.1603
R3126 cap_res_Y.t77 cap_res_Y.t42 0.1603
R3127 cap_res_Y.t57 cap_res_Y.t93 0.1603
R3128 cap_res_Y.t115 cap_res_Y.t82 0.1603
R3129 cap_res_Y.t96 cap_res_Y.t2 0.1603
R3130 cap_res_Y.t15 cap_res_Y.t124 0.1603
R3131 cap_res_Y.t64 cap_res_Y.t98 0.1603
R3132 cap_res_Y.t126 cap_res_Y.t85 0.1603
R3133 cap_res_Y.t105 cap_res_Y.t5 0.1603
R3134 cap_res_Y.t22 cap_res_Y.t130 0.1603
R3135 cap_res_Y.t122 cap_res_Y.t69 0.1603
R3136 cap_res_Y.t133 cap_res_Y.t40 0.1603
R3137 cap_res_Y.t117 cap_res_Y.t67 0.1603
R3138 cap_res_Y.t76 cap_res_Y.t88 0.1603
R3139 cap_res_Y.t29 cap_res_Y.t128 0.1603
R3140 cap_res_Y.t120 cap_res_Y.t19 0.1603
R3141 cap_res_Y.t103 cap_res_Y.t68 0.1603
R3142 cap_res_Y.t55 cap_res_Y.t100 0.1603
R3143 cap_res_Y.t52 cap_res_Y.t56 0.1603
R3144 cap_res_Y.t44 cap_res_Y.t108 0.1603
R3145 cap_res_Y.t137 cap_res_Y.t7 0.1603
R3146 cap_res_Y.t87 cap_res_Y.t41 0.1603
R3147 cap_res_Y.t39 cap_res_Y.t74 0.1603
R3148 cap_res_Y.t21 cap_res_Y.t51 0.1603
R3149 cap_res_Y.t16 cap_res_Y.t50 0.1603
R3150 cap_res_Y.t46 cap_res_Y.t16 0.1603
R3151 cap_res_Y.t12 cap_res_Y.t46 0.1603
R3152 cap_res_Y.t60 cap_res_Y.t136 0.1603
R3153 cap_res_Y.t99 cap_res_Y.t31 0.1603
R3154 cap_res_Y.t4 cap_res_Y.t59 0.1603
R3155 cap_res_Y.t121 cap_res_Y.t113 0.1603
R3156 cap_res_Y.t114 cap_res_Y.t13 0.1603
R3157 cap_res_Y.t9 cap_res_Y.t114 0.1603
R3158 cap_res_Y.t18 cap_res_Y.t9 0.1603
R3159 cap_res_Y.t70 cap_res_Y.t107 0.1603
R3160 cap_res_Y.t102 cap_res_Y.t70 0.1603
R3161 cap_res_Y.t3 cap_res_Y.t102 0.1603
R3162 cap_res_Y.t14 cap_res_Y.t116 0.1603
R3163 cap_res_Y.t123 cap_res_Y.t14 0.1603
R3164 cap_res_Y.t20 cap_res_Y.t123 0.1603
R3165 cap_res_Y.n31 cap_res_Y.t30 0.159278
R3166 cap_res_Y.t25 cap_res_Y.n15 0.159278
R3167 cap_res_Y.t32 cap_res_Y.n16 0.159278
R3168 cap_res_Y.t73 cap_res_Y.n17 0.159278
R3169 cap_res_Y.t36 cap_res_Y.n18 0.159278
R3170 cap_res_Y.t62 cap_res_Y.n19 0.159278
R3171 cap_res_Y.t28 cap_res_Y.n20 0.159278
R3172 cap_res_Y.t132 cap_res_Y.n21 0.159278
R3173 cap_res_Y.t23 cap_res_Y.n22 0.159278
R3174 cap_res_Y.t127 cap_res_Y.n23 0.159278
R3175 cap_res_Y.t83 cap_res_Y.n24 0.159278
R3176 cap_res_Y.t43 cap_res_Y.n25 0.159278
R3177 cap_res_Y.t79 cap_res_Y.n26 0.159278
R3178 cap_res_Y.t38 cap_res_Y.n27 0.159278
R3179 cap_res_Y.t1 cap_res_Y.n28 0.159278
R3180 cap_res_Y.t34 cap_res_Y.n29 0.159278
R3181 cap_res_Y.t66 cap_res_Y.n30 0.159278
R3182 cap_res_Y.n32 cap_res_Y.t45 0.159278
R3183 cap_res_Y.n33 cap_res_Y.t11 0.159278
R3184 cap_res_Y.n34 cap_res_Y.t112 0.159278
R3185 cap_res_Y.n0 cap_res_Y.t26 0.159278
R3186 cap_res_Y.n1 cap_res_Y.t58 0.159278
R3187 cap_res_Y.n2 cap_res_Y.t95 0.159278
R3188 cap_res_Y.n3 cap_res_Y.t81 0.159278
R3189 cap_res_Y.n4 cap_res_Y.t119 0.159278
R3190 cap_res_Y.n5 cap_res_Y.t94 0.159278
R3191 cap_res_Y.n35 cap_res_Y.t78 0.159278
R3192 cap_res_Y.t30 cap_res_Y.t61 0.137822
R3193 cap_res_Y.n31 cap_res_Y.t104 0.1368
R3194 cap_res_Y.n30 cap_res_Y.t63 0.1368
R3195 cap_res_Y.n30 cap_res_Y.t125 0.1368
R3196 cap_res_Y.n29 cap_res_Y.t35 0.1368
R3197 cap_res_Y.n29 cap_res_Y.t86 0.1368
R3198 cap_res_Y.n28 cap_res_Y.t72 0.1368
R3199 cap_res_Y.n28 cap_res_Y.t131 0.1368
R3200 cap_res_Y.n27 cap_res_Y.t110 0.1368
R3201 cap_res_Y.n27 cap_res_Y.t27 0.1368
R3202 cap_res_Y.n26 cap_res_Y.t80 0.1368
R3203 cap_res_Y.n26 cap_res_Y.t135 0.1368
R3204 cap_res_Y.n25 cap_res_Y.t118 0.1368
R3205 cap_res_Y.n25 cap_res_Y.t33 0.1368
R3206 cap_res_Y.n24 cap_res_Y.t17 0.1368
R3207 cap_res_Y.n24 cap_res_Y.t71 0.1368
R3208 cap_res_Y.n23 cap_res_Y.t53 0.1368
R3209 cap_res_Y.n23 cap_res_Y.t109 0.1368
R3210 cap_res_Y.n22 cap_res_Y.t24 0.1368
R3211 cap_res_Y.n22 cap_res_Y.t77 0.1368
R3212 cap_res_Y.n21 cap_res_Y.t57 0.1368
R3213 cap_res_Y.n21 cap_res_Y.t115 0.1368
R3214 cap_res_Y.n20 cap_res_Y.t96 0.1368
R3215 cap_res_Y.n20 cap_res_Y.t15 0.1368
R3216 cap_res_Y.n19 cap_res_Y.t64 0.1368
R3217 cap_res_Y.n19 cap_res_Y.t126 0.1368
R3218 cap_res_Y.n18 cap_res_Y.t105 0.1368
R3219 cap_res_Y.n18 cap_res_Y.t22 0.1368
R3220 cap_res_Y.n17 cap_res_Y.t122 0.1368
R3221 cap_res_Y.n17 cap_res_Y.t133 0.1368
R3222 cap_res_Y.n16 cap_res_Y.t117 0.1368
R3223 cap_res_Y.n15 cap_res_Y.t21 0.1368
R3224 cap_res_Y.n6 cap_res_Y.t76 0.114322
R3225 cap_res_Y.n7 cap_res_Y.n6 0.1133
R3226 cap_res_Y.n8 cap_res_Y.n7 0.1133
R3227 cap_res_Y.n9 cap_res_Y.n8 0.1133
R3228 cap_res_Y.n10 cap_res_Y.n9 0.1133
R3229 cap_res_Y.n11 cap_res_Y.n10 0.1133
R3230 cap_res_Y.n12 cap_res_Y.n11 0.1133
R3231 cap_res_Y.n13 cap_res_Y.n12 0.1133
R3232 cap_res_Y.n14 cap_res_Y.n13 0.1133
R3233 cap_res_Y.n16 cap_res_Y.n14 0.1133
R3234 cap_res_Y.n32 cap_res_Y.n31 0.1133
R3235 cap_res_Y.n33 cap_res_Y.n32 0.1133
R3236 cap_res_Y.n34 cap_res_Y.n33 0.1133
R3237 cap_res_Y.n1 cap_res_Y.n0 0.1133
R3238 cap_res_Y.n2 cap_res_Y.n1 0.1133
R3239 cap_res_Y.n3 cap_res_Y.n2 0.1133
R3240 cap_res_Y.n4 cap_res_Y.n3 0.1133
R3241 cap_res_Y.n5 cap_res_Y.n4 0.1133
R3242 cap_res_Y.n35 cap_res_Y.n5 0.1133
R3243 cap_res_Y.n35 cap_res_Y.n34 0.1133
R3244 cap_res_Y.n6 cap_res_Y.t29 0.00152174
R3245 cap_res_Y.n7 cap_res_Y.t120 0.00152174
R3246 cap_res_Y.n8 cap_res_Y.t103 0.00152174
R3247 cap_res_Y.n9 cap_res_Y.t55 0.00152174
R3248 cap_res_Y.n10 cap_res_Y.t52 0.00152174
R3249 cap_res_Y.n11 cap_res_Y.t44 0.00152174
R3250 cap_res_Y.n12 cap_res_Y.t137 0.00152174
R3251 cap_res_Y.n13 cap_res_Y.t87 0.00152174
R3252 cap_res_Y.n14 cap_res_Y.t39 0.00152174
R3253 cap_res_Y.n15 cap_res_Y.t129 0.00152174
R3254 cap_res_Y.n16 cap_res_Y.t25 0.00152174
R3255 cap_res_Y.n17 cap_res_Y.t32 0.00152174
R3256 cap_res_Y.n18 cap_res_Y.t73 0.00152174
R3257 cap_res_Y.n19 cap_res_Y.t36 0.00152174
R3258 cap_res_Y.n20 cap_res_Y.t62 0.00152174
R3259 cap_res_Y.n21 cap_res_Y.t28 0.00152174
R3260 cap_res_Y.n22 cap_res_Y.t132 0.00152174
R3261 cap_res_Y.n23 cap_res_Y.t23 0.00152174
R3262 cap_res_Y.n24 cap_res_Y.t127 0.00152174
R3263 cap_res_Y.n25 cap_res_Y.t83 0.00152174
R3264 cap_res_Y.n26 cap_res_Y.t43 0.00152174
R3265 cap_res_Y.n27 cap_res_Y.t79 0.00152174
R3266 cap_res_Y.n28 cap_res_Y.t38 0.00152174
R3267 cap_res_Y.n29 cap_res_Y.t1 0.00152174
R3268 cap_res_Y.n30 cap_res_Y.t34 0.00152174
R3269 cap_res_Y.n31 cap_res_Y.t66 0.00152174
R3270 cap_res_Y.n32 cap_res_Y.t89 0.00152174
R3271 cap_res_Y.n33 cap_res_Y.t49 0.00152174
R3272 cap_res_Y.n34 cap_res_Y.t12 0.00152174
R3273 cap_res_Y.n0 cap_res_Y.t60 0.00152174
R3274 cap_res_Y.n1 cap_res_Y.t99 0.00152174
R3275 cap_res_Y.n2 cap_res_Y.t4 0.00152174
R3276 cap_res_Y.n3 cap_res_Y.t121 0.00152174
R3277 cap_res_Y.n4 cap_res_Y.t18 0.00152174
R3278 cap_res_Y.n5 cap_res_Y.t3 0.00152174
R3279 cap_res_Y.t116 cap_res_Y.n35 0.00152174
R3280 V_tail_gate.n11 V_tail_gate.t11 610.534
R3281 V_tail_gate.n2 V_tail_gate.t8 610.534
R3282 V_tail_gate.n11 V_tail_gate.t21 433.8
R3283 V_tail_gate.n12 V_tail_gate.t9 433.8
R3284 V_tail_gate.n13 V_tail_gate.t18 433.8
R3285 V_tail_gate.n14 V_tail_gate.t14 433.8
R3286 V_tail_gate.n15 V_tail_gate.t23 433.8
R3287 V_tail_gate.n16 V_tail_gate.t12 433.8
R3288 V_tail_gate.n17 V_tail_gate.t16 433.8
R3289 V_tail_gate.n18 V_tail_gate.t5 433.8
R3290 V_tail_gate.n19 V_tail_gate.t15 433.8
R3291 V_tail_gate.n10 V_tail_gate.t4 433.8
R3292 V_tail_gate.n9 V_tail_gate.t13 433.8
R3293 V_tail_gate.n8 V_tail_gate.t22 433.8
R3294 V_tail_gate.n7 V_tail_gate.t19 433.8
R3295 V_tail_gate.n6 V_tail_gate.t7 433.8
R3296 V_tail_gate.n5 V_tail_gate.t17 433.8
R3297 V_tail_gate.n4 V_tail_gate.t6 433.8
R3298 V_tail_gate.n3 V_tail_gate.t10 433.8
R3299 V_tail_gate.n2 V_tail_gate.t20 433.8
R3300 V_tail_gate.n21 V_tail_gate.n20 221.356
R3301 V_tail_gate.n19 V_tail_gate.n18 176.733
R3302 V_tail_gate.n18 V_tail_gate.n17 176.733
R3303 V_tail_gate.n17 V_tail_gate.n16 176.733
R3304 V_tail_gate.n16 V_tail_gate.n15 176.733
R3305 V_tail_gate.n15 V_tail_gate.n14 176.733
R3306 V_tail_gate.n14 V_tail_gate.n13 176.733
R3307 V_tail_gate.n13 V_tail_gate.n12 176.733
R3308 V_tail_gate.n12 V_tail_gate.n11 176.733
R3309 V_tail_gate.n3 V_tail_gate.n2 176.733
R3310 V_tail_gate.n4 V_tail_gate.n3 176.733
R3311 V_tail_gate.n5 V_tail_gate.n4 176.733
R3312 V_tail_gate.n6 V_tail_gate.n5 176.733
R3313 V_tail_gate.n7 V_tail_gate.n6 176.733
R3314 V_tail_gate.n8 V_tail_gate.n7 176.733
R3315 V_tail_gate.n9 V_tail_gate.n8 176.733
R3316 V_tail_gate.n10 V_tail_gate.n9 176.733
R3317 V_tail_gate.n22 V_tail_gate.n0 113.261
R3318 V_tail_gate.n22 V_tail_gate.n21 69.7049
R3319 V_tail_gate.n20 V_tail_gate.n19 56.2338
R3320 V_tail_gate.n20 V_tail_gate.n10 56.2338
R3321 V_tail_gate.n21 V_tail_gate.n1 53.2453
R3322 V_tail_gate.n0 V_tail_gate.t3 16.0005
R3323 V_tail_gate.n0 V_tail_gate.t0 16.0005
R3324 V_tail_gate.n1 V_tail_gate.t1 16.0005
R3325 V_tail_gate.n1 V_tail_gate.t2 16.0005
R3326 V_tail_gate V_tail_gate.n22 0.063
R3327 err_amp_out.n0 err_amp_out.t12 669.486
R3328 err_amp_out err_amp_out.n1 631.982
R3329 err_amp_out err_amp_out.n3 627.128
R3330 err_amp_out err_amp_out.n2 627.128
R3331 err_amp_out.n0 err_amp_out.n6 226.534
R3332 err_amp_out.n0 err_amp_out.n5 226.534
R3333 err_amp_out.n7 err_amp_out.n4 222.034
R3334 err_amp_out.n3 err_amp_out.t5 78.8005
R3335 err_amp_out.n3 err_amp_out.t4 78.8005
R3336 err_amp_out.n2 err_amp_out.t0 78.8005
R3337 err_amp_out.n2 err_amp_out.t3 78.8005
R3338 err_amp_out.n1 err_amp_out.t6 78.8005
R3339 err_amp_out.n1 err_amp_out.t9 78.8005
R3340 err_amp_out.n6 err_amp_out.t8 48.0005
R3341 err_amp_out.n6 err_amp_out.t2 48.0005
R3342 err_amp_out.n4 err_amp_out.t11 48.0005
R3343 err_amp_out.n4 err_amp_out.t7 48.0005
R3344 err_amp_out.n5 err_amp_out.t10 48.0005
R3345 err_amp_out.n5 err_amp_out.t1 48.0005
R3346 err_amp_out err_amp_out.n7 10.2505
R3347 err_amp_out.n7 err_amp_out.n0 7.0005
R3348 V_CMFB_S2.n11 V_CMFB_S2.t0 120.66
R3349 V_CMFB_S2.n4 V_CMFB_S2.n3 96.8384
R3350 V_CMFB_S2.n6 V_CMFB_S2.n5 96.8384
R3351 V_CMFB_S2.n8 V_CMFB_S2.n7 96.8384
R3352 V_CMFB_S2.n10 V_CMFB_S2.n9 96.8384
R3353 V_CMFB_S2.n2 V_CMFB_S2.n1 92.3384
R3354 V_CMFB_S2.n1 V_CMFB_S2.t6 8.0005
R3355 V_CMFB_S2.n1 V_CMFB_S2.t1 8.0005
R3356 V_CMFB_S2.n3 V_CMFB_S2.t10 8.0005
R3357 V_CMFB_S2.n3 V_CMFB_S2.t4 8.0005
R3358 V_CMFB_S2.n5 V_CMFB_S2.t7 8.0005
R3359 V_CMFB_S2.n5 V_CMFB_S2.t5 8.0005
R3360 V_CMFB_S2.n7 V_CMFB_S2.t8 8.0005
R3361 V_CMFB_S2.n7 V_CMFB_S2.t2 8.0005
R3362 V_CMFB_S2.n9 V_CMFB_S2.t9 8.0005
R3363 V_CMFB_S2.n9 V_CMFB_S2.t3 8.0005
R3364 V_CMFB_S2.n11 V_CMFB_S2.n10 5.938
R3365 V_CMFB_S2.n4 V_CMFB_S2.n2 5.063
R3366 V_CMFB_S2.n2 V_CMFB_S2.n0 2.15675
R3367 V_CMFB_S2.n10 V_CMFB_S2.n8 0.563
R3368 V_CMFB_S2.n8 V_CMFB_S2.n6 0.563
R3369 V_CMFB_S2.n6 V_CMFB_S2.n4 0.563
R3370 V_CMFB_S2 V_CMFB_S2.n11 0.063
R3371 V_CMFB_S4.n9 V_CMFB_S4.t0 120.66
R3372 V_CMFB_S4.n2 V_CMFB_S4.n0 97.4009
R3373 V_CMFB_S4.n8 V_CMFB_S4.n7 96.8384
R3374 V_CMFB_S4.n6 V_CMFB_S4.n5 96.8384
R3375 V_CMFB_S4.n4 V_CMFB_S4.n3 96.8384
R3376 V_CMFB_S4.n2 V_CMFB_S4.n1 96.8384
R3377 V_CMFB_S4.n7 V_CMFB_S4.t10 8.0005
R3378 V_CMFB_S4.n7 V_CMFB_S4.t4 8.0005
R3379 V_CMFB_S4.n5 V_CMFB_S4.t1 8.0005
R3380 V_CMFB_S4.n5 V_CMFB_S4.t5 8.0005
R3381 V_CMFB_S4.n3 V_CMFB_S4.t2 8.0005
R3382 V_CMFB_S4.n3 V_CMFB_S4.t6 8.0005
R3383 V_CMFB_S4.n1 V_CMFB_S4.t3 8.0005
R3384 V_CMFB_S4.n1 V_CMFB_S4.t7 8.0005
R3385 V_CMFB_S4.n0 V_CMFB_S4.t9 8.0005
R3386 V_CMFB_S4.n0 V_CMFB_S4.t8 8.0005
R3387 V_CMFB_S4.n9 V_CMFB_S4.n8 5.938
R3388 V_CMFB_S4.n4 V_CMFB_S4.n2 0.563
R3389 V_CMFB_S4.n6 V_CMFB_S4.n4 0.563
R3390 V_CMFB_S4.n8 V_CMFB_S4.n6 0.563
R3391 V_CMFB_S4 V_CMFB_S4.n9 0.063
R3392 V_err_gate.n21 V_err_gate.n19 630.857
R3393 V_err_gate.n24 V_err_gate.n22 627.316
R3394 V_err_gate.n26 V_err_gate.n25 626.784
R3395 V_err_gate.n24 V_err_gate.n23 626.784
R3396 V_err_gate.n21 V_err_gate.n20 626.784
R3397 V_err_gate.n29 V_err_gate.n28 585
R3398 V_err_gate.n16 V_err_gate.t19 289.2
R3399 V_err_gate.n0 V_err_gate.t15 289.2
R3400 V_err_gate.n17 V_err_gate.n16 176.733
R3401 V_err_gate.n1 V_err_gate.n0 176.733
R3402 V_err_gate.n2 V_err_gate.n1 176.733
R3403 V_err_gate.n3 V_err_gate.n2 176.733
R3404 V_err_gate.n4 V_err_gate.n3 176.733
R3405 V_err_gate.n5 V_err_gate.n4 176.733
R3406 V_err_gate.n6 V_err_gate.n5 176.733
R3407 V_err_gate.n7 V_err_gate.n6 176.733
R3408 V_err_gate.n8 V_err_gate.n7 176.733
R3409 V_err_gate.n9 V_err_gate.n8 176.733
R3410 V_err_gate.n10 V_err_gate.n9 176.733
R3411 V_err_gate.n11 V_err_gate.n10 176.733
R3412 V_err_gate.n12 V_err_gate.n11 176.733
R3413 V_err_gate.n13 V_err_gate.n12 176.733
R3414 V_err_gate.n14 V_err_gate.n13 176.733
R3415 V_err_gate.n15 V_err_gate.n14 176.733
R3416 V_err_gate V_err_gate.n18 162.494
R3417 V_err_gate.n17 V_err_gate.t16 112.468
R3418 V_err_gate.n16 V_err_gate.t27 112.468
R3419 V_err_gate.n0 V_err_gate.t26 112.468
R3420 V_err_gate.n1 V_err_gate.t18 112.468
R3421 V_err_gate.n2 V_err_gate.t28 112.468
R3422 V_err_gate.n3 V_err_gate.t24 112.468
R3423 V_err_gate.n4 V_err_gate.t14 112.468
R3424 V_err_gate.n5 V_err_gate.t25 112.468
R3425 V_err_gate.n6 V_err_gate.t17 112.468
R3426 V_err_gate.n7 V_err_gate.t20 112.468
R3427 V_err_gate.n8 V_err_gate.t30 112.468
R3428 V_err_gate.n9 V_err_gate.t22 112.468
R3429 V_err_gate.n10 V_err_gate.t12 112.468
R3430 V_err_gate.n11 V_err_gate.t23 112.468
R3431 V_err_gate.n12 V_err_gate.t13 112.468
R3432 V_err_gate.n13 V_err_gate.t29 112.468
R3433 V_err_gate.n14 V_err_gate.t21 112.468
R3434 V_err_gate.n15 V_err_gate.t31 112.468
R3435 V_err_gate.n28 V_err_gate.t8 78.8005
R3436 V_err_gate.n28 V_err_gate.t0 78.8005
R3437 V_err_gate.n25 V_err_gate.t4 78.8005
R3438 V_err_gate.n25 V_err_gate.t9 78.8005
R3439 V_err_gate.n23 V_err_gate.t5 78.8005
R3440 V_err_gate.n23 V_err_gate.t7 78.8005
R3441 V_err_gate.n22 V_err_gate.t1 78.8005
R3442 V_err_gate.n22 V_err_gate.t11 78.8005
R3443 V_err_gate.n20 V_err_gate.t2 78.8005
R3444 V_err_gate.n20 V_err_gate.t6 78.8005
R3445 V_err_gate.n19 V_err_gate.t10 78.8005
R3446 V_err_gate.n19 V_err_gate.t3 78.8005
R3447 V_err_gate.n18 V_err_gate.n17 49.8072
R3448 V_err_gate.n18 V_err_gate.n15 49.8072
R3449 V_err_gate.n29 V_err_gate.n27 41.7838
R3450 V_err_gate V_err_gate.n29 39.8443
R3451 V_err_gate.n26 V_err_gate.n24 0.59425
R3452 V_err_gate.n27 V_err_gate.n21 0.59425
R3453 V_err_gate.n27 V_err_gate.n26 0.53175
R3454 V_err_p.n5 V_err_p.n3 630.827
R3455 V_err_p.n9 V_err_p.n8 630.264
R3456 V_err_p.n7 V_err_p.n6 630.264
R3457 V_err_p.n5 V_err_p.n4 630.264
R3458 V_err_p.n17 V_err_p.n15 627.784
R3459 V_err_p.n12 V_err_p.n0 627.784
R3460 V_err_p.n10 V_err_p.n2 627.168
R3461 V_err_p.n17 V_err_p.n16 626.534
R3462 V_err_p.n14 V_err_p.n13 626.534
R3463 V_err_p.n19 V_err_p.n18 626.534
R3464 V_err_p.n11 V_err_p.n1 622.034
R3465 V_err_p.n16 V_err_p.t15 78.8005
R3466 V_err_p.n16 V_err_p.t11 78.8005
R3467 V_err_p.n15 V_err_p.t17 78.8005
R3468 V_err_p.n15 V_err_p.t9 78.8005
R3469 V_err_p.n13 V_err_p.t18 78.8005
R3470 V_err_p.n13 V_err_p.t16 78.8005
R3471 V_err_p.n1 V_err_p.t12 78.8005
R3472 V_err_p.n1 V_err_p.t13 78.8005
R3473 V_err_p.n8 V_err_p.t8 78.8005
R3474 V_err_p.n8 V_err_p.t6 78.8005
R3475 V_err_p.n6 V_err_p.t4 78.8005
R3476 V_err_p.n6 V_err_p.t7 78.8005
R3477 V_err_p.n4 V_err_p.t3 78.8005
R3478 V_err_p.n4 V_err_p.t0 78.8005
R3479 V_err_p.n3 V_err_p.t21 78.8005
R3480 V_err_p.n3 V_err_p.t2 78.8005
R3481 V_err_p.n2 V_err_p.t5 78.8005
R3482 V_err_p.n2 V_err_p.t1 78.8005
R3483 V_err_p.n0 V_err_p.t10 78.8005
R3484 V_err_p.n0 V_err_p.t19 78.8005
R3485 V_err_p.t20 V_err_p.n19 78.8005
R3486 V_err_p.n19 V_err_p.t14 78.8005
R3487 V_err_p.n10 V_err_p.n9 5.0005
R3488 V_err_p.n12 V_err_p.n11 4.5005
R3489 V_err_p.n11 V_err_p.n10 1.60845
R3490 V_err_p.n18 V_err_p.n17 1.2505
R3491 V_err_p.n14 V_err_p.n12 1.2505
R3492 V_err_p.n18 V_err_p.n14 1.2505
R3493 V_err_p.n7 V_err_p.n5 0.563
R3494 V_err_p.n9 V_err_p.n7 0.563
R3495 Vb2_Vb3.n1 Vb2_Vb3.t0 720.312
R3496 Vb2_Vb3.n2 Vb2_Vb3.t3 720.312
R3497 Vb2_Vb3.t1 Vb2_Vb3.n1 207.362
R3498 Vb2_Vb3.n2 Vb2_Vb3.t4 207.362
R3499 Vb2_Vb3 Vb2_Vb3.n5 179.933
R3500 Vb2_Vb3.n4 Vb2_Vb3.n0 170.3
R3501 Vb2_Vb3.t9 Vb2_Vb3.t1 142.5
R3502 Vb2_Vb3.t4 Vb2_Vb3.t9 142.5
R3503 Vb2_Vb3.n1 Vb2_Vb3.t2 75.9449
R3504 Vb2_Vb3.n2 Vb2_Vb3.t6 75.9449
R3505 Vb2_Vb3.n3 Vb2_Vb3.n1 66.5398
R3506 Vb2_Vb3.n3 Vb2_Vb3.n2 66.1648
R3507 Vb2_Vb3.n5 Vb2_Vb3.t7 11.0991
R3508 Vb2_Vb3.n5 Vb2_Vb3.t8 11.0991
R3509 Vb2_Vb3.n0 Vb2_Vb3.t10 10.9449
R3510 Vb2_Vb3.n0 Vb2_Vb3.t5 10.9449
R3511 Vb2_Vb3 Vb2_Vb3.n4 6.21925
R3512 Vb2_Vb3.n4 Vb2_Vb3.n3 4.5005
R3513 Vb1.n14 Vb1.t3 449.868
R3514 Vb1.n10 Vb1.t5 449.868
R3515 Vb1.n5 Vb1.t4 449.868
R3516 Vb1.n1 Vb1.t6 449.868
R3517 Vb1.n14 Vb1.t13 273.134
R3518 Vb1.n15 Vb1.t21 273.134
R3519 Vb1.n16 Vb1.t11 273.134
R3520 Vb1.n17 Vb1.t18 273.134
R3521 Vb1.n13 Vb1.t7 273.134
R3522 Vb1.n12 Vb1.t19 273.134
R3523 Vb1.n11 Vb1.t8 273.134
R3524 Vb1.n10 Vb1.t16 273.134
R3525 Vb1.n5 Vb1.t14 273.134
R3526 Vb1.n6 Vb1.t2 273.134
R3527 Vb1.n7 Vb1.t12 273.134
R3528 Vb1.n8 Vb1.t20 273.134
R3529 Vb1.n4 Vb1.t9 273.134
R3530 Vb1.n3 Vb1.t15 273.134
R3531 Vb1.n2 Vb1.t10 273.134
R3532 Vb1.n1 Vb1.t17 273.134
R3533 Vb1.n0 Vb1.t1 184.625
R3534 Vb1.n17 Vb1.n16 176.733
R3535 Vb1.n16 Vb1.n15 176.733
R3536 Vb1.n15 Vb1.n14 176.733
R3537 Vb1.n11 Vb1.n10 176.733
R3538 Vb1.n12 Vb1.n11 176.733
R3539 Vb1.n13 Vb1.n12 176.733
R3540 Vb1.n8 Vb1.n7 176.733
R3541 Vb1.n7 Vb1.n6 176.733
R3542 Vb1.n6 Vb1.n5 176.733
R3543 Vb1.n2 Vb1.n1 176.733
R3544 Vb1.n3 Vb1.n2 176.733
R3545 Vb1.n4 Vb1.n3 176.733
R3546 Vb1.n19 Vb1.n9 171.644
R3547 Vb1.n19 Vb1.n18 165.8
R3548 Vb1.n0 Vb1.t0 61.1914
R3549 Vb1.n18 Vb1.n17 56.2338
R3550 Vb1.n18 Vb1.n13 56.2338
R3551 Vb1.n9 Vb1.n8 56.2338
R3552 Vb1.n9 Vb1.n4 56.2338
R3553 Vb1.n20 Vb1.n0 23.6235
R3554 Vb1.n20 Vb1.n19 7.98488
R3555 Vb1 Vb1.n20 0.063
R3556 V_tot.n6 V_tot.t13 327.623
R3557 V_tot.n4 V_tot.t12 326.365
R3558 V_tot.n5 V_tot.t6 168.701
R3559 V_tot.n5 V_tot.t11 168.701
R3560 V_tot.n3 V_tot.n1 167.05
R3561 V_tot.n8 V_tot.n7 165.8
R3562 V_tot.n6 V_tot.n5 165.8
R3563 V_tot.n3 V_tot.n2 165.8
R3564 V_tot.n7 V_tot.t8 157.989
R3565 V_tot.n7 V_tot.t10 157.989
R3566 V_tot.n2 V_tot.t5 157.989
R3567 V_tot.n2 V_tot.t7 157.989
R3568 V_tot.n1 V_tot.t4 157.989
R3569 V_tot.n1 V_tot.t9 157.989
R3570 V_tot.n0 V_tot.t1 117.591
R3571 V_tot.t0 V_tot.n11 117.591
R3572 V_tot.n11 V_tot.t2 108.424
R3573 V_tot.n0 V_tot.t3 108.424
R3574 V_tot.n11 V_tot.n10 36.3621
R3575 V_tot.n10 V_tot.n0 35.9871
R3576 V_tot.n10 V_tot.n9 10.6255
R3577 V_tot.n9 V_tot.n8 2.063
R3578 V_tot.n8 V_tot.n6 1.26612
R3579 V_tot.n4 V_tot.n3 1.15363
R3580 V_tot.n9 V_tot.n4 1.12862
R3581 err_amp_mir.n4 err_amp_mir.n2 628.034
R3582 err_amp_mir.n4 err_amp_mir.n3 626.784
R3583 err_amp_mir.n5 err_amp_mir.n1 622.284
R3584 err_amp_mir.n18 err_amp_mir.t19 289.2
R3585 err_amp_mir.n8 err_amp_mir.t2 289.2
R3586 err_amp_mir.n6 err_amp_mir.n0 227.252
R3587 err_amp_mir.n12 err_amp_mir.n11 212.733
R3588 err_amp_mir.n21 err_amp_mir.n20 212.733
R3589 err_amp_mir.n15 err_amp_mir.n14 176.733
R3590 err_amp_mir.n16 err_amp_mir.n15 176.733
R3591 err_amp_mir.n17 err_amp_mir.n16 176.733
R3592 err_amp_mir.n9 err_amp_mir.n8 176.733
R3593 err_amp_mir.n10 err_amp_mir.n9 176.733
R3594 err_amp_mir.n13 err_amp_mir.n12 152
R3595 err_amp_mir.n20 err_amp_mir.n19 152
R3596 err_amp_mir.n18 err_amp_mir.t4 112.468
R3597 err_amp_mir.n17 err_amp_mir.t8 112.468
R3598 err_amp_mir.n16 err_amp_mir.t20 112.468
R3599 err_amp_mir.n15 err_amp_mir.t17 112.468
R3600 err_amp_mir.n14 err_amp_mir.t6 112.468
R3601 err_amp_mir.n10 err_amp_mir.t0 112.468
R3602 err_amp_mir.n9 err_amp_mir.t21 112.468
R3603 err_amp_mir.n8 err_amp_mir.t18 112.468
R3604 err_amp_mir.n3 err_amp_mir.t14 78.8005
R3605 err_amp_mir.n3 err_amp_mir.t15 78.8005
R3606 err_amp_mir.n2 err_amp_mir.t13 78.8005
R3607 err_amp_mir.n2 err_amp_mir.t16 78.8005
R3608 err_amp_mir.n1 err_amp_mir.t12 78.8005
R3609 err_amp_mir.n1 err_amp_mir.t10 78.8005
R3610 err_amp_mir.n11 err_amp_mir.t1 48.0005
R3611 err_amp_mir.n11 err_amp_mir.t7 48.0005
R3612 err_amp_mir.n0 err_amp_mir.t11 48.0005
R3613 err_amp_mir.n0 err_amp_mir.t3 48.0005
R3614 err_amp_mir.t9 err_amp_mir.n21 48.0005
R3615 err_amp_mir.n21 err_amp_mir.t5 48.0005
R3616 err_amp_mir.n19 err_amp_mir.n18 45.5227
R3617 err_amp_mir.n19 err_amp_mir.n17 45.5227
R3618 err_amp_mir.n14 err_amp_mir.n13 45.5227
R3619 err_amp_mir.n13 err_amp_mir.n10 45.5227
R3620 err_amp_mir.n20 err_amp_mir.n7 15.488
R3621 err_amp_mir.n12 err_amp_mir.n7 14.1755
R3622 err_amp_mir.n5 err_amp_mir.n4 5.7505
R3623 err_amp_mir.n6 err_amp_mir.n5 5.28175
R3624 err_amp_mir.n7 err_amp_mir.n6 0.84425
R3625 V_CMFB_S1.n4 V_CMFB_S1.n3 205.488
R3626 V_CMFB_S1.n6 V_CMFB_S1.n5 205.488
R3627 V_CMFB_S1.n8 V_CMFB_S1.n7 205.488
R3628 V_CMFB_S1.n10 V_CMFB_S1.n9 205.488
R3629 V_CMFB_S1.n2 V_CMFB_S1.n1 200.988
R3630 V_CMFB_S1.n11 V_CMFB_S1.t0 122.504
R3631 V_CMFB_S1.n1 V_CMFB_S1.t8 19.7005
R3632 V_CMFB_S1.n1 V_CMFB_S1.t3 19.7005
R3633 V_CMFB_S1.n3 V_CMFB_S1.t2 19.7005
R3634 V_CMFB_S1.n3 V_CMFB_S1.t6 19.7005
R3635 V_CMFB_S1.n5 V_CMFB_S1.t9 19.7005
R3636 V_CMFB_S1.n5 V_CMFB_S1.t7 19.7005
R3637 V_CMFB_S1.n7 V_CMFB_S1.t10 19.7005
R3638 V_CMFB_S1.n7 V_CMFB_S1.t4 19.7005
R3639 V_CMFB_S1.n9 V_CMFB_S1.t1 19.7005
R3640 V_CMFB_S1.n9 V_CMFB_S1.t5 19.7005
R3641 V_CMFB_S1.n11 V_CMFB_S1.n10 6.21925
R3642 V_CMFB_S1.n4 V_CMFB_S1.n2 5.063
R3643 V_CMFB_S1.n2 V_CMFB_S1.n0 2.29738
R3644 V_CMFB_S1.n10 V_CMFB_S1.n8 0.563
R3645 V_CMFB_S1.n8 V_CMFB_S1.n6 0.563
R3646 V_CMFB_S1.n6 V_CMFB_S1.n4 0.563
R3647 V_CMFB_S1 V_CMFB_S1.n11 0.063
R3648 VD2.n2 VD2.n0 114.719
R3649 VD2.n19 VD2.n18 114.719
R3650 VD2.n4 VD2.n3 114.156
R3651 VD2.n2 VD2.n1 114.156
R3652 VD2.n14 VD2.n12 112.456
R3653 VD2.n9 VD2.n7 112.456
R3654 VD2.n14 VD2.n13 111.206
R3655 VD2.n11 VD2.n10 111.206
R3656 VD2.n9 VD2.n8 111.206
R3657 VD2.n17 VD2.n5 109.656
R3658 VD2.n16 VD2.n6 106.706
R3659 VD2.n5 VD2.t18 16.0005
R3660 VD2.n5 VD2.t13 16.0005
R3661 VD2.n13 VD2.t6 16.0005
R3662 VD2.n13 VD2.t4 16.0005
R3663 VD2.n12 VD2.t5 16.0005
R3664 VD2.n12 VD2.t11 16.0005
R3665 VD2.n10 VD2.t9 16.0005
R3666 VD2.n10 VD2.t10 16.0005
R3667 VD2.n8 VD2.t2 16.0005
R3668 VD2.n8 VD2.t1 16.0005
R3669 VD2.n7 VD2.t0 16.0005
R3670 VD2.n7 VD2.t7 16.0005
R3671 VD2.n6 VD2.t3 16.0005
R3672 VD2.n6 VD2.t8 16.0005
R3673 VD2.n3 VD2.t19 16.0005
R3674 VD2.n3 VD2.t14 16.0005
R3675 VD2.n1 VD2.t17 16.0005
R3676 VD2.n1 VD2.t12 16.0005
R3677 VD2.n0 VD2.t16 16.0005
R3678 VD2.n0 VD2.t21 16.0005
R3679 VD2.t20 VD2.n19 16.0005
R3680 VD2.n19 VD2.t15 16.0005
R3681 VD2.n16 VD2.n15 4.5005
R3682 VD2.n18 VD2.n17 4.5005
R3683 VD2.n15 VD2.n11 3.6255
R3684 VD2.n15 VD2.n14 1.2505
R3685 VD2.n11 VD2.n9 1.2505
R3686 VD2.n17 VD2.n16 0.78175
R3687 VD2.n4 VD2.n2 0.563
R3688 VD2.n18 VD2.n4 0.563
R3689 V_CMFB_S3.n2 V_CMFB_S3.n0 206.052
R3690 V_CMFB_S3.n8 V_CMFB_S3.n7 205.488
R3691 V_CMFB_S3.n6 V_CMFB_S3.n5 205.488
R3692 V_CMFB_S3.n4 V_CMFB_S3.n3 205.488
R3693 V_CMFB_S3.n2 V_CMFB_S3.n1 205.488
R3694 V_CMFB_S3.n9 V_CMFB_S3.t0 122.504
R3695 V_CMFB_S3.n7 V_CMFB_S3.t2 19.7005
R3696 V_CMFB_S3.n7 V_CMFB_S3.t6 19.7005
R3697 V_CMFB_S3.n5 V_CMFB_S3.t3 19.7005
R3698 V_CMFB_S3.n5 V_CMFB_S3.t7 19.7005
R3699 V_CMFB_S3.n3 V_CMFB_S3.t4 19.7005
R3700 V_CMFB_S3.n3 V_CMFB_S3.t8 19.7005
R3701 V_CMFB_S3.n1 V_CMFB_S3.t5 19.7005
R3702 V_CMFB_S3.n1 V_CMFB_S3.t9 19.7005
R3703 V_CMFB_S3.n0 V_CMFB_S3.t1 19.7005
R3704 V_CMFB_S3.n0 V_CMFB_S3.t10 19.7005
R3705 V_CMFB_S3.n9 V_CMFB_S3.n8 6.21925
R3706 V_CMFB_S3.n4 V_CMFB_S3.n2 0.563
R3707 V_CMFB_S3.n6 V_CMFB_S3.n4 0.563
R3708 V_CMFB_S3.n8 V_CMFB_S3.n6 0.563
R3709 V_CMFB_S3 V_CMFB_S3.n9 0.063
R3710 V_err_amp_ref.n1 V_err_amp_ref.t9 323.491
R3711 V_err_amp_ref.n4 V_err_amp_ref.t0 322.692
R3712 V_err_amp_ref.n7 V_err_amp_ref.t4 270.591
R3713 V_err_amp_ref.n5 V_err_amp_ref.t1 270.591
R3714 V_err_amp_ref.n2 V_err_amp_ref.t2 270.591
R3715 V_err_amp_ref.n0 V_err_amp_ref.t7 270.591
R3716 V_err_amp_ref.n8 V_err_amp_ref.n7 233.374
R3717 V_err_amp_ref.n6 V_err_amp_ref.n5 233.374
R3718 V_err_amp_ref.n3 V_err_amp_ref.n2 233.374
R3719 V_err_amp_ref.n1 V_err_amp_ref.n0 233.374
R3720 V_err_amp_ref.n7 V_err_amp_ref.t8 129.24
R3721 V_err_amp_ref.n5 V_err_amp_ref.t5 129.24
R3722 V_err_amp_ref.n2 V_err_amp_ref.t6 129.24
R3723 V_err_amp_ref.n0 V_err_amp_ref.t3 129.24
R3724 V_err_amp_ref.n4 V_err_amp_ref.n3 3.688
R3725 V_err_amp_ref V_err_amp_ref.n8 2.0005
R3726 V_err_amp_ref.n3 V_err_amp_ref.n1 1.2755
R3727 V_err_amp_ref.n8 V_err_amp_ref.n6 1.2755
R3728 V_err_amp_ref.n6 V_err_amp_ref.n4 0.8005
R3729 V_err_mir_p.n3 V_err_mir_p.n1 632.186
R3730 V_err_mir_p.n7 V_err_mir_p.n6 630.264
R3731 V_err_mir_p.n5 V_err_mir_p.n4 630.264
R3732 V_err_mir_p.n3 V_err_mir_p.n2 630.264
R3733 V_err_mir_p.n15 V_err_mir_p.n14 628.003
R3734 V_err_mir_p.n11 V_err_mir_p.n9 628.003
R3735 V_err_mir_p.n13 V_err_mir_p.n12 626.753
R3736 V_err_mir_p.n11 V_err_mir_p.n10 626.753
R3737 V_err_mir_p.n8 V_err_mir_p.n0 625.756
R3738 V_err_mir_p.n17 V_err_mir_p.n16 622.231
R3739 V_err_mir_p.n14 V_err_mir_p.t12 78.8005
R3740 V_err_mir_p.n14 V_err_mir_p.t7 78.8005
R3741 V_err_mir_p.n12 V_err_mir_p.t5 78.8005
R3742 V_err_mir_p.n12 V_err_mir_p.t10 78.8005
R3743 V_err_mir_p.n10 V_err_mir_p.t13 78.8005
R3744 V_err_mir_p.n10 V_err_mir_p.t9 78.8005
R3745 V_err_mir_p.n9 V_err_mir_p.t8 78.8005
R3746 V_err_mir_p.n9 V_err_mir_p.t11 78.8005
R3747 V_err_mir_p.n6 V_err_mir_p.t18 78.8005
R3748 V_err_mir_p.n6 V_err_mir_p.t1 78.8005
R3749 V_err_mir_p.n4 V_err_mir_p.t3 78.8005
R3750 V_err_mir_p.n4 V_err_mir_p.t16 78.8005
R3751 V_err_mir_p.n2 V_err_mir_p.t19 78.8005
R3752 V_err_mir_p.n2 V_err_mir_p.t0 78.8005
R3753 V_err_mir_p.n1 V_err_mir_p.t2 78.8005
R3754 V_err_mir_p.n1 V_err_mir_p.t15 78.8005
R3755 V_err_mir_p.n0 V_err_mir_p.t4 78.8005
R3756 V_err_mir_p.n0 V_err_mir_p.t17 78.8005
R3757 V_err_mir_p.t14 V_err_mir_p.n17 78.8005
R3758 V_err_mir_p.n17 V_err_mir_p.t6 78.8005
R3759 V_err_mir_p.n8 V_err_mir_p.n7 5.063
R3760 V_err_mir_p.n16 V_err_mir_p.n15 4.5005
R3761 V_err_mir_p.n13 V_err_mir_p.n11 1.2505
R3762 V_err_mir_p.n15 V_err_mir_p.n13 1.2505
R3763 V_err_mir_p.n16 V_err_mir_p.n8 1.22272
R3764 V_err_mir_p.n5 V_err_mir_p.n3 0.563
R3765 V_err_mir_p.n7 V_err_mir_p.n5 0.563
R3766 V_b_2nd_stage.n4 V_b_2nd_stage.t7 525.38
R3767 V_b_2nd_stage.n0 V_b_2nd_stage.t2 525.38
R3768 V_b_2nd_stage.n6 V_b_2nd_stage.t4 366.856
R3769 V_b_2nd_stage.n2 V_b_2nd_stage.t5 366.856
R3770 V_b_2nd_stage.n4 V_b_2nd_stage.t3 281.168
R3771 V_b_2nd_stage.n5 V_b_2nd_stage.t8 281.168
R3772 V_b_2nd_stage.n0 V_b_2nd_stage.t6 281.168
R3773 V_b_2nd_stage.n1 V_b_2nd_stage.t9 281.168
R3774 V_b_2nd_stage.n5 V_b_2nd_stage.n4 244.214
R3775 V_b_2nd_stage.n1 V_b_2nd_stage.n0 244.214
R3776 V_b_2nd_stage.n7 V_b_2nd_stage.n6 166.03
R3777 V_b_2nd_stage.n3 V_b_2nd_stage.n2 166.03
R3778 V_b_2nd_stage.t0 V_b_2nd_stage.n7 117.974
R3779 V_b_2nd_stage.n3 V_b_2nd_stage.t1 117.849
R3780 V_b_2nd_stage.n6 V_b_2nd_stage.n5 85.6894
R3781 V_b_2nd_stage.n2 V_b_2nd_stage.n1 85.6894
R3782 V_b_2nd_stage.n7 V_b_2nd_stage.n3 36.813
R3783 VIN+.n9 VIN+.t9 485.127
R3784 VIN+.n4 VIN+.t5 485.127
R3785 VIN+.n3 VIN+.t0 485.127
R3786 VIN+.n7 VIN+.t2 318.656
R3787 VIN+.n7 VIN+.t7 318.656
R3788 VIN+.n5 VIN+.t1 318.656
R3789 VIN+.n5 VIN+.t6 318.656
R3790 VIN+.n1 VIN+.t4 318.656
R3791 VIN+.n1 VIN+.t10 318.656
R3792 VIN+.n0 VIN+.t3 318.656
R3793 VIN+.n0 VIN+.t8 318.656
R3794 VIN+.n2 VIN+.n0 167.05
R3795 VIN+.n8 VIN+.n7 165.8
R3796 VIN+.n6 VIN+.n5 165.8
R3797 VIN+.n2 VIN+.n1 165.8
R3798 VIN+.n6 VIN+.n4 2.34425
R3799 VIN+.n4 VIN+.n3 1.3005
R3800 VIN+.n8 VIN+.n6 1.2505
R3801 VIN+.n3 VIN+.n2 1.15675
R3802 VIN+.n9 VIN+.n8 1.15675
R3803 VIN+ VIN+.n9 0.963
R3804 V_p_mir.n1 V_p_mir.n0 219.99
R3805 V_p_mir.n0 V_p_mir.t0 16.0005
R3806 V_p_mir.n0 V_p_mir.t3 16.0005
R3807 V_p_mir.n1 V_p_mir.t1 9.6005
R3808 V_p_mir.t2 V_p_mir.n1 9.6005
R3809 a_109420_966.t0 a_109420_966.t1 169.905
R3810 a_109020_3958.t0 a_109020_3958.t1 169.905
R3811 a_117950_966.t0 a_117950_966.t1 169.905
R3812 a_118270_3958.t0 a_118270_3958.t1 294.339
R3813 a_118390_3958.t0 a_118390_3958.t1 169.905
R3814 a_108900_3958.t0 a_108900_3958.t1 294.339
C0 X V_CMFB_S1 0.624653f
C1 a_109990_5430# VOUT+ 0.054387f
C2 cap_res_Y VOUT- 0.028842f
C3 V_err_gate V_err_amp_ref 1.2227f
C4 V_CMFB_S4 V_CMFB_S3 1.24433f
C5 a_111200_5430# VDDA 0.087006f
C6 X VIN- 0.012706f
C7 V_CMFB_S2 X 0.711653f
C8 V_tail_gate Vb1 0.018702f
C9 Vb2 V_err_gate 0.031005f
C10 a_116370_5430# X 0.0255f
C11 VOUT+ VDDA 5.80669f
C12 err_amp_out VDDA 0.208638f
C13 Vb2_Vb3 VDDA 0.870514f
C14 VIN- Vb1 0.034729f
C15 VD1 X 0.986893f
C16 X VDDA 4.25983f
C17 VOUT+ VOUT- 0.305434f
C18 V_err_amp_ref VDDA 0.60945f
C19 V_CMFB_S3 VDDA 0.170191f
C20 Vb2_Vb3 VOUT- 0.026323f
C21 VD4 VDDA 3.82421f
C22 Vb3 VDDA 3.39276f
C23 VIN+ Vb1 0.011575f
C24 V_CMFB_S2 V_CMFB_S1 1.24433f
C25 V_tail_gate VIN- 0.230783f
C26 VD1 Vb1 0.27266f
C27 X VOUT- 2.15923f
C28 Vb1 VDDA 0.652968f
C29 Vb2 VDDA 1.24599f
C30 cap_res_Y VOUT+ 50.841f
C31 a_117580_5430# VDDA 0.086667f
C32 V_tail_gate VIN+ 0.107958f
C33 V_CMFB_S1 VDDA 0.169887f
C34 V_tail_gate VD1 0.21454f
C35 V_CMFB_S4 VDDA 2.21677f
C36 V_err_gate VDDA 1.34743f
C37 a_117580_5430# VOUT- 0.054387f
C38 VD4 cap_res_Y 0.037866f
C39 VIN- VIN+ 0.559567f
C40 Vb3 cap_res_Y 0.057312f
C41 VD1 VIN- 0.889f
C42 V_CMFB_S1 VOUT- 0.060463f
C43 a_111200_5430# VOUT+ 0.054329f
C44 a_109990_5430# VDDA 0.086666f
C45 V_CMFB_S2 VDDA 2.21711f
C46 cap_res_Y Vb1 0.016415f
C47 a_116370_5430# VDDA 0.087029f
C48 VD1 VIN+ 0.06006f
C49 a_116370_5430# VOUT- 0.054329f
C50 err_amp_out X 0.284856f
C51 V_CMFB_S3 VOUT+ 0.064245f
C52 err_amp_out V_err_amp_ref 0.596514f
C53 Vb2_Vb3 Vb3 0.717641f
C54 VOUT- VDDA 5.7703f
C55 Vb3 X 0.236637f
C56 VD4 Vb3 1.13534f
C57 Vb2_Vb3 Vb2 0.194352f
C58 X Vb1 0.837472f
C59 Vb1 V_err_amp_ref 0.011274f
C60 Vb2 X 1.09875f
C61 cap_res_Y VDDA 0.811299f
C62 a_117580_5430# X 0.015758f
C63 err_amp_out V_err_gate 0.105132f
C64 err_amp_out V_tail_gate 0.025573f
C65 VD4 Vb2 1.23863f
C66 Vb3 Vb2 1.95154f
C67 V_CMFB_S2 GNDA 1.017056f
C68 V_tail_gate GNDA 3.47641f
C69 VIN+ GNDA 2.019015f
C70 VIN- GNDA 1.933225f
C71 V_CMFB_S4 GNDA 1.019446f
C72 V_CMFB_S1 GNDA 2.42512f
C73 Vb1 GNDA 5.94722f
C74 V_CMFB_S3 GNDA 2.42066f
C75 VOUT- GNDA 17.95247f
C76 V_err_amp_ref GNDA 1.14478f
C77 VOUT+ GNDA 17.94547f
C78 V_err_gate GNDA 1.97686f
C79 Vb2 GNDA 2.72127f
C80 Vb3 GNDA 3.364983f
C81 VDDA GNDA 55.78524f
C82 m2_115460_3030# GNDA 0.054912f $ **FLOATING
C83 VD1 GNDA 2.58595f
C84 err_amp_out GNDA 4.361154f
C85 cap_res_Y GNDA 33.860977f
C86 a_117580_5430# GNDA 0.035194f
C87 a_116370_5430# GNDA 0.034748f
C88 a_111200_5430# GNDA 0.034748f
C89 a_109990_5430# GNDA 0.035194f
C90 X GNDA 6.590617f
C91 VD4 GNDA 4.994748f
C92 Vb2_Vb3 GNDA 2.77375f
C93 VIN+.t8 GNDA 0.042153f
C94 VIN+.t3 GNDA 0.042153f
C95 VIN+.n0 GNDA 0.087115f
C96 VIN+.t10 GNDA 0.042153f
C97 VIN+.t4 GNDA 0.042153f
C98 VIN+.n1 GNDA 0.085908f
C99 VIN+.n2 GNDA 0.362773f
C100 VIN+.t0 GNDA 0.059304f
C101 VIN+.n3 GNDA 0.217138f
C102 VIN+.t5 GNDA 0.059304f
C103 VIN+.n4 GNDA 0.264788f
C104 VIN+.t6 GNDA 0.042153f
C105 VIN+.t1 GNDA 0.042153f
C106 VIN+.n5 GNDA 0.085908f
C107 VIN+.n6 GNDA 0.250437f
C108 VIN+.t7 GNDA 0.042153f
C109 VIN+.t2 GNDA 0.042153f
C110 VIN+.n7 GNDA 0.085908f
C111 VIN+.n8 GNDA 0.202639f
C112 VIN+.t9 GNDA 0.059304f
C113 VIN+.n9 GNDA 0.203261f
C114 V_b_2nd_stage.t1 GNDA 0.107702f
C115 V_b_2nd_stage.t9 GNDA 0.269049f
C116 V_b_2nd_stage.t6 GNDA 0.269049f
C117 V_b_2nd_stage.t2 GNDA 0.319319f
C118 V_b_2nd_stage.n0 GNDA 0.168662f
C119 V_b_2nd_stage.n1 GNDA 0.106742f
C120 V_b_2nd_stage.t5 GNDA 0.293365f
C121 V_b_2nd_stage.n2 GNDA 0.098647f
C122 V_b_2nd_stage.n3 GNDA 0.565881f
C123 V_b_2nd_stage.t4 GNDA 0.293365f
C124 V_b_2nd_stage.t8 GNDA 0.269049f
C125 V_b_2nd_stage.t3 GNDA 0.269049f
C126 V_b_2nd_stage.t7 GNDA 0.319319f
C127 V_b_2nd_stage.n4 GNDA 0.168662f
C128 V_b_2nd_stage.n5 GNDA 0.106742f
C129 V_b_2nd_stage.n6 GNDA 0.098647f
C130 V_b_2nd_stage.n7 GNDA 0.568835f
C131 V_b_2nd_stage.t0 GNDA 0.107918f
C132 VD2.t15 GNDA 0.013877f
C133 VD2.t16 GNDA 0.013877f
C134 VD2.t21 GNDA 0.013877f
C135 VD2.n0 GNDA 0.050131f
C136 VD2.t17 GNDA 0.013877f
C137 VD2.t12 GNDA 0.013877f
C138 VD2.n1 GNDA 0.04969f
C139 VD2.n2 GNDA 0.186051f
C140 VD2.t19 GNDA 0.013877f
C141 VD2.t14 GNDA 0.013877f
C142 VD2.n3 GNDA 0.04969f
C143 VD2.n4 GNDA 0.096484f
C144 VD2.t18 GNDA 0.013877f
C145 VD2.t13 GNDA 0.013877f
C146 VD2.n5 GNDA 0.04687f
C147 VD2.t3 GNDA 0.013877f
C148 VD2.t8 GNDA 0.013877f
C149 VD2.n6 GNDA 0.045463f
C150 VD2.t0 GNDA 0.013877f
C151 VD2.t7 GNDA 0.013877f
C152 VD2.n7 GNDA 0.048872f
C153 VD2.t2 GNDA 0.013877f
C154 VD2.t1 GNDA 0.013877f
C155 VD2.n8 GNDA 0.047884f
C156 VD2.n9 GNDA 0.193373f
C157 VD2.t9 GNDA 0.013877f
C158 VD2.t10 GNDA 0.013877f
C159 VD2.n10 GNDA 0.047884f
C160 VD2.n11 GNDA 0.140662f
C161 VD2.t5 GNDA 0.013877f
C162 VD2.t11 GNDA 0.013877f
C163 VD2.n12 GNDA 0.048872f
C164 VD2.t6 GNDA 0.013877f
C165 VD2.t4 GNDA 0.013877f
C166 VD2.n13 GNDA 0.047884f
C167 VD2.n14 GNDA 0.193373f
C168 VD2.n15 GNDA 0.083264f
C169 VD2.n16 GNDA 0.069533f
C170 VD2.n17 GNDA 0.081264f
C171 VD2.n18 GNDA 0.117321f
C172 VD2.n19 GNDA 0.050132f
C173 VD2.t20 GNDA 0.013877f
C174 V_tot.t2 GNDA 0.080458f
C175 V_tot.t1 GNDA 0.085707f
C176 V_tot.t3 GNDA 0.080458f
C177 V_tot.n0 GNDA 0.400236f
C178 V_tot.n1 GNDA 0.018935f
C179 V_tot.n2 GNDA 0.018591f
C180 V_tot.n3 GNDA 0.103225f
C181 V_tot.n4 GNDA 0.05423f
C182 V_tot.n5 GNDA 0.015822f
C183 V_tot.n6 GNDA 0.092524f
C184 V_tot.n7 GNDA 0.018591f
C185 V_tot.n8 GNDA 0.068227f
C186 V_tot.n9 GNDA 0.073631f
C187 V_tot.n10 GNDA 0.64879f
C188 V_tot.n11 GNDA 0.401534f
C189 V_tot.t0 GNDA 0.085717f
C190 V_CMFB_S4.t0 GNDA 0.156142f
C191 V_CMFB_S4.t9 GNDA 0.037623f
C192 V_CMFB_S4.t8 GNDA 0.037623f
C193 V_CMFB_S4.n0 GNDA 0.155586f
C194 V_CMFB_S4.t3 GNDA 0.037623f
C195 V_CMFB_S4.t7 GNDA 0.037623f
C196 V_CMFB_S4.n1 GNDA 0.154989f
C197 V_CMFB_S4.n2 GNDA 0.214892f
C198 V_CMFB_S4.t2 GNDA 0.037623f
C199 V_CMFB_S4.t6 GNDA 0.037623f
C200 V_CMFB_S4.n3 GNDA 0.154989f
C201 V_CMFB_S4.n4 GNDA 0.112134f
C202 V_CMFB_S4.t1 GNDA 0.037623f
C203 V_CMFB_S4.t5 GNDA 0.037623f
C204 V_CMFB_S4.n5 GNDA 0.154989f
C205 V_CMFB_S4.n6 GNDA 0.112134f
C206 V_CMFB_S4.t10 GNDA 0.037623f
C207 V_CMFB_S4.t4 GNDA 0.037623f
C208 V_CMFB_S4.n7 GNDA 0.154989f
C209 V_CMFB_S4.n8 GNDA 0.164859f
C210 V_CMFB_S4.n9 GNDA 0.283052f
C211 V_CMFB_S2.t0 GNDA 0.156142f
C212 V_CMFB_S2.n0 GNDA -0.163033f
C213 V_CMFB_S2.t6 GNDA 0.037623f
C214 V_CMFB_S2.t1 GNDA 0.037623f
C215 V_CMFB_S2.n1 GNDA 0.151358f
C216 V_CMFB_S2.n2 GNDA 0.24438f
C217 V_CMFB_S2.t10 GNDA 0.037623f
C218 V_CMFB_S2.t4 GNDA 0.037623f
C219 V_CMFB_S2.n3 GNDA 0.154989f
C220 V_CMFB_S2.n4 GNDA 0.137773f
C221 V_CMFB_S2.t7 GNDA 0.037623f
C222 V_CMFB_S2.t5 GNDA 0.037623f
C223 V_CMFB_S2.n5 GNDA 0.154989f
C224 V_CMFB_S2.n6 GNDA 0.112134f
C225 V_CMFB_S2.t8 GNDA 0.037623f
C226 V_CMFB_S2.t2 GNDA 0.037623f
C227 V_CMFB_S2.n7 GNDA 0.154989f
C228 V_CMFB_S2.n8 GNDA 0.112134f
C229 V_CMFB_S2.t9 GNDA 0.037623f
C230 V_CMFB_S2.t3 GNDA 0.037623f
C231 V_CMFB_S2.n9 GNDA 0.154989f
C232 V_CMFB_S2.n10 GNDA 0.164859f
C233 V_CMFB_S2.n11 GNDA 0.283052f
C234 err_amp_out.n0 GNDA 1.19233f
C235 err_amp_out.n1 GNDA 0.017541f
C236 err_amp_out.n2 GNDA 0.017349f
C237 err_amp_out.n3 GNDA 0.017349f
C238 err_amp_out.n4 GNDA 0.01937f
C239 err_amp_out.t12 GNDA 0.06858f
C240 err_amp_out.n5 GNDA 0.020693f
C241 err_amp_out.n6 GNDA 0.020693f
C242 err_amp_out.n7 GNDA 0.177079f
C243 cap_res_Y.t26 GNDA 0.343734f
C244 cap_res_Y.t136 GNDA 0.344881f
C245 cap_res_Y.t60 GNDA 0.185242f
C246 cap_res_Y.n0 GNDA 0.197802f
C247 cap_res_Y.t58 GNDA 0.343734f
C248 cap_res_Y.t31 GNDA 0.344881f
C249 cap_res_Y.t99 GNDA 0.185242f
C250 cap_res_Y.n1 GNDA 0.216311f
C251 cap_res_Y.t95 GNDA 0.343734f
C252 cap_res_Y.t59 GNDA 0.344881f
C253 cap_res_Y.t4 GNDA 0.185242f
C254 cap_res_Y.n2 GNDA 0.216311f
C255 cap_res_Y.t81 GNDA 0.343734f
C256 cap_res_Y.t113 GNDA 0.344881f
C257 cap_res_Y.t121 GNDA 0.185242f
C258 cap_res_Y.n3 GNDA 0.216311f
C259 cap_res_Y.t119 GNDA 0.343734f
C260 cap_res_Y.t13 GNDA 0.344881f
C261 cap_res_Y.t114 GNDA 0.36339f
C262 cap_res_Y.t9 GNDA 0.36339f
C263 cap_res_Y.t18 GNDA 0.185242f
C264 cap_res_Y.n4 GNDA 0.216311f
C265 cap_res_Y.t94 GNDA 0.343734f
C266 cap_res_Y.t107 GNDA 0.344881f
C267 cap_res_Y.t70 GNDA 0.36339f
C268 cap_res_Y.t102 GNDA 0.36339f
C269 cap_res_Y.t3 GNDA 0.185242f
C270 cap_res_Y.n5 GNDA 0.216311f
C271 cap_res_Y.t6 GNDA 0.344881f
C272 cap_res_Y.t104 GNDA 0.346131f
C273 cap_res_Y.t101 GNDA 0.344881f
C274 cap_res_Y.t61 GNDA 0.347585f
C275 cap_res_Y.t30 GNDA 0.378048f
C276 cap_res_Y.t84 GNDA 0.344881f
C277 cap_res_Y.t125 GNDA 0.346131f
C278 cap_res_Y.t97 GNDA 0.344881f
C279 cap_res_Y.t63 GNDA 0.346131f
C280 cap_res_Y.t47 GNDA 0.344881f
C281 cap_res_Y.t86 GNDA 0.346131f
C282 cap_res_Y.t65 GNDA 0.344881f
C283 cap_res_Y.t35 GNDA 0.346131f
C284 cap_res_Y.t90 GNDA 0.344881f
C285 cap_res_Y.t131 GNDA 0.346131f
C286 cap_res_Y.t106 GNDA 0.344881f
C287 cap_res_Y.t72 GNDA 0.346131f
C288 cap_res_Y.t134 GNDA 0.344881f
C289 cap_res_Y.t27 GNDA 0.346131f
C290 cap_res_Y.t8 GNDA 0.344881f
C291 cap_res_Y.t110 GNDA 0.346131f
C292 cap_res_Y.t92 GNDA 0.344881f
C293 cap_res_Y.t135 GNDA 0.346131f
C294 cap_res_Y.t111 GNDA 0.344881f
C295 cap_res_Y.t80 GNDA 0.346131f
C296 cap_res_Y.t138 GNDA 0.344881f
C297 cap_res_Y.t33 GNDA 0.346131f
C298 cap_res_Y.t10 GNDA 0.344881f
C299 cap_res_Y.t118 GNDA 0.346131f
C300 cap_res_Y.t37 GNDA 0.344881f
C301 cap_res_Y.t71 GNDA 0.346131f
C302 cap_res_Y.t48 GNDA 0.344881f
C303 cap_res_Y.t17 GNDA 0.346131f
C304 cap_res_Y.t75 GNDA 0.344881f
C305 cap_res_Y.t109 GNDA 0.346131f
C306 cap_res_Y.t91 GNDA 0.344881f
C307 cap_res_Y.t53 GNDA 0.346131f
C308 cap_res_Y.t42 GNDA 0.344881f
C309 cap_res_Y.t77 GNDA 0.346131f
C310 cap_res_Y.t54 GNDA 0.344881f
C311 cap_res_Y.t24 GNDA 0.346131f
C312 cap_res_Y.t82 GNDA 0.344881f
C313 cap_res_Y.t115 GNDA 0.346131f
C314 cap_res_Y.t93 GNDA 0.344881f
C315 cap_res_Y.t57 GNDA 0.346131f
C316 cap_res_Y.t124 GNDA 0.344881f
C317 cap_res_Y.t15 GNDA 0.346131f
C318 cap_res_Y.t2 GNDA 0.344881f
C319 cap_res_Y.t96 GNDA 0.346131f
C320 cap_res_Y.t85 GNDA 0.344881f
C321 cap_res_Y.t126 GNDA 0.346131f
C322 cap_res_Y.t98 GNDA 0.344881f
C323 cap_res_Y.t64 GNDA 0.346131f
C324 cap_res_Y.t130 GNDA 0.344881f
C325 cap_res_Y.t22 GNDA 0.346131f
C326 cap_res_Y.t5 GNDA 0.344881f
C327 cap_res_Y.t105 GNDA 0.346131f
C328 cap_res_Y.t40 GNDA 0.344881f
C329 cap_res_Y.t133 GNDA 0.346131f
C330 cap_res_Y.t69 GNDA 0.344881f
C331 cap_res_Y.t122 GNDA 0.346131f
C332 cap_res_Y.t88 GNDA 0.344881f
C333 cap_res_Y.t76 GNDA 0.36179f
C334 cap_res_Y.t128 GNDA 0.344881f
C335 cap_res_Y.t29 GNDA 0.185242f
C336 cap_res_Y.n6 GNDA 0.198255f
C337 cap_res_Y.t19 GNDA 0.344881f
C338 cap_res_Y.t120 GNDA 0.185242f
C339 cap_res_Y.n7 GNDA 0.196656f
C340 cap_res_Y.t68 GNDA 0.344881f
C341 cap_res_Y.t103 GNDA 0.185242f
C342 cap_res_Y.n8 GNDA 0.196656f
C343 cap_res_Y.t100 GNDA 0.344881f
C344 cap_res_Y.t55 GNDA 0.185242f
C345 cap_res_Y.n9 GNDA 0.196656f
C346 cap_res_Y.t56 GNDA 0.344881f
C347 cap_res_Y.t52 GNDA 0.185242f
C348 cap_res_Y.n10 GNDA 0.196656f
C349 cap_res_Y.t108 GNDA 0.344881f
C350 cap_res_Y.t44 GNDA 0.185242f
C351 cap_res_Y.n11 GNDA 0.196656f
C352 cap_res_Y.t7 GNDA 0.344881f
C353 cap_res_Y.t137 GNDA 0.185242f
C354 cap_res_Y.n12 GNDA 0.196656f
C355 cap_res_Y.t41 GNDA 0.344881f
C356 cap_res_Y.t87 GNDA 0.185242f
C357 cap_res_Y.n13 GNDA 0.196656f
C358 cap_res_Y.t74 GNDA 0.344881f
C359 cap_res_Y.t39 GNDA 0.185242f
C360 cap_res_Y.n14 GNDA 0.196656f
C361 cap_res_Y.t67 GNDA 0.344881f
C362 cap_res_Y.t117 GNDA 0.346131f
C363 cap_res_Y.t51 GNDA 0.344881f
C364 cap_res_Y.t21 GNDA 0.346131f
C365 cap_res_Y.t129 GNDA 0.166734f
C366 cap_res_Y.n15 GNDA 0.215061f
C367 cap_res_Y.t25 GNDA 0.184096f
C368 cap_res_Y.n16 GNDA 0.23357f
C369 cap_res_Y.t32 GNDA 0.184096f
C370 cap_res_Y.n17 GNDA 0.250829f
C371 cap_res_Y.t73 GNDA 0.184096f
C372 cap_res_Y.n18 GNDA 0.250829f
C373 cap_res_Y.t36 GNDA 0.184096f
C374 cap_res_Y.n19 GNDA 0.250829f
C375 cap_res_Y.t62 GNDA 0.184096f
C376 cap_res_Y.n20 GNDA 0.250829f
C377 cap_res_Y.t28 GNDA 0.184096f
C378 cap_res_Y.n21 GNDA 0.250829f
C379 cap_res_Y.t132 GNDA 0.184096f
C380 cap_res_Y.n22 GNDA 0.250829f
C381 cap_res_Y.t23 GNDA 0.184096f
C382 cap_res_Y.n23 GNDA 0.250829f
C383 cap_res_Y.t127 GNDA 0.184096f
C384 cap_res_Y.n24 GNDA 0.250829f
C385 cap_res_Y.t83 GNDA 0.184096f
C386 cap_res_Y.n25 GNDA 0.250829f
C387 cap_res_Y.t43 GNDA 0.184096f
C388 cap_res_Y.n26 GNDA 0.250829f
C389 cap_res_Y.t79 GNDA 0.184096f
C390 cap_res_Y.n27 GNDA 0.250829f
C391 cap_res_Y.t38 GNDA 0.184096f
C392 cap_res_Y.n28 GNDA 0.250829f
C393 cap_res_Y.t1 GNDA 0.184096f
C394 cap_res_Y.n29 GNDA 0.250829f
C395 cap_res_Y.t34 GNDA 0.184096f
C396 cap_res_Y.n30 GNDA 0.250829f
C397 cap_res_Y.t66 GNDA 0.184096f
C398 cap_res_Y.n31 GNDA 0.23357f
C399 cap_res_Y.t45 GNDA 0.343734f
C400 cap_res_Y.t89 GNDA 0.166734f
C401 cap_res_Y.n32 GNDA 0.216311f
C402 cap_res_Y.t11 GNDA 0.343734f
C403 cap_res_Y.t49 GNDA 0.166734f
C404 cap_res_Y.n33 GNDA 0.216311f
C405 cap_res_Y.t112 GNDA 0.343734f
C406 cap_res_Y.t50 GNDA 0.344881f
C407 cap_res_Y.t16 GNDA 0.36339f
C408 cap_res_Y.t46 GNDA 0.36339f
C409 cap_res_Y.t12 GNDA 0.185242f
C410 cap_res_Y.n34 GNDA 0.216311f
C411 cap_res_Y.t78 GNDA 0.343734f
C412 cap_res_Y.n35 GNDA 0.216311f
C413 cap_res_Y.t116 GNDA 0.185242f
C414 cap_res_Y.t14 GNDA 0.36339f
C415 cap_res_Y.t123 GNDA 0.36339f
C416 cap_res_Y.t20 GNDA 0.434792f
C417 cap_res_Y.t0 GNDA 0.291879f
C418 VOUT+.t3 GNDA 0.043062f
C419 VOUT+.t4 GNDA 0.043062f
C420 VOUT+.n0 GNDA 0.173078f
C421 VOUT+.t9 GNDA 0.043062f
C422 VOUT+.t14 GNDA 0.043062f
C423 VOUT+.n1 GNDA 0.173078f
C424 VOUT+.t10 GNDA 0.043062f
C425 VOUT+.t5 GNDA 0.043062f
C426 VOUT+.n2 GNDA 0.17276f
C427 VOUT+.n3 GNDA 0.170189f
C428 VOUT+.t11 GNDA 0.043062f
C429 VOUT+.t6 GNDA 0.043062f
C430 VOUT+.n4 GNDA 0.17276f
C431 VOUT+.n5 GNDA 0.087765f
C432 VOUT+.t12 GNDA 0.043062f
C433 VOUT+.t7 GNDA 0.043062f
C434 VOUT+.n6 GNDA 0.17276f
C435 VOUT+.n7 GNDA 0.087765f
C436 VOUT+.n8 GNDA 0.103954f
C437 VOUT+.t13 GNDA 0.043062f
C438 VOUT+.t8 GNDA 0.043062f
C439 VOUT+.n9 GNDA 0.170645f
C440 VOUT+.n10 GNDA 0.211034f
C441 VOUT+.t28 GNDA 0.28708f
C442 VOUT+.t106 GNDA 0.29197f
C443 VOUT+.t136 GNDA 0.28708f
C444 VOUT+.n11 GNDA 0.192478f
C445 VOUT+.n12 GNDA 0.125597f
C446 VOUT+.t83 GNDA 0.291357f
C447 VOUT+.t116 GNDA 0.291357f
C448 VOUT+.t150 GNDA 0.291357f
C449 VOUT+.t49 GNDA 0.291357f
C450 VOUT+.t101 GNDA 0.291357f
C451 VOUT+.t57 GNDA 0.291357f
C452 VOUT+.t89 GNDA 0.291357f
C453 VOUT+.t138 GNDA 0.291357f
C454 VOUT+.t29 GNDA 0.291357f
C455 VOUT+.t69 GNDA 0.291357f
C456 VOUT+.t81 GNDA 0.28708f
C457 VOUT+.n13 GNDA 0.19309f
C458 VOUT+.t128 GNDA 0.28708f
C459 VOUT+.n14 GNDA 0.246917f
C460 VOUT+.t37 GNDA 0.28708f
C461 VOUT+.n15 GNDA 0.246917f
C462 VOUT+.t54 GNDA 0.28708f
C463 VOUT+.n16 GNDA 0.246917f
C464 VOUT+.t102 GNDA 0.28708f
C465 VOUT+.n17 GNDA 0.246917f
C466 VOUT+.t105 GNDA 0.28708f
C467 VOUT+.n18 GNDA 0.246917f
C468 VOUT+.t113 GNDA 0.28708f
C469 VOUT+.n19 GNDA 0.246917f
C470 VOUT+.t20 GNDA 0.28708f
C471 VOUT+.n20 GNDA 0.246917f
C472 VOUT+.t70 GNDA 0.28708f
C473 VOUT+.n21 GNDA 0.246917f
C474 VOUT+.t118 GNDA 0.28708f
C475 VOUT+.n22 GNDA 0.246917f
C476 VOUT+.t132 GNDA 0.28708f
C477 VOUT+.t90 GNDA 0.29197f
C478 VOUT+.t40 GNDA 0.28708f
C479 VOUT+.n23 GNDA 0.192478f
C480 VOUT+.n24 GNDA 0.233252f
C481 VOUT+.t117 GNDA 0.29197f
C482 VOUT+.t24 GNDA 0.28708f
C483 VOUT+.n25 GNDA 0.192478f
C484 VOUT+.t125 GNDA 0.28708f
C485 VOUT+.t88 GNDA 0.29197f
C486 VOUT+.t35 GNDA 0.28708f
C487 VOUT+.n26 GNDA 0.192478f
C488 VOUT+.n27 GNDA 0.233252f
C489 VOUT+.t27 GNDA 0.29197f
C490 VOUT+.t135 GNDA 0.28708f
C491 VOUT+.n28 GNDA 0.192478f
C492 VOUT+.t84 GNDA 0.28708f
C493 VOUT+.t152 GNDA 0.29197f
C494 VOUT+.t52 GNDA 0.28708f
C495 VOUT+.n29 GNDA 0.192478f
C496 VOUT+.n30 GNDA 0.233252f
C497 VOUT+.t72 GNDA 0.29197f
C498 VOUT+.t31 GNDA 0.28708f
C499 VOUT+.n31 GNDA 0.192478f
C500 VOUT+.t121 GNDA 0.28708f
C501 VOUT+.t59 GNDA 0.29197f
C502 VOUT+.t93 GNDA 0.28708f
C503 VOUT+.n32 GNDA 0.192478f
C504 VOUT+.n33 GNDA 0.233252f
C505 VOUT+.t33 GNDA 0.29197f
C506 VOUT+.t142 GNDA 0.28708f
C507 VOUT+.n34 GNDA 0.192478f
C508 VOUT+.t95 GNDA 0.28708f
C509 VOUT+.t155 GNDA 0.29197f
C510 VOUT+.t61 GNDA 0.28708f
C511 VOUT+.n35 GNDA 0.192478f
C512 VOUT+.n36 GNDA 0.233252f
C513 VOUT+.t127 GNDA 0.28708f
C514 VOUT+.t56 GNDA 0.29197f
C515 VOUT+.t96 GNDA 0.28708f
C516 VOUT+.n37 GNDA 0.192478f
C517 VOUT+.n38 GNDA 0.125597f
C518 VOUT+.t112 GNDA 0.291357f
C519 VOUT+.t146 GNDA 0.291357f
C520 VOUT+.t107 GNDA 0.29197f
C521 VOUT+.t141 GNDA 0.28708f
C522 VOUT+.n39 GNDA 0.192478f
C523 VOUT+.t111 GNDA 0.28708f
C524 VOUT+.n40 GNDA 0.121112f
C525 VOUT+.t45 GNDA 0.291357f
C526 VOUT+.t137 GNDA 0.29197f
C527 VOUT+.t34 GNDA 0.28708f
C528 VOUT+.n41 GNDA 0.192478f
C529 VOUT+.t143 GNDA 0.28708f
C530 VOUT+.n42 GNDA 0.121112f
C531 VOUT+.t79 GNDA 0.291357f
C532 VOUT+.t50 GNDA 0.29197f
C533 VOUT+.t87 GNDA 0.28708f
C534 VOUT+.n43 GNDA 0.192478f
C535 VOUT+.t55 GNDA 0.28708f
C536 VOUT+.n44 GNDA 0.121112f
C537 VOUT+.t63 GNDA 0.291357f
C538 VOUT+.t144 GNDA 0.29197f
C539 VOUT+.t43 GNDA 0.28708f
C540 VOUT+.n45 GNDA 0.192478f
C541 VOUT+.t148 GNDA 0.28708f
C542 VOUT+.n46 GNDA 0.121112f
C543 VOUT+.t38 GNDA 0.291357f
C544 VOUT+.t44 GNDA 0.291598f
C545 VOUT+.t76 GNDA 0.291357f
C546 VOUT+.t98 GNDA 0.291598f
C547 VOUT+.t62 GNDA 0.291357f
C548 VOUT+.t126 GNDA 0.291598f
C549 VOUT+.t99 GNDA 0.291357f
C550 VOUT+.t21 GNDA 0.291598f
C551 VOUT+.t131 GNDA 0.291357f
C552 VOUT+.t97 GNDA 0.28708f
C553 VOUT+.n47 GNDA 0.317758f
C554 VOUT+.t58 GNDA 0.28708f
C555 VOUT+.n48 GNDA 0.371586f
C556 VOUT+.t153 GNDA 0.28708f
C557 VOUT+.n49 GNDA 0.371586f
C558 VOUT+.t36 GNDA 0.28708f
C559 VOUT+.n50 GNDA 0.371586f
C560 VOUT+.t139 GNDA 0.28708f
C561 VOUT+.n51 GNDA 0.305231f
C562 VOUT+.t154 GNDA 0.28708f
C563 VOUT+.n52 GNDA 0.305231f
C564 VOUT+.t41 GNDA 0.28708f
C565 VOUT+.n53 GNDA 0.305231f
C566 VOUT+.t145 GNDA 0.28708f
C567 VOUT+.n54 GNDA 0.305231f
C568 VOUT+.t108 GNDA 0.28708f
C569 VOUT+.n55 GNDA 0.246917f
C570 VOUT+.t68 GNDA 0.28708f
C571 VOUT+.n56 GNDA 0.246917f
C572 VOUT+.t91 GNDA 0.28708f
C573 VOUT+.t151 GNDA 0.29197f
C574 VOUT+.t53 GNDA 0.28708f
C575 VOUT+.n57 GNDA 0.192478f
C576 VOUT+.n58 GNDA 0.233252f
C577 VOUT+.t73 GNDA 0.29197f
C578 VOUT+.t32 GNDA 0.28708f
C579 VOUT+.n59 GNDA 0.192478f
C580 VOUT+.t123 GNDA 0.28708f
C581 VOUT+.t60 GNDA 0.29197f
C582 VOUT+.t94 GNDA 0.28708f
C583 VOUT+.n60 GNDA 0.192478f
C584 VOUT+.n61 GNDA 0.233252f
C585 VOUT+.t110 GNDA 0.29197f
C586 VOUT+.t71 GNDA 0.28708f
C587 VOUT+.n62 GNDA 0.192478f
C588 VOUT+.t156 GNDA 0.28708f
C589 VOUT+.t92 GNDA 0.29197f
C590 VOUT+.t122 GNDA 0.28708f
C591 VOUT+.n63 GNDA 0.192478f
C592 VOUT+.n64 GNDA 0.233252f
C593 VOUT+.t67 GNDA 0.29197f
C594 VOUT+.t26 GNDA 0.28708f
C595 VOUT+.n65 GNDA 0.192478f
C596 VOUT+.t119 GNDA 0.28708f
C597 VOUT+.t51 GNDA 0.29197f
C598 VOUT+.t85 GNDA 0.28708f
C599 VOUT+.n66 GNDA 0.192478f
C600 VOUT+.n67 GNDA 0.233252f
C601 VOUT+.t23 GNDA 0.29197f
C602 VOUT+.t130 GNDA 0.28708f
C603 VOUT+.n68 GNDA 0.192478f
C604 VOUT+.t78 GNDA 0.28708f
C605 VOUT+.t149 GNDA 0.29197f
C606 VOUT+.t47 GNDA 0.28708f
C607 VOUT+.n69 GNDA 0.192478f
C608 VOUT+.n70 GNDA 0.233252f
C609 VOUT+.t65 GNDA 0.29197f
C610 VOUT+.t22 GNDA 0.28708f
C611 VOUT+.n71 GNDA 0.192478f
C612 VOUT+.t114 GNDA 0.28708f
C613 VOUT+.t46 GNDA 0.29197f
C614 VOUT+.t77 GNDA 0.28708f
C615 VOUT+.n72 GNDA 0.192478f
C616 VOUT+.n73 GNDA 0.233252f
C617 VOUT+.t19 GNDA 0.29197f
C618 VOUT+.t124 GNDA 0.28708f
C619 VOUT+.n74 GNDA 0.192478f
C620 VOUT+.t74 GNDA 0.28708f
C621 VOUT+.t147 GNDA 0.29197f
C622 VOUT+.t39 GNDA 0.28708f
C623 VOUT+.n75 GNDA 0.192478f
C624 VOUT+.n76 GNDA 0.233252f
C625 VOUT+.t120 GNDA 0.29197f
C626 VOUT+.t86 GNDA 0.28708f
C627 VOUT+.n77 GNDA 0.192478f
C628 VOUT+.t30 GNDA 0.28708f
C629 VOUT+.t109 GNDA 0.29197f
C630 VOUT+.t140 GNDA 0.28708f
C631 VOUT+.n78 GNDA 0.192478f
C632 VOUT+.n79 GNDA 0.233252f
C633 VOUT+.t82 GNDA 0.29197f
C634 VOUT+.t48 GNDA 0.28708f
C635 VOUT+.n80 GNDA 0.192478f
C636 VOUT+.t134 GNDA 0.28708f
C637 VOUT+.t66 GNDA 0.29197f
C638 VOUT+.t104 GNDA 0.28708f
C639 VOUT+.n81 GNDA 0.192478f
C640 VOUT+.n82 GNDA 0.233252f
C641 VOUT+.t115 GNDA 0.29197f
C642 VOUT+.t80 GNDA 0.28708f
C643 VOUT+.n83 GNDA 0.192478f
C644 VOUT+.t25 GNDA 0.28708f
C645 VOUT+.t103 GNDA 0.29197f
C646 VOUT+.t133 GNDA 0.28708f
C647 VOUT+.n84 GNDA 0.192478f
C648 VOUT+.n85 GNDA 0.233252f
C649 VOUT+.t64 GNDA 0.29197f
C650 VOUT+.t100 GNDA 0.28708f
C651 VOUT+.n86 GNDA 0.192478f
C652 VOUT+.t129 GNDA 0.28708f
C653 VOUT+.n87 GNDA 0.233252f
C654 VOUT+.t42 GNDA 0.28708f
C655 VOUT+.n88 GNDA 0.125597f
C656 VOUT+.t75 GNDA 0.28708f
C657 VOUT+.n89 GNDA 0.228298f
C658 VOUT+.n90 GNDA 0.245854f
C659 VOUT+.t16 GNDA 0.050239f
C660 VOUT+.t18 GNDA 0.050239f
C661 VOUT+.n91 GNDA 0.232408f
C662 VOUT+.t2 GNDA 0.050239f
C663 VOUT+.t0 GNDA 0.050239f
C664 VOUT+.n92 GNDA 0.23163f
C665 VOUT+.n93 GNDA 0.143136f
C666 VOUT+.t17 GNDA 0.050239f
C667 VOUT+.t15 GNDA 0.050239f
C668 VOUT+.n94 GNDA 0.23163f
C669 VOUT+.n95 GNDA 0.089541f
C670 VOUT+.t1 GNDA 0.083063f
C671 VOUT+.n96 GNDA 0.145316f
C672 VOUT+.n97 GNDA 0.067878f
C673 cap_res_X.t18 GNDA 0.344881f
C674 cap_res_X.t55 GNDA 0.346131f
C675 cap_res_X.t121 GNDA 0.344881f
C676 cap_res_X.t17 GNDA 0.347585f
C677 cap_res_X.t48 GNDA 0.378048f
C678 cap_res_X.t126 GNDA 0.344881f
C679 cap_res_X.t21 GNDA 0.346131f
C680 cap_res_X.t63 GNDA 0.344881f
C681 cap_res_X.t105 GNDA 0.346131f
C682 cap_res_X.t86 GNDA 0.344881f
C683 cap_res_X.t128 GNDA 0.346131f
C684 cap_res_X.t29 GNDA 0.344881f
C685 cap_res_X.t74 GNDA 0.346131f
C686 cap_res_X.t130 GNDA 0.344881f
C687 cap_res_X.t27 GNDA 0.346131f
C688 cap_res_X.t69 GNDA 0.344881f
C689 cap_res_X.t112 GNDA 0.346131f
C690 cap_res_X.t31 GNDA 0.344881f
C691 cap_res_X.t67 GNDA 0.346131f
C692 cap_res_X.t106 GNDA 0.344881f
C693 cap_res_X.t8 GNDA 0.346131f
C694 cap_res_X.t131 GNDA 0.344881f
C695 cap_res_X.t33 GNDA 0.346131f
C696 cap_res_X.t75 GNDA 0.344881f
C697 cap_res_X.t118 GNDA 0.346131f
C698 cap_res_X.t36 GNDA 0.344881f
C699 cap_res_X.t73 GNDA 0.346131f
C700 cap_res_X.t113 GNDA 0.344881f
C701 cap_res_X.t15 GNDA 0.346131f
C702 cap_res_X.t78 GNDA 0.344881f
C703 cap_res_X.t110 GNDA 0.346131f
C704 cap_res_X.t9 GNDA 0.344881f
C705 cap_res_X.t53 GNDA 0.346131f
C706 cap_res_X.t116 GNDA 0.344881f
C707 cap_res_X.t6 GNDA 0.346131f
C708 cap_res_X.t45 GNDA 0.344881f
C709 cap_res_X.t92 GNDA 0.346131f
C710 cap_res_X.t81 GNDA 0.344881f
C711 cap_res_X.t117 GNDA 0.346131f
C712 cap_res_X.t16 GNDA 0.344881f
C713 cap_res_X.t65 GNDA 0.346131f
C714 cap_res_X.t123 GNDA 0.344881f
C715 cap_res_X.t14 GNDA 0.346131f
C716 cap_res_X.t54 GNDA 0.344881f
C717 cap_res_X.t101 GNDA 0.346131f
C718 cap_res_X.t20 GNDA 0.344881f
C719 cap_res_X.t51 GNDA 0.346131f
C720 cap_res_X.t93 GNDA 0.344881f
C721 cap_res_X.t135 GNDA 0.346131f
C722 cap_res_X.t127 GNDA 0.344881f
C723 cap_res_X.t22 GNDA 0.346131f
C724 cap_res_X.t66 GNDA 0.344881f
C725 cap_res_X.t107 GNDA 0.346131f
C726 cap_res_X.t26 GNDA 0.344881f
C727 cap_res_X.t61 GNDA 0.346131f
C728 cap_res_X.t100 GNDA 0.344881f
C729 cap_res_X.t138 GNDA 0.346131f
C730 cap_res_X.t32 GNDA 0.344881f
C731 cap_res_X.t122 GNDA 0.346131f
C732 cap_res_X.t39 GNDA 0.344881f
C733 cap_res_X.t111 GNDA 0.346131f
C734 cap_res_X.t108 GNDA 0.344881f
C735 cap_res_X.t57 GNDA 0.346131f
C736 cap_res_X.t42 GNDA 0.344881f
C737 cap_res_X.t96 GNDA 0.361791f
C738 cap_res_X.t11 GNDA 0.344881f
C739 cap_res_X.t3 GNDA 0.185242f
C740 cap_res_X.n0 GNDA 0.198255f
C741 cap_res_X.t119 GNDA 0.344881f
C742 cap_res_X.t52 GNDA 0.185242f
C743 cap_res_X.n1 GNDA 0.196656f
C744 cap_res_X.t82 GNDA 0.344881f
C745 cap_res_X.t102 GNDA 0.185242f
C746 cap_res_X.n2 GNDA 0.196656f
C747 cap_res_X.t34 GNDA 0.344881f
C748 cap_res_X.t120 GNDA 0.185242f
C749 cap_res_X.n3 GNDA 0.196656f
C750 cap_res_X.t133 GNDA 0.344881f
C751 cap_res_X.t28 GNDA 0.185242f
C752 cap_res_X.n4 GNDA 0.196656f
C753 cap_res_X.t99 GNDA 0.344881f
C754 cap_res_X.t77 GNDA 0.185242f
C755 cap_res_X.n5 GNDA 0.196656f
C756 cap_res_X.t43 GNDA 0.344881f
C757 cap_res_X.t85 GNDA 0.185242f
C758 cap_res_X.n6 GNDA 0.196656f
C759 cap_res_X.t13 GNDA 0.344881f
C760 cap_res_X.t132 GNDA 0.185242f
C761 cap_res_X.n7 GNDA 0.196656f
C762 cap_res_X.t60 GNDA 0.344881f
C763 cap_res_X.t134 GNDA 0.185242f
C764 cap_res_X.n8 GNDA 0.196656f
C765 cap_res_X.t80 GNDA 0.344881f
C766 cap_res_X.t115 GNDA 0.346131f
C767 cap_res_X.t4 GNDA 0.166734f
C768 cap_res_X.n9 GNDA 0.215061f
C769 cap_res_X.t5 GNDA 0.184096f
C770 cap_res_X.n10 GNDA 0.23357f
C771 cap_res_X.t71 GNDA 0.184096f
C772 cap_res_X.n11 GNDA 0.250829f
C773 cap_res_X.t91 GNDA 0.184096f
C774 cap_res_X.n12 GNDA 0.250829f
C775 cap_res_X.t50 GNDA 0.184096f
C776 cap_res_X.n13 GNDA 0.250829f
C777 cap_res_X.t87 GNDA 0.184096f
C778 cap_res_X.n14 GNDA 0.250829f
C779 cap_res_X.t44 GNDA 0.184096f
C780 cap_res_X.n15 GNDA 0.250829f
C781 cap_res_X.t7 GNDA 0.184096f
C782 cap_res_X.n16 GNDA 0.250829f
C783 cap_res_X.t40 GNDA 0.184096f
C784 cap_res_X.n17 GNDA 0.250829f
C785 cap_res_X.t136 GNDA 0.184096f
C786 cap_res_X.n18 GNDA 0.250829f
C787 cap_res_X.t103 GNDA 0.184096f
C788 cap_res_X.n19 GNDA 0.250829f
C789 cap_res_X.t68 GNDA 0.184096f
C790 cap_res_X.n20 GNDA 0.250829f
C791 cap_res_X.t97 GNDA 0.184096f
C792 cap_res_X.n21 GNDA 0.250829f
C793 cap_res_X.t62 GNDA 0.184096f
C794 cap_res_X.n22 GNDA 0.250829f
C795 cap_res_X.t23 GNDA 0.184096f
C796 cap_res_X.n23 GNDA 0.250829f
C797 cap_res_X.t49 GNDA 0.184096f
C798 cap_res_X.n24 GNDA 0.250829f
C799 cap_res_X.t90 GNDA 0.184096f
C800 cap_res_X.n25 GNDA 0.23357f
C801 cap_res_X.t35 GNDA 0.343735f
C802 cap_res_X.t76 GNDA 0.166734f
C803 cap_res_X.n26 GNDA 0.216311f
C804 cap_res_X.t12 GNDA 0.343735f
C805 cap_res_X.t47 GNDA 0.166734f
C806 cap_res_X.n27 GNDA 0.216311f
C807 cap_res_X.t46 GNDA 0.343735f
C808 cap_res_X.t98 GNDA 0.344881f
C809 cap_res_X.t64 GNDA 0.36339f
C810 cap_res_X.t94 GNDA 0.36339f
C811 cap_res_X.t88 GNDA 0.185242f
C812 cap_res_X.n28 GNDA 0.216311f
C813 cap_res_X.t56 GNDA 0.343735f
C814 cap_res_X.t89 GNDA 0.344881f
C815 cap_res_X.t95 GNDA 0.185242f
C816 cap_res_X.n29 GNDA 0.197803f
C817 cap_res_X.t19 GNDA 0.343735f
C818 cap_res_X.t58 GNDA 0.344881f
C819 cap_res_X.t59 GNDA 0.185242f
C820 cap_res_X.n30 GNDA 0.216311f
C821 cap_res_X.t124 GNDA 0.343735f
C822 cap_res_X.t25 GNDA 0.344881f
C823 cap_res_X.t24 GNDA 0.185242f
C824 cap_res_X.n31 GNDA 0.216311f
C825 cap_res_X.t84 GNDA 0.343735f
C826 cap_res_X.t129 GNDA 0.344881f
C827 cap_res_X.t125 GNDA 0.185242f
C828 cap_res_X.n32 GNDA 0.216311f
C829 cap_res_X.t104 GNDA 0.343735f
C830 cap_res_X.t83 GNDA 0.344881f
C831 cap_res_X.t38 GNDA 0.36339f
C832 cap_res_X.t79 GNDA 0.36339f
C833 cap_res_X.t137 GNDA 0.185242f
C834 cap_res_X.n33 GNDA 0.216311f
C835 cap_res_X.t70 GNDA 0.343735f
C836 cap_res_X.t41 GNDA 0.344881f
C837 cap_res_X.t2 GNDA 0.36339f
C838 cap_res_X.t37 GNDA 0.36339f
C839 cap_res_X.t109 GNDA 0.185242f
C840 cap_res_X.n34 GNDA 0.216311f
C841 cap_res_X.t30 GNDA 0.343735f
C842 cap_res_X.n35 GNDA 0.216311f
C843 cap_res_X.t72 GNDA 0.185242f
C844 cap_res_X.t1 GNDA 0.36339f
C845 cap_res_X.t114 GNDA 0.36339f
C846 cap_res_X.t10 GNDA 0.736617f
C847 cap_res_X.t0 GNDA 0.297532f
C848 VOUT-.t5 GNDA 0.043062f
C849 VOUT-.t16 GNDA 0.043062f
C850 VOUT-.n0 GNDA 0.173079f
C851 VOUT-.t10 GNDA 0.043062f
C852 VOUT-.t15 GNDA 0.043062f
C853 VOUT-.n1 GNDA 0.17276f
C854 VOUT-.n2 GNDA 0.170188f
C855 VOUT-.t9 GNDA 0.043062f
C856 VOUT-.t14 GNDA 0.043062f
C857 VOUT-.n3 GNDA 0.17276f
C858 VOUT-.n4 GNDA 0.087765f
C859 VOUT-.t12 GNDA 0.043062f
C860 VOUT-.t7 GNDA 0.043062f
C861 VOUT-.n5 GNDA 0.17276f
C862 VOUT-.n6 GNDA 0.087765f
C863 VOUT-.t8 GNDA 0.043062f
C864 VOUT-.t4 GNDA 0.043062f
C865 VOUT-.n7 GNDA 0.173078f
C866 VOUT-.n8 GNDA 0.103954f
C867 VOUT-.t11 GNDA 0.043062f
C868 VOUT-.t13 GNDA 0.043062f
C869 VOUT-.n9 GNDA 0.170645f
C870 VOUT-.n10 GNDA 0.211034f
C871 VOUT-.t77 GNDA 0.29197f
C872 VOUT-.t42 GNDA 0.28708f
C873 VOUT-.n11 GNDA 0.192478f
C874 VOUT-.t153 GNDA 0.28708f
C875 VOUT-.n12 GNDA 0.125597f
C876 VOUT-.t49 GNDA 0.29197f
C877 VOUT-.t100 GNDA 0.28708f
C878 VOUT-.n13 GNDA 0.192478f
C879 VOUT-.t152 GNDA 0.28708f
C880 VOUT-.t97 GNDA 0.291357f
C881 VOUT-.t144 GNDA 0.291357f
C882 VOUT-.t114 GNDA 0.291357f
C883 VOUT-.t58 GNDA 0.291357f
C884 VOUT-.t24 GNDA 0.291357f
C885 VOUT-.t123 GNDA 0.291357f
C886 VOUT-.t75 GNDA 0.291357f
C887 VOUT-.t38 GNDA 0.291357f
C888 VOUT-.t146 GNDA 0.291357f
C889 VOUT-.t115 GNDA 0.291357f
C890 VOUT-.t61 GNDA 0.28708f
C891 VOUT-.n14 GNDA 0.19309f
C892 VOUT-.t154 GNDA 0.28708f
C893 VOUT-.n15 GNDA 0.246917f
C894 VOUT-.t105 GNDA 0.28708f
C895 VOUT-.n16 GNDA 0.246917f
C896 VOUT-.t55 GNDA 0.28708f
C897 VOUT-.n17 GNDA 0.246917f
C898 VOUT-.t37 GNDA 0.28708f
C899 VOUT-.n18 GNDA 0.246917f
C900 VOUT-.t129 GNDA 0.28708f
C901 VOUT-.n19 GNDA 0.246917f
C902 VOUT-.t80 GNDA 0.28708f
C903 VOUT-.n20 GNDA 0.246917f
C904 VOUT-.t72 GNDA 0.28708f
C905 VOUT-.n21 GNDA 0.246917f
C906 VOUT-.t25 GNDA 0.28708f
C907 VOUT-.n22 GNDA 0.246917f
C908 VOUT-.t23 GNDA 0.28708f
C909 VOUT-.n23 GNDA 0.246917f
C910 VOUT-.n24 GNDA 0.233252f
C911 VOUT-.t125 GNDA 0.29197f
C912 VOUT-.t35 GNDA 0.28708f
C913 VOUT-.n25 GNDA 0.192478f
C914 VOUT-.t86 GNDA 0.28708f
C915 VOUT-.t118 GNDA 0.29197f
C916 VOUT-.t46 GNDA 0.28708f
C917 VOUT-.n26 GNDA 0.192478f
C918 VOUT-.n27 GNDA 0.233252f
C919 VOUT-.t131 GNDA 0.29197f
C920 VOUT-.t96 GNDA 0.28708f
C921 VOUT-.n28 GNDA 0.192478f
C922 VOUT-.t66 GNDA 0.28708f
C923 VOUT-.t57 GNDA 0.29197f
C924 VOUT-.t19 GNDA 0.28708f
C925 VOUT-.n29 GNDA 0.192478f
C926 VOUT-.n30 GNDA 0.233252f
C927 VOUT-.t30 GNDA 0.29197f
C928 VOUT-.t135 GNDA 0.28708f
C929 VOUT-.n31 GNDA 0.192478f
C930 VOUT-.t107 GNDA 0.28708f
C931 VOUT-.t91 GNDA 0.29197f
C932 VOUT-.t50 GNDA 0.28708f
C933 VOUT-.n32 GNDA 0.192478f
C934 VOUT-.n33 GNDA 0.233252f
C935 VOUT-.t137 GNDA 0.29197f
C936 VOUT-.t106 GNDA 0.28708f
C937 VOUT-.n34 GNDA 0.192478f
C938 VOUT-.t70 GNDA 0.28708f
C939 VOUT-.t64 GNDA 0.29197f
C940 VOUT-.t22 GNDA 0.28708f
C941 VOUT-.n35 GNDA 0.192478f
C942 VOUT-.n36 GNDA 0.233252f
C943 VOUT-.t36 GNDA 0.29197f
C944 VOUT-.t140 GNDA 0.28708f
C945 VOUT-.n37 GNDA 0.192478f
C946 VOUT-.t109 GNDA 0.28708f
C947 VOUT-.n38 GNDA 0.125597f
C948 VOUT-.t139 GNDA 0.29197f
C949 VOUT-.t102 GNDA 0.28708f
C950 VOUT-.n39 GNDA 0.192478f
C951 VOUT-.t67 GNDA 0.28708f
C952 VOUT-.t122 GNDA 0.291357f
C953 VOUT-.t145 GNDA 0.291357f
C954 VOUT-.t59 GNDA 0.29197f
C955 VOUT-.t93 GNDA 0.28708f
C956 VOUT-.n40 GNDA 0.192478f
C957 VOUT-.t63 GNDA 0.28708f
C958 VOUT-.n41 GNDA 0.121112f
C959 VOUT-.t111 GNDA 0.291357f
C960 VOUT-.t147 GNDA 0.29197f
C961 VOUT-.t43 GNDA 0.28708f
C962 VOUT-.n42 GNDA 0.192478f
C963 VOUT-.t156 GNDA 0.28708f
C964 VOUT-.n43 GNDA 0.121112f
C965 VOUT-.t127 GNDA 0.291357f
C966 VOUT-.t116 GNDA 0.29197f
C967 VOUT-.t155 GNDA 0.28708f
C968 VOUT-.n44 GNDA 0.192478f
C969 VOUT-.t120 GNDA 0.28708f
C970 VOUT-.n45 GNDA 0.121112f
C971 VOUT-.t87 GNDA 0.291357f
C972 VOUT-.t74 GNDA 0.29197f
C973 VOUT-.t119 GNDA 0.28708f
C974 VOUT-.n46 GNDA 0.192478f
C975 VOUT-.t78 GNDA 0.28708f
C976 VOUT-.n47 GNDA 0.121112f
C977 VOUT-.t53 GNDA 0.291357f
C978 VOUT-.t28 GNDA 0.291598f
C979 VOUT-.t73 GNDA 0.291357f
C980 VOUT-.t132 GNDA 0.291598f
C981 VOUT-.t33 GNDA 0.291357f
C982 VOUT-.t99 GNDA 0.291598f
C983 VOUT-.t138 GNDA 0.291357f
C984 VOUT-.t68 GNDA 0.291598f
C985 VOUT-.t101 GNDA 0.291357f
C986 VOUT-.t62 GNDA 0.28708f
C987 VOUT-.n48 GNDA 0.317758f
C988 VOUT-.t98 GNDA 0.28708f
C989 VOUT-.n49 GNDA 0.371586f
C990 VOUT-.t133 GNDA 0.28708f
C991 VOUT-.n50 GNDA 0.371586f
C992 VOUT-.t32 GNDA 0.28708f
C993 VOUT-.n51 GNDA 0.371586f
C994 VOUT-.t20 GNDA 0.28708f
C995 VOUT-.n52 GNDA 0.305231f
C996 VOUT-.t48 GNDA 0.28708f
C997 VOUT-.n53 GNDA 0.305231f
C998 VOUT-.t85 GNDA 0.28708f
C999 VOUT-.n54 GNDA 0.305231f
C1000 VOUT-.t69 GNDA 0.28708f
C1001 VOUT-.n55 GNDA 0.305231f
C1002 VOUT-.t110 GNDA 0.28708f
C1003 VOUT-.n56 GNDA 0.246917f
C1004 VOUT-.t81 GNDA 0.28708f
C1005 VOUT-.n57 GNDA 0.246917f
C1006 VOUT-.n58 GNDA 0.233252f
C1007 VOUT-.t31 GNDA 0.29197f
C1008 VOUT-.t136 GNDA 0.28708f
C1009 VOUT-.n59 GNDA 0.192478f
C1010 VOUT-.t108 GNDA 0.28708f
C1011 VOUT-.t94 GNDA 0.29197f
C1012 VOUT-.t52 GNDA 0.28708f
C1013 VOUT-.n60 GNDA 0.192478f
C1014 VOUT-.n61 GNDA 0.233252f
C1015 VOUT-.t71 GNDA 0.29197f
C1016 VOUT-.t29 GNDA 0.28708f
C1017 VOUT-.n62 GNDA 0.192478f
C1018 VOUT-.t134 GNDA 0.28708f
C1019 VOUT-.t128 GNDA 0.29197f
C1020 VOUT-.t83 GNDA 0.28708f
C1021 VOUT-.n63 GNDA 0.192478f
C1022 VOUT-.n64 GNDA 0.233252f
C1023 VOUT-.t27 GNDA 0.29197f
C1024 VOUT-.t130 GNDA 0.28708f
C1025 VOUT-.n65 GNDA 0.192478f
C1026 VOUT-.t95 GNDA 0.28708f
C1027 VOUT-.t88 GNDA 0.29197f
C1028 VOUT-.t45 GNDA 0.28708f
C1029 VOUT-.n66 GNDA 0.192478f
C1030 VOUT-.n67 GNDA 0.233252f
C1031 VOUT-.t126 GNDA 0.29197f
C1032 VOUT-.t90 GNDA 0.28708f
C1033 VOUT-.n68 GNDA 0.192478f
C1034 VOUT-.t60 GNDA 0.28708f
C1035 VOUT-.t51 GNDA 0.29197f
C1036 VOUT-.t149 GNDA 0.28708f
C1037 VOUT-.n69 GNDA 0.192478f
C1038 VOUT-.n70 GNDA 0.233252f
C1039 VOUT-.t26 GNDA 0.29197f
C1040 VOUT-.t124 GNDA 0.28708f
C1041 VOUT-.n71 GNDA 0.192478f
C1042 VOUT-.t89 GNDA 0.28708f
C1043 VOUT-.t82 GNDA 0.29197f
C1044 VOUT-.t39 GNDA 0.28708f
C1045 VOUT-.n72 GNDA 0.192478f
C1046 VOUT-.n73 GNDA 0.233252f
C1047 VOUT-.t121 GNDA 0.29197f
C1048 VOUT-.t84 GNDA 0.28708f
C1049 VOUT-.n74 GNDA 0.192478f
C1050 VOUT-.t54 GNDA 0.28708f
C1051 VOUT-.t44 GNDA 0.29197f
C1052 VOUT-.t142 GNDA 0.28708f
C1053 VOUT-.n75 GNDA 0.192478f
C1054 VOUT-.n76 GNDA 0.233252f
C1055 VOUT-.t79 GNDA 0.29197f
C1056 VOUT-.t47 GNDA 0.28708f
C1057 VOUT-.n77 GNDA 0.192478f
C1058 VOUT-.t21 GNDA 0.28708f
C1059 VOUT-.t148 GNDA 0.29197f
C1060 VOUT-.t104 GNDA 0.28708f
C1061 VOUT-.n78 GNDA 0.192478f
C1062 VOUT-.n79 GNDA 0.233252f
C1063 VOUT-.t41 GNDA 0.29197f
C1064 VOUT-.t151 GNDA 0.28708f
C1065 VOUT-.n80 GNDA 0.192478f
C1066 VOUT-.t117 GNDA 0.28708f
C1067 VOUT-.t112 GNDA 0.29197f
C1068 VOUT-.t65 GNDA 0.28708f
C1069 VOUT-.n81 GNDA 0.192478f
C1070 VOUT-.n82 GNDA 0.233252f
C1071 VOUT-.t76 GNDA 0.29197f
C1072 VOUT-.t40 GNDA 0.28708f
C1073 VOUT-.n83 GNDA 0.192478f
C1074 VOUT-.t150 GNDA 0.28708f
C1075 VOUT-.t141 GNDA 0.29197f
C1076 VOUT-.t92 GNDA 0.28708f
C1077 VOUT-.n84 GNDA 0.192478f
C1078 VOUT-.n85 GNDA 0.233252f
C1079 VOUT-.t34 GNDA 0.29197f
C1080 VOUT-.t143 GNDA 0.28708f
C1081 VOUT-.n86 GNDA 0.192478f
C1082 VOUT-.t113 GNDA 0.28708f
C1083 VOUT-.n87 GNDA 0.233252f
C1084 VOUT-.t56 GNDA 0.28708f
C1085 VOUT-.n88 GNDA 0.125597f
C1086 VOUT-.t103 GNDA 0.28708f
C1087 VOUT-.n89 GNDA 0.228298f
C1088 VOUT-.n90 GNDA 0.245854f
C1089 VOUT-.t1 GNDA 0.050239f
C1090 VOUT-.t17 GNDA 0.050239f
C1091 VOUT-.n91 GNDA 0.232408f
C1092 VOUT-.t3 GNDA 0.050239f
C1093 VOUT-.t0 GNDA 0.050239f
C1094 VOUT-.n92 GNDA 0.23163f
C1095 VOUT-.n93 GNDA 0.143136f
C1096 VOUT-.t18 GNDA 0.050239f
C1097 VOUT-.t2 GNDA 0.050239f
C1098 VOUT-.n94 GNDA 0.23163f
C1099 VOUT-.n95 GNDA 0.088105f
C1100 VOUT-.t6 GNDA 0.083063f
C1101 VOUT-.n96 GNDA 0.145743f
C1102 VOUT-.n97 GNDA 0.068886f
C1103 X.t3 GNDA 0.021176f
C1104 X.t2 GNDA 0.021176f
C1105 X.n0 GNDA 0.071494f
C1106 X.t23 GNDA 0.021176f
C1107 X.t7 GNDA 0.021176f
C1108 X.n1 GNDA 0.076412f
C1109 X.t4 GNDA 0.021176f
C1110 X.t24 GNDA 0.021176f
C1111 X.n2 GNDA 0.076412f
C1112 X.t0 GNDA 0.021176f
C1113 X.t8 GNDA 0.021176f
C1114 X.n3 GNDA 0.075745f
C1115 X.n4 GNDA 0.281241f
C1116 X.t6 GNDA 0.021176f
C1117 X.t1 GNDA 0.021176f
C1118 X.n5 GNDA 0.075745f
C1119 X.n6 GNDA 0.145895f
C1120 X.t10 GNDA 0.021176f
C1121 X.t5 GNDA 0.021176f
C1122 X.n7 GNDA 0.075745f
C1123 X.n8 GNDA 0.145895f
C1124 X.n9 GNDA 0.177697f
C1125 X.n10 GNDA 0.143638f
C1126 X.t9 GNDA 0.676735f
C1127 X.t28 GNDA 0.093173f
C1128 X.t43 GNDA 0.093173f
C1129 X.t25 GNDA 0.099236f
C1130 X.n11 GNDA 0.07864f
C1131 X.n12 GNDA 0.04204f
C1132 X.t46 GNDA 0.093173f
C1133 X.t31 GNDA 0.093173f
C1134 X.t38 GNDA 0.093173f
C1135 X.t53 GNDA 0.093173f
C1136 X.t40 GNDA 0.093173f
C1137 X.t34 GNDA 0.093173f
C1138 X.t50 GNDA 0.099236f
C1139 X.n13 GNDA 0.07864f
C1140 X.n14 GNDA 0.044469f
C1141 X.n15 GNDA 0.044469f
C1142 X.n16 GNDA 0.044469f
C1143 X.n17 GNDA 0.044469f
C1144 X.n18 GNDA 0.04204f
C1145 X.n19 GNDA 0.022779f
C1146 X.n20 GNDA 0.753199f
C1147 X.t18 GNDA 0.04941f
C1148 X.t22 GNDA 0.04941f
C1149 X.n21 GNDA 0.171837f
C1150 X.t17 GNDA 0.04941f
C1151 X.t15 GNDA 0.04941f
C1152 X.n22 GNDA 0.171229f
C1153 X.n23 GNDA 0.323263f
C1154 X.t12 GNDA 0.04941f
C1155 X.t14 GNDA 0.04941f
C1156 X.n24 GNDA 0.171229f
C1157 X.n25 GNDA 0.167583f
C1158 X.t20 GNDA 0.04941f
C1159 X.t11 GNDA 0.04941f
C1160 X.n26 GNDA 0.171229f
C1161 X.n27 GNDA 0.167583f
C1162 X.t16 GNDA 0.04941f
C1163 X.t19 GNDA 0.04941f
C1164 X.n28 GNDA 0.171229f
C1165 X.n29 GNDA 0.197332f
C1166 X.t21 GNDA 0.04941f
C1167 X.t13 GNDA 0.04941f
C1168 X.n30 GNDA 0.167682f
C1169 X.n31 GNDA 0.334482f
C1170 X.t39 GNDA 0.029646f
C1171 X.t51 GNDA 0.029646f
C1172 X.t36 GNDA 0.029646f
C1173 X.t30 GNDA 0.029646f
C1174 X.t45 GNDA 0.029646f
C1175 X.t27 GNDA 0.029646f
C1176 X.t42 GNDA 0.029646f
C1177 X.t54 GNDA 0.035999f
C1178 X.n32 GNDA 0.035999f
C1179 X.n33 GNDA 0.023293f
C1180 X.n34 GNDA 0.023293f
C1181 X.n35 GNDA 0.023293f
C1182 X.n36 GNDA 0.023293f
C1183 X.n37 GNDA 0.023293f
C1184 X.n38 GNDA 0.020864f
C1185 X.t33 GNDA 0.029646f
C1186 X.t49 GNDA 0.035999f
C1187 X.n39 GNDA 0.033569f
C1188 X.n40 GNDA 0.02052f
C1189 X.t44 GNDA 0.045528f
C1190 X.t26 GNDA 0.045528f
C1191 X.t41 GNDA 0.045528f
C1192 X.t35 GNDA 0.045528f
C1193 X.t48 GNDA 0.045528f
C1194 X.t32 GNDA 0.045528f
C1195 X.t47 GNDA 0.045528f
C1196 X.t29 GNDA 0.051757f
C1197 X.n41 GNDA 0.04671f
C1198 X.n42 GNDA 0.028587f
C1199 X.n43 GNDA 0.028587f
C1200 X.n44 GNDA 0.028587f
C1201 X.n45 GNDA 0.028587f
C1202 X.n46 GNDA 0.028587f
C1203 X.n47 GNDA 0.026158f
C1204 X.t37 GNDA 0.045528f
C1205 X.t52 GNDA 0.051757f
C1206 X.n48 GNDA 0.04428f
C1207 X.n49 GNDA 0.020477f
C1208 X.n50 GNDA 0.220698f
C1209 X.n51 GNDA 0.459548f
C1210 X.n52 GNDA 0.214361f
C1211 X.n53 GNDA 0.091429f
C1212 VDDA.t199 GNDA 0.018811f
C1213 VDDA.t227 GNDA 0.018811f
C1214 VDDA.n0 GNDA 0.077794f
C1215 VDDA.t197 GNDA 0.018811f
C1216 VDDA.t219 GNDA 0.018811f
C1217 VDDA.n1 GNDA 0.077496f
C1218 VDDA.n2 GNDA 0.107444f
C1219 VDDA.t203 GNDA 0.018811f
C1220 VDDA.t182 GNDA 0.018811f
C1221 VDDA.n3 GNDA 0.077496f
C1222 VDDA.n4 GNDA 0.056066f
C1223 VDDA.t207 GNDA 0.018811f
C1224 VDDA.t188 GNDA 0.018811f
C1225 VDDA.n5 GNDA 0.077496f
C1226 VDDA.n6 GNDA 0.056066f
C1227 VDDA.t211 GNDA 0.018811f
C1228 VDDA.t187 GNDA 0.018811f
C1229 VDDA.n7 GNDA 0.077496f
C1230 VDDA.n8 GNDA 0.056066f
C1231 VDDA.t226 GNDA 0.018811f
C1232 VDDA.t218 GNDA 0.018811f
C1233 VDDA.n9 GNDA 0.077496f
C1234 VDDA.n10 GNDA 0.0976f
C1235 VDDA.n12 GNDA 0.012541f
C1236 VDDA.n15 GNDA 0.012541f
C1237 VDDA.n16 GNDA 0.021947f
C1238 VDDA.t125 GNDA 0.018905f
C1239 VDDA.n17 GNDA 0.047345f
C1240 VDDA.n18 GNDA 0.012541f
C1241 VDDA.n19 GNDA 0.021947f
C1242 VDDA.t127 GNDA 0.033064f
C1243 VDDA.n21 GNDA 0.030535f
C1244 VDDA.n22 GNDA 0.010308f
C1245 VDDA.n23 GNDA 0.110988f
C1246 VDDA.t126 GNDA 0.092176f
C1247 VDDA.t202 GNDA 0.082771f
C1248 VDDA.t190 GNDA 0.082771f
C1249 VDDA.t206 GNDA 0.082771f
C1250 VDDA.t191 GNDA 0.082771f
C1251 VDDA.t210 GNDA 0.082771f
C1252 VDDA.t194 GNDA 0.082771f
C1253 VDDA.t214 GNDA 0.082771f
C1254 VDDA.t198 GNDA 0.082771f
C1255 VDDA.t217 GNDA 0.082771f
C1256 VDDA.t189 GNDA 0.082771f
C1257 VDDA.t178 GNDA 0.092176f
C1258 VDDA.n24 GNDA 0.012541f
C1259 VDDA.t179 GNDA 0.033064f
C1260 VDDA.n25 GNDA 0.021947f
C1261 VDDA.n26 GNDA 0.021947f
C1262 VDDA.n27 GNDA 0.027645f
C1263 VDDA.n28 GNDA 0.013198f
C1264 VDDA.n29 GNDA 0.110988f
C1265 VDDA.n30 GNDA 0.012541f
C1266 VDDA.n31 GNDA 0.025626f
C1267 VDDA.t177 GNDA 0.018228f
C1268 VDDA.n32 GNDA 0.036672f
C1269 VDDA.n33 GNDA 0.14674f
C1270 VDDA.t148 GNDA 0.011424f
C1271 VDDA.n34 GNDA 0.026145f
C1272 VDDA.t145 GNDA 0.011424f
C1273 VDDA.n35 GNDA 0.051619f
C1274 VDDA.t144 GNDA 0.04695f
C1275 VDDA.t27 GNDA 0.031039f
C1276 VDDA.t21 GNDA 0.031039f
C1277 VDDA.t71 GNDA 0.031039f
C1278 VDDA.t74 GNDA 0.031039f
C1279 VDDA.t19 GNDA 0.031039f
C1280 VDDA.t28 GNDA 0.031039f
C1281 VDDA.t80 GNDA 0.031039f
C1282 VDDA.t48 GNDA 0.031039f
C1283 VDDA.t73 GNDA 0.031039f
C1284 VDDA.t20 GNDA 0.031039f
C1285 VDDA.t147 GNDA 0.046649f
C1286 VDDA.n36 GNDA 0.044224f
C1287 VDDA.n37 GNDA 0.12013f
C1288 VDDA.t184 GNDA 0.037623f
C1289 VDDA.t216 GNDA 0.037623f
C1290 VDDA.n38 GNDA 0.150938f
C1291 VDDA.n39 GNDA 0.076681f
C1292 VDDA.n41 GNDA 0.012541f
C1293 VDDA.n46 GNDA 0.013198f
C1294 VDDA.n52 GNDA 0.013198f
C1295 VDDA.n53 GNDA 0.012541f
C1296 VDDA.t196 GNDA 0.037623f
C1297 VDDA.t213 GNDA 0.037623f
C1298 VDDA.n54 GNDA 0.150938f
C1299 VDDA.n55 GNDA 0.076681f
C1300 VDDA.t193 GNDA 0.037623f
C1301 VDDA.t209 GNDA 0.037623f
C1302 VDDA.n56 GNDA 0.150938f
C1303 VDDA.n57 GNDA 0.076681f
C1304 VDDA.t181 GNDA 0.037623f
C1305 VDDA.t205 GNDA 0.037623f
C1306 VDDA.n58 GNDA 0.150938f
C1307 VDDA.n59 GNDA 0.076681f
C1308 VDDA.t186 GNDA 0.037623f
C1309 VDDA.t201 GNDA 0.037623f
C1310 VDDA.n60 GNDA 0.150938f
C1311 VDDA.n61 GNDA 0.106392f
C1312 VDDA.n62 GNDA 0.021947f
C1313 VDDA.n63 GNDA 0.012541f
C1314 VDDA.n64 GNDA 0.012541f
C1315 VDDA.n67 GNDA 0.012541f
C1316 VDDA.n68 GNDA 0.012541f
C1317 VDDA.n69 GNDA 0.024951f
C1318 VDDA.n70 GNDA 0.031767f
C1319 VDDA.n71 GNDA 0.012541f
C1320 VDDA.n72 GNDA 0.021947f
C1321 VDDA.n73 GNDA 0.021947f
C1322 VDDA.n74 GNDA 0.012541f
C1323 VDDA.n75 GNDA 0.012541f
C1324 VDDA.n76 GNDA 0.021947f
C1325 VDDA.n77 GNDA 0.021947f
C1326 VDDA.n78 GNDA 0.012541f
C1327 VDDA.n79 GNDA 0.012541f
C1328 VDDA.n80 GNDA 0.021947f
C1329 VDDA.n81 GNDA 0.021947f
C1330 VDDA.n82 GNDA 0.012541f
C1331 VDDA.n83 GNDA 0.012541f
C1332 VDDA.n84 GNDA 0.021947f
C1333 VDDA.n85 GNDA 0.021947f
C1334 VDDA.n86 GNDA 0.012541f
C1335 VDDA.n87 GNDA 0.012541f
C1336 VDDA.n88 GNDA 0.021947f
C1337 VDDA.n89 GNDA 0.024951f
C1338 VDDA.n91 GNDA 0.030752f
C1339 VDDA.n92 GNDA 0.012541f
C1340 VDDA.n93 GNDA 0.295967f
C1341 VDDA.t220 GNDA 0.245803f
C1342 VDDA.t200 GNDA 0.220721f
C1343 VDDA.t185 GNDA 0.220721f
C1344 VDDA.t204 GNDA 0.220721f
C1345 VDDA.t180 GNDA 0.220721f
C1346 VDDA.t208 GNDA 0.220721f
C1347 VDDA.t192 GNDA 0.220721f
C1348 VDDA.t212 GNDA 0.220721f
C1349 VDDA.t195 GNDA 0.220721f
C1350 VDDA.t215 GNDA 0.220721f
C1351 VDDA.t183 GNDA 0.220721f
C1352 VDDA.t81 GNDA 0.245803f
C1353 VDDA.n94 GNDA 0.012541f
C1354 VDDA.n95 GNDA 0.021947f
C1355 VDDA.n96 GNDA 0.024951f
C1356 VDDA.n97 GNDA 0.012541f
C1357 VDDA.n98 GNDA 0.012541f
C1358 VDDA.n101 GNDA 0.012541f
C1359 VDDA.n102 GNDA 0.012541f
C1360 VDDA.n103 GNDA 0.024951f
C1361 VDDA.n104 GNDA 0.031767f
C1362 VDDA.n105 GNDA 0.012541f
C1363 VDDA.n106 GNDA 0.021947f
C1364 VDDA.n107 GNDA 0.021947f
C1365 VDDA.n108 GNDA 0.012541f
C1366 VDDA.n109 GNDA 0.012541f
C1367 VDDA.n110 GNDA 0.021947f
C1368 VDDA.n111 GNDA 0.021947f
C1369 VDDA.n112 GNDA 0.012541f
C1370 VDDA.n113 GNDA 0.012541f
C1371 VDDA.n114 GNDA 0.021947f
C1372 VDDA.n115 GNDA 0.021947f
C1373 VDDA.n116 GNDA 0.012541f
C1374 VDDA.n117 GNDA 0.012541f
C1375 VDDA.n118 GNDA 0.021947f
C1376 VDDA.n119 GNDA 0.021947f
C1377 VDDA.n120 GNDA 0.021947f
C1378 VDDA.n121 GNDA 0.012541f
C1379 VDDA.n122 GNDA 0.295967f
C1380 VDDA.n124 GNDA 0.033104f
C1381 VDDA.n125 GNDA 0.053368f
C1382 VDDA.n126 GNDA 0.091863f
C1383 VDDA.t90 GNDA 0.021947f
C1384 VDDA.t124 GNDA 0.021947f
C1385 VDDA.n127 GNDA 0.076056f
C1386 VDDA.n128 GNDA 0.074436f
C1387 VDDA.t136 GNDA 0.021947f
C1388 VDDA.n129 GNDA 0.06584f
C1389 VDDA.n130 GNDA 0.021947f
C1390 VDDA.n131 GNDA 0.012541f
C1391 VDDA.n135 GNDA 0.012541f
C1392 VDDA.t110 GNDA 0.021947f
C1393 VDDA.t120 GNDA 0.021947f
C1394 VDDA.n136 GNDA 0.076056f
C1395 VDDA.n137 GNDA 0.104714f
C1396 VDDA.n138 GNDA 0.021947f
C1397 VDDA.n140 GNDA 0.021947f
C1398 VDDA.n141 GNDA 0.012541f
C1399 VDDA.n142 GNDA 0.012541f
C1400 VDDA.n143 GNDA 0.021947f
C1401 VDDA.n145 GNDA 0.021947f
C1402 VDDA.n146 GNDA 0.012541f
C1403 VDDA.n147 GNDA 0.012541f
C1404 VDDA.n148 GNDA 0.021947f
C1405 VDDA.t155 GNDA 0.038972f
C1406 VDDA.n149 GNDA 0.048957f
C1407 VDDA.t157 GNDA 0.021947f
C1408 VDDA.n151 GNDA 0.06584f
C1409 VDDA.n152 GNDA 0.027097f
C1410 VDDA.n153 GNDA 0.012541f
C1411 VDDA.n154 GNDA 0.183412f
C1412 VDDA.t156 GNDA 0.158957f
C1413 VDDA.t109 GNDA 0.14673f
C1414 VDDA.t119 GNDA 0.14673f
C1415 VDDA.t89 GNDA 0.14673f
C1416 VDDA.t123 GNDA 0.14673f
C1417 VDDA.t95 GNDA 0.14673f
C1418 VDDA.t101 GNDA 0.14673f
C1419 VDDA.t111 GNDA 0.14673f
C1420 VDDA.t121 GNDA 0.14673f
C1421 VDDA.t115 GNDA 0.14673f
C1422 VDDA.t85 GNDA 0.14673f
C1423 VDDA.t135 GNDA 0.158957f
C1424 VDDA.n157 GNDA 0.012541f
C1425 VDDA.t134 GNDA 0.038972f
C1426 VDDA.n159 GNDA 0.048957f
C1427 VDDA.n161 GNDA 0.021947f
C1428 VDDA.n162 GNDA 0.012541f
C1429 VDDA.n163 GNDA 0.012541f
C1430 VDDA.n164 GNDA 0.021947f
C1431 VDDA.n166 GNDA 0.021947f
C1432 VDDA.n167 GNDA 0.021947f
C1433 VDDA.n168 GNDA 0.012541f
C1434 VDDA.n169 GNDA 0.183412f
C1435 VDDA.n171 GNDA 0.029905f
C1436 VDDA.t116 GNDA 0.021947f
C1437 VDDA.t86 GNDA 0.021947f
C1438 VDDA.n172 GNDA 0.076056f
C1439 VDDA.n173 GNDA 0.104714f
C1440 VDDA.t112 GNDA 0.021947f
C1441 VDDA.t122 GNDA 0.021947f
C1442 VDDA.n174 GNDA 0.076056f
C1443 VDDA.n175 GNDA 0.074436f
C1444 VDDA.n176 GNDA 0.020066f
C1445 VDDA.t96 GNDA 0.021947f
C1446 VDDA.t102 GNDA 0.021947f
C1447 VDDA.n177 GNDA 0.07448f
C1448 VDDA.n178 GNDA 0.08673f
C1449 VDDA.t224 GNDA 0.018811f
C1450 VDDA.t29 GNDA 0.018811f
C1451 VDDA.n179 GNDA 0.077794f
C1452 VDDA.t60 GNDA 0.018811f
C1453 VDDA.t14 GNDA 0.018811f
C1454 VDDA.n180 GNDA 0.077496f
C1455 VDDA.n181 GNDA 0.107444f
C1456 VDDA.t35 GNDA 0.018811f
C1457 VDDA.t0 GNDA 0.018811f
C1458 VDDA.n182 GNDA 0.077496f
C1459 VDDA.n183 GNDA 0.056066f
C1460 VDDA.t235 GNDA 0.018811f
C1461 VDDA.t54 GNDA 0.018811f
C1462 VDDA.n184 GNDA 0.077496f
C1463 VDDA.n185 GNDA 0.056066f
C1464 VDDA.t33 GNDA 0.018811f
C1465 VDDA.t231 GNDA 0.018811f
C1466 VDDA.n186 GNDA 0.077496f
C1467 VDDA.n187 GNDA 0.056066f
C1468 VDDA.t244 GNDA 0.018811f
C1469 VDDA.t225 GNDA 0.018811f
C1470 VDDA.n188 GNDA 0.077496f
C1471 VDDA.n189 GNDA 0.097133f
C1472 VDDA.n191 GNDA 0.012541f
C1473 VDDA.n193 GNDA 0.012541f
C1474 VDDA.n194 GNDA 0.021947f
C1475 VDDA.t149 GNDA 0.018905f
C1476 VDDA.n195 GNDA 0.047345f
C1477 VDDA.n196 GNDA 0.012541f
C1478 VDDA.n197 GNDA 0.021947f
C1479 VDDA.t151 GNDA 0.033064f
C1480 VDDA.n199 GNDA 0.030535f
C1481 VDDA.n200 GNDA 0.010308f
C1482 VDDA.n201 GNDA 0.110988f
C1483 VDDA.t150 GNDA 0.092176f
C1484 VDDA.t79 GNDA 0.082771f
C1485 VDDA.t30 GNDA 0.082771f
C1486 VDDA.t240 GNDA 0.082771f
C1487 VDDA.t34 GNDA 0.082771f
C1488 VDDA.t68 GNDA 0.082771f
C1489 VDDA.t230 GNDA 0.082771f
C1490 VDDA.t7 GNDA 0.082771f
C1491 VDDA.t232 GNDA 0.082771f
C1492 VDDA.t12 GNDA 0.082771f
C1493 VDDA.t24 GNDA 0.082771f
C1494 VDDA.t162 GNDA 0.092176f
C1495 VDDA.n203 GNDA 0.012541f
C1496 VDDA.n204 GNDA 0.021947f
C1497 VDDA.n205 GNDA 0.021947f
C1498 VDDA.t163 GNDA 0.033064f
C1499 VDDA.n206 GNDA 0.027645f
C1500 VDDA.n207 GNDA 0.013198f
C1501 VDDA.n208 GNDA 0.110988f
C1502 VDDA.n209 GNDA 0.012541f
C1503 VDDA.n210 GNDA 0.025791f
C1504 VDDA.t161 GNDA 0.018228f
C1505 VDDA.n211 GNDA 0.033815f
C1506 VDDA.n212 GNDA 0.146137f
C1507 VDDA.t166 GNDA 0.011424f
C1508 VDDA.n213 GNDA 0.051619f
C1509 VDDA.t165 GNDA 0.04695f
C1510 VDDA.t6 GNDA 0.031039f
C1511 VDDA.t61 GNDA 0.031039f
C1512 VDDA.t62 GNDA 0.031039f
C1513 VDDA.t72 GNDA 0.031039f
C1514 VDDA.t65 GNDA 0.031039f
C1515 VDDA.t57 GNDA 0.031039f
C1516 VDDA.t1 GNDA 0.031039f
C1517 VDDA.t51 GNDA 0.031039f
C1518 VDDA.t13 GNDA 0.031039f
C1519 VDDA.t243 GNDA 0.031039f
C1520 VDDA.t153 GNDA 0.046649f
C1521 VDDA.t154 GNDA 0.011424f
C1522 VDDA.n214 GNDA 0.026145f
C1523 VDDA.n215 GNDA 0.044414f
C1524 VDDA.n216 GNDA 0.120567f
C1525 VDDA.t76 GNDA 0.037623f
C1526 VDDA.t53 GNDA 0.037623f
C1527 VDDA.n217 GNDA 0.150938f
C1528 VDDA.n218 GNDA 0.076681f
C1529 VDDA.n220 GNDA 0.012541f
C1530 VDDA.n226 GNDA 0.013198f
C1531 VDDA.n227 GNDA 0.012541f
C1532 VDDA.t37 GNDA 0.037623f
C1533 VDDA.t234 GNDA 0.037623f
C1534 VDDA.n228 GNDA 0.150938f
C1535 VDDA.n229 GNDA 0.076681f
C1536 VDDA.t9 GNDA 0.037623f
C1537 VDDA.t229 GNDA 0.037623f
C1538 VDDA.n230 GNDA 0.150938f
C1539 VDDA.n231 GNDA 0.076681f
C1540 VDDA.t39 GNDA 0.037623f
C1541 VDDA.t59 GNDA 0.037623f
C1542 VDDA.n232 GNDA 0.150938f
C1543 VDDA.n233 GNDA 0.076681f
C1544 VDDA.t11 GNDA 0.037623f
C1545 VDDA.t32 GNDA 0.037623f
C1546 VDDA.n234 GNDA 0.150938f
C1547 VDDA.n235 GNDA 0.106392f
C1548 VDDA.n236 GNDA 0.024951f
C1549 VDDA.n237 GNDA 0.012541f
C1550 VDDA.n238 GNDA 0.012541f
C1551 VDDA.n239 GNDA 0.021947f
C1552 VDDA.n240 GNDA 0.012541f
C1553 VDDA.n241 GNDA 0.012541f
C1554 VDDA.n242 GNDA 0.012541f
C1555 VDDA.n243 GNDA 0.012541f
C1556 VDDA.n244 GNDA 0.021947f
C1557 VDDA.n245 GNDA 0.024951f
C1558 VDDA.n246 GNDA 0.012541f
C1559 VDDA.n247 GNDA 0.012541f
C1560 VDDA.n248 GNDA 0.012541f
C1561 VDDA.n249 GNDA 0.031767f
C1562 VDDA.n250 GNDA 0.021947f
C1563 VDDA.n251 GNDA 0.021947f
C1564 VDDA.n252 GNDA 0.021947f
C1565 VDDA.n253 GNDA 0.012541f
C1566 VDDA.n254 GNDA 0.012541f
C1567 VDDA.n256 GNDA 0.021947f
C1568 VDDA.n257 GNDA 0.021947f
C1569 VDDA.n259 GNDA 0.012541f
C1570 VDDA.n260 GNDA 0.012541f
C1571 VDDA.n261 GNDA 0.021947f
C1572 VDDA.n262 GNDA 0.021947f
C1573 VDDA.n263 GNDA 0.021947f
C1574 VDDA.n265 GNDA 0.030752f
C1575 VDDA.n266 GNDA 0.012541f
C1576 VDDA.n267 GNDA 0.295967f
C1577 VDDA.t77 GNDA 0.245803f
C1578 VDDA.t10 GNDA 0.220721f
C1579 VDDA.t31 GNDA 0.220721f
C1580 VDDA.t38 GNDA 0.220721f
C1581 VDDA.t58 GNDA 0.220721f
C1582 VDDA.t8 GNDA 0.220721f
C1583 VDDA.t228 GNDA 0.220721f
C1584 VDDA.t36 GNDA 0.220721f
C1585 VDDA.t233 GNDA 0.220721f
C1586 VDDA.t75 GNDA 0.220721f
C1587 VDDA.t52 GNDA 0.220721f
C1588 VDDA.t66 GNDA 0.245803f
C1589 VDDA.n272 GNDA 0.013198f
C1590 VDDA.n273 GNDA 0.012541f
C1591 VDDA.n274 GNDA 0.021947f
C1592 VDDA.n275 GNDA 0.024951f
C1593 VDDA.n276 GNDA 0.012541f
C1594 VDDA.n277 GNDA 0.012541f
C1595 VDDA.n280 GNDA 0.012541f
C1596 VDDA.n281 GNDA 0.012541f
C1597 VDDA.n282 GNDA 0.024951f
C1598 VDDA.n283 GNDA 0.031767f
C1599 VDDA.n284 GNDA 0.012541f
C1600 VDDA.n285 GNDA 0.021947f
C1601 VDDA.n286 GNDA 0.021947f
C1602 VDDA.n287 GNDA 0.012541f
C1603 VDDA.n288 GNDA 0.012541f
C1604 VDDA.n289 GNDA 0.021947f
C1605 VDDA.n290 GNDA 0.021947f
C1606 VDDA.n291 GNDA 0.012541f
C1607 VDDA.n292 GNDA 0.012541f
C1608 VDDA.n293 GNDA 0.021947f
C1609 VDDA.n294 GNDA 0.021947f
C1610 VDDA.n295 GNDA 0.012541f
C1611 VDDA.n296 GNDA 0.012541f
C1612 VDDA.n297 GNDA 0.021947f
C1613 VDDA.n298 GNDA 0.021947f
C1614 VDDA.n299 GNDA 0.021947f
C1615 VDDA.n300 GNDA 0.012541f
C1616 VDDA.n301 GNDA 0.295967f
C1617 VDDA.n303 GNDA 0.033104f
C1618 VDDA.n304 GNDA 0.038005f
C1619 VDDA.n306 GNDA 0.048012f
C1620 VDDA.t130 GNDA 0.011424f
C1621 VDDA.n308 GNDA 0.048012f
C1622 VDDA.n310 GNDA 0.048012f
C1623 VDDA.n312 GNDA 0.048012f
C1624 VDDA.n314 GNDA 0.048012f
C1625 VDDA.n316 GNDA 0.048012f
C1626 VDDA.n318 GNDA 0.048012f
C1627 VDDA.n320 GNDA 0.048012f
C1628 VDDA.n322 GNDA 0.048012f
C1629 VDDA.n324 GNDA 0.076451f
C1630 VDDA.n325 GNDA 0.060176f
C1631 VDDA.t129 GNDA 0.04695f
C1632 VDDA.t63 GNDA 0.031039f
C1633 VDDA.t2 GNDA 0.031039f
C1634 VDDA.t25 GNDA 0.031039f
C1635 VDDA.t49 GNDA 0.031039f
C1636 VDDA.t241 GNDA 0.031039f
C1637 VDDA.t15 GNDA 0.031039f
C1638 VDDA.t46 GNDA 0.031039f
C1639 VDDA.t247 GNDA 0.031039f
C1640 VDDA.t42 GNDA 0.031039f
C1641 VDDA.t245 GNDA 0.031039f
C1642 VDDA.t55 GNDA 0.031039f
C1643 VDDA.t249 GNDA 0.031039f
C1644 VDDA.t22 GNDA 0.031039f
C1645 VDDA.t44 GNDA 0.031039f
C1646 VDDA.t238 GNDA 0.031039f
C1647 VDDA.t40 GNDA 0.031039f
C1648 VDDA.t4 GNDA 0.031039f
C1649 VDDA.t69 GNDA 0.031039f
C1650 VDDA.t236 GNDA 0.031039f
C1651 VDDA.t17 GNDA 0.031039f
C1652 VDDA.t141 GNDA 0.04695f
C1653 VDDA.t142 GNDA 0.011424f
C1654 VDDA.n326 GNDA 0.059691f
C1655 VDDA.n327 GNDA 0.057455f
C1656 VDDA.n328 GNDA 0.046402f
C1657 VDDA.n329 GNDA 0.116648f
C1658 VDDA.n330 GNDA 0.227544f
C1659 VDDA.t94 GNDA 0.021947f
C1660 VDDA.t98 GNDA 0.021947f
C1661 VDDA.n331 GNDA 0.076056f
C1662 VDDA.n332 GNDA 0.074436f
C1663 VDDA.t139 GNDA 0.021947f
C1664 VDDA.n333 GNDA 0.06584f
C1665 VDDA.n334 GNDA 0.021947f
C1666 VDDA.n335 GNDA 0.012541f
C1667 VDDA.n339 GNDA 0.012541f
C1668 VDDA.t104 GNDA 0.021947f
C1669 VDDA.t114 GNDA 0.021947f
C1670 VDDA.n340 GNDA 0.076056f
C1671 VDDA.n341 GNDA 0.104666f
C1672 VDDA.n342 GNDA 0.023514f
C1673 VDDA.n344 GNDA 0.023514f
C1674 VDDA.n345 GNDA 0.012541f
C1675 VDDA.n346 GNDA 0.012541f
C1676 VDDA.n347 GNDA 0.023514f
C1677 VDDA.n349 GNDA 0.023514f
C1678 VDDA.n350 GNDA 0.012541f
C1679 VDDA.n351 GNDA 0.012541f
C1680 VDDA.n352 GNDA 0.023514f
C1681 VDDA.t171 GNDA 0.038963f
C1682 VDDA.n353 GNDA 0.050377f
C1683 VDDA.t173 GNDA 0.021947f
C1684 VDDA.n355 GNDA 0.076814f
C1685 VDDA.n356 GNDA 0.028556f
C1686 VDDA.n357 GNDA 0.012541f
C1687 VDDA.n358 GNDA 0.189526f
C1688 VDDA.t172 GNDA 0.165071f
C1689 VDDA.t103 GNDA 0.14673f
C1690 VDDA.t113 GNDA 0.14673f
C1691 VDDA.t93 GNDA 0.14673f
C1692 VDDA.t97 GNDA 0.14673f
C1693 VDDA.t105 GNDA 0.14673f
C1694 VDDA.t99 GNDA 0.14673f
C1695 VDDA.t107 GNDA 0.14673f
C1696 VDDA.t117 GNDA 0.14673f
C1697 VDDA.t87 GNDA 0.14673f
C1698 VDDA.t91 GNDA 0.14673f
C1699 VDDA.t138 GNDA 0.158957f
C1700 VDDA.n361 GNDA 0.012541f
C1701 VDDA.t137 GNDA 0.038972f
C1702 VDDA.n363 GNDA 0.048957f
C1703 VDDA.n365 GNDA 0.021947f
C1704 VDDA.n366 GNDA 0.012541f
C1705 VDDA.n367 GNDA 0.012541f
C1706 VDDA.n368 GNDA 0.021947f
C1707 VDDA.n370 GNDA 0.021947f
C1708 VDDA.n371 GNDA 0.021947f
C1709 VDDA.n372 GNDA 0.012541f
C1710 VDDA.n373 GNDA 0.183412f
C1711 VDDA.n375 GNDA 0.029905f
C1712 VDDA.t88 GNDA 0.021947f
C1713 VDDA.t92 GNDA 0.021947f
C1714 VDDA.n376 GNDA 0.076056f
C1715 VDDA.n377 GNDA 0.104714f
C1716 VDDA.t108 GNDA 0.021947f
C1717 VDDA.t118 GNDA 0.021947f
C1718 VDDA.n378 GNDA 0.076056f
C1719 VDDA.n379 GNDA 0.074436f
C1720 VDDA.n380 GNDA 0.020066f
C1721 VDDA.t106 GNDA 0.021947f
C1722 VDDA.t100 GNDA 0.021947f
C1723 VDDA.n381 GNDA 0.07448f
C1724 VDDA.n382 GNDA 0.08694f
C1725 VDDA.n383 GNDA 0.196938f
C1726 VDDA.n384 GNDA 0.077315f
C1727 VDDA.n386 GNDA 0.061522f
C1728 VDDA.t170 GNDA 0.014657f
C1729 VDDA.t167 GNDA 0.013265f
C1730 VDDA.n387 GNDA 0.117824f
C1731 VDDA.t133 GNDA 0.079301f
C1732 VDDA.t131 GNDA 0.041991f
C1733 VDDA.t174 GNDA 0.041991f
C1734 VDDA.t84 GNDA 0.02226f
C1735 VDDA.n388 GNDA 0.079394f
C1736 VDDA.t176 GNDA 0.101562f
C1737 VDDA.n389 GNDA 0.256336f
C1738 VDDA.t175 GNDA 0.219783f
C1739 VDDA.t83 GNDA 0.169303f
C1740 VDDA.t132 GNDA 0.219783f
C1741 VDDA.n390 GNDA 0.256149f
C1742 VDDA.n391 GNDA 0.113353f
C1743 VDDA.n392 GNDA 0.070486f
C1744 VDDA.t158 GNDA 0.013265f
C1745 VDDA.t160 GNDA 0.014657f
C1746 VDDA.n393 GNDA 0.062854f
C1747 VDDA.t159 GNDA 0.058092f
C1748 VDDA.t222 GNDA 0.039504f
C1749 VDDA.t168 GNDA 0.058092f
C1750 VDDA.n394 GNDA 0.06493f
C1751 VDDA.n395 GNDA 0.06887f
C1752 VDDA.n396 GNDA 0.56988f
C1753 VD3.t35 GNDA 0.050359f
C1754 VD3.n1 GNDA 0.059633f
C1755 VD3.n3 GNDA 0.028359f
C1756 VD3.n4 GNDA 0.028359f
C1757 VD3.n5 GNDA 0.016205f
C1758 VD3.n6 GNDA 0.016205f
C1759 VD3.t36 GNDA 0.205398f
C1760 VD3.t0 GNDA 0.028359f
C1761 VD3.t8 GNDA 0.028359f
C1762 VD3.n7 GNDA 0.098626f
C1763 VD3.t4 GNDA 0.028359f
C1764 VD3.t10 GNDA 0.028359f
C1765 VD3.n8 GNDA 0.098276f
C1766 VD3.n9 GNDA 0.185535f
C1767 VD3.t9 GNDA 0.028359f
C1768 VD3.t6 GNDA 0.028359f
C1769 VD3.n10 GNDA 0.098276f
C1770 VD3.n11 GNDA 0.096183f
C1771 VD3.t5 GNDA 0.028359f
C1772 VD3.t3 GNDA 0.028359f
C1773 VD3.n12 GNDA 0.098276f
C1774 VD3.n13 GNDA 0.096183f
C1775 VD3.t7 GNDA 0.028359f
C1776 VD3.t2 GNDA 0.028359f
C1777 VD3.n14 GNDA 0.098276f
C1778 VD3.n15 GNDA 0.096183f
C1779 VD3.t11 GNDA 0.028359f
C1780 VD3.t1 GNDA 0.028359f
C1781 VD3.n16 GNDA 0.098276f
C1782 VD3.n17 GNDA 0.18012f
C1783 VD3.n18 GNDA 0.016205f
C1784 VD3.n19 GNDA 0.028359f
C1785 VD3.n22 GNDA 0.028359f
C1786 VD3.n23 GNDA 0.016205f
C1787 VD3.n24 GNDA 0.016205f
C1788 VD3.n26 GNDA 0.016205f
C1789 VD3.n27 GNDA 0.028359f
C1790 VD3.n28 GNDA 0.028359f
C1791 VD3.n29 GNDA 0.016205f
C1792 VD3.n30 GNDA 0.028359f
C1793 VD3.n31 GNDA 0.016205f
C1794 VD3.t26 GNDA 0.189598f
C1795 VD3.t20 GNDA 0.189598f
C1796 VD3.t24 GNDA 0.189598f
C1797 VD3.t18 GNDA 0.189598f
C1798 VD3.t14 GNDA 0.189598f
C1799 VD3.t12 GNDA 0.189598f
C1800 VD3.t30 GNDA 0.189598f
C1801 VD3.t28 GNDA 0.189598f
C1802 VD3.t22 GNDA 0.189598f
C1803 VD3.t16 GNDA 0.189598f
C1804 VD3.t33 GNDA 0.205398f
C1805 VD3.n33 GNDA 0.236997f
C1806 VD3.n34 GNDA 0.012577f
C1807 VD3.t32 GNDA 0.050359f
C1808 VD3.n35 GNDA 0.063261f
C1809 VD3.t34 GNDA 0.028359f
C1810 VD3.n37 GNDA 0.085076f
C1811 VD3.n38 GNDA 0.034347f
C1812 VD3.n39 GNDA 0.113043f
C1813 VD3.t17 GNDA 0.028359f
C1814 VD3.t23 GNDA 0.028359f
C1815 VD3.n40 GNDA 0.098276f
C1816 VD3.n41 GNDA 0.096184f
C1817 VD3.t29 GNDA 0.028359f
C1818 VD3.t31 GNDA 0.028359f
C1819 VD3.n42 GNDA 0.098276f
C1820 VD3.n43 GNDA 0.096184f
C1821 VD3.t13 GNDA 0.028359f
C1822 VD3.t15 GNDA 0.028359f
C1823 VD3.n44 GNDA 0.098276f
C1824 VD3.n45 GNDA 0.096184f
C1825 VD3.t19 GNDA 0.028359f
C1826 VD3.t25 GNDA 0.028359f
C1827 VD3.n46 GNDA 0.098276f
C1828 VD3.n47 GNDA 0.096184f
C1829 VD3.t21 GNDA 0.028359f
C1830 VD3.t27 GNDA 0.028359f
C1831 VD3.n48 GNDA 0.098276f
C1832 VD3.n49 GNDA 0.135308f
C1833 VD3.n50 GNDA 0.038641f
C1834 VD3.n51 GNDA 0.012577f
C1835 VD3.n52 GNDA 0.016205f
C1836 VD3.n53 GNDA 0.028359f
C1837 VD3.n54 GNDA 0.016205f
C1838 VD3.n55 GNDA 0.028359f
C1839 VD3.n56 GNDA 0.016205f
C1840 VD3.n58 GNDA 0.236997f
C1841 VD3.n60 GNDA 0.016205f
C1842 VD3.n61 GNDA 0.028359f
C1843 VD3.n63 GNDA 0.085076f
C1844 VD3.t37 GNDA 0.028359f
C1845 Vb3.t16 GNDA 0.054986f
C1846 Vb3.t2 GNDA 0.054986f
C1847 Vb3.t19 GNDA 0.054986f
C1848 Vb3.t4 GNDA 0.054986f
C1849 Vb3.t9 GNDA 0.063453f
C1850 Vb3.n0 GNDA 0.051517f
C1851 Vb3.n1 GNDA 0.031658f
C1852 Vb3.n2 GNDA 0.031658f
C1853 Vb3.n3 GNDA 0.029644f
C1854 Vb3.t13 GNDA 0.054986f
C1855 Vb3.t8 GNDA 0.054986f
C1856 Vb3.t3 GNDA 0.054986f
C1857 Vb3.t6 GNDA 0.054986f
C1858 Vb3.t21 GNDA 0.063453f
C1859 Vb3.n4 GNDA 0.051517f
C1860 Vb3.n5 GNDA 0.031658f
C1861 Vb3.n6 GNDA 0.031658f
C1862 Vb3.n7 GNDA 0.029644f
C1863 Vb3.n8 GNDA 0.02992f
C1864 Vb3.t12 GNDA 0.054986f
C1865 Vb3.t15 GNDA 0.054986f
C1866 Vb3.t17 GNDA 0.054986f
C1867 Vb3.t7 GNDA 0.054986f
C1868 Vb3.t11 GNDA 0.063453f
C1869 Vb3.n9 GNDA 0.051517f
C1870 Vb3.n10 GNDA 0.031658f
C1871 Vb3.n11 GNDA 0.031658f
C1872 Vb3.n12 GNDA 0.029644f
C1873 Vb3.t14 GNDA 0.054986f
C1874 Vb3.t10 GNDA 0.054986f
C1875 Vb3.t5 GNDA 0.054986f
C1876 Vb3.t20 GNDA 0.054986f
C1877 Vb3.t18 GNDA 0.063453f
C1878 Vb3.n13 GNDA 0.051517f
C1879 Vb3.n14 GNDA 0.031658f
C1880 Vb3.n15 GNDA 0.031658f
C1881 Vb3.n16 GNDA 0.029644f
C1882 Vb3.n17 GNDA 0.032121f
C1883 Vb3.t1 GNDA 0.03999f
C1884 Vb3.t0 GNDA 0.03999f
C1885 Vb3.n18 GNDA 0.153569f
C1886 Vb3.t22 GNDA 0.068937f
C1887 Vb3.n19 GNDA 0.451236f
C1888 Vb3.n20 GNDA 0.485892f
C1889 V_source.n0 GNDA 0.083087f
C1890 V_source.t6 GNDA 0.012033f
C1891 V_source.t9 GNDA 0.012033f
C1892 V_source.t10 GNDA 0.012033f
C1893 V_source.n1 GNDA 0.047997f
C1894 V_source.t38 GNDA 0.012033f
C1895 V_source.t15 GNDA 0.012033f
C1896 V_source.n2 GNDA 0.047775f
C1897 V_source.n3 GNDA 0.08183f
C1898 V_source.t36 GNDA 0.012033f
C1899 V_source.t39 GNDA 0.012033f
C1900 V_source.n4 GNDA 0.047775f
C1901 V_source.n5 GNDA 0.042711f
C1902 V_source.t20 GNDA 0.049521f
C1903 V_source.t16 GNDA 0.012033f
C1904 V_source.t37 GNDA 0.012033f
C1905 V_source.n6 GNDA 0.04643f
C1906 V_source.n7 GNDA 0.325194f
C1907 V_source.n8 GNDA 0.014439f
C1908 V_source.t13 GNDA 0.012033f
C1909 V_source.t14 GNDA 0.012033f
C1910 V_source.n9 GNDA 0.047775f
C1911 V_source.n10 GNDA 0.042711f
C1912 V_source.t8 GNDA 0.012033f
C1913 V_source.t40 GNDA 0.012033f
C1914 V_source.n11 GNDA 0.047775f
C1915 V_source.n12 GNDA 0.042711f
C1916 V_source.t7 GNDA 0.012033f
C1917 V_source.t25 GNDA 0.012033f
C1918 V_source.n13 GNDA 0.047775f
C1919 V_source.n14 GNDA 0.042711f
C1920 V_source.t17 GNDA 0.012033f
C1921 V_source.t11 GNDA 0.012033f
C1922 V_source.n15 GNDA 0.04643f
C1923 V_source.n16 GNDA 0.024528f
C1924 V_source.n17 GNDA 0.025938f
C1925 V_source.n18 GNDA 0.025737f
C1926 V_source.n19 GNDA 0.087039f
C1927 V_source.n20 GNDA 0.025737f
C1928 V_source.n21 GNDA 0.045304f
C1929 V_source.n22 GNDA 0.025737f
C1930 V_source.n23 GNDA 0.025926f
C1931 V_source.n24 GNDA 0.025737f
C1932 V_source.n25 GNDA 0.086183f
C1933 V_source.n26 GNDA 0.025737f
C1934 V_source.n27 GNDA 0.045304f
C1935 V_source.n28 GNDA 0.025737f
C1936 V_source.n29 GNDA 0.045304f
C1937 V_source.n30 GNDA 0.025737f
C1938 V_source.n31 GNDA 0.069129f
C1939 V_source.n32 GNDA 0.041164f
C1940 V_source.n33 GNDA 0.040838f
C1941 V_source.n34 GNDA 0.014439f
C1942 V_source.t21 GNDA 0.012033f
C1943 V_source.t24 GNDA 0.012033f
C1944 V_source.n35 GNDA 0.047775f
C1945 V_source.n36 GNDA 0.083233f
C1946 V_source.n37 GNDA 0.048039f
C1947 V_source.t0 GNDA 0.012033f
C1948 VIN-.t4 GNDA 0.051074f
C1949 VIN-.t10 GNDA 0.033698f
C1950 VIN-.t6 GNDA 0.041603f
C1951 VIN-.n0 GNDA 0.059781f
C1952 VIN-.n1 GNDA 0.282874f
C1953 VIN-.t1 GNDA 0.033144f
C1954 VIN-.t8 GNDA 0.041618f
C1955 VIN-.n2 GNDA 0.065446f
C1956 VIN-.n3 GNDA 0.202595f
C1957 VIN-.t3 GNDA 0.050506f
C1958 VIN-.n4 GNDA 0.238259f
C1959 VIN-.t2 GNDA 0.050856f
C1960 VIN-.n5 GNDA 0.182164f
C1961 VIN-.t7 GNDA 0.033698f
C1962 VIN-.t0 GNDA 0.041603f
C1963 VIN-.n6 GNDA 0.059781f
C1964 VIN-.n7 GNDA 0.150907f
C1965 VIN-.t9 GNDA 0.033144f
C1966 VIN-.t5 GNDA 0.041618f
C1967 VIN-.n8 GNDA 0.065446f
C1968 VIN-.n9 GNDA 0.17917f
C1969 VD4.t30 GNDA 0.028359f
C1970 VD4.t32 GNDA 0.028359f
C1971 VD4.n0 GNDA 0.098276f
C1972 VD4.n1 GNDA 0.096184f
C1973 VD4.t16 GNDA 0.028359f
C1974 VD4.n2 GNDA 0.085076f
C1975 VD4.n3 GNDA 0.028359f
C1976 VD4.n4 GNDA 0.016205f
C1977 VD4.n7 GNDA 0.012577f
C1978 VD4.n8 GNDA 0.016205f
C1979 VD4.t22 GNDA 0.028359f
C1980 VD4.t26 GNDA 0.028359f
C1981 VD4.n9 GNDA 0.098276f
C1982 VD4.n10 GNDA 0.096183f
C1983 VD4.t18 GNDA 0.028359f
C1984 VD4.t36 GNDA 0.028359f
C1985 VD4.n11 GNDA 0.098276f
C1986 VD4.n12 GNDA 0.096184f
C1987 VD4.t28 GNDA 0.028359f
C1988 VD4.t34 GNDA 0.028359f
C1989 VD4.n13 GNDA 0.098276f
C1990 VD4.n14 GNDA 0.096184f
C1991 VD4.t20 GNDA 0.028359f
C1992 VD4.t24 GNDA 0.028359f
C1993 VD4.n15 GNDA 0.098276f
C1994 VD4.n16 GNDA 0.135308f
C1995 VD4.n17 GNDA 0.028359f
C1996 VD4.n19 GNDA 0.028359f
C1997 VD4.n20 GNDA 0.016205f
C1998 VD4.n21 GNDA 0.016205f
C1999 VD4.n22 GNDA 0.028359f
C2000 VD4.n24 GNDA 0.028359f
C2001 VD4.n25 GNDA 0.016205f
C2002 VD4.n26 GNDA 0.016205f
C2003 VD4.n27 GNDA 0.028359f
C2004 VD4.t11 GNDA 0.050359f
C2005 VD4.n28 GNDA 0.06326f
C2006 VD4.t13 GNDA 0.028359f
C2007 VD4.n30 GNDA 0.085076f
C2008 VD4.n31 GNDA 0.035014f
C2009 VD4.n32 GNDA 0.016205f
C2010 VD4.n33 GNDA 0.236997f
C2011 VD4.t12 GNDA 0.205398f
C2012 VD4.t19 GNDA 0.189598f
C2013 VD4.t23 GNDA 0.189598f
C2014 VD4.t27 GNDA 0.189598f
C2015 VD4.t33 GNDA 0.189598f
C2016 VD4.t17 GNDA 0.189598f
C2017 VD4.t35 GNDA 0.189598f
C2018 VD4.t21 GNDA 0.189598f
C2019 VD4.t25 GNDA 0.189598f
C2020 VD4.t29 GNDA 0.189598f
C2021 VD4.t31 GNDA 0.189598f
C2022 VD4.t15 GNDA 0.205398f
C2023 VD4.n35 GNDA 0.012577f
C2024 VD4.n36 GNDA 0.016205f
C2025 VD4.t14 GNDA 0.050359f
C2026 VD4.n38 GNDA 0.06326f
C2027 VD4.n40 GNDA 0.028359f
C2028 VD4.n41 GNDA 0.016205f
C2029 VD4.n42 GNDA 0.016205f
C2030 VD4.n43 GNDA 0.028359f
C2031 VD4.n45 GNDA 0.028359f
C2032 VD4.n46 GNDA 0.028359f
C2033 VD4.n47 GNDA 0.016205f
C2034 VD4.n48 GNDA 0.236997f
C2035 VD4.n49 GNDA 0.012577f
C2036 VD4.n50 GNDA 0.037974f
C2037 VD4.n51 GNDA 0.060662f
C2038 VD4.t8 GNDA 0.028359f
C2039 VD4.t3 GNDA 0.028359f
C2040 VD4.n52 GNDA 0.098625f
C2041 VD4.t4 GNDA 0.028359f
C2042 VD4.t1 GNDA 0.028359f
C2043 VD4.n53 GNDA 0.098276f
C2044 VD4.n54 GNDA 0.185535f
C2045 VD4.t2 GNDA 0.028359f
C2046 VD4.t9 GNDA 0.028359f
C2047 VD4.n55 GNDA 0.098276f
C2048 VD4.n56 GNDA 0.096183f
C2049 VD4.t7 GNDA 0.028359f
C2050 VD4.t6 GNDA 0.028359f
C2051 VD4.n57 GNDA 0.098276f
C2052 VD4.n58 GNDA 0.096183f
C2053 VD4.t10 GNDA 0.028359f
C2054 VD4.t5 GNDA 0.028359f
C2055 VD4.n59 GNDA 0.098276f
C2056 VD4.n60 GNDA 0.096183f
C2057 VD4.t37 GNDA 0.028359f
C2058 VD4.t0 GNDA 0.028359f
C2059 VD4.n61 GNDA 0.098276f
C2060 VD4.n62 GNDA 0.148152f
C2061 Y.t11 GNDA 0.020284f
C2062 Y.t5 GNDA 0.020284f
C2063 Y.n0 GNDA 0.068484f
C2064 Y.t12 GNDA 0.020284f
C2065 Y.t10 GNDA 0.020284f
C2066 Y.n1 GNDA 0.073194f
C2067 Y.t7 GNDA 0.020284f
C2068 Y.t1 GNDA 0.020284f
C2069 Y.n2 GNDA 0.072555f
C2070 Y.n3 GNDA 0.269399f
C2071 Y.t6 GNDA 0.020284f
C2072 Y.t0 GNDA 0.020284f
C2073 Y.n4 GNDA 0.072555f
C2074 Y.n5 GNDA 0.139752f
C2075 Y.t2 GNDA 0.020284f
C2076 Y.t23 GNDA 0.020284f
C2077 Y.n6 GNDA 0.072555f
C2078 Y.n7 GNDA 0.139752f
C2079 Y.t24 GNDA 0.020284f
C2080 Y.t4 GNDA 0.020284f
C2081 Y.n8 GNDA 0.073194f
C2082 Y.n9 GNDA 0.170215f
C2083 Y.n10 GNDA 0.21308f
C2084 Y.t9 GNDA 0.04733f
C2085 Y.t18 GNDA 0.04733f
C2086 Y.n11 GNDA 0.164603f
C2087 Y.t14 GNDA 0.04733f
C2088 Y.t17 GNDA 0.04733f
C2089 Y.n12 GNDA 0.164019f
C2090 Y.n13 GNDA 0.309652f
C2091 Y.t19 GNDA 0.04733f
C2092 Y.t22 GNDA 0.04733f
C2093 Y.n14 GNDA 0.164019f
C2094 Y.n15 GNDA 0.160527f
C2095 Y.t13 GNDA 0.04733f
C2096 Y.t21 GNDA 0.04733f
C2097 Y.n16 GNDA 0.164019f
C2098 Y.n17 GNDA 0.160527f
C2099 Y.t15 GNDA 0.04733f
C2100 Y.t20 GNDA 0.04733f
C2101 Y.n18 GNDA 0.164019f
C2102 Y.n19 GNDA 0.189023f
C2103 Y.t16 GNDA 0.04733f
C2104 Y.t3 GNDA 0.04733f
C2105 Y.n20 GNDA 0.160621f
C2106 Y.n21 GNDA 0.320399f
C2107 Y.t27 GNDA 0.028398f
C2108 Y.t51 GNDA 0.034483f
C2109 Y.n22 GNDA 0.032156f
C2110 Y.t42 GNDA 0.028398f
C2111 Y.t29 GNDA 0.028398f
C2112 Y.t44 GNDA 0.028398f
C2113 Y.t32 GNDA 0.028398f
C2114 Y.t47 GNDA 0.028398f
C2115 Y.t35 GNDA 0.028398f
C2116 Y.t50 GNDA 0.028398f
C2117 Y.t38 GNDA 0.034483f
C2118 Y.n23 GNDA 0.034483f
C2119 Y.n24 GNDA 0.022313f
C2120 Y.n25 GNDA 0.022313f
C2121 Y.n26 GNDA 0.022313f
C2122 Y.n27 GNDA 0.022313f
C2123 Y.n28 GNDA 0.022313f
C2124 Y.n29 GNDA 0.019986f
C2125 Y.n30 GNDA 0.019656f
C2126 Y.t31 GNDA 0.043611f
C2127 Y.t26 GNDA 0.049578f
C2128 Y.n31 GNDA 0.042416f
C2129 Y.t46 GNDA 0.043611f
C2130 Y.t34 GNDA 0.043611f
C2131 Y.t49 GNDA 0.043611f
C2132 Y.t37 GNDA 0.043611f
C2133 Y.t54 GNDA 0.043611f
C2134 Y.t40 GNDA 0.043611f
C2135 Y.t25 GNDA 0.043611f
C2136 Y.t41 GNDA 0.049578f
C2137 Y.n32 GNDA 0.044743f
C2138 Y.n33 GNDA 0.027384f
C2139 Y.n34 GNDA 0.027384f
C2140 Y.n35 GNDA 0.027384f
C2141 Y.n36 GNDA 0.027384f
C2142 Y.n37 GNDA 0.027384f
C2143 Y.n38 GNDA 0.025057f
C2144 Y.n39 GNDA 0.019615f
C2145 Y.n40 GNDA 0.211405f
C2146 Y.n41 GNDA 0.440199f
C2147 Y.n42 GNDA 0.222835f
C2148 Y.t48 GNDA 0.08925f
C2149 Y.t33 GNDA 0.08925f
C2150 Y.t45 GNDA 0.08925f
C2151 Y.t30 GNDA 0.08925f
C2152 Y.t43 GNDA 0.08925f
C2153 Y.t28 GNDA 0.08925f
C2154 Y.t53 GNDA 0.095058f
C2155 Y.n43 GNDA 0.075329f
C2156 Y.n44 GNDA 0.042597f
C2157 Y.n45 GNDA 0.042597f
C2158 Y.n46 GNDA 0.042597f
C2159 Y.n47 GNDA 0.042597f
C2160 Y.n48 GNDA 0.04027f
C2161 Y.t36 GNDA 0.08925f
C2162 Y.t52 GNDA 0.08925f
C2163 Y.t39 GNDA 0.095058f
C2164 Y.n49 GNDA 0.075329f
C2165 Y.n50 GNDA 0.04027f
C2166 Y.n51 GNDA 0.02182f
C2167 Y.n52 GNDA 0.721482f
C2168 Y.t8 GNDA 0.648245f
.ends

