magic
tech sky130A
timestamp 1738172952
<< nwell >>
rect -3570 220 -1745 460
rect -695 215 5 1055
<< pwell >>
rect -3030 5 -2825 115
rect -2575 5 -2370 115
rect -2115 5 -1910 115
<< nmos >>
rect -3500 10 -3485 110
rect -3350 10 -3335 110
rect -3200 10 -3185 110
rect -2975 10 -2960 110
rect -2750 10 -2735 110
rect -2520 10 -2505 110
rect -2290 10 -2275 110
rect -2060 10 -2045 110
rect -1830 10 -1815 110
rect -1125 -265 -1065 135
rect -625 -265 -565 135
rect -125 -265 -65 135
<< pmos >>
rect -3500 240 -3485 440
rect -3350 240 -3335 440
rect -3200 240 -3185 440
rect -2975 240 -2960 440
rect -2750 240 -2735 440
rect -2520 240 -2505 440
rect -2290 240 -2275 440
rect -2060 240 -2045 440
rect -1830 240 -1815 440
rect -625 235 -565 1035
rect -125 235 -65 1035
<< ndiff >>
rect -3550 95 -3500 110
rect -3550 25 -3535 95
rect -3515 25 -3500 95
rect -3550 10 -3500 25
rect -3485 95 -3435 110
rect -3485 25 -3470 95
rect -3450 25 -3435 95
rect -3485 10 -3435 25
rect -3400 95 -3350 110
rect -3400 25 -3385 95
rect -3365 25 -3350 95
rect -3400 10 -3350 25
rect -3335 95 -3285 110
rect -3335 25 -3320 95
rect -3300 25 -3285 95
rect -3335 10 -3285 25
rect -3250 95 -3200 110
rect -3250 25 -3235 95
rect -3215 25 -3200 95
rect -3250 10 -3200 25
rect -3185 95 -3135 110
rect -3185 25 -3170 95
rect -3150 25 -3135 95
rect -3025 95 -2975 110
rect -3185 10 -3135 25
rect -3025 25 -3010 95
rect -2990 25 -2975 95
rect -3025 10 -2975 25
rect -2960 95 -2910 110
rect -2960 25 -2945 95
rect -2925 25 -2910 95
rect -2960 10 -2910 25
rect -2800 95 -2750 110
rect -2800 25 -2785 95
rect -2765 25 -2750 95
rect -2800 10 -2750 25
rect -2735 95 -2685 110
rect -2735 25 -2720 95
rect -2700 25 -2685 95
rect -2570 95 -2520 110
rect -2735 10 -2685 25
rect -2570 25 -2555 95
rect -2535 25 -2520 95
rect -2570 10 -2520 25
rect -2505 95 -2455 110
rect -2505 25 -2490 95
rect -2470 25 -2455 95
rect -2505 10 -2455 25
rect -2340 95 -2290 110
rect -2340 25 -2325 95
rect -2305 25 -2290 95
rect -2340 10 -2290 25
rect -2275 95 -2225 110
rect -2275 25 -2260 95
rect -2240 25 -2225 95
rect -2110 95 -2060 110
rect -2275 10 -2225 25
rect -2110 25 -2095 95
rect -2075 25 -2060 95
rect -2110 10 -2060 25
rect -2045 95 -1995 110
rect -2045 25 -2030 95
rect -2010 25 -1995 95
rect -2045 10 -1995 25
rect -1880 95 -1830 110
rect -1880 25 -1865 95
rect -1845 25 -1830 95
rect -1880 10 -1830 25
rect -1815 95 -1765 110
rect -1815 25 -1800 95
rect -1780 25 -1765 95
rect -1815 10 -1765 25
rect -1175 120 -1125 135
rect -1175 -250 -1160 120
rect -1140 -250 -1125 120
rect -1175 -265 -1125 -250
rect -1065 120 -1015 135
rect -1065 -250 -1050 120
rect -1030 -250 -1015 120
rect -1065 -265 -1015 -250
rect -675 120 -625 135
rect -675 -250 -660 120
rect -640 -250 -625 120
rect -675 -265 -625 -250
rect -565 120 -515 135
rect -565 -250 -550 120
rect -530 -250 -515 120
rect -565 -265 -515 -250
rect -175 120 -125 135
rect -175 -250 -160 120
rect -140 -250 -125 120
rect -175 -265 -125 -250
rect -65 120 -15 135
rect -65 -250 -50 120
rect -30 -250 -15 120
rect -65 -265 -15 -250
<< pdiff >>
rect -675 1020 -625 1035
rect -3550 425 -3500 440
rect -3550 255 -3535 425
rect -3515 255 -3500 425
rect -3550 240 -3500 255
rect -3485 425 -3435 440
rect -3485 255 -3470 425
rect -3450 255 -3435 425
rect -3485 240 -3435 255
rect -3400 425 -3350 440
rect -3400 255 -3385 425
rect -3365 255 -3350 425
rect -3400 240 -3350 255
rect -3335 425 -3285 440
rect -3335 255 -3320 425
rect -3300 255 -3285 425
rect -3335 240 -3285 255
rect -3250 425 -3200 440
rect -3250 255 -3235 425
rect -3215 255 -3200 425
rect -3250 240 -3200 255
rect -3185 425 -3135 440
rect -3185 255 -3170 425
rect -3150 255 -3135 425
rect -3185 240 -3135 255
rect -3025 425 -2975 440
rect -3025 255 -3010 425
rect -2990 255 -2975 425
rect -3025 240 -2975 255
rect -2960 425 -2910 440
rect -2960 255 -2945 425
rect -2925 255 -2910 425
rect -2800 425 -2750 440
rect -2960 240 -2910 255
rect -2800 255 -2785 425
rect -2765 255 -2750 425
rect -2800 240 -2750 255
rect -2735 425 -2685 440
rect -2735 255 -2720 425
rect -2700 255 -2685 425
rect -2735 240 -2685 255
rect -2570 425 -2520 440
rect -2570 255 -2555 425
rect -2535 255 -2520 425
rect -2570 240 -2520 255
rect -2505 425 -2455 440
rect -2505 255 -2490 425
rect -2470 255 -2455 425
rect -2340 425 -2290 440
rect -2505 240 -2455 255
rect -2340 255 -2325 425
rect -2305 255 -2290 425
rect -2340 240 -2290 255
rect -2275 425 -2225 440
rect -2275 255 -2260 425
rect -2240 255 -2225 425
rect -2275 240 -2225 255
rect -2110 425 -2060 440
rect -2110 255 -2095 425
rect -2075 255 -2060 425
rect -2110 240 -2060 255
rect -2045 425 -1995 440
rect -2045 255 -2030 425
rect -2010 255 -1995 425
rect -1880 425 -1830 440
rect -2045 240 -1995 255
rect -1880 255 -1865 425
rect -1845 255 -1830 425
rect -1880 240 -1830 255
rect -1815 425 -1765 440
rect -1815 255 -1800 425
rect -1780 255 -1765 425
rect -1815 240 -1765 255
rect -675 250 -660 1020
rect -640 250 -625 1020
rect -675 235 -625 250
rect -565 1020 -515 1035
rect -565 250 -550 1020
rect -530 250 -515 1020
rect -565 235 -515 250
rect -175 1020 -125 1035
rect -175 250 -160 1020
rect -140 250 -125 1020
rect -175 235 -125 250
rect -65 1020 -15 1035
rect -65 250 -50 1020
rect -30 250 -15 1020
rect -65 235 -15 250
<< ndiffc >>
rect -3535 25 -3515 95
rect -3470 25 -3450 95
rect -3385 25 -3365 95
rect -3320 25 -3300 95
rect -3235 25 -3215 95
rect -3170 25 -3150 95
rect -3010 25 -2990 95
rect -2945 25 -2925 95
rect -2785 25 -2765 95
rect -2720 25 -2700 95
rect -2555 25 -2535 95
rect -2490 25 -2470 95
rect -2325 25 -2305 95
rect -2260 25 -2240 95
rect -2095 25 -2075 95
rect -2030 25 -2010 95
rect -1865 25 -1845 95
rect -1800 25 -1780 95
rect -1160 -250 -1140 120
rect -1050 -250 -1030 120
rect -660 -250 -640 120
rect -550 -250 -530 120
rect -160 -250 -140 120
rect -50 -250 -30 120
<< pdiffc >>
rect -3535 255 -3515 425
rect -3470 255 -3450 425
rect -3385 255 -3365 425
rect -3320 255 -3300 425
rect -3235 255 -3215 425
rect -3170 255 -3150 425
rect -3010 255 -2990 425
rect -2945 255 -2925 425
rect -2785 255 -2765 425
rect -2720 255 -2700 425
rect -2555 255 -2535 425
rect -2490 255 -2470 425
rect -2325 255 -2305 425
rect -2260 255 -2240 425
rect -2095 255 -2075 425
rect -2030 255 -2010 425
rect -1865 255 -1845 425
rect -1800 255 -1780 425
rect -660 250 -640 1020
rect -550 250 -530 1020
rect -160 250 -140 1020
rect -50 250 -30 1020
<< psubdiff >>
rect -2880 95 -2830 110
rect -2880 25 -2865 95
rect -2845 25 -2830 95
rect -2880 10 -2830 25
rect -2425 95 -2375 110
rect -2425 25 -2410 95
rect -2390 25 -2375 95
rect -2425 10 -2375 25
rect -1965 95 -1915 110
rect -1965 25 -1950 95
rect -1930 25 -1915 95
rect -1965 10 -1915 25
rect -1015 120 -965 135
rect -1015 -250 -1000 120
rect -980 -250 -965 120
rect -1015 -265 -965 -250
rect -515 120 -465 135
rect -515 -250 -500 120
rect -480 -250 -465 120
rect -515 -265 -465 -250
rect -225 120 -175 135
rect -225 -250 -210 120
rect -190 -250 -175 120
rect -225 -265 -175 -250
<< nsubdiff >>
rect -3105 425 -3055 440
rect -3105 255 -3090 425
rect -3070 255 -3055 425
rect -3105 240 -3055 255
rect -2650 425 -2600 440
rect -2650 255 -2635 425
rect -2615 255 -2600 425
rect -2650 240 -2600 255
rect -2190 425 -2140 440
rect -2190 255 -2175 425
rect -2155 255 -2140 425
rect -2190 240 -2140 255
rect -515 1020 -465 1035
rect -515 250 -500 1020
rect -480 250 -465 1020
rect -515 235 -465 250
rect -225 1020 -175 1035
rect -225 250 -210 1020
rect -190 250 -175 1020
rect -225 235 -175 250
<< psubdiffcont >>
rect -2865 25 -2845 95
rect -2410 25 -2390 95
rect -1950 25 -1930 95
rect -1000 -250 -980 120
rect -500 -250 -480 120
rect -210 -250 -190 120
<< nsubdiffcont >>
rect -3090 255 -3070 425
rect -2635 255 -2615 425
rect -2175 255 -2155 425
rect -500 250 -480 1020
rect -210 250 -190 1020
<< poly >>
rect -1560 1235 495 1250
rect -1560 875 -1545 1235
rect -625 1035 -565 1050
rect -125 1035 -65 1050
rect -3160 860 -1545 875
rect -3160 740 -3145 860
rect -1695 740 -1680 860
rect -3160 730 -3120 740
rect -3160 710 -3150 730
rect -3130 710 -3120 730
rect -3160 700 -3120 710
rect -3020 730 -1680 740
rect -3020 710 -3010 730
rect -2990 725 -1680 730
rect -2990 710 -2980 725
rect -3020 700 -2980 710
rect -2940 690 -1720 700
rect -2940 670 -2930 690
rect -2910 685 -1720 690
rect -2910 670 -2900 685
rect -2940 660 -2900 670
rect -3200 620 -1815 635
rect -3500 440 -3485 455
rect -3350 440 -3335 455
rect -3200 440 -3185 620
rect -3160 585 -3120 595
rect -3160 565 -3150 585
rect -3130 570 -3120 585
rect -3130 565 -2960 570
rect -3160 555 -2960 565
rect -2975 440 -2960 555
rect -2520 455 -2415 470
rect -2750 440 -2735 455
rect -2520 440 -2505 455
rect -2430 445 -2415 455
rect -2885 430 -2845 440
rect -2885 410 -2875 430
rect -2855 410 -2845 430
rect -2885 400 -2845 410
rect -2430 435 -2390 445
rect -2290 440 -2275 455
rect -2060 440 -2045 455
rect -1830 440 -1815 620
rect -2430 415 -2420 435
rect -2400 415 -2390 435
rect -2430 405 -2390 415
rect -1970 425 -1930 435
rect -1970 405 -1960 425
rect -1940 405 -1930 425
rect -1970 395 -1930 405
rect -3500 185 -3485 240
rect -3350 200 -3335 240
rect -3200 200 -3185 240
rect -2975 225 -2960 240
rect -3565 170 -3485 185
rect -3500 110 -3485 170
rect -3375 190 -3335 200
rect -3375 170 -3365 190
rect -3345 170 -3335 190
rect -3375 160 -3335 170
rect -3225 190 -3185 200
rect -3225 170 -3215 190
rect -3195 170 -3185 190
rect -3225 160 -3185 170
rect -3020 190 -2980 200
rect -3020 170 -3010 190
rect -2990 170 -2980 190
rect -3020 160 -2980 170
rect -2955 190 -2915 200
rect -2955 170 -2945 190
rect -2925 170 -2915 190
rect -2955 160 -2915 170
rect -3350 110 -3335 160
rect -3200 135 -3185 160
rect -3200 120 -2960 135
rect -3200 110 -3185 120
rect -2975 110 -2960 120
rect -2750 110 -2735 240
rect -2520 225 -2505 240
rect -2290 215 -2275 240
rect -2060 215 -2045 240
rect -1830 225 -1815 240
rect -2290 200 -1850 215
rect -2710 190 -2670 200
rect -2710 170 -2700 190
rect -2680 185 -2670 190
rect -2565 190 -2525 200
rect -2565 185 -2555 190
rect -2680 170 -2555 185
rect -2535 170 -2525 190
rect -2710 160 -2670 170
rect -2565 160 -2525 170
rect -2500 190 -2460 200
rect -2500 170 -2490 190
rect -2470 185 -2460 190
rect -2315 190 -2275 200
rect -2315 185 -2305 190
rect -2470 170 -2305 185
rect -2285 170 -2275 190
rect -2500 160 -2460 170
rect -2315 160 -2275 170
rect -2520 110 -2505 125
rect -2290 110 -2275 160
rect -1865 135 -1850 200
rect -1735 200 -1720 685
rect -1210 225 -1090 240
rect 480 875 495 1235
rect 480 860 590 875
rect 590 240 605 250
rect -625 225 -565 235
rect -1445 210 -1195 225
rect -1105 210 -565 225
rect -125 225 -65 235
rect 465 225 605 240
rect -125 210 480 225
rect -1445 200 -1430 210
rect -1735 185 -1430 200
rect -1170 180 -1130 190
rect -1170 165 -1160 180
rect -1400 160 -1160 165
rect -1140 165 -1130 180
rect -1140 160 -565 165
rect -1400 150 -565 160
rect -2060 110 -2045 125
rect -1865 120 -1815 135
rect -1830 110 -1815 120
rect -3090 40 -3050 50
rect -3090 20 -3080 40
rect -3060 20 -3050 40
rect -3090 10 -3050 20
rect -2635 40 -2595 50
rect -2635 20 -2625 40
rect -2605 20 -2595 40
rect -2635 10 -2595 20
rect -2175 40 -2135 50
rect -2175 20 -2165 40
rect -2145 20 -2135 40
rect -2175 10 -2135 20
rect -3500 -5 -3485 10
rect -3350 -5 -3335 10
rect -3200 -5 -3185 10
rect -2975 -5 -2960 10
rect -2750 -120 -2735 10
rect -2610 0 -2595 10
rect -2520 0 -2505 10
rect -2610 -15 -2505 0
rect -2290 -5 -2275 10
rect -3565 -135 -2735 -120
rect -2250 -55 -2210 -50
rect -2060 -55 -2045 10
rect -1830 -5 -1815 10
rect -2250 -60 -2045 -55
rect -2250 -80 -2240 -60
rect -2220 -70 -2045 -60
rect -2020 -65 -1980 -55
rect -2220 -80 -2210 -70
rect -2250 -90 -2210 -80
rect -2020 -85 -2010 -65
rect -1990 -80 -1980 -65
rect -1400 -80 -1385 150
rect -1125 145 -565 150
rect -1125 135 -1065 145
rect -625 135 -565 145
rect -125 145 170 160
rect -125 135 -65 145
rect -1990 -85 -1385 -80
rect -2250 -160 -2235 -90
rect -2020 -95 -1385 -85
rect -2105 -105 -2065 -95
rect -2105 -125 -2095 -105
rect -2075 -120 -2065 -105
rect -2075 -125 -1625 -120
rect -2105 -135 -1625 -125
rect -1640 -160 -1625 -135
rect -2250 -175 -1545 -160
rect -1560 -475 -1545 -175
rect 155 125 170 145
rect 155 110 605 125
rect 590 100 605 110
rect 480 -175 590 -160
rect -1125 -280 -1065 -265
rect -625 -280 -565 -265
rect -125 -280 -65 -265
rect 480 -475 495 -175
rect -1560 -490 495 -475
<< polycont >>
rect -3150 710 -3130 730
rect -3010 710 -2990 730
rect -2930 670 -2910 690
rect -3150 565 -3130 585
rect -2875 410 -2855 430
rect -2420 415 -2400 435
rect -1960 405 -1940 425
rect -3365 170 -3345 190
rect -3215 170 -3195 190
rect -3010 170 -2990 190
rect -2945 170 -2925 190
rect -2700 170 -2680 190
rect -2555 170 -2535 190
rect -2490 170 -2470 190
rect -2305 170 -2285 190
rect -1160 160 -1140 180
rect -3080 20 -3060 40
rect -2625 20 -2605 40
rect -2165 20 -2145 40
rect -2240 -80 -2220 -60
rect -2010 -85 -1990 -65
rect -2095 -125 -2075 -105
<< locali >>
rect -670 1020 -630 1030
rect -3310 760 -1855 780
rect -3310 435 -3290 760
rect -3160 730 -3120 740
rect -3160 710 -3150 730
rect -3130 710 -3120 730
rect -3160 700 -3120 710
rect -3020 730 -2980 740
rect -3020 710 -3010 730
rect -2990 710 -2980 730
rect -3020 700 -2980 710
rect -3160 595 -3140 700
rect -3160 585 -3120 595
rect -3160 565 -3150 585
rect -3130 565 -3120 585
rect -3160 555 -3120 565
rect -3160 435 -3140 555
rect -3020 435 -3000 700
rect -2940 690 -2900 700
rect -2940 670 -2930 690
rect -2910 670 -2900 690
rect -2940 660 -2900 670
rect -2940 435 -2920 660
rect -3545 425 -3505 435
rect -3545 255 -3535 425
rect -3515 255 -3505 425
rect -3545 245 -3505 255
rect -3480 425 -3440 435
rect -3480 255 -3470 425
rect -3450 255 -3440 425
rect -3480 245 -3440 255
rect -3395 425 -3355 435
rect -3395 255 -3385 425
rect -3365 255 -3355 425
rect -3395 245 -3355 255
rect -3330 425 -3290 435
rect -3330 255 -3320 425
rect -3300 255 -3290 425
rect -3330 245 -3290 255
rect -3245 425 -3205 435
rect -3245 255 -3235 425
rect -3215 255 -3205 425
rect -3245 245 -3205 255
rect -3180 425 -3140 435
rect -3180 255 -3170 425
rect -3150 255 -3140 425
rect -3180 245 -3140 255
rect -3100 425 -3060 435
rect -3100 255 -3090 425
rect -3070 255 -3060 425
rect -3100 245 -3060 255
rect -3020 425 -2980 435
rect -3020 255 -3010 425
rect -2990 255 -2980 425
rect -3020 245 -2980 255
rect -2955 425 -2915 435
rect -2955 255 -2945 425
rect -2925 255 -2915 425
rect -2885 430 -2845 440
rect -2430 435 -2390 445
rect -1875 435 -1855 760
rect -2885 410 -2875 430
rect -2855 410 -2845 430
rect -2885 400 -2845 410
rect -2955 245 -2915 255
rect -3460 190 -3440 245
rect -3375 190 -3335 200
rect -3460 170 -3365 190
rect -3345 170 -3335 190
rect -3460 105 -3440 170
rect -3375 160 -3335 170
rect -3310 190 -3290 245
rect -3225 190 -3185 200
rect -3310 170 -3215 190
rect -3195 170 -3185 190
rect -3310 105 -3290 170
rect -3225 160 -3185 170
rect -3160 105 -3140 245
rect -3545 95 -3505 105
rect -3545 25 -3535 95
rect -3515 25 -3505 95
rect -3545 15 -3505 25
rect -3480 95 -3440 105
rect -3480 25 -3470 95
rect -3450 25 -3440 95
rect -3480 15 -3440 25
rect -3395 95 -3355 105
rect -3395 25 -3385 95
rect -3365 25 -3355 95
rect -3395 15 -3355 25
rect -3330 95 -3290 105
rect -3330 25 -3320 95
rect -3300 25 -3290 95
rect -3330 15 -3290 25
rect -3245 95 -3205 105
rect -3245 25 -3235 95
rect -3215 25 -3205 95
rect -3245 15 -3205 25
rect -3180 95 -3140 105
rect -3180 25 -3170 95
rect -3150 25 -3140 95
rect -3180 15 -3140 25
rect -3090 50 -3070 245
rect -3010 200 -2990 245
rect -2945 200 -2925 245
rect -3020 190 -2980 200
rect -3020 170 -3010 190
rect -2990 170 -2980 190
rect -3020 160 -2980 170
rect -2955 190 -2915 200
rect -2955 170 -2945 190
rect -2925 170 -2915 190
rect -2955 160 -2915 170
rect -3010 105 -2990 160
rect -2945 105 -2925 160
rect -2865 105 -2845 400
rect -2795 425 -2755 435
rect -2795 255 -2785 425
rect -2765 255 -2755 425
rect -2795 245 -2755 255
rect -2730 425 -2690 435
rect -2730 255 -2720 425
rect -2700 255 -2690 425
rect -2730 245 -2690 255
rect -2645 425 -2605 435
rect -2645 255 -2635 425
rect -2615 255 -2605 425
rect -2645 245 -2605 255
rect -2565 425 -2525 435
rect -2565 255 -2555 425
rect -2535 255 -2525 425
rect -2565 245 -2525 255
rect -2500 425 -2460 435
rect -2500 255 -2490 425
rect -2470 255 -2460 425
rect -2430 415 -2420 435
rect -2400 415 -2390 435
rect -2430 405 -2390 415
rect -2500 245 -2460 255
rect -2710 200 -2690 245
rect -2710 190 -2670 200
rect -2710 170 -2700 190
rect -2680 170 -2670 190
rect -2710 160 -2670 170
rect -2710 105 -2690 160
rect -3020 95 -2980 105
rect -3090 40 -3050 50
rect -3090 20 -3080 40
rect -3060 20 -3050 40
rect -3090 10 -3050 20
rect -3020 25 -3010 95
rect -2990 25 -2980 95
rect -3020 15 -2980 25
rect -2955 95 -2915 105
rect -2955 25 -2945 95
rect -2925 25 -2915 95
rect -2955 15 -2915 25
rect -2875 95 -2835 105
rect -2875 25 -2865 95
rect -2845 25 -2835 95
rect -2875 15 -2835 25
rect -2795 95 -2755 105
rect -2795 25 -2785 95
rect -2765 25 -2755 95
rect -2795 15 -2755 25
rect -2730 95 -2690 105
rect -2730 25 -2720 95
rect -2700 25 -2690 95
rect -2730 15 -2690 25
rect -2635 50 -2615 245
rect -2555 200 -2535 245
rect -2490 200 -2470 245
rect -2565 190 -2525 200
rect -2565 170 -2555 190
rect -2535 170 -2525 190
rect -2565 160 -2525 170
rect -2500 190 -2460 200
rect -2500 170 -2490 190
rect -2470 170 -2460 190
rect -2500 160 -2460 170
rect -2555 105 -2535 160
rect -2490 105 -2470 160
rect -2410 105 -2390 405
rect -2335 425 -2295 435
rect -2335 255 -2325 425
rect -2305 255 -2295 425
rect -2335 245 -2295 255
rect -2270 425 -2230 435
rect -2270 255 -2260 425
rect -2240 255 -2230 425
rect -2270 245 -2230 255
rect -2185 425 -2145 435
rect -2185 255 -2175 425
rect -2155 255 -2145 425
rect -2185 245 -2145 255
rect -2105 425 -2065 435
rect -2105 255 -2095 425
rect -2075 255 -2065 425
rect -2105 245 -2065 255
rect -2040 425 -2000 435
rect -2040 255 -2030 425
rect -2010 255 -2000 425
rect -1970 425 -1930 435
rect -1970 405 -1960 425
rect -1940 405 -1930 425
rect -1970 395 -1930 405
rect -2040 245 -2000 255
rect -2315 190 -2275 200
rect -2315 170 -2305 190
rect -2285 170 -2275 190
rect -2315 160 -2275 170
rect -2250 105 -2230 245
rect -2565 95 -2525 105
rect -2635 40 -2595 50
rect -2635 20 -2625 40
rect -2605 20 -2595 40
rect -2635 10 -2595 20
rect -2565 25 -2555 95
rect -2535 25 -2525 95
rect -2565 15 -2525 25
rect -2500 95 -2460 105
rect -2500 25 -2490 95
rect -2470 25 -2460 95
rect -2500 15 -2460 25
rect -2420 95 -2380 105
rect -2420 25 -2410 95
rect -2390 25 -2380 95
rect -2420 15 -2380 25
rect -2335 95 -2295 105
rect -2335 25 -2325 95
rect -2305 25 -2295 95
rect -2335 15 -2295 25
rect -2270 95 -2230 105
rect -2270 25 -2260 95
rect -2240 25 -2230 95
rect -2270 15 -2230 25
rect -2250 -50 -2230 15
rect -2175 50 -2155 245
rect -2095 105 -2075 245
rect -2030 105 -2010 245
rect -1950 105 -1930 395
rect -1875 425 -1835 435
rect -1875 255 -1865 425
rect -1845 255 -1835 425
rect -1875 245 -1835 255
rect -1810 425 -1770 435
rect -1810 255 -1800 425
rect -1780 255 -1770 425
rect -1810 245 -1770 255
rect -670 250 -660 1020
rect -640 250 -630 1020
rect -670 240 -630 250
rect -560 1020 -470 1030
rect -560 250 -550 1020
rect -530 250 -500 1020
rect -480 250 -470 1020
rect -560 240 -470 250
rect -220 1020 -130 1030
rect -220 250 -210 1020
rect -190 250 -160 1020
rect -140 250 -130 1020
rect -220 240 -130 250
rect -60 1020 -20 1030
rect -60 250 -50 1020
rect -30 250 -20 1020
rect 590 890 645 900
rect 590 855 600 890
rect 635 855 645 890
rect 590 845 645 855
rect 590 295 645 305
rect 590 260 600 295
rect 635 260 645 295
rect 590 250 645 260
rect -60 240 -20 250
rect -1170 180 -1130 190
rect -1170 160 -1160 180
rect -1140 160 -1130 180
rect -1170 150 -1130 160
rect -1160 130 -1140 150
rect -660 130 -640 240
rect -50 185 -30 240
rect -50 165 1325 185
rect -50 130 -30 165
rect -1170 120 -1130 130
rect -2105 95 -2065 105
rect -2175 40 -2135 50
rect -2175 20 -2165 40
rect -2145 20 -2135 40
rect -2175 10 -2135 20
rect -2105 25 -2095 95
rect -2075 25 -2065 95
rect -2105 15 -2065 25
rect -2040 95 -1995 105
rect -2040 25 -2030 95
rect -2010 25 -1995 95
rect -2040 15 -1995 25
rect -1965 95 -1920 105
rect -1965 25 -1950 95
rect -1930 25 -1920 95
rect -1965 15 -1920 25
rect -1875 95 -1835 105
rect -1875 25 -1865 95
rect -1845 25 -1835 95
rect -1875 15 -1835 25
rect -1810 95 -1770 105
rect -1810 25 -1800 95
rect -1780 25 -1770 95
rect -1810 15 -1770 25
rect -2250 -60 -2210 -50
rect -2250 -80 -2240 -60
rect -2220 -80 -2210 -60
rect -2250 -90 -2210 -80
rect -2095 -95 -2075 15
rect -2020 -5 -2000 15
rect -1865 -5 -1845 15
rect -2020 -25 -1845 -5
rect -2020 -55 -2000 -25
rect -2020 -65 -1980 -55
rect -2020 -85 -2010 -65
rect -1990 -85 -1980 -65
rect -2020 -95 -1980 -85
rect -2105 -105 -2065 -95
rect -2105 -125 -2095 -105
rect -2075 -125 -2065 -105
rect -2105 -135 -2065 -125
rect -1170 -210 -1160 120
rect -3565 -230 -1160 -210
rect -1170 -250 -1160 -230
rect -1140 -250 -1130 120
rect -1170 -260 -1130 -250
rect -1060 120 -970 130
rect -1060 -250 -1050 120
rect -1030 -250 -1000 120
rect -980 -250 -970 120
rect -1060 -260 -970 -250
rect -670 120 -630 130
rect -670 -250 -660 120
rect -640 -250 -630 120
rect -670 -260 -630 -250
rect -560 120 -470 130
rect -560 -250 -550 120
rect -530 -250 -500 120
rect -480 -250 -470 120
rect -560 -260 -470 -250
rect -220 120 -130 130
rect -220 -250 -210 120
rect -190 -250 -160 120
rect -140 -250 -130 120
rect -220 -260 -130 -250
rect -60 120 -20 130
rect -60 -250 -50 120
rect -30 -250 -20 120
rect 590 90 645 100
rect 590 55 600 90
rect 635 55 645 90
rect 590 45 645 55
rect 590 -130 645 -120
rect 590 -165 600 -130
rect 635 -165 645 -130
rect 590 -175 645 -165
rect -60 -260 -20 -250
<< viali >>
rect -3535 255 -3515 425
rect -3385 255 -3365 425
rect -3235 255 -3215 425
rect -2875 410 -2855 430
rect -3535 25 -3515 95
rect -3385 25 -3365 95
rect -3235 25 -3215 95
rect -2785 255 -2765 425
rect -2420 415 -2400 435
rect -3080 20 -3060 40
rect -2785 25 -2765 95
rect -2325 255 -2305 425
rect -1960 405 -1940 425
rect -2625 20 -2605 40
rect -2325 25 -2305 95
rect -1800 255 -1780 425
rect -550 250 -530 1020
rect -500 250 -480 1020
rect -210 250 -190 1020
rect -160 250 -140 1020
rect 600 855 635 890
rect 600 260 635 295
rect -2165 20 -2145 40
rect -1800 25 -1780 95
rect -1050 -250 -1030 120
rect -1000 -250 -980 120
rect -550 -250 -530 120
rect -500 -250 -480 120
rect -210 -250 -190 120
rect -160 -250 -140 120
rect 600 55 635 90
rect 600 -165 635 -130
<< metal1 >>
rect -1550 1020 -15 1035
rect -1550 440 -550 1020
rect -3600 435 -550 440
rect -3600 430 -2420 435
rect -3600 425 -2875 430
rect -3600 255 -3535 425
rect -3515 255 -3385 425
rect -3365 255 -3235 425
rect -3215 410 -2875 425
rect -2855 425 -2420 430
rect -2855 410 -2785 425
rect -3215 255 -2785 410
rect -2765 415 -2420 425
rect -2400 425 -550 435
rect -2400 415 -2325 425
rect -2765 255 -2325 415
rect -2305 405 -1960 425
rect -1940 405 -1800 425
rect -2305 255 -1800 405
rect -1780 255 -550 425
rect -3600 250 -550 255
rect -530 250 -500 1020
rect -480 250 -210 1020
rect -190 250 -160 1020
rect -140 250 -15 1020
rect 590 890 645 900
rect 590 855 600 890
rect 635 855 645 890
rect 590 845 645 855
rect 590 295 645 305
rect 590 260 600 295
rect 635 260 645 295
rect 590 250 645 260
rect -3600 240 -15 250
rect -1555 235 -15 240
rect -1545 120 -15 135
rect -1545 110 -1050 120
rect -3600 95 -1050 110
rect -3600 25 -3535 95
rect -3515 25 -3385 95
rect -3365 25 -3235 95
rect -3215 40 -2785 95
rect -3215 25 -3080 40
rect -3600 20 -3080 25
rect -3060 25 -2785 40
rect -2765 40 -2325 95
rect -2765 25 -2625 40
rect -3060 20 -2625 25
rect -2605 25 -2325 40
rect -2305 40 -1800 95
rect -2305 25 -2165 40
rect -2605 20 -2165 25
rect -2145 25 -1800 40
rect -1780 25 -1050 95
rect -2145 20 -1050 25
rect -3600 0 -1050 20
rect -1545 -250 -1050 0
rect -1030 -250 -1000 120
rect -980 -250 -550 120
rect -530 -250 -500 120
rect -480 -250 -210 120
rect -190 -250 -160 120
rect -140 -250 -15 120
rect 590 90 645 100
rect 590 55 600 90
rect 635 55 645 90
rect 590 45 645 55
rect 590 -130 645 -120
rect 590 -165 600 -130
rect 635 -165 645 -130
rect 590 -175 645 -165
rect -1545 -265 -15 -250
<< via1 >>
rect 600 855 635 890
rect 600 260 635 295
rect 600 55 635 90
rect 600 -165 635 -130
<< metal2 >>
rect 590 890 645 900
rect 590 855 600 890
rect 635 855 645 890
rect 590 845 645 855
rect 590 295 645 305
rect 590 260 600 295
rect 635 260 645 295
rect 590 250 645 260
rect 590 90 645 100
rect 590 55 600 90
rect 635 55 645 90
rect 590 45 645 55
rect 590 -130 645 -120
rect 590 -165 600 -130
rect 635 -165 645 -130
rect 590 -175 645 -165
<< via2 >>
rect 600 855 635 890
rect 600 260 635 295
rect 600 55 635 90
rect 600 -165 635 -130
<< metal3 >>
rect 765 900 1215 925
rect 590 890 1215 900
rect 590 855 600 890
rect 635 855 1215 890
rect 590 845 1215 855
rect 765 305 1215 845
rect 590 295 1215 305
rect 590 260 600 295
rect 635 260 1215 295
rect 590 250 1215 260
rect 765 235 1215 250
rect 765 100 1055 115
rect 590 90 1055 100
rect 590 55 600 90
rect 635 55 1055 90
rect 590 45 1055 55
rect 765 -120 1055 45
rect 590 -130 1055 -120
rect 590 -165 600 -130
rect 635 -165 1055 -130
rect 590 -175 1055 -165
<< via3 >>
rect 600 260 635 295
rect 600 55 635 90
<< mimcap >>
rect 780 295 1200 910
rect 780 260 790 295
rect 825 260 1200 295
rect 780 250 1200 260
rect 780 90 1040 100
rect 780 55 790 90
rect 825 55 1040 90
rect 780 -160 1040 55
<< mimcapcontact >>
rect 790 260 825 295
rect 790 55 825 90
<< metal4 >>
rect 590 295 645 305
rect 590 260 600 295
rect 635 260 645 295
rect 590 250 645 260
rect 780 295 835 305
rect 780 260 790 295
rect 825 260 835 295
rect 780 250 835 260
rect 590 90 645 100
rect 590 55 600 90
rect 635 55 645 90
rect 590 45 645 55
rect 780 90 835 100
rect 780 55 790 90
rect 825 55 835 90
rect 780 45 835 55
<< labels >>
flabel locali 1325 175 1325 175 3 FreeSans 400 0 80 0 VOUT
flabel locali -3565 -220 -3565 -220 7 FreeSans 400 0 -200 0 I_IN
flabel poly -3565 -125 -3565 -125 7 FreeSans 400 0 -200 0 DOWN_PFD
flabel poly -3565 175 -3565 175 7 FreeSans 400 0 -200 0 UP_PFD
flabel metal1 -3600 340 -3600 340 7 FreeSans 400 0 -200 0 VDDA
flabel metal1 -3600 60 -3600 60 7 FreeSans 400 0 -200 0 GNDA
<< end >>
