* SPICE3 file created from pnp.ext - technology: sky130A

X0 GND GND EMITTER sky130_fd_pr__pnp_05v5_W0p68L0p68
X1 GND GND EMITTER sky130_fd_pr__pnp_05v5_W0p68L0p68
