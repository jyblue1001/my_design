magic
tech sky130A
timestamp 1748714285
<< error_p >>
rect -975 -940 -972 -937
rect -970 -940 -964 -939
rect -978 -943 -975 -940
rect -976 -951 -975 -945
rect -976 -970 -975 -964
rect -978 -975 -975 -972
rect -975 -978 -972 -975
rect -970 -976 -964 -975
<< pwell >>
rect 4545 2790 4765 2890
rect 4795 2790 6635 2890
rect 4400 2400 6780 2700
rect 4155 1850 4305 1950
rect 4335 1850 5575 1950
rect 5605 1850 6845 1950
rect -45 1685 130 1725
rect 4755 1565 5395 1615
rect 5785 1565 6425 1615
rect 4425 1160 5545 1410
rect 5635 1160 6755 1410
rect 4530 965 6650 1065
rect 4680 810 4810 910
rect 4840 810 6590 910
<< nmos >>
rect 4585 2790 4635 2890
rect 4675 2790 4725 2890
rect 4835 2790 4885 2890
rect 4925 2790 4975 2890
rect 5015 2790 5065 2890
rect 5105 2790 5155 2890
rect 5195 2790 5245 2890
rect 5285 2790 5335 2890
rect 5375 2790 5425 2890
rect 5465 2790 5515 2890
rect 5555 2790 5605 2890
rect 5645 2790 5695 2890
rect 5735 2790 5785 2890
rect 5825 2790 5875 2890
rect 5915 2790 5965 2890
rect 6005 2790 6055 2890
rect 6095 2790 6145 2890
rect 6185 2790 6235 2890
rect 6275 2790 6325 2890
rect 6365 2790 6415 2890
rect 6455 2790 6505 2890
rect 6545 2790 6595 2890
rect 4440 2400 4490 2700
rect 4530 2400 4580 2700
rect 4620 2400 4670 2700
rect 4710 2400 4760 2700
rect 4800 2400 4850 2700
rect 4890 2400 4940 2700
rect 4980 2400 5030 2700
rect 5070 2400 5120 2700
rect 5160 2400 5210 2700
rect 5250 2400 5300 2700
rect 5340 2400 5390 2700
rect 5430 2400 5480 2700
rect 5520 2400 5570 2700
rect 5610 2400 5660 2700
rect 5700 2400 5750 2700
rect 5790 2400 5840 2700
rect 5880 2400 5930 2700
rect 5970 2400 6020 2700
rect 6060 2400 6110 2700
rect 6150 2400 6200 2700
rect 6240 2400 6290 2700
rect 6330 2400 6380 2700
rect 6420 2400 6470 2700
rect 6510 2400 6560 2700
rect 6600 2400 6650 2700
rect 6690 2400 6740 2700
rect 4195 1850 4210 1950
rect 4250 1850 4265 1950
rect 4375 1850 4395 1950
rect 4435 1850 4455 1950
rect 4495 1850 4515 1950
rect 4555 1850 4575 1950
rect 4615 1850 4635 1950
rect 4675 1850 4695 1950
rect 4735 1850 4755 1950
rect 4795 1850 4815 1950
rect 4855 1850 4875 1950
rect 4915 1850 4935 1950
rect 4975 1850 4995 1950
rect 5035 1850 5055 1950
rect 5095 1850 5115 1950
rect 5155 1850 5175 1950
rect 5215 1850 5235 1950
rect 5275 1850 5295 1950
rect 5335 1850 5355 1950
rect 5395 1850 5415 1950
rect 5455 1850 5475 1950
rect 5515 1850 5535 1950
rect 5645 1850 5665 1950
rect 5705 1850 5725 1950
rect 5765 1850 5785 1950
rect 5825 1850 5845 1950
rect 5885 1850 5905 1950
rect 5945 1850 5965 1950
rect 6005 1850 6025 1950
rect 6065 1850 6085 1950
rect 6125 1850 6145 1950
rect 6185 1850 6205 1950
rect 6245 1850 6265 1950
rect 6305 1850 6325 1950
rect 6365 1850 6385 1950
rect 6425 1850 6445 1950
rect 6485 1850 6505 1950
rect 6545 1850 6565 1950
rect 6605 1850 6625 1950
rect 6665 1850 6685 1950
rect 6725 1850 6745 1950
rect 6785 1850 6805 1950
rect 4795 1565 4815 1615
rect 4855 1565 4875 1615
rect 4915 1565 4935 1615
rect 4975 1565 4995 1615
rect 5035 1565 5055 1615
rect 5095 1565 5115 1615
rect 5155 1565 5175 1615
rect 5215 1565 5235 1615
rect 5275 1565 5295 1615
rect 5335 1565 5355 1615
rect 5825 1565 5845 1615
rect 5885 1565 5905 1615
rect 5945 1565 5965 1615
rect 6005 1565 6025 1615
rect 6065 1565 6085 1615
rect 6125 1565 6145 1615
rect 6185 1565 6205 1615
rect 6245 1565 6265 1615
rect 6305 1565 6325 1615
rect 6365 1565 6385 1615
rect 4465 1160 4965 1410
rect 5005 1160 5505 1410
rect 5675 1160 6175 1410
rect 6215 1160 6715 1410
rect 4570 965 5570 1065
rect 5610 965 6610 1065
rect 4720 810 4770 910
rect 4880 810 4930 910
rect 4970 810 5020 910
rect 5060 810 5110 910
rect 5150 810 5200 910
rect 5240 810 5290 910
rect 5330 810 5380 910
rect 5420 810 5470 910
rect 5510 810 5560 910
rect 5600 810 5650 910
rect 5690 810 5740 910
rect 5780 810 5830 910
rect 5870 810 5920 910
rect 5960 810 6010 910
rect 6050 810 6100 910
rect 6140 810 6190 910
rect 6230 810 6280 910
rect 6320 810 6370 910
rect 6410 810 6460 910
rect 6500 810 6550 910
<< ndiff >>
rect 4545 2875 4585 2890
rect 4545 2855 4555 2875
rect 4575 2855 4585 2875
rect 4545 2825 4585 2855
rect 4545 2805 4555 2825
rect 4575 2805 4585 2825
rect 4545 2790 4585 2805
rect 4635 2875 4675 2890
rect 4635 2855 4645 2875
rect 4665 2855 4675 2875
rect 4635 2825 4675 2855
rect 4635 2805 4645 2825
rect 4665 2805 4675 2825
rect 4635 2790 4675 2805
rect 4725 2875 4765 2890
rect 4725 2855 4735 2875
rect 4755 2855 4765 2875
rect 4725 2825 4765 2855
rect 4725 2805 4735 2825
rect 4755 2805 4765 2825
rect 4725 2790 4765 2805
rect 4795 2875 4835 2890
rect 4795 2855 4805 2875
rect 4825 2855 4835 2875
rect 4795 2825 4835 2855
rect 4795 2805 4805 2825
rect 4825 2805 4835 2825
rect 4795 2790 4835 2805
rect 4885 2875 4925 2890
rect 4885 2855 4895 2875
rect 4915 2855 4925 2875
rect 4885 2825 4925 2855
rect 4885 2805 4895 2825
rect 4915 2805 4925 2825
rect 4885 2790 4925 2805
rect 4975 2875 5015 2890
rect 4975 2855 4985 2875
rect 5005 2855 5015 2875
rect 4975 2825 5015 2855
rect 4975 2805 4985 2825
rect 5005 2805 5015 2825
rect 4975 2790 5015 2805
rect 5065 2875 5105 2890
rect 5065 2855 5075 2875
rect 5095 2855 5105 2875
rect 5065 2825 5105 2855
rect 5065 2805 5075 2825
rect 5095 2805 5105 2825
rect 5065 2790 5105 2805
rect 5155 2875 5195 2890
rect 5155 2855 5165 2875
rect 5185 2855 5195 2875
rect 5155 2825 5195 2855
rect 5155 2805 5165 2825
rect 5185 2805 5195 2825
rect 5155 2790 5195 2805
rect 5245 2875 5285 2890
rect 5245 2855 5255 2875
rect 5275 2855 5285 2875
rect 5245 2825 5285 2855
rect 5245 2805 5255 2825
rect 5275 2805 5285 2825
rect 5245 2790 5285 2805
rect 5335 2875 5375 2890
rect 5335 2855 5345 2875
rect 5365 2855 5375 2875
rect 5335 2825 5375 2855
rect 5335 2805 5345 2825
rect 5365 2805 5375 2825
rect 5335 2790 5375 2805
rect 5425 2875 5465 2890
rect 5425 2855 5435 2875
rect 5455 2855 5465 2875
rect 5425 2825 5465 2855
rect 5425 2805 5435 2825
rect 5455 2805 5465 2825
rect 5425 2790 5465 2805
rect 5515 2875 5555 2890
rect 5515 2855 5525 2875
rect 5545 2855 5555 2875
rect 5515 2825 5555 2855
rect 5515 2805 5525 2825
rect 5545 2805 5555 2825
rect 5515 2790 5555 2805
rect 5605 2875 5645 2890
rect 5605 2855 5615 2875
rect 5635 2855 5645 2875
rect 5605 2825 5645 2855
rect 5605 2805 5615 2825
rect 5635 2805 5645 2825
rect 5605 2790 5645 2805
rect 5695 2875 5735 2890
rect 5695 2855 5705 2875
rect 5725 2855 5735 2875
rect 5695 2825 5735 2855
rect 5695 2805 5705 2825
rect 5725 2805 5735 2825
rect 5695 2790 5735 2805
rect 5785 2875 5825 2890
rect 5785 2855 5795 2875
rect 5815 2855 5825 2875
rect 5785 2825 5825 2855
rect 5785 2805 5795 2825
rect 5815 2805 5825 2825
rect 5785 2790 5825 2805
rect 5875 2875 5915 2890
rect 5875 2855 5885 2875
rect 5905 2855 5915 2875
rect 5875 2825 5915 2855
rect 5875 2805 5885 2825
rect 5905 2805 5915 2825
rect 5875 2790 5915 2805
rect 5965 2875 6005 2890
rect 5965 2855 5975 2875
rect 5995 2855 6005 2875
rect 5965 2825 6005 2855
rect 5965 2805 5975 2825
rect 5995 2805 6005 2825
rect 5965 2790 6005 2805
rect 6055 2875 6095 2890
rect 6055 2855 6065 2875
rect 6085 2855 6095 2875
rect 6055 2825 6095 2855
rect 6055 2805 6065 2825
rect 6085 2805 6095 2825
rect 6055 2790 6095 2805
rect 6145 2875 6185 2890
rect 6145 2855 6155 2875
rect 6175 2855 6185 2875
rect 6145 2825 6185 2855
rect 6145 2805 6155 2825
rect 6175 2805 6185 2825
rect 6145 2790 6185 2805
rect 6235 2875 6275 2890
rect 6235 2855 6245 2875
rect 6265 2855 6275 2875
rect 6235 2825 6275 2855
rect 6235 2805 6245 2825
rect 6265 2805 6275 2825
rect 6235 2790 6275 2805
rect 6325 2875 6365 2890
rect 6325 2855 6335 2875
rect 6355 2855 6365 2875
rect 6325 2825 6365 2855
rect 6325 2805 6335 2825
rect 6355 2805 6365 2825
rect 6325 2790 6365 2805
rect 6415 2875 6455 2890
rect 6415 2855 6425 2875
rect 6445 2855 6455 2875
rect 6415 2825 6455 2855
rect 6415 2805 6425 2825
rect 6445 2805 6455 2825
rect 6415 2790 6455 2805
rect 6505 2875 6545 2890
rect 6505 2855 6515 2875
rect 6535 2855 6545 2875
rect 6505 2825 6545 2855
rect 6505 2805 6515 2825
rect 6535 2805 6545 2825
rect 6505 2790 6545 2805
rect 6595 2875 6635 2890
rect 6595 2855 6605 2875
rect 6625 2855 6635 2875
rect 6595 2825 6635 2855
rect 6595 2805 6605 2825
rect 6625 2805 6635 2825
rect 6595 2790 6635 2805
rect 4400 2685 4440 2700
rect 4400 2665 4410 2685
rect 4430 2665 4440 2685
rect 4400 2635 4440 2665
rect 4400 2615 4410 2635
rect 4430 2615 4440 2635
rect 4400 2585 4440 2615
rect 4400 2565 4410 2585
rect 4430 2565 4440 2585
rect 4400 2535 4440 2565
rect 4400 2515 4410 2535
rect 4430 2515 4440 2535
rect 4400 2485 4440 2515
rect 4400 2465 4410 2485
rect 4430 2465 4440 2485
rect 4400 2435 4440 2465
rect 4400 2415 4410 2435
rect 4430 2415 4440 2435
rect 4400 2400 4440 2415
rect 4490 2685 4530 2700
rect 4490 2665 4500 2685
rect 4520 2665 4530 2685
rect 4490 2635 4530 2665
rect 4490 2615 4500 2635
rect 4520 2615 4530 2635
rect 4490 2585 4530 2615
rect 4490 2565 4500 2585
rect 4520 2565 4530 2585
rect 4490 2535 4530 2565
rect 4490 2515 4500 2535
rect 4520 2515 4530 2535
rect 4490 2485 4530 2515
rect 4490 2465 4500 2485
rect 4520 2465 4530 2485
rect 4490 2435 4530 2465
rect 4490 2415 4500 2435
rect 4520 2415 4530 2435
rect 4490 2400 4530 2415
rect 4580 2685 4620 2700
rect 4580 2665 4590 2685
rect 4610 2665 4620 2685
rect 4580 2635 4620 2665
rect 4580 2615 4590 2635
rect 4610 2615 4620 2635
rect 4580 2585 4620 2615
rect 4580 2565 4590 2585
rect 4610 2565 4620 2585
rect 4580 2535 4620 2565
rect 4580 2515 4590 2535
rect 4610 2515 4620 2535
rect 4580 2485 4620 2515
rect 4580 2465 4590 2485
rect 4610 2465 4620 2485
rect 4580 2435 4620 2465
rect 4580 2415 4590 2435
rect 4610 2415 4620 2435
rect 4580 2400 4620 2415
rect 4670 2685 4710 2700
rect 4670 2665 4680 2685
rect 4700 2665 4710 2685
rect 4670 2635 4710 2665
rect 4670 2615 4680 2635
rect 4700 2615 4710 2635
rect 4670 2585 4710 2615
rect 4670 2565 4680 2585
rect 4700 2565 4710 2585
rect 4670 2535 4710 2565
rect 4670 2515 4680 2535
rect 4700 2515 4710 2535
rect 4670 2485 4710 2515
rect 4670 2465 4680 2485
rect 4700 2465 4710 2485
rect 4670 2435 4710 2465
rect 4670 2415 4680 2435
rect 4700 2415 4710 2435
rect 4670 2400 4710 2415
rect 4760 2685 4800 2700
rect 4760 2665 4770 2685
rect 4790 2665 4800 2685
rect 4760 2635 4800 2665
rect 4760 2615 4770 2635
rect 4790 2615 4800 2635
rect 4760 2585 4800 2615
rect 4760 2565 4770 2585
rect 4790 2565 4800 2585
rect 4760 2535 4800 2565
rect 4760 2515 4770 2535
rect 4790 2515 4800 2535
rect 4760 2485 4800 2515
rect 4760 2465 4770 2485
rect 4790 2465 4800 2485
rect 4760 2435 4800 2465
rect 4760 2415 4770 2435
rect 4790 2415 4800 2435
rect 4760 2400 4800 2415
rect 4850 2685 4890 2700
rect 4850 2665 4860 2685
rect 4880 2665 4890 2685
rect 4850 2635 4890 2665
rect 4850 2615 4860 2635
rect 4880 2615 4890 2635
rect 4850 2585 4890 2615
rect 4850 2565 4860 2585
rect 4880 2565 4890 2585
rect 4850 2535 4890 2565
rect 4850 2515 4860 2535
rect 4880 2515 4890 2535
rect 4850 2485 4890 2515
rect 4850 2465 4860 2485
rect 4880 2465 4890 2485
rect 4850 2435 4890 2465
rect 4850 2415 4860 2435
rect 4880 2415 4890 2435
rect 4850 2400 4890 2415
rect 4940 2685 4980 2700
rect 4940 2665 4950 2685
rect 4970 2665 4980 2685
rect 4940 2635 4980 2665
rect 4940 2615 4950 2635
rect 4970 2615 4980 2635
rect 4940 2585 4980 2615
rect 4940 2565 4950 2585
rect 4970 2565 4980 2585
rect 4940 2535 4980 2565
rect 4940 2515 4950 2535
rect 4970 2515 4980 2535
rect 4940 2485 4980 2515
rect 4940 2465 4950 2485
rect 4970 2465 4980 2485
rect 4940 2435 4980 2465
rect 4940 2415 4950 2435
rect 4970 2415 4980 2435
rect 4940 2400 4980 2415
rect 5030 2685 5070 2700
rect 5030 2665 5040 2685
rect 5060 2665 5070 2685
rect 5030 2635 5070 2665
rect 5030 2615 5040 2635
rect 5060 2615 5070 2635
rect 5030 2585 5070 2615
rect 5030 2565 5040 2585
rect 5060 2565 5070 2585
rect 5030 2535 5070 2565
rect 5030 2515 5040 2535
rect 5060 2515 5070 2535
rect 5030 2485 5070 2515
rect 5030 2465 5040 2485
rect 5060 2465 5070 2485
rect 5030 2435 5070 2465
rect 5030 2415 5040 2435
rect 5060 2415 5070 2435
rect 5030 2400 5070 2415
rect 5120 2685 5160 2700
rect 5120 2665 5130 2685
rect 5150 2665 5160 2685
rect 5120 2635 5160 2665
rect 5120 2615 5130 2635
rect 5150 2615 5160 2635
rect 5120 2585 5160 2615
rect 5120 2565 5130 2585
rect 5150 2565 5160 2585
rect 5120 2535 5160 2565
rect 5120 2515 5130 2535
rect 5150 2515 5160 2535
rect 5120 2485 5160 2515
rect 5120 2465 5130 2485
rect 5150 2465 5160 2485
rect 5120 2435 5160 2465
rect 5120 2415 5130 2435
rect 5150 2415 5160 2435
rect 5120 2400 5160 2415
rect 5210 2685 5250 2700
rect 5210 2665 5220 2685
rect 5240 2665 5250 2685
rect 5210 2635 5250 2665
rect 5210 2615 5220 2635
rect 5240 2615 5250 2635
rect 5210 2585 5250 2615
rect 5210 2565 5220 2585
rect 5240 2565 5250 2585
rect 5210 2535 5250 2565
rect 5210 2515 5220 2535
rect 5240 2515 5250 2535
rect 5210 2485 5250 2515
rect 5210 2465 5220 2485
rect 5240 2465 5250 2485
rect 5210 2435 5250 2465
rect 5210 2415 5220 2435
rect 5240 2415 5250 2435
rect 5210 2400 5250 2415
rect 5300 2685 5340 2700
rect 5300 2665 5310 2685
rect 5330 2665 5340 2685
rect 5300 2635 5340 2665
rect 5300 2615 5310 2635
rect 5330 2615 5340 2635
rect 5300 2585 5340 2615
rect 5300 2565 5310 2585
rect 5330 2565 5340 2585
rect 5300 2535 5340 2565
rect 5300 2515 5310 2535
rect 5330 2515 5340 2535
rect 5300 2485 5340 2515
rect 5300 2465 5310 2485
rect 5330 2465 5340 2485
rect 5300 2435 5340 2465
rect 5300 2415 5310 2435
rect 5330 2415 5340 2435
rect 5300 2400 5340 2415
rect 5390 2685 5430 2700
rect 5390 2665 5400 2685
rect 5420 2665 5430 2685
rect 5390 2635 5430 2665
rect 5390 2615 5400 2635
rect 5420 2615 5430 2635
rect 5390 2585 5430 2615
rect 5390 2565 5400 2585
rect 5420 2565 5430 2585
rect 5390 2535 5430 2565
rect 5390 2515 5400 2535
rect 5420 2515 5430 2535
rect 5390 2485 5430 2515
rect 5390 2465 5400 2485
rect 5420 2465 5430 2485
rect 5390 2435 5430 2465
rect 5390 2415 5400 2435
rect 5420 2415 5430 2435
rect 5390 2400 5430 2415
rect 5480 2685 5520 2700
rect 5480 2665 5490 2685
rect 5510 2665 5520 2685
rect 5480 2635 5520 2665
rect 5480 2615 5490 2635
rect 5510 2615 5520 2635
rect 5480 2585 5520 2615
rect 5480 2565 5490 2585
rect 5510 2565 5520 2585
rect 5480 2535 5520 2565
rect 5480 2515 5490 2535
rect 5510 2515 5520 2535
rect 5480 2485 5520 2515
rect 5480 2465 5490 2485
rect 5510 2465 5520 2485
rect 5480 2435 5520 2465
rect 5480 2415 5490 2435
rect 5510 2415 5520 2435
rect 5480 2400 5520 2415
rect 5570 2685 5610 2700
rect 5570 2665 5580 2685
rect 5600 2665 5610 2685
rect 5570 2635 5610 2665
rect 5570 2615 5580 2635
rect 5600 2615 5610 2635
rect 5570 2585 5610 2615
rect 5570 2565 5580 2585
rect 5600 2565 5610 2585
rect 5570 2535 5610 2565
rect 5570 2515 5580 2535
rect 5600 2515 5610 2535
rect 5570 2485 5610 2515
rect 5570 2465 5580 2485
rect 5600 2465 5610 2485
rect 5570 2435 5610 2465
rect 5570 2415 5580 2435
rect 5600 2415 5610 2435
rect 5570 2400 5610 2415
rect 5660 2685 5700 2700
rect 5660 2665 5670 2685
rect 5690 2665 5700 2685
rect 5660 2635 5700 2665
rect 5660 2615 5670 2635
rect 5690 2615 5700 2635
rect 5660 2585 5700 2615
rect 5660 2565 5670 2585
rect 5690 2565 5700 2585
rect 5660 2535 5700 2565
rect 5660 2515 5670 2535
rect 5690 2515 5700 2535
rect 5660 2485 5700 2515
rect 5660 2465 5670 2485
rect 5690 2465 5700 2485
rect 5660 2435 5700 2465
rect 5660 2415 5670 2435
rect 5690 2415 5700 2435
rect 5660 2400 5700 2415
rect 5750 2685 5790 2700
rect 5750 2665 5760 2685
rect 5780 2665 5790 2685
rect 5750 2635 5790 2665
rect 5750 2615 5760 2635
rect 5780 2615 5790 2635
rect 5750 2585 5790 2615
rect 5750 2565 5760 2585
rect 5780 2565 5790 2585
rect 5750 2535 5790 2565
rect 5750 2515 5760 2535
rect 5780 2515 5790 2535
rect 5750 2485 5790 2515
rect 5750 2465 5760 2485
rect 5780 2465 5790 2485
rect 5750 2435 5790 2465
rect 5750 2415 5760 2435
rect 5780 2415 5790 2435
rect 5750 2400 5790 2415
rect 5840 2685 5880 2700
rect 5840 2665 5850 2685
rect 5870 2665 5880 2685
rect 5840 2635 5880 2665
rect 5840 2615 5850 2635
rect 5870 2615 5880 2635
rect 5840 2585 5880 2615
rect 5840 2565 5850 2585
rect 5870 2565 5880 2585
rect 5840 2535 5880 2565
rect 5840 2515 5850 2535
rect 5870 2515 5880 2535
rect 5840 2485 5880 2515
rect 5840 2465 5850 2485
rect 5870 2465 5880 2485
rect 5840 2435 5880 2465
rect 5840 2415 5850 2435
rect 5870 2415 5880 2435
rect 5840 2400 5880 2415
rect 5930 2685 5970 2700
rect 5930 2665 5940 2685
rect 5960 2665 5970 2685
rect 5930 2635 5970 2665
rect 5930 2615 5940 2635
rect 5960 2615 5970 2635
rect 5930 2585 5970 2615
rect 5930 2565 5940 2585
rect 5960 2565 5970 2585
rect 5930 2535 5970 2565
rect 5930 2515 5940 2535
rect 5960 2515 5970 2535
rect 5930 2485 5970 2515
rect 5930 2465 5940 2485
rect 5960 2465 5970 2485
rect 5930 2435 5970 2465
rect 5930 2415 5940 2435
rect 5960 2415 5970 2435
rect 5930 2400 5970 2415
rect 6020 2685 6060 2700
rect 6020 2665 6030 2685
rect 6050 2665 6060 2685
rect 6020 2635 6060 2665
rect 6020 2615 6030 2635
rect 6050 2615 6060 2635
rect 6020 2585 6060 2615
rect 6020 2565 6030 2585
rect 6050 2565 6060 2585
rect 6020 2535 6060 2565
rect 6020 2515 6030 2535
rect 6050 2515 6060 2535
rect 6020 2485 6060 2515
rect 6020 2465 6030 2485
rect 6050 2465 6060 2485
rect 6020 2435 6060 2465
rect 6020 2415 6030 2435
rect 6050 2415 6060 2435
rect 6020 2400 6060 2415
rect 6110 2685 6150 2700
rect 6110 2665 6120 2685
rect 6140 2665 6150 2685
rect 6110 2635 6150 2665
rect 6110 2615 6120 2635
rect 6140 2615 6150 2635
rect 6110 2585 6150 2615
rect 6110 2565 6120 2585
rect 6140 2565 6150 2585
rect 6110 2535 6150 2565
rect 6110 2515 6120 2535
rect 6140 2515 6150 2535
rect 6110 2485 6150 2515
rect 6110 2465 6120 2485
rect 6140 2465 6150 2485
rect 6110 2435 6150 2465
rect 6110 2415 6120 2435
rect 6140 2415 6150 2435
rect 6110 2400 6150 2415
rect 6200 2685 6240 2700
rect 6200 2665 6210 2685
rect 6230 2665 6240 2685
rect 6200 2635 6240 2665
rect 6200 2615 6210 2635
rect 6230 2615 6240 2635
rect 6200 2585 6240 2615
rect 6200 2565 6210 2585
rect 6230 2565 6240 2585
rect 6200 2535 6240 2565
rect 6200 2515 6210 2535
rect 6230 2515 6240 2535
rect 6200 2485 6240 2515
rect 6200 2465 6210 2485
rect 6230 2465 6240 2485
rect 6200 2435 6240 2465
rect 6200 2415 6210 2435
rect 6230 2415 6240 2435
rect 6200 2400 6240 2415
rect 6290 2685 6330 2700
rect 6290 2665 6300 2685
rect 6320 2665 6330 2685
rect 6290 2635 6330 2665
rect 6290 2615 6300 2635
rect 6320 2615 6330 2635
rect 6290 2585 6330 2615
rect 6290 2565 6300 2585
rect 6320 2565 6330 2585
rect 6290 2535 6330 2565
rect 6290 2515 6300 2535
rect 6320 2515 6330 2535
rect 6290 2485 6330 2515
rect 6290 2465 6300 2485
rect 6320 2465 6330 2485
rect 6290 2435 6330 2465
rect 6290 2415 6300 2435
rect 6320 2415 6330 2435
rect 6290 2400 6330 2415
rect 6380 2685 6420 2700
rect 6380 2665 6390 2685
rect 6410 2665 6420 2685
rect 6380 2635 6420 2665
rect 6380 2615 6390 2635
rect 6410 2615 6420 2635
rect 6380 2585 6420 2615
rect 6380 2565 6390 2585
rect 6410 2565 6420 2585
rect 6380 2535 6420 2565
rect 6380 2515 6390 2535
rect 6410 2515 6420 2535
rect 6380 2485 6420 2515
rect 6380 2465 6390 2485
rect 6410 2465 6420 2485
rect 6380 2435 6420 2465
rect 6380 2415 6390 2435
rect 6410 2415 6420 2435
rect 6380 2400 6420 2415
rect 6470 2685 6510 2700
rect 6470 2665 6480 2685
rect 6500 2665 6510 2685
rect 6470 2635 6510 2665
rect 6470 2615 6480 2635
rect 6500 2615 6510 2635
rect 6470 2585 6510 2615
rect 6470 2565 6480 2585
rect 6500 2565 6510 2585
rect 6470 2535 6510 2565
rect 6470 2515 6480 2535
rect 6500 2515 6510 2535
rect 6470 2485 6510 2515
rect 6470 2465 6480 2485
rect 6500 2465 6510 2485
rect 6470 2435 6510 2465
rect 6470 2415 6480 2435
rect 6500 2415 6510 2435
rect 6470 2400 6510 2415
rect 6560 2685 6600 2700
rect 6560 2665 6570 2685
rect 6590 2665 6600 2685
rect 6560 2635 6600 2665
rect 6560 2615 6570 2635
rect 6590 2615 6600 2635
rect 6560 2585 6600 2615
rect 6560 2565 6570 2585
rect 6590 2565 6600 2585
rect 6560 2535 6600 2565
rect 6560 2515 6570 2535
rect 6590 2515 6600 2535
rect 6560 2485 6600 2515
rect 6560 2465 6570 2485
rect 6590 2465 6600 2485
rect 6560 2435 6600 2465
rect 6560 2415 6570 2435
rect 6590 2415 6600 2435
rect 6560 2400 6600 2415
rect 6650 2685 6690 2700
rect 6650 2665 6660 2685
rect 6680 2665 6690 2685
rect 6650 2635 6690 2665
rect 6650 2615 6660 2635
rect 6680 2615 6690 2635
rect 6650 2585 6690 2615
rect 6650 2565 6660 2585
rect 6680 2565 6690 2585
rect 6650 2535 6690 2565
rect 6650 2515 6660 2535
rect 6680 2515 6690 2535
rect 6650 2485 6690 2515
rect 6650 2465 6660 2485
rect 6680 2465 6690 2485
rect 6650 2435 6690 2465
rect 6650 2415 6660 2435
rect 6680 2415 6690 2435
rect 6650 2400 6690 2415
rect 6740 2685 6780 2700
rect 6740 2665 6750 2685
rect 6770 2665 6780 2685
rect 6740 2635 6780 2665
rect 6740 2615 6750 2635
rect 6770 2615 6780 2635
rect 6740 2585 6780 2615
rect 6740 2565 6750 2585
rect 6770 2565 6780 2585
rect 6740 2535 6780 2565
rect 6740 2515 6750 2535
rect 6770 2515 6780 2535
rect 6740 2485 6780 2515
rect 6740 2465 6750 2485
rect 6770 2465 6780 2485
rect 6740 2435 6780 2465
rect 6740 2415 6750 2435
rect 6770 2415 6780 2435
rect 6740 2400 6780 2415
rect 4155 1935 4195 1950
rect 4155 1915 4165 1935
rect 4185 1915 4195 1935
rect 4155 1885 4195 1915
rect 4155 1865 4165 1885
rect 4185 1865 4195 1885
rect 4155 1850 4195 1865
rect 4210 1935 4250 1950
rect 4210 1915 4220 1935
rect 4240 1915 4250 1935
rect 4210 1885 4250 1915
rect 4210 1865 4220 1885
rect 4240 1865 4250 1885
rect 4210 1850 4250 1865
rect 4265 1935 4305 1950
rect 4265 1915 4275 1935
rect 4295 1915 4305 1935
rect 4265 1885 4305 1915
rect 4265 1865 4275 1885
rect 4295 1865 4305 1885
rect 4265 1850 4305 1865
rect 4335 1935 4375 1950
rect 4335 1915 4345 1935
rect 4365 1915 4375 1935
rect 4335 1885 4375 1915
rect 4335 1865 4345 1885
rect 4365 1865 4375 1885
rect 4335 1850 4375 1865
rect 4395 1935 4435 1950
rect 4395 1915 4405 1935
rect 4425 1915 4435 1935
rect 4395 1885 4435 1915
rect 4395 1865 4405 1885
rect 4425 1865 4435 1885
rect 4395 1850 4435 1865
rect 4455 1935 4495 1950
rect 4455 1915 4465 1935
rect 4485 1915 4495 1935
rect 4455 1885 4495 1915
rect 4455 1865 4465 1885
rect 4485 1865 4495 1885
rect 4455 1850 4495 1865
rect 4515 1935 4555 1950
rect 4515 1915 4525 1935
rect 4545 1915 4555 1935
rect 4515 1885 4555 1915
rect 4515 1865 4525 1885
rect 4545 1865 4555 1885
rect 4515 1850 4555 1865
rect 4575 1935 4615 1950
rect 4575 1915 4585 1935
rect 4605 1915 4615 1935
rect 4575 1885 4615 1915
rect 4575 1865 4585 1885
rect 4605 1865 4615 1885
rect 4575 1850 4615 1865
rect 4635 1935 4675 1950
rect 4635 1915 4645 1935
rect 4665 1915 4675 1935
rect 4635 1885 4675 1915
rect 4635 1865 4645 1885
rect 4665 1865 4675 1885
rect 4635 1850 4675 1865
rect 4695 1935 4735 1950
rect 4695 1915 4705 1935
rect 4725 1915 4735 1935
rect 4695 1885 4735 1915
rect 4695 1865 4705 1885
rect 4725 1865 4735 1885
rect 4695 1850 4735 1865
rect 4755 1935 4795 1950
rect 4755 1915 4765 1935
rect 4785 1915 4795 1935
rect 4755 1885 4795 1915
rect 4755 1865 4765 1885
rect 4785 1865 4795 1885
rect 4755 1850 4795 1865
rect 4815 1935 4855 1950
rect 4815 1915 4825 1935
rect 4845 1915 4855 1935
rect 4815 1885 4855 1915
rect 4815 1865 4825 1885
rect 4845 1865 4855 1885
rect 4815 1850 4855 1865
rect 4875 1935 4915 1950
rect 4875 1915 4885 1935
rect 4905 1915 4915 1935
rect 4875 1885 4915 1915
rect 4875 1865 4885 1885
rect 4905 1865 4915 1885
rect 4875 1850 4915 1865
rect 4935 1935 4975 1950
rect 4935 1915 4945 1935
rect 4965 1915 4975 1935
rect 4935 1885 4975 1915
rect 4935 1865 4945 1885
rect 4965 1865 4975 1885
rect 4935 1850 4975 1865
rect 4995 1935 5035 1950
rect 4995 1915 5005 1935
rect 5025 1915 5035 1935
rect 4995 1885 5035 1915
rect 4995 1865 5005 1885
rect 5025 1865 5035 1885
rect 4995 1850 5035 1865
rect 5055 1935 5095 1950
rect 5055 1915 5065 1935
rect 5085 1915 5095 1935
rect 5055 1885 5095 1915
rect 5055 1865 5065 1885
rect 5085 1865 5095 1885
rect 5055 1850 5095 1865
rect 5115 1935 5155 1950
rect 5115 1915 5125 1935
rect 5145 1915 5155 1935
rect 5115 1885 5155 1915
rect 5115 1865 5125 1885
rect 5145 1865 5155 1885
rect 5115 1850 5155 1865
rect 5175 1935 5215 1950
rect 5175 1915 5185 1935
rect 5205 1915 5215 1935
rect 5175 1885 5215 1915
rect 5175 1865 5185 1885
rect 5205 1865 5215 1885
rect 5175 1850 5215 1865
rect 5235 1935 5275 1950
rect 5235 1915 5245 1935
rect 5265 1915 5275 1935
rect 5235 1885 5275 1915
rect 5235 1865 5245 1885
rect 5265 1865 5275 1885
rect 5235 1850 5275 1865
rect 5295 1935 5335 1950
rect 5295 1915 5305 1935
rect 5325 1915 5335 1935
rect 5295 1885 5335 1915
rect 5295 1865 5305 1885
rect 5325 1865 5335 1885
rect 5295 1850 5335 1865
rect 5355 1935 5395 1950
rect 5355 1915 5365 1935
rect 5385 1915 5395 1935
rect 5355 1885 5395 1915
rect 5355 1865 5365 1885
rect 5385 1865 5395 1885
rect 5355 1850 5395 1865
rect 5415 1935 5455 1950
rect 5415 1915 5425 1935
rect 5445 1915 5455 1935
rect 5415 1885 5455 1915
rect 5415 1865 5425 1885
rect 5445 1865 5455 1885
rect 5415 1850 5455 1865
rect 5475 1935 5515 1950
rect 5475 1915 5485 1935
rect 5505 1915 5515 1935
rect 5475 1885 5515 1915
rect 5475 1865 5485 1885
rect 5505 1865 5515 1885
rect 5475 1850 5515 1865
rect 5535 1935 5575 1950
rect 5535 1915 5545 1935
rect 5565 1915 5575 1935
rect 5535 1885 5575 1915
rect 5535 1865 5545 1885
rect 5565 1865 5575 1885
rect 5535 1850 5575 1865
rect 5605 1935 5645 1950
rect 5605 1915 5615 1935
rect 5635 1915 5645 1935
rect 5605 1885 5645 1915
rect 5605 1865 5615 1885
rect 5635 1865 5645 1885
rect 5605 1850 5645 1865
rect 5665 1935 5705 1950
rect 5665 1915 5675 1935
rect 5695 1915 5705 1935
rect 5665 1885 5705 1915
rect 5665 1865 5675 1885
rect 5695 1865 5705 1885
rect 5665 1850 5705 1865
rect 5725 1935 5765 1950
rect 5725 1915 5735 1935
rect 5755 1915 5765 1935
rect 5725 1885 5765 1915
rect 5725 1865 5735 1885
rect 5755 1865 5765 1885
rect 5725 1850 5765 1865
rect 5785 1935 5825 1950
rect 5785 1915 5795 1935
rect 5815 1915 5825 1935
rect 5785 1885 5825 1915
rect 5785 1865 5795 1885
rect 5815 1865 5825 1885
rect 5785 1850 5825 1865
rect 5845 1935 5885 1950
rect 5845 1915 5855 1935
rect 5875 1915 5885 1935
rect 5845 1885 5885 1915
rect 5845 1865 5855 1885
rect 5875 1865 5885 1885
rect 5845 1850 5885 1865
rect 5905 1935 5945 1950
rect 5905 1915 5915 1935
rect 5935 1915 5945 1935
rect 5905 1885 5945 1915
rect 5905 1865 5915 1885
rect 5935 1865 5945 1885
rect 5905 1850 5945 1865
rect 5965 1935 6005 1950
rect 5965 1915 5975 1935
rect 5995 1915 6005 1935
rect 5965 1885 6005 1915
rect 5965 1865 5975 1885
rect 5995 1865 6005 1885
rect 5965 1850 6005 1865
rect 6025 1935 6065 1950
rect 6025 1915 6035 1935
rect 6055 1915 6065 1935
rect 6025 1885 6065 1915
rect 6025 1865 6035 1885
rect 6055 1865 6065 1885
rect 6025 1850 6065 1865
rect 6085 1935 6125 1950
rect 6085 1915 6095 1935
rect 6115 1915 6125 1935
rect 6085 1885 6125 1915
rect 6085 1865 6095 1885
rect 6115 1865 6125 1885
rect 6085 1850 6125 1865
rect 6145 1935 6185 1950
rect 6145 1915 6155 1935
rect 6175 1915 6185 1935
rect 6145 1885 6185 1915
rect 6145 1865 6155 1885
rect 6175 1865 6185 1885
rect 6145 1850 6185 1865
rect 6205 1935 6245 1950
rect 6205 1915 6215 1935
rect 6235 1915 6245 1935
rect 6205 1885 6245 1915
rect 6205 1865 6215 1885
rect 6235 1865 6245 1885
rect 6205 1850 6245 1865
rect 6265 1935 6305 1950
rect 6265 1915 6275 1935
rect 6295 1915 6305 1935
rect 6265 1885 6305 1915
rect 6265 1865 6275 1885
rect 6295 1865 6305 1885
rect 6265 1850 6305 1865
rect 6325 1935 6365 1950
rect 6325 1915 6335 1935
rect 6355 1915 6365 1935
rect 6325 1885 6365 1915
rect 6325 1865 6335 1885
rect 6355 1865 6365 1885
rect 6325 1850 6365 1865
rect 6385 1935 6425 1950
rect 6385 1915 6395 1935
rect 6415 1915 6425 1935
rect 6385 1885 6425 1915
rect 6385 1865 6395 1885
rect 6415 1865 6425 1885
rect 6385 1850 6425 1865
rect 6445 1935 6485 1950
rect 6445 1915 6455 1935
rect 6475 1915 6485 1935
rect 6445 1885 6485 1915
rect 6445 1865 6455 1885
rect 6475 1865 6485 1885
rect 6445 1850 6485 1865
rect 6505 1935 6545 1950
rect 6505 1915 6515 1935
rect 6535 1915 6545 1935
rect 6505 1885 6545 1915
rect 6505 1865 6515 1885
rect 6535 1865 6545 1885
rect 6505 1850 6545 1865
rect 6565 1935 6605 1950
rect 6565 1915 6575 1935
rect 6595 1915 6605 1935
rect 6565 1885 6605 1915
rect 6565 1865 6575 1885
rect 6595 1865 6605 1885
rect 6565 1850 6605 1865
rect 6625 1935 6665 1950
rect 6625 1915 6635 1935
rect 6655 1915 6665 1935
rect 6625 1885 6665 1915
rect 6625 1865 6635 1885
rect 6655 1865 6665 1885
rect 6625 1850 6665 1865
rect 6685 1935 6725 1950
rect 6685 1915 6695 1935
rect 6715 1915 6725 1935
rect 6685 1885 6725 1915
rect 6685 1865 6695 1885
rect 6715 1865 6725 1885
rect 6685 1850 6725 1865
rect 6745 1935 6785 1950
rect 6745 1915 6755 1935
rect 6775 1915 6785 1935
rect 6745 1885 6785 1915
rect 6745 1865 6755 1885
rect 6775 1865 6785 1885
rect 6745 1850 6785 1865
rect 6805 1935 6845 1950
rect 6805 1915 6815 1935
rect 6835 1915 6845 1935
rect 6805 1885 6845 1915
rect 6805 1865 6815 1885
rect 6835 1865 6845 1885
rect 6805 1850 6845 1865
rect 4755 1600 4795 1615
rect 4755 1580 4765 1600
rect 4785 1580 4795 1600
rect 4755 1565 4795 1580
rect 4815 1600 4855 1615
rect 4815 1580 4825 1600
rect 4845 1580 4855 1600
rect 4815 1565 4855 1580
rect 4875 1600 4915 1615
rect 4875 1580 4885 1600
rect 4905 1580 4915 1600
rect 4875 1565 4915 1580
rect 4935 1600 4975 1615
rect 4935 1580 4945 1600
rect 4965 1580 4975 1600
rect 4935 1565 4975 1580
rect 4995 1600 5035 1615
rect 4995 1580 5005 1600
rect 5025 1580 5035 1600
rect 4995 1565 5035 1580
rect 5055 1600 5095 1615
rect 5055 1580 5065 1600
rect 5085 1580 5095 1600
rect 5055 1565 5095 1580
rect 5115 1600 5155 1615
rect 5115 1580 5125 1600
rect 5145 1580 5155 1600
rect 5115 1565 5155 1580
rect 5175 1600 5215 1615
rect 5175 1580 5185 1600
rect 5205 1580 5215 1600
rect 5175 1565 5215 1580
rect 5235 1600 5275 1615
rect 5235 1580 5245 1600
rect 5265 1580 5275 1600
rect 5235 1565 5275 1580
rect 5295 1600 5335 1615
rect 5295 1580 5305 1600
rect 5325 1580 5335 1600
rect 5295 1565 5335 1580
rect 5355 1600 5395 1615
rect 5355 1580 5365 1600
rect 5385 1580 5395 1600
rect 5355 1565 5395 1580
rect 5785 1600 5825 1615
rect 5785 1580 5795 1600
rect 5815 1580 5825 1600
rect 5785 1565 5825 1580
rect 5845 1600 5885 1615
rect 5845 1580 5855 1600
rect 5875 1580 5885 1600
rect 5845 1565 5885 1580
rect 5905 1600 5945 1615
rect 5905 1580 5915 1600
rect 5935 1580 5945 1600
rect 5905 1565 5945 1580
rect 5965 1600 6005 1615
rect 5965 1580 5975 1600
rect 5995 1580 6005 1600
rect 5965 1565 6005 1580
rect 6025 1600 6065 1615
rect 6025 1580 6035 1600
rect 6055 1580 6065 1600
rect 6025 1565 6065 1580
rect 6085 1600 6125 1615
rect 6085 1580 6095 1600
rect 6115 1580 6125 1600
rect 6085 1565 6125 1580
rect 6145 1600 6185 1615
rect 6145 1580 6155 1600
rect 6175 1580 6185 1600
rect 6145 1565 6185 1580
rect 6205 1600 6245 1615
rect 6205 1580 6215 1600
rect 6235 1580 6245 1600
rect 6205 1565 6245 1580
rect 6265 1600 6305 1615
rect 6265 1580 6275 1600
rect 6295 1580 6305 1600
rect 6265 1565 6305 1580
rect 6325 1600 6365 1615
rect 6325 1580 6335 1600
rect 6355 1580 6365 1600
rect 6325 1565 6365 1580
rect 6385 1600 6425 1615
rect 6385 1580 6395 1600
rect 6415 1580 6425 1600
rect 6385 1565 6425 1580
rect 4425 1395 4465 1410
rect 4425 1375 4435 1395
rect 4455 1375 4465 1395
rect 4425 1345 4465 1375
rect 4425 1325 4435 1345
rect 4455 1325 4465 1345
rect 4425 1295 4465 1325
rect 4425 1275 4435 1295
rect 4455 1275 4465 1295
rect 4425 1245 4465 1275
rect 4425 1225 4435 1245
rect 4455 1225 4465 1245
rect 4425 1195 4465 1225
rect 4425 1175 4435 1195
rect 4455 1175 4465 1195
rect 4425 1160 4465 1175
rect 4965 1395 5005 1410
rect 4965 1375 4975 1395
rect 4995 1375 5005 1395
rect 4965 1345 5005 1375
rect 4965 1325 4975 1345
rect 4995 1325 5005 1345
rect 4965 1295 5005 1325
rect 4965 1275 4975 1295
rect 4995 1275 5005 1295
rect 4965 1245 5005 1275
rect 4965 1225 4975 1245
rect 4995 1225 5005 1245
rect 4965 1195 5005 1225
rect 4965 1175 4975 1195
rect 4995 1175 5005 1195
rect 4965 1160 5005 1175
rect 5505 1395 5545 1410
rect 5505 1375 5515 1395
rect 5535 1375 5545 1395
rect 5505 1345 5545 1375
rect 5505 1325 5515 1345
rect 5535 1325 5545 1345
rect 5505 1295 5545 1325
rect 5505 1275 5515 1295
rect 5535 1275 5545 1295
rect 5505 1245 5545 1275
rect 5505 1225 5515 1245
rect 5535 1225 5545 1245
rect 5505 1195 5545 1225
rect 5505 1175 5515 1195
rect 5535 1175 5545 1195
rect 5505 1160 5545 1175
rect 5635 1395 5675 1410
rect 5635 1375 5645 1395
rect 5665 1375 5675 1395
rect 5635 1345 5675 1375
rect 5635 1325 5645 1345
rect 5665 1325 5675 1345
rect 5635 1295 5675 1325
rect 5635 1275 5645 1295
rect 5665 1275 5675 1295
rect 5635 1245 5675 1275
rect 5635 1225 5645 1245
rect 5665 1225 5675 1245
rect 5635 1195 5675 1225
rect 5635 1175 5645 1195
rect 5665 1175 5675 1195
rect 5635 1160 5675 1175
rect 6175 1395 6215 1410
rect 6175 1375 6185 1395
rect 6205 1375 6215 1395
rect 6175 1345 6215 1375
rect 6175 1325 6185 1345
rect 6205 1325 6215 1345
rect 6175 1295 6215 1325
rect 6175 1275 6185 1295
rect 6205 1275 6215 1295
rect 6175 1245 6215 1275
rect 6175 1225 6185 1245
rect 6205 1225 6215 1245
rect 6175 1195 6215 1225
rect 6175 1175 6185 1195
rect 6205 1175 6215 1195
rect 6175 1160 6215 1175
rect 6715 1395 6755 1410
rect 6715 1375 6725 1395
rect 6745 1375 6755 1395
rect 6715 1345 6755 1375
rect 6715 1325 6725 1345
rect 6745 1325 6755 1345
rect 6715 1295 6755 1325
rect 6715 1275 6725 1295
rect 6745 1275 6755 1295
rect 6715 1245 6755 1275
rect 6715 1225 6725 1245
rect 6745 1225 6755 1245
rect 6715 1195 6755 1225
rect 6715 1175 6725 1195
rect 6745 1175 6755 1195
rect 6715 1160 6755 1175
rect 4530 1050 4570 1065
rect 4530 1030 4540 1050
rect 4560 1030 4570 1050
rect 4530 1000 4570 1030
rect 4530 980 4540 1000
rect 4560 980 4570 1000
rect 4530 965 4570 980
rect 5570 1050 5610 1065
rect 5570 1030 5580 1050
rect 5600 1030 5610 1050
rect 5570 1000 5610 1030
rect 5570 980 5580 1000
rect 5600 980 5610 1000
rect 5570 965 5610 980
rect 6610 1050 6650 1065
rect 6610 1030 6620 1050
rect 6640 1030 6650 1050
rect 6610 1000 6650 1030
rect 6610 980 6620 1000
rect 6640 980 6650 1000
rect 6610 965 6650 980
rect 4680 895 4720 910
rect 4680 875 4690 895
rect 4710 875 4720 895
rect 4680 845 4720 875
rect 4680 825 4690 845
rect 4710 825 4720 845
rect 4680 810 4720 825
rect 4770 895 4810 910
rect 4770 875 4780 895
rect 4800 875 4810 895
rect 4770 845 4810 875
rect 4770 825 4780 845
rect 4800 825 4810 845
rect 4770 810 4810 825
rect 4840 895 4880 910
rect 4840 875 4850 895
rect 4870 875 4880 895
rect 4840 845 4880 875
rect 4840 825 4850 845
rect 4870 825 4880 845
rect 4840 810 4880 825
rect 4930 895 4970 910
rect 4930 875 4940 895
rect 4960 875 4970 895
rect 4930 845 4970 875
rect 4930 825 4940 845
rect 4960 825 4970 845
rect 4930 810 4970 825
rect 5020 895 5060 910
rect 5020 875 5030 895
rect 5050 875 5060 895
rect 5020 845 5060 875
rect 5020 825 5030 845
rect 5050 825 5060 845
rect 5020 810 5060 825
rect 5110 895 5150 910
rect 5110 875 5120 895
rect 5140 875 5150 895
rect 5110 845 5150 875
rect 5110 825 5120 845
rect 5140 825 5150 845
rect 5110 810 5150 825
rect 5200 895 5240 910
rect 5200 875 5210 895
rect 5230 875 5240 895
rect 5200 845 5240 875
rect 5200 825 5210 845
rect 5230 825 5240 845
rect 5200 810 5240 825
rect 5290 895 5330 910
rect 5290 875 5300 895
rect 5320 875 5330 895
rect 5290 845 5330 875
rect 5290 825 5300 845
rect 5320 825 5330 845
rect 5290 810 5330 825
rect 5380 895 5420 910
rect 5380 875 5390 895
rect 5410 875 5420 895
rect 5380 845 5420 875
rect 5380 825 5390 845
rect 5410 825 5420 845
rect 5380 810 5420 825
rect 5470 895 5510 910
rect 5470 875 5480 895
rect 5500 875 5510 895
rect 5470 845 5510 875
rect 5470 825 5480 845
rect 5500 825 5510 845
rect 5470 810 5510 825
rect 5560 895 5600 910
rect 5560 875 5570 895
rect 5590 875 5600 895
rect 5560 845 5600 875
rect 5560 825 5570 845
rect 5590 825 5600 845
rect 5560 810 5600 825
rect 5650 895 5690 910
rect 5650 875 5660 895
rect 5680 875 5690 895
rect 5650 845 5690 875
rect 5650 825 5660 845
rect 5680 825 5690 845
rect 5650 810 5690 825
rect 5740 895 5780 910
rect 5740 875 5750 895
rect 5770 875 5780 895
rect 5740 845 5780 875
rect 5740 825 5750 845
rect 5770 825 5780 845
rect 5740 810 5780 825
rect 5830 895 5870 910
rect 5830 875 5840 895
rect 5860 875 5870 895
rect 5830 845 5870 875
rect 5830 825 5840 845
rect 5860 825 5870 845
rect 5830 810 5870 825
rect 5920 895 5960 910
rect 5920 875 5930 895
rect 5950 875 5960 895
rect 5920 845 5960 875
rect 5920 825 5930 845
rect 5950 825 5960 845
rect 5920 810 5960 825
rect 6010 895 6050 910
rect 6010 875 6020 895
rect 6040 875 6050 895
rect 6010 845 6050 875
rect 6010 825 6020 845
rect 6040 825 6050 845
rect 6010 810 6050 825
rect 6100 895 6140 910
rect 6100 875 6110 895
rect 6130 875 6140 895
rect 6100 845 6140 875
rect 6100 825 6110 845
rect 6130 825 6140 845
rect 6100 810 6140 825
rect 6190 895 6230 910
rect 6190 875 6200 895
rect 6220 875 6230 895
rect 6190 845 6230 875
rect 6190 825 6200 845
rect 6220 825 6230 845
rect 6190 810 6230 825
rect 6280 895 6320 910
rect 6280 875 6290 895
rect 6310 875 6320 895
rect 6280 845 6320 875
rect 6280 825 6290 845
rect 6310 825 6320 845
rect 6280 810 6320 825
rect 6370 895 6410 910
rect 6370 875 6380 895
rect 6400 875 6410 895
rect 6370 845 6410 875
rect 6370 825 6380 845
rect 6400 825 6410 845
rect 6370 810 6410 825
rect 6460 895 6500 910
rect 6460 875 6470 895
rect 6490 875 6500 895
rect 6460 845 6500 875
rect 6460 825 6470 845
rect 6490 825 6500 845
rect 6460 810 6500 825
rect 6550 895 6590 910
rect 6550 875 6560 895
rect 6580 875 6590 895
rect 6550 845 6590 875
rect 6550 825 6560 845
rect 6580 825 6590 845
rect 6550 810 6590 825
<< ndiffc >>
rect 4555 2855 4575 2875
rect 4555 2805 4575 2825
rect 4645 2855 4665 2875
rect 4645 2805 4665 2825
rect 4735 2855 4755 2875
rect 4735 2805 4755 2825
rect 4805 2855 4825 2875
rect 4805 2805 4825 2825
rect 4895 2855 4915 2875
rect 4895 2805 4915 2825
rect 4985 2855 5005 2875
rect 4985 2805 5005 2825
rect 5075 2855 5095 2875
rect 5075 2805 5095 2825
rect 5165 2855 5185 2875
rect 5165 2805 5185 2825
rect 5255 2855 5275 2875
rect 5255 2805 5275 2825
rect 5345 2855 5365 2875
rect 5345 2805 5365 2825
rect 5435 2855 5455 2875
rect 5435 2805 5455 2825
rect 5525 2855 5545 2875
rect 5525 2805 5545 2825
rect 5615 2855 5635 2875
rect 5615 2805 5635 2825
rect 5705 2855 5725 2875
rect 5705 2805 5725 2825
rect 5795 2855 5815 2875
rect 5795 2805 5815 2825
rect 5885 2855 5905 2875
rect 5885 2805 5905 2825
rect 5975 2855 5995 2875
rect 5975 2805 5995 2825
rect 6065 2855 6085 2875
rect 6065 2805 6085 2825
rect 6155 2855 6175 2875
rect 6155 2805 6175 2825
rect 6245 2855 6265 2875
rect 6245 2805 6265 2825
rect 6335 2855 6355 2875
rect 6335 2805 6355 2825
rect 6425 2855 6445 2875
rect 6425 2805 6445 2825
rect 6515 2855 6535 2875
rect 6515 2805 6535 2825
rect 6605 2855 6625 2875
rect 6605 2805 6625 2825
rect 4410 2665 4430 2685
rect 4410 2615 4430 2635
rect 4410 2565 4430 2585
rect 4410 2515 4430 2535
rect 4410 2465 4430 2485
rect 4410 2415 4430 2435
rect 4500 2665 4520 2685
rect 4500 2615 4520 2635
rect 4500 2565 4520 2585
rect 4500 2515 4520 2535
rect 4500 2465 4520 2485
rect 4500 2415 4520 2435
rect 4590 2665 4610 2685
rect 4590 2615 4610 2635
rect 4590 2565 4610 2585
rect 4590 2515 4610 2535
rect 4590 2465 4610 2485
rect 4590 2415 4610 2435
rect 4680 2665 4700 2685
rect 4680 2615 4700 2635
rect 4680 2565 4700 2585
rect 4680 2515 4700 2535
rect 4680 2465 4700 2485
rect 4680 2415 4700 2435
rect 4770 2665 4790 2685
rect 4770 2615 4790 2635
rect 4770 2565 4790 2585
rect 4770 2515 4790 2535
rect 4770 2465 4790 2485
rect 4770 2415 4790 2435
rect 4860 2665 4880 2685
rect 4860 2615 4880 2635
rect 4860 2565 4880 2585
rect 4860 2515 4880 2535
rect 4860 2465 4880 2485
rect 4860 2415 4880 2435
rect 4950 2665 4970 2685
rect 4950 2615 4970 2635
rect 4950 2565 4970 2585
rect 4950 2515 4970 2535
rect 4950 2465 4970 2485
rect 4950 2415 4970 2435
rect 5040 2665 5060 2685
rect 5040 2615 5060 2635
rect 5040 2565 5060 2585
rect 5040 2515 5060 2535
rect 5040 2465 5060 2485
rect 5040 2415 5060 2435
rect 5130 2665 5150 2685
rect 5130 2615 5150 2635
rect 5130 2565 5150 2585
rect 5130 2515 5150 2535
rect 5130 2465 5150 2485
rect 5130 2415 5150 2435
rect 5220 2665 5240 2685
rect 5220 2615 5240 2635
rect 5220 2565 5240 2585
rect 5220 2515 5240 2535
rect 5220 2465 5240 2485
rect 5220 2415 5240 2435
rect 5310 2665 5330 2685
rect 5310 2615 5330 2635
rect 5310 2565 5330 2585
rect 5310 2515 5330 2535
rect 5310 2465 5330 2485
rect 5310 2415 5330 2435
rect 5400 2665 5420 2685
rect 5400 2615 5420 2635
rect 5400 2565 5420 2585
rect 5400 2515 5420 2535
rect 5400 2465 5420 2485
rect 5400 2415 5420 2435
rect 5490 2665 5510 2685
rect 5490 2615 5510 2635
rect 5490 2565 5510 2585
rect 5490 2515 5510 2535
rect 5490 2465 5510 2485
rect 5490 2415 5510 2435
rect 5580 2665 5600 2685
rect 5580 2615 5600 2635
rect 5580 2565 5600 2585
rect 5580 2515 5600 2535
rect 5580 2465 5600 2485
rect 5580 2415 5600 2435
rect 5670 2665 5690 2685
rect 5670 2615 5690 2635
rect 5670 2565 5690 2585
rect 5670 2515 5690 2535
rect 5670 2465 5690 2485
rect 5670 2415 5690 2435
rect 5760 2665 5780 2685
rect 5760 2615 5780 2635
rect 5760 2565 5780 2585
rect 5760 2515 5780 2535
rect 5760 2465 5780 2485
rect 5760 2415 5780 2435
rect 5850 2665 5870 2685
rect 5850 2615 5870 2635
rect 5850 2565 5870 2585
rect 5850 2515 5870 2535
rect 5850 2465 5870 2485
rect 5850 2415 5870 2435
rect 5940 2665 5960 2685
rect 5940 2615 5960 2635
rect 5940 2565 5960 2585
rect 5940 2515 5960 2535
rect 5940 2465 5960 2485
rect 5940 2415 5960 2435
rect 6030 2665 6050 2685
rect 6030 2615 6050 2635
rect 6030 2565 6050 2585
rect 6030 2515 6050 2535
rect 6030 2465 6050 2485
rect 6030 2415 6050 2435
rect 6120 2665 6140 2685
rect 6120 2615 6140 2635
rect 6120 2565 6140 2585
rect 6120 2515 6140 2535
rect 6120 2465 6140 2485
rect 6120 2415 6140 2435
rect 6210 2665 6230 2685
rect 6210 2615 6230 2635
rect 6210 2565 6230 2585
rect 6210 2515 6230 2535
rect 6210 2465 6230 2485
rect 6210 2415 6230 2435
rect 6300 2665 6320 2685
rect 6300 2615 6320 2635
rect 6300 2565 6320 2585
rect 6300 2515 6320 2535
rect 6300 2465 6320 2485
rect 6300 2415 6320 2435
rect 6390 2665 6410 2685
rect 6390 2615 6410 2635
rect 6390 2565 6410 2585
rect 6390 2515 6410 2535
rect 6390 2465 6410 2485
rect 6390 2415 6410 2435
rect 6480 2665 6500 2685
rect 6480 2615 6500 2635
rect 6480 2565 6500 2585
rect 6480 2515 6500 2535
rect 6480 2465 6500 2485
rect 6480 2415 6500 2435
rect 6570 2665 6590 2685
rect 6570 2615 6590 2635
rect 6570 2565 6590 2585
rect 6570 2515 6590 2535
rect 6570 2465 6590 2485
rect 6570 2415 6590 2435
rect 6660 2665 6680 2685
rect 6660 2615 6680 2635
rect 6660 2565 6680 2585
rect 6660 2515 6680 2535
rect 6660 2465 6680 2485
rect 6660 2415 6680 2435
rect 6750 2665 6770 2685
rect 6750 2615 6770 2635
rect 6750 2565 6770 2585
rect 6750 2515 6770 2535
rect 6750 2465 6770 2485
rect 6750 2415 6770 2435
rect 4165 1915 4185 1935
rect 4165 1865 4185 1885
rect 4220 1915 4240 1935
rect 4220 1865 4240 1885
rect 4275 1915 4295 1935
rect 4275 1865 4295 1885
rect 4345 1915 4365 1935
rect 4345 1865 4365 1885
rect 4405 1915 4425 1935
rect 4405 1865 4425 1885
rect 4465 1915 4485 1935
rect 4465 1865 4485 1885
rect 4525 1915 4545 1935
rect 4525 1865 4545 1885
rect 4585 1915 4605 1935
rect 4585 1865 4605 1885
rect 4645 1915 4665 1935
rect 4645 1865 4665 1885
rect 4705 1915 4725 1935
rect 4705 1865 4725 1885
rect 4765 1915 4785 1935
rect 4765 1865 4785 1885
rect 4825 1915 4845 1935
rect 4825 1865 4845 1885
rect 4885 1915 4905 1935
rect 4885 1865 4905 1885
rect 4945 1915 4965 1935
rect 4945 1865 4965 1885
rect 5005 1915 5025 1935
rect 5005 1865 5025 1885
rect 5065 1915 5085 1935
rect 5065 1865 5085 1885
rect 5125 1915 5145 1935
rect 5125 1865 5145 1885
rect 5185 1915 5205 1935
rect 5185 1865 5205 1885
rect 5245 1915 5265 1935
rect 5245 1865 5265 1885
rect 5305 1915 5325 1935
rect 5305 1865 5325 1885
rect 5365 1915 5385 1935
rect 5365 1865 5385 1885
rect 5425 1915 5445 1935
rect 5425 1865 5445 1885
rect 5485 1915 5505 1935
rect 5485 1865 5505 1885
rect 5545 1915 5565 1935
rect 5545 1865 5565 1885
rect 5615 1915 5635 1935
rect 5615 1865 5635 1885
rect 5675 1915 5695 1935
rect 5675 1865 5695 1885
rect 5735 1915 5755 1935
rect 5735 1865 5755 1885
rect 5795 1915 5815 1935
rect 5795 1865 5815 1885
rect 5855 1915 5875 1935
rect 5855 1865 5875 1885
rect 5915 1915 5935 1935
rect 5915 1865 5935 1885
rect 5975 1915 5995 1935
rect 5975 1865 5995 1885
rect 6035 1915 6055 1935
rect 6035 1865 6055 1885
rect 6095 1915 6115 1935
rect 6095 1865 6115 1885
rect 6155 1915 6175 1935
rect 6155 1865 6175 1885
rect 6215 1915 6235 1935
rect 6215 1865 6235 1885
rect 6275 1915 6295 1935
rect 6275 1865 6295 1885
rect 6335 1915 6355 1935
rect 6335 1865 6355 1885
rect 6395 1915 6415 1935
rect 6395 1865 6415 1885
rect 6455 1915 6475 1935
rect 6455 1865 6475 1885
rect 6515 1915 6535 1935
rect 6515 1865 6535 1885
rect 6575 1915 6595 1935
rect 6575 1865 6595 1885
rect 6635 1915 6655 1935
rect 6635 1865 6655 1885
rect 6695 1915 6715 1935
rect 6695 1865 6715 1885
rect 6755 1915 6775 1935
rect 6755 1865 6775 1885
rect 6815 1915 6835 1935
rect 6815 1865 6835 1885
rect 4765 1580 4785 1600
rect 4825 1580 4845 1600
rect 4885 1580 4905 1600
rect 4945 1580 4965 1600
rect 5005 1580 5025 1600
rect 5065 1580 5085 1600
rect 5125 1580 5145 1600
rect 5185 1580 5205 1600
rect 5245 1580 5265 1600
rect 5305 1580 5325 1600
rect 5365 1580 5385 1600
rect 5795 1580 5815 1600
rect 5855 1580 5875 1600
rect 5915 1580 5935 1600
rect 5975 1580 5995 1600
rect 6035 1580 6055 1600
rect 6095 1580 6115 1600
rect 6155 1580 6175 1600
rect 6215 1580 6235 1600
rect 6275 1580 6295 1600
rect 6335 1580 6355 1600
rect 6395 1580 6415 1600
rect 4435 1375 4455 1395
rect 4435 1325 4455 1345
rect 4435 1275 4455 1295
rect 4435 1225 4455 1245
rect 4435 1175 4455 1195
rect 4975 1375 4995 1395
rect 4975 1325 4995 1345
rect 4975 1275 4995 1295
rect 4975 1225 4995 1245
rect 4975 1175 4995 1195
rect 5515 1375 5535 1395
rect 5515 1325 5535 1345
rect 5515 1275 5535 1295
rect 5515 1225 5535 1245
rect 5515 1175 5535 1195
rect 5645 1375 5665 1395
rect 5645 1325 5665 1345
rect 5645 1275 5665 1295
rect 5645 1225 5665 1245
rect 5645 1175 5665 1195
rect 6185 1375 6205 1395
rect 6185 1325 6205 1345
rect 6185 1275 6205 1295
rect 6185 1225 6205 1245
rect 6185 1175 6205 1195
rect 6725 1375 6745 1395
rect 6725 1325 6745 1345
rect 6725 1275 6745 1295
rect 6725 1225 6745 1245
rect 6725 1175 6745 1195
rect 4540 1030 4560 1050
rect 4540 980 4560 1000
rect 5580 1030 5600 1050
rect 5580 980 5600 1000
rect 6620 1030 6640 1050
rect 6620 980 6640 1000
rect 4690 875 4710 895
rect 4690 825 4710 845
rect 4780 875 4800 895
rect 4780 825 4800 845
rect 4850 875 4870 895
rect 4850 825 4870 845
rect 4940 875 4960 895
rect 4940 825 4960 845
rect 5030 875 5050 895
rect 5030 825 5050 845
rect 5120 875 5140 895
rect 5120 825 5140 845
rect 5210 875 5230 895
rect 5210 825 5230 845
rect 5300 875 5320 895
rect 5300 825 5320 845
rect 5390 875 5410 895
rect 5390 825 5410 845
rect 5480 875 5500 895
rect 5480 825 5500 845
rect 5570 875 5590 895
rect 5570 825 5590 845
rect 5660 875 5680 895
rect 5660 825 5680 845
rect 5750 875 5770 895
rect 5750 825 5770 845
rect 5840 875 5860 895
rect 5840 825 5860 845
rect 5930 875 5950 895
rect 5930 825 5950 845
rect 6020 875 6040 895
rect 6020 825 6040 845
rect 6110 875 6130 895
rect 6110 825 6130 845
rect 6200 875 6220 895
rect 6200 825 6220 845
rect 6290 875 6310 895
rect 6290 825 6310 845
rect 6380 875 6400 895
rect 6380 825 6400 845
rect 6470 875 6490 895
rect 6470 825 6490 845
rect 6560 875 6580 895
rect 6560 825 6580 845
<< psubdiff >>
rect -50 1715 100 1730
rect -50 1695 -35 1715
rect -15 1695 15 1715
rect 35 1695 65 1715
rect 85 1695 100 1715
rect -50 1680 100 1695
<< psubdiffcont >>
rect -35 1695 -15 1715
rect 15 1695 35 1715
rect 65 1695 85 1715
<< poly >>
rect 4585 2890 4635 2905
rect 4675 2890 4725 2905
rect 4835 2890 4885 2905
rect 4925 2890 4975 2905
rect 5015 2890 5065 2905
rect 5105 2890 5155 2905
rect 5195 2890 5245 2905
rect 5285 2890 5335 2905
rect 5375 2890 5425 2905
rect 5465 2890 5515 2905
rect 5555 2890 5605 2905
rect 5645 2890 5695 2905
rect 5735 2890 5785 2905
rect 5825 2890 5875 2905
rect 5915 2890 5965 2905
rect 6005 2890 6055 2905
rect 6095 2890 6145 2905
rect 6185 2890 6235 2905
rect 6275 2890 6325 2905
rect 6365 2890 6415 2905
rect 6455 2890 6505 2905
rect 6545 2890 6595 2905
rect 4585 2775 4635 2790
rect 4675 2775 4725 2790
rect 4835 2775 4885 2790
rect 4925 2775 4975 2790
rect 5015 2775 5065 2790
rect 5105 2775 5155 2790
rect 5195 2775 5245 2790
rect 5285 2775 5335 2790
rect 5375 2775 5425 2790
rect 5465 2775 5515 2790
rect 5555 2775 5605 2790
rect 5645 2775 5695 2790
rect 5735 2775 5785 2790
rect 5825 2775 5875 2790
rect 5915 2775 5965 2790
rect 6005 2775 6055 2790
rect 6095 2775 6145 2790
rect 6185 2775 6235 2790
rect 6275 2775 6325 2790
rect 6365 2775 6415 2790
rect 6455 2775 6505 2790
rect 6545 2775 6595 2790
rect 4440 2700 4490 2715
rect 4530 2700 4580 2715
rect 4620 2700 4670 2715
rect 4710 2700 4760 2715
rect 4800 2700 4850 2715
rect 4890 2700 4940 2715
rect 4980 2700 5030 2715
rect 5070 2700 5120 2715
rect 5160 2700 5210 2715
rect 5250 2700 5300 2715
rect 5340 2700 5390 2715
rect 5430 2700 5480 2715
rect 5520 2700 5570 2715
rect 5610 2700 5660 2715
rect 5700 2700 5750 2715
rect 5790 2700 5840 2715
rect 5880 2700 5930 2715
rect 5970 2700 6020 2715
rect 6060 2700 6110 2715
rect 6150 2700 6200 2715
rect 6240 2700 6290 2715
rect 6330 2700 6380 2715
rect 6420 2700 6470 2715
rect 6510 2700 6560 2715
rect 6600 2700 6650 2715
rect 6690 2700 6740 2715
rect 4440 2390 4490 2400
rect 4400 2375 4490 2390
rect 4530 2390 4580 2400
rect 4620 2390 4670 2400
rect 4710 2390 4760 2400
rect 4800 2390 4850 2400
rect 4890 2390 4940 2400
rect 4980 2390 5030 2400
rect 5070 2390 5120 2400
rect 5160 2390 5210 2400
rect 5250 2390 5300 2400
rect 5340 2390 5390 2400
rect 5430 2390 5480 2400
rect 5520 2390 5570 2400
rect 5610 2390 5660 2400
rect 5700 2390 5750 2400
rect 5790 2390 5840 2400
rect 5880 2390 5930 2400
rect 5970 2390 6020 2400
rect 6060 2390 6110 2400
rect 6150 2390 6200 2400
rect 6240 2390 6290 2400
rect 6330 2390 6380 2400
rect 6420 2390 6470 2400
rect 6510 2390 6560 2400
rect 6600 2390 6650 2400
rect 4530 2375 6650 2390
rect 6690 2390 6740 2400
rect 6690 2375 6780 2390
rect 4400 2355 4410 2375
rect 4430 2355 4440 2375
rect 4400 2345 4440 2355
rect 4580 2370 4620 2375
rect 4580 2350 4590 2370
rect 4610 2350 4620 2370
rect 4580 2340 4620 2350
rect 5335 2355 5345 2375
rect 5365 2355 5375 2375
rect 5335 2345 5375 2355
rect 6740 2355 6750 2375
rect 6770 2355 6780 2375
rect 6740 2345 6780 2355
rect 4335 1995 4375 2005
rect 4335 1975 4345 1995
rect 4365 1980 4375 1995
rect 5535 1995 5575 2005
rect 5535 1980 5545 1995
rect 4365 1975 4395 1980
rect 4335 1965 4395 1975
rect 5515 1975 5545 1980
rect 5565 1975 5575 1995
rect 5515 1965 5575 1975
rect 5605 1995 5645 2005
rect 5605 1975 5615 1995
rect 5635 1980 5645 1995
rect 6805 1995 6845 2005
rect 6805 1980 6815 1995
rect 5635 1975 5665 1980
rect 5605 1965 5665 1975
rect 6785 1975 6815 1980
rect 6835 1975 6845 1995
rect 6785 1965 6845 1975
rect 4195 1950 4210 1965
rect 4250 1950 4265 1965
rect 4375 1950 4395 1965
rect 4435 1950 4455 1965
rect 4495 1950 4515 1965
rect 4555 1950 4575 1965
rect 4615 1950 4635 1965
rect 4675 1950 4695 1965
rect 4735 1950 4755 1965
rect 4795 1950 4815 1965
rect 4855 1950 4875 1965
rect 4915 1950 4935 1965
rect 4975 1950 4995 1965
rect 5035 1950 5055 1965
rect 5095 1950 5115 1965
rect 5155 1950 5175 1965
rect 5215 1950 5235 1965
rect 5275 1950 5295 1965
rect 5335 1950 5355 1965
rect 5395 1950 5415 1965
rect 5455 1950 5475 1965
rect 5515 1950 5535 1965
rect 5645 1950 5665 1965
rect 5705 1950 5725 1965
rect 5765 1950 5785 1965
rect 5825 1950 5845 1965
rect 5885 1950 5905 1965
rect 5945 1950 5965 1965
rect 6005 1950 6025 1965
rect 6065 1950 6085 1965
rect 6125 1950 6145 1965
rect 6185 1950 6205 1965
rect 6245 1950 6265 1965
rect 6305 1950 6325 1965
rect 6365 1950 6385 1965
rect 6425 1950 6445 1965
rect 6485 1950 6505 1965
rect 6545 1950 6565 1965
rect 6605 1950 6625 1965
rect 6665 1950 6685 1965
rect 6725 1950 6745 1965
rect 6785 1950 6805 1965
rect 4195 1840 4210 1850
rect 4250 1840 4265 1850
rect 4195 1825 4265 1840
rect 4375 1835 4395 1850
rect 4435 1835 4455 1850
rect 4495 1840 4515 1850
rect 4555 1840 4575 1850
rect 4615 1840 4635 1850
rect 4675 1840 4695 1850
rect 4425 1825 4465 1835
rect 4495 1825 4695 1840
rect 4735 1840 4755 1850
rect 4795 1840 4815 1850
rect 4735 1825 4815 1840
rect 4855 1840 4875 1850
rect 4915 1840 4935 1850
rect 4975 1840 4995 1850
rect 5035 1840 5055 1850
rect 4855 1825 5055 1840
rect 5095 1840 5115 1850
rect 5155 1840 5175 1850
rect 5095 1825 5175 1840
rect 5215 1840 5235 1850
rect 5275 1840 5295 1850
rect 5335 1840 5355 1850
rect 5395 1840 5415 1850
rect 5215 1825 5415 1840
rect 5455 1835 5475 1850
rect 5515 1835 5535 1850
rect 5645 1835 5665 1850
rect 5705 1835 5725 1850
rect 5765 1840 5785 1850
rect 5825 1840 5845 1850
rect 5885 1840 5905 1850
rect 5945 1840 5965 1850
rect 5445 1825 5485 1835
rect 4210 1805 4220 1825
rect 4240 1805 4250 1825
rect 4210 1795 4250 1805
rect 4425 1805 4435 1825
rect 4455 1805 4465 1825
rect 4425 1795 4465 1805
rect 4515 1805 4525 1825
rect 4545 1805 4555 1825
rect 4515 1795 4555 1805
rect 4755 1805 4765 1825
rect 4785 1805 4795 1825
rect 4755 1795 4795 1805
rect 4875 1805 4885 1825
rect 4905 1805 4915 1825
rect 4875 1795 4915 1805
rect 5115 1805 5125 1825
rect 5145 1805 5155 1825
rect 5115 1795 5155 1805
rect 5235 1805 5245 1825
rect 5265 1805 5275 1825
rect 5235 1795 5275 1805
rect 5445 1805 5455 1825
rect 5475 1805 5485 1825
rect 5445 1795 5485 1805
rect 5695 1825 5735 1835
rect 5765 1825 5965 1840
rect 6005 1840 6025 1850
rect 6065 1840 6085 1850
rect 6005 1825 6085 1840
rect 6125 1840 6145 1850
rect 6185 1840 6205 1850
rect 6245 1840 6265 1850
rect 6305 1840 6325 1850
rect 6125 1825 6325 1840
rect 6365 1840 6385 1850
rect 6425 1840 6445 1850
rect 6365 1825 6445 1840
rect 6485 1840 6505 1850
rect 6545 1840 6565 1850
rect 6605 1840 6625 1850
rect 6665 1840 6685 1850
rect 6485 1825 6685 1840
rect 6725 1835 6745 1850
rect 6785 1835 6805 1850
rect 6715 1825 6755 1835
rect 5695 1805 5705 1825
rect 5725 1805 5735 1825
rect 5695 1795 5735 1805
rect 5905 1805 5915 1825
rect 5935 1805 5945 1825
rect 5905 1795 5945 1805
rect 6025 1805 6035 1825
rect 6055 1805 6065 1825
rect 6025 1795 6065 1805
rect 6265 1805 6275 1825
rect 6295 1805 6305 1825
rect 6265 1795 6305 1805
rect 6385 1805 6395 1825
rect 6415 1805 6425 1825
rect 6385 1795 6425 1805
rect 6625 1805 6635 1825
rect 6655 1805 6665 1825
rect 6625 1795 6665 1805
rect 6715 1805 6725 1825
rect 6745 1805 6755 1825
rect 6715 1795 6755 1805
rect 4815 1705 4855 1715
rect 4815 1685 4825 1705
rect 4845 1685 4855 1705
rect 4815 1670 4855 1685
rect 6325 1705 6365 1715
rect 6325 1685 6335 1705
rect 6355 1685 6365 1705
rect 6325 1670 6365 1685
rect 4815 1655 5355 1670
rect 4795 1615 4815 1630
rect 4855 1615 4875 1655
rect 4915 1615 4935 1655
rect 4975 1615 4995 1630
rect 5035 1615 5055 1630
rect 5095 1615 5115 1655
rect 5155 1615 5175 1655
rect 5215 1615 5235 1630
rect 5275 1615 5295 1630
rect 5335 1615 5355 1655
rect 5825 1655 6365 1670
rect 5825 1615 5845 1655
rect 5885 1615 5905 1630
rect 5945 1615 5965 1630
rect 6005 1615 6025 1655
rect 6065 1615 6085 1655
rect 6125 1615 6145 1630
rect 6185 1615 6205 1630
rect 6245 1615 6265 1655
rect 6305 1615 6325 1655
rect 6365 1615 6385 1630
rect 4795 1550 4815 1565
rect 4855 1550 4875 1565
rect 4915 1550 4935 1565
rect 4755 1540 4815 1550
rect 4755 1520 4765 1540
rect 4785 1525 4815 1540
rect 4975 1525 4995 1565
rect 5035 1525 5055 1565
rect 5095 1550 5115 1565
rect 5155 1550 5175 1565
rect 5215 1525 5235 1565
rect 5275 1525 5295 1565
rect 5335 1550 5355 1565
rect 5825 1550 5845 1565
rect 4785 1520 5295 1525
rect 4755 1510 5295 1520
rect 5885 1525 5905 1565
rect 5945 1525 5965 1565
rect 6005 1550 6025 1565
rect 6065 1550 6085 1565
rect 6125 1525 6145 1565
rect 6185 1525 6205 1565
rect 6245 1550 6265 1565
rect 6305 1550 6325 1565
rect 6365 1550 6385 1565
rect 6365 1540 6425 1550
rect 6365 1525 6395 1540
rect 5885 1520 6395 1525
rect 6415 1520 6425 1540
rect 5885 1510 6425 1520
rect 4465 1410 4965 1425
rect 5005 1410 5505 1425
rect 5675 1410 6175 1425
rect 6215 1410 6715 1425
rect 4465 1145 4965 1160
rect 5005 1145 5505 1160
rect 5675 1145 6175 1160
rect 6215 1145 6715 1160
rect 4610 1080 4650 1120
rect 4690 1080 4730 1120
rect 4770 1080 4810 1120
rect 4850 1080 4890 1120
rect 4930 1080 4970 1120
rect 5010 1080 5050 1120
rect 5090 1080 5130 1120
rect 5170 1080 5210 1120
rect 5250 1080 5290 1120
rect 5330 1080 5370 1120
rect 5410 1080 5450 1120
rect 5490 1080 5530 1120
rect 5650 1080 5690 1120
rect 5730 1080 5770 1120
rect 5810 1080 5850 1120
rect 5890 1080 5930 1120
rect 5970 1080 6010 1120
rect 6050 1080 6090 1120
rect 6130 1080 6170 1120
rect 6210 1080 6250 1120
rect 6290 1080 6330 1120
rect 6370 1080 6410 1120
rect 6450 1080 6490 1120
rect 6530 1080 6570 1120
rect 4570 1065 5570 1080
rect 5610 1065 6610 1080
rect 4570 950 5570 965
rect 5610 950 6610 965
rect 4720 910 4770 925
rect 4880 910 4930 925
rect 4970 910 5020 925
rect 5060 910 5110 925
rect 5150 910 5200 925
rect 5240 910 5290 925
rect 5330 910 5380 925
rect 5420 910 5470 925
rect 5510 910 5560 925
rect 5600 910 5650 925
rect 5690 910 5740 925
rect 5780 910 5830 925
rect 5870 910 5920 925
rect 5960 910 6010 925
rect 6050 910 6100 925
rect 6140 910 6190 925
rect 6230 910 6280 925
rect 6320 910 6370 925
rect 6410 910 6460 925
rect 6500 910 6550 925
rect 4720 795 4770 810
rect 4880 795 4930 810
rect 4970 795 5020 810
rect 5060 795 5110 810
rect 5150 795 5200 810
rect 5240 795 5290 810
rect 5330 795 5380 810
rect 5420 795 5470 810
rect 5510 795 5560 810
rect 5600 795 5650 810
rect 5690 795 5740 810
rect 5780 795 5830 810
rect 5870 795 5920 810
rect 5960 795 6010 810
rect 6050 795 6100 810
rect 6140 795 6190 810
rect 6230 795 6280 810
rect 6320 795 6370 810
rect 6410 795 6460 810
rect 6500 795 6550 810
<< polycont >>
rect 4410 2355 4430 2375
rect 4590 2350 4610 2370
rect 5345 2355 5365 2375
rect 6750 2355 6770 2375
rect 4345 1975 4365 1995
rect 5545 1975 5565 1995
rect 5615 1975 5635 1995
rect 6815 1975 6835 1995
rect 4220 1805 4240 1825
rect 4435 1805 4455 1825
rect 4525 1805 4545 1825
rect 4765 1805 4785 1825
rect 4885 1805 4905 1825
rect 5125 1805 5145 1825
rect 5245 1805 5265 1825
rect 5455 1805 5475 1825
rect 5705 1805 5725 1825
rect 5915 1805 5935 1825
rect 6035 1805 6055 1825
rect 6275 1805 6295 1825
rect 6395 1805 6415 1825
rect 6635 1805 6655 1825
rect 6725 1805 6745 1825
rect 4825 1685 4845 1705
rect 6335 1685 6355 1705
rect 4765 1520 4785 1540
rect 6395 1520 6415 1540
<< xpolycontact >>
rect 2385 1570 2605 1605
rect 3205 1570 3425 1605
rect 2385 1510 2605 1545
rect 3205 1510 3425 1545
rect 2385 1450 2605 1485
rect 3205 1450 3425 1485
rect 2385 1390 2605 1425
rect 3205 1390 3425 1425
rect 2385 1330 2605 1365
rect 3205 1330 3425 1365
rect 2385 1270 2605 1305
rect 3205 1270 3425 1305
rect 2390 995 2610 1030
rect 2840 995 3060 1030
rect 2505 935 2725 970
rect 3330 935 3550 970
rect 2505 875 2725 910
rect 3330 875 3550 910
rect 2505 795 2725 830
rect 3325 795 3545 830
rect 2505 735 2725 770
rect 3325 735 3545 770
rect -795 -435 -575 -400
rect -31 -435 189 -400
rect -795 -495 -575 -460
rect -31 -495 189 -460
rect -795 -555 -575 -520
rect -31 -555 189 -520
rect -795 -615 -575 -580
rect -31 -615 189 -580
rect -795 -675 -575 -640
rect -31 -675 189 -640
rect -795 -735 -575 -700
rect -31 -735 189 -700
rect -795 -795 -575 -760
rect -31 -795 189 -760
rect -795 -855 -575 -820
rect -31 -855 189 -820
rect -795 -915 -575 -880
rect -31 -915 189 -880
rect -795 -975 -575 -940
rect -241 -975 -21 -940
rect -795 -1035 -575 -1000
rect -31 -1035 189 -1000
rect -795 -1095 -575 -1060
rect -31 -1095 189 -1060
rect -795 -1155 -575 -1120
rect -31 -1155 189 -1120
rect -795 -1215 -575 -1180
rect -31 -1215 189 -1180
rect -795 -1275 -575 -1240
rect -31 -1275 189 -1240
rect -795 -1335 -575 -1300
rect -31 -1335 189 -1300
rect -795 -1395 -575 -1360
rect -31 -1395 189 -1360
rect -795 -1455 -575 -1420
rect -31 -1455 189 -1420
rect -795 -1515 -575 -1480
rect -31 -1515 189 -1480
<< xpolyres >>
rect 2605 1570 3205 1605
rect 2605 1510 3205 1545
rect 2605 1450 3205 1485
rect 2605 1390 3205 1425
rect 2605 1330 3205 1365
rect 2605 1270 3205 1305
rect 2610 995 2840 1030
rect 2725 935 3330 970
rect 2725 875 3330 910
rect 2725 795 3325 830
rect 2725 735 3325 770
rect -575 -435 -31 -400
rect -575 -495 -31 -460
rect -575 -555 -31 -520
rect -575 -615 -31 -580
rect -575 -675 -31 -640
rect -575 -735 -31 -700
rect -575 -795 -31 -760
rect -575 -855 -31 -820
rect -575 -915 -31 -880
rect -575 -975 -241 -940
rect -575 -1035 -31 -1000
rect -575 -1095 -31 -1060
rect -575 -1155 -31 -1120
rect -575 -1215 -31 -1180
rect -575 -1275 -31 -1240
rect -575 -1335 -31 -1300
rect -575 -1395 -31 -1360
rect -575 -1455 -31 -1420
rect -575 -1515 -31 -1480
<< locali >>
rect 4550 3045 4580 3075
rect 7040 3045 7070 3075
rect 4545 2935 4585 2945
rect 4545 2915 4555 2935
rect 4575 2915 4585 2935
rect 4545 2905 4585 2915
rect 4555 2885 4575 2905
rect 4550 2875 4580 2885
rect 4550 2855 4555 2875
rect 4575 2855 4580 2875
rect 4550 2825 4580 2855
rect 4550 2805 4555 2825
rect 4575 2805 4580 2825
rect 4550 2795 4580 2805
rect 4640 2875 4670 2885
rect 4640 2855 4645 2875
rect 4665 2855 4670 2875
rect 4640 2825 4670 2855
rect 4640 2805 4645 2825
rect 4665 2805 4670 2825
rect 4640 2795 4670 2805
rect 4730 2875 4760 2885
rect 4730 2855 4735 2875
rect 4755 2855 4760 2875
rect 4730 2825 4760 2855
rect 4730 2805 4735 2825
rect 4755 2805 4760 2825
rect 4730 2795 4760 2805
rect 4800 2875 4830 2885
rect 4800 2855 4805 2875
rect 4825 2855 4830 2875
rect 4800 2825 4830 2855
rect 4800 2805 4805 2825
rect 4825 2805 4830 2825
rect 4800 2795 4830 2805
rect 4890 2875 4920 2885
rect 4890 2855 4895 2875
rect 4915 2855 4920 2875
rect 4890 2825 4920 2855
rect 4890 2805 4895 2825
rect 4915 2805 4920 2825
rect 4890 2795 4920 2805
rect 4980 2875 5010 2885
rect 4980 2855 4985 2875
rect 5005 2855 5010 2875
rect 4980 2825 5010 2855
rect 4980 2805 4985 2825
rect 5005 2805 5010 2825
rect 4980 2795 5010 2805
rect 5070 2875 5100 2885
rect 5070 2855 5075 2875
rect 5095 2855 5100 2875
rect 5070 2825 5100 2855
rect 5070 2805 5075 2825
rect 5095 2805 5100 2825
rect 5070 2795 5100 2805
rect 5160 2875 5190 2885
rect 5160 2855 5165 2875
rect 5185 2855 5190 2875
rect 5160 2825 5190 2855
rect 5160 2805 5165 2825
rect 5185 2805 5190 2825
rect 5160 2795 5190 2805
rect 5250 2875 5280 2885
rect 5250 2855 5255 2875
rect 5275 2855 5280 2875
rect 5250 2825 5280 2855
rect 5250 2805 5255 2825
rect 5275 2805 5280 2825
rect 5250 2795 5280 2805
rect 5340 2875 5370 2885
rect 5340 2855 5345 2875
rect 5365 2855 5370 2875
rect 5340 2825 5370 2855
rect 5340 2805 5345 2825
rect 5365 2805 5370 2825
rect 5340 2795 5370 2805
rect 5430 2875 5460 2885
rect 5430 2855 5435 2875
rect 5455 2855 5460 2875
rect 5430 2825 5460 2855
rect 5430 2805 5435 2825
rect 5455 2805 5460 2825
rect 5430 2795 5460 2805
rect 5520 2875 5550 2885
rect 5520 2855 5525 2875
rect 5545 2855 5550 2875
rect 5520 2825 5550 2855
rect 5520 2805 5525 2825
rect 5545 2805 5550 2825
rect 5520 2795 5550 2805
rect 5610 2875 5640 2885
rect 5610 2855 5615 2875
rect 5635 2855 5640 2875
rect 5610 2825 5640 2855
rect 5610 2805 5615 2825
rect 5635 2805 5640 2825
rect 5610 2795 5640 2805
rect 5700 2875 5730 2885
rect 5700 2855 5705 2875
rect 5725 2855 5730 2875
rect 5700 2825 5730 2855
rect 5700 2805 5705 2825
rect 5725 2805 5730 2825
rect 5700 2795 5730 2805
rect 5790 2875 5820 2885
rect 5790 2855 5795 2875
rect 5815 2855 5820 2875
rect 5790 2825 5820 2855
rect 5790 2805 5795 2825
rect 5815 2805 5820 2825
rect 5790 2795 5820 2805
rect 5880 2875 5910 2885
rect 5880 2855 5885 2875
rect 5905 2855 5910 2875
rect 5880 2825 5910 2855
rect 5880 2805 5885 2825
rect 5905 2805 5910 2825
rect 5880 2795 5910 2805
rect 5970 2875 6000 2885
rect 5970 2855 5975 2875
rect 5995 2855 6000 2875
rect 5970 2825 6000 2855
rect 5970 2805 5975 2825
rect 5995 2805 6000 2825
rect 5970 2795 6000 2805
rect 6060 2875 6090 2885
rect 6060 2855 6065 2875
rect 6085 2855 6090 2875
rect 6060 2825 6090 2855
rect 6060 2805 6065 2825
rect 6085 2805 6090 2825
rect 6060 2795 6090 2805
rect 6150 2875 6180 2885
rect 6150 2855 6155 2875
rect 6175 2855 6180 2875
rect 6150 2825 6180 2855
rect 6150 2805 6155 2825
rect 6175 2805 6180 2825
rect 6150 2795 6180 2805
rect 6240 2875 6270 2885
rect 6240 2855 6245 2875
rect 6265 2855 6270 2875
rect 6240 2825 6270 2855
rect 6240 2805 6245 2825
rect 6265 2805 6270 2825
rect 6240 2795 6270 2805
rect 6330 2875 6360 2885
rect 6330 2855 6335 2875
rect 6355 2855 6360 2875
rect 6330 2825 6360 2855
rect 6330 2805 6335 2825
rect 6355 2805 6360 2825
rect 6330 2795 6360 2805
rect 6420 2875 6450 2885
rect 6420 2855 6425 2875
rect 6445 2855 6450 2875
rect 6420 2825 6450 2855
rect 6420 2805 6425 2825
rect 6445 2805 6450 2825
rect 6420 2795 6450 2805
rect 6510 2875 6540 2885
rect 6510 2855 6515 2875
rect 6535 2855 6540 2875
rect 6510 2825 6540 2855
rect 6510 2805 6515 2825
rect 6535 2805 6540 2825
rect 6510 2795 6540 2805
rect 6600 2875 6630 2885
rect 6600 2855 6605 2875
rect 6625 2855 6630 2875
rect 6600 2825 6630 2855
rect 6600 2805 6605 2825
rect 6625 2805 6630 2825
rect 6600 2795 6630 2805
rect 4580 2745 4620 2755
rect 4580 2725 4590 2745
rect 4610 2725 4620 2745
rect 4580 2715 4620 2725
rect 4760 2745 4800 2755
rect 4760 2725 4770 2745
rect 4790 2725 4800 2745
rect 4760 2715 4800 2725
rect 4940 2745 4980 2755
rect 4940 2725 4950 2745
rect 4970 2725 4980 2745
rect 4940 2715 4980 2725
rect 5120 2745 5160 2755
rect 5120 2725 5130 2745
rect 5150 2725 5160 2745
rect 5120 2715 5160 2725
rect 5300 2745 5340 2755
rect 5300 2725 5310 2745
rect 5330 2725 5340 2745
rect 5300 2715 5340 2725
rect 5480 2745 5520 2755
rect 5480 2725 5490 2745
rect 5510 2725 5520 2745
rect 5480 2715 5520 2725
rect 5660 2745 5700 2755
rect 5660 2725 5670 2745
rect 5690 2725 5700 2745
rect 5660 2715 5700 2725
rect 5840 2745 5880 2755
rect 5840 2725 5850 2745
rect 5870 2725 5880 2745
rect 5840 2715 5880 2725
rect 6020 2745 6060 2755
rect 6020 2725 6030 2745
rect 6050 2725 6060 2745
rect 6020 2715 6060 2725
rect 6200 2745 6240 2755
rect 6200 2725 6210 2745
rect 6230 2725 6240 2745
rect 6200 2715 6240 2725
rect 6380 2745 6420 2755
rect 6380 2725 6390 2745
rect 6410 2725 6420 2745
rect 6380 2715 6420 2725
rect 6560 2745 6600 2755
rect 6560 2725 6570 2745
rect 6590 2725 6600 2745
rect 6560 2715 6600 2725
rect 650 2055 775 2700
rect 1330 2055 1455 2700
rect 2010 2055 2135 2700
rect 4590 2695 4610 2715
rect 4770 2695 4790 2715
rect 4950 2695 4970 2715
rect 5130 2695 5150 2715
rect 5310 2695 5330 2715
rect 5490 2695 5510 2715
rect 5670 2695 5690 2715
rect 5850 2695 5870 2715
rect 6030 2695 6050 2715
rect 6210 2695 6230 2715
rect 6390 2695 6410 2715
rect 6570 2695 6590 2715
rect 4405 2685 4435 2695
rect 4405 2665 4410 2685
rect 4430 2665 4435 2685
rect 4405 2635 4435 2665
rect 4405 2615 4410 2635
rect 4430 2615 4435 2635
rect 4405 2585 4435 2615
rect 4405 2565 4410 2585
rect 4430 2565 4435 2585
rect 4405 2535 4435 2565
rect 4405 2515 4410 2535
rect 4430 2515 4435 2535
rect 4405 2485 4435 2515
rect 4405 2465 4410 2485
rect 4430 2465 4435 2485
rect 4405 2435 4435 2465
rect 4405 2415 4410 2435
rect 4430 2415 4435 2435
rect 4405 2405 4435 2415
rect 4495 2685 4525 2695
rect 4495 2665 4500 2685
rect 4520 2665 4525 2685
rect 4495 2635 4525 2665
rect 4495 2615 4500 2635
rect 4520 2615 4525 2635
rect 4495 2585 4525 2615
rect 4495 2565 4500 2585
rect 4520 2565 4525 2585
rect 4495 2535 4525 2565
rect 4495 2515 4500 2535
rect 4520 2515 4525 2535
rect 4495 2485 4525 2515
rect 4495 2465 4500 2485
rect 4520 2465 4525 2485
rect 4495 2435 4525 2465
rect 4495 2415 4500 2435
rect 4520 2415 4525 2435
rect 4495 2405 4525 2415
rect 4585 2685 4615 2695
rect 4585 2665 4590 2685
rect 4610 2665 4615 2685
rect 4585 2635 4615 2665
rect 4585 2615 4590 2635
rect 4610 2615 4615 2635
rect 4585 2585 4615 2615
rect 4585 2565 4590 2585
rect 4610 2565 4615 2585
rect 4585 2535 4615 2565
rect 4585 2515 4590 2535
rect 4610 2515 4615 2535
rect 4585 2485 4615 2515
rect 4585 2465 4590 2485
rect 4610 2465 4615 2485
rect 4585 2435 4615 2465
rect 4585 2415 4590 2435
rect 4610 2415 4615 2435
rect 4585 2405 4615 2415
rect 4675 2685 4705 2695
rect 4675 2665 4680 2685
rect 4700 2665 4705 2685
rect 4675 2635 4705 2665
rect 4675 2615 4680 2635
rect 4700 2615 4705 2635
rect 4675 2585 4705 2615
rect 4675 2565 4680 2585
rect 4700 2565 4705 2585
rect 4675 2535 4705 2565
rect 4675 2515 4680 2535
rect 4700 2515 4705 2535
rect 4675 2485 4705 2515
rect 4675 2465 4680 2485
rect 4700 2465 4705 2485
rect 4675 2435 4705 2465
rect 4675 2415 4680 2435
rect 4700 2415 4705 2435
rect 4675 2405 4705 2415
rect 4765 2685 4795 2695
rect 4765 2665 4770 2685
rect 4790 2665 4795 2685
rect 4765 2635 4795 2665
rect 4765 2615 4770 2635
rect 4790 2615 4795 2635
rect 4765 2585 4795 2615
rect 4765 2565 4770 2585
rect 4790 2565 4795 2585
rect 4765 2535 4795 2565
rect 4765 2515 4770 2535
rect 4790 2515 4795 2535
rect 4765 2485 4795 2515
rect 4765 2465 4770 2485
rect 4790 2465 4795 2485
rect 4765 2435 4795 2465
rect 4765 2415 4770 2435
rect 4790 2415 4795 2435
rect 4765 2405 4795 2415
rect 4855 2685 4885 2695
rect 4855 2665 4860 2685
rect 4880 2665 4885 2685
rect 4855 2635 4885 2665
rect 4855 2615 4860 2635
rect 4880 2615 4885 2635
rect 4855 2585 4885 2615
rect 4855 2565 4860 2585
rect 4880 2565 4885 2585
rect 4855 2535 4885 2565
rect 4855 2515 4860 2535
rect 4880 2515 4885 2535
rect 4855 2485 4885 2515
rect 4855 2465 4860 2485
rect 4880 2465 4885 2485
rect 4855 2435 4885 2465
rect 4855 2415 4860 2435
rect 4880 2415 4885 2435
rect 4855 2405 4885 2415
rect 4945 2685 4975 2695
rect 4945 2665 4950 2685
rect 4970 2665 4975 2685
rect 4945 2635 4975 2665
rect 4945 2615 4950 2635
rect 4970 2615 4975 2635
rect 4945 2585 4975 2615
rect 4945 2565 4950 2585
rect 4970 2565 4975 2585
rect 4945 2535 4975 2565
rect 4945 2515 4950 2535
rect 4970 2515 4975 2535
rect 4945 2485 4975 2515
rect 4945 2465 4950 2485
rect 4970 2465 4975 2485
rect 4945 2435 4975 2465
rect 4945 2415 4950 2435
rect 4970 2415 4975 2435
rect 4945 2405 4975 2415
rect 5035 2685 5065 2695
rect 5035 2665 5040 2685
rect 5060 2665 5065 2685
rect 5035 2635 5065 2665
rect 5035 2615 5040 2635
rect 5060 2615 5065 2635
rect 5035 2585 5065 2615
rect 5035 2565 5040 2585
rect 5060 2565 5065 2585
rect 5035 2535 5065 2565
rect 5035 2515 5040 2535
rect 5060 2515 5065 2535
rect 5035 2485 5065 2515
rect 5035 2465 5040 2485
rect 5060 2465 5065 2485
rect 5035 2435 5065 2465
rect 5035 2415 5040 2435
rect 5060 2415 5065 2435
rect 5035 2405 5065 2415
rect 5125 2685 5155 2695
rect 5125 2665 5130 2685
rect 5150 2665 5155 2685
rect 5125 2635 5155 2665
rect 5125 2615 5130 2635
rect 5150 2615 5155 2635
rect 5125 2585 5155 2615
rect 5125 2565 5130 2585
rect 5150 2565 5155 2585
rect 5125 2535 5155 2565
rect 5125 2515 5130 2535
rect 5150 2515 5155 2535
rect 5125 2485 5155 2515
rect 5125 2465 5130 2485
rect 5150 2465 5155 2485
rect 5125 2435 5155 2465
rect 5125 2415 5130 2435
rect 5150 2415 5155 2435
rect 5125 2405 5155 2415
rect 5215 2685 5245 2695
rect 5215 2665 5220 2685
rect 5240 2665 5245 2685
rect 5215 2635 5245 2665
rect 5215 2615 5220 2635
rect 5240 2615 5245 2635
rect 5215 2585 5245 2615
rect 5215 2565 5220 2585
rect 5240 2565 5245 2585
rect 5215 2535 5245 2565
rect 5215 2515 5220 2535
rect 5240 2515 5245 2535
rect 5215 2485 5245 2515
rect 5215 2465 5220 2485
rect 5240 2465 5245 2485
rect 5215 2435 5245 2465
rect 5215 2415 5220 2435
rect 5240 2415 5245 2435
rect 5215 2405 5245 2415
rect 5305 2685 5335 2695
rect 5305 2665 5310 2685
rect 5330 2665 5335 2685
rect 5305 2635 5335 2665
rect 5305 2615 5310 2635
rect 5330 2615 5335 2635
rect 5305 2585 5335 2615
rect 5305 2565 5310 2585
rect 5330 2565 5335 2585
rect 5305 2535 5335 2565
rect 5305 2515 5310 2535
rect 5330 2515 5335 2535
rect 5305 2485 5335 2515
rect 5305 2465 5310 2485
rect 5330 2465 5335 2485
rect 5305 2435 5335 2465
rect 5305 2415 5310 2435
rect 5330 2415 5335 2435
rect 5305 2405 5335 2415
rect 5395 2685 5425 2695
rect 5395 2665 5400 2685
rect 5420 2665 5425 2685
rect 5395 2635 5425 2665
rect 5395 2615 5400 2635
rect 5420 2615 5425 2635
rect 5395 2585 5425 2615
rect 5395 2565 5400 2585
rect 5420 2565 5425 2585
rect 5395 2535 5425 2565
rect 5395 2515 5400 2535
rect 5420 2515 5425 2535
rect 5395 2485 5425 2515
rect 5395 2465 5400 2485
rect 5420 2465 5425 2485
rect 5395 2435 5425 2465
rect 5395 2415 5400 2435
rect 5420 2415 5425 2435
rect 5395 2405 5425 2415
rect 5485 2685 5515 2695
rect 5485 2665 5490 2685
rect 5510 2665 5515 2685
rect 5485 2635 5515 2665
rect 5485 2615 5490 2635
rect 5510 2615 5515 2635
rect 5485 2585 5515 2615
rect 5485 2565 5490 2585
rect 5510 2565 5515 2585
rect 5485 2535 5515 2565
rect 5485 2515 5490 2535
rect 5510 2515 5515 2535
rect 5485 2485 5515 2515
rect 5485 2465 5490 2485
rect 5510 2465 5515 2485
rect 5485 2435 5515 2465
rect 5485 2415 5490 2435
rect 5510 2415 5515 2435
rect 5485 2405 5515 2415
rect 5575 2685 5605 2695
rect 5575 2665 5580 2685
rect 5600 2665 5605 2685
rect 5575 2635 5605 2665
rect 5575 2615 5580 2635
rect 5600 2615 5605 2635
rect 5575 2585 5605 2615
rect 5575 2565 5580 2585
rect 5600 2565 5605 2585
rect 5575 2535 5605 2565
rect 5575 2515 5580 2535
rect 5600 2515 5605 2535
rect 5575 2485 5605 2515
rect 5575 2465 5580 2485
rect 5600 2465 5605 2485
rect 5575 2435 5605 2465
rect 5575 2415 5580 2435
rect 5600 2415 5605 2435
rect 5575 2405 5605 2415
rect 5665 2685 5695 2695
rect 5665 2665 5670 2685
rect 5690 2665 5695 2685
rect 5665 2635 5695 2665
rect 5665 2615 5670 2635
rect 5690 2615 5695 2635
rect 5665 2585 5695 2615
rect 5665 2565 5670 2585
rect 5690 2565 5695 2585
rect 5665 2535 5695 2565
rect 5665 2515 5670 2535
rect 5690 2515 5695 2535
rect 5665 2485 5695 2515
rect 5665 2465 5670 2485
rect 5690 2465 5695 2485
rect 5665 2435 5695 2465
rect 5665 2415 5670 2435
rect 5690 2415 5695 2435
rect 5665 2405 5695 2415
rect 5755 2685 5785 2695
rect 5755 2665 5760 2685
rect 5780 2665 5785 2685
rect 5755 2635 5785 2665
rect 5755 2615 5760 2635
rect 5780 2615 5785 2635
rect 5755 2585 5785 2615
rect 5755 2565 5760 2585
rect 5780 2565 5785 2585
rect 5755 2535 5785 2565
rect 5755 2515 5760 2535
rect 5780 2515 5785 2535
rect 5755 2485 5785 2515
rect 5755 2465 5760 2485
rect 5780 2465 5785 2485
rect 5755 2435 5785 2465
rect 5755 2415 5760 2435
rect 5780 2415 5785 2435
rect 5755 2405 5785 2415
rect 5845 2685 5875 2695
rect 5845 2665 5850 2685
rect 5870 2665 5875 2685
rect 5845 2635 5875 2665
rect 5845 2615 5850 2635
rect 5870 2615 5875 2635
rect 5845 2585 5875 2615
rect 5845 2565 5850 2585
rect 5870 2565 5875 2585
rect 5845 2535 5875 2565
rect 5845 2515 5850 2535
rect 5870 2515 5875 2535
rect 5845 2485 5875 2515
rect 5845 2465 5850 2485
rect 5870 2465 5875 2485
rect 5845 2435 5875 2465
rect 5845 2415 5850 2435
rect 5870 2415 5875 2435
rect 5845 2405 5875 2415
rect 5935 2685 5965 2695
rect 5935 2665 5940 2685
rect 5960 2665 5965 2685
rect 5935 2635 5965 2665
rect 5935 2615 5940 2635
rect 5960 2615 5965 2635
rect 5935 2585 5965 2615
rect 5935 2565 5940 2585
rect 5960 2565 5965 2585
rect 5935 2535 5965 2565
rect 5935 2515 5940 2535
rect 5960 2515 5965 2535
rect 5935 2485 5965 2515
rect 5935 2465 5940 2485
rect 5960 2465 5965 2485
rect 5935 2435 5965 2465
rect 5935 2415 5940 2435
rect 5960 2415 5965 2435
rect 5935 2405 5965 2415
rect 6025 2685 6055 2695
rect 6025 2665 6030 2685
rect 6050 2665 6055 2685
rect 6025 2635 6055 2665
rect 6025 2615 6030 2635
rect 6050 2615 6055 2635
rect 6025 2585 6055 2615
rect 6025 2565 6030 2585
rect 6050 2565 6055 2585
rect 6025 2535 6055 2565
rect 6025 2515 6030 2535
rect 6050 2515 6055 2535
rect 6025 2485 6055 2515
rect 6025 2465 6030 2485
rect 6050 2465 6055 2485
rect 6025 2435 6055 2465
rect 6025 2415 6030 2435
rect 6050 2415 6055 2435
rect 6025 2405 6055 2415
rect 6115 2685 6145 2695
rect 6115 2665 6120 2685
rect 6140 2665 6145 2685
rect 6115 2635 6145 2665
rect 6115 2615 6120 2635
rect 6140 2615 6145 2635
rect 6115 2585 6145 2615
rect 6115 2565 6120 2585
rect 6140 2565 6145 2585
rect 6115 2535 6145 2565
rect 6115 2515 6120 2535
rect 6140 2515 6145 2535
rect 6115 2485 6145 2515
rect 6115 2465 6120 2485
rect 6140 2465 6145 2485
rect 6115 2435 6145 2465
rect 6115 2415 6120 2435
rect 6140 2415 6145 2435
rect 6115 2405 6145 2415
rect 6205 2685 6235 2695
rect 6205 2665 6210 2685
rect 6230 2665 6235 2685
rect 6205 2635 6235 2665
rect 6205 2615 6210 2635
rect 6230 2615 6235 2635
rect 6205 2585 6235 2615
rect 6205 2565 6210 2585
rect 6230 2565 6235 2585
rect 6205 2535 6235 2565
rect 6205 2515 6210 2535
rect 6230 2515 6235 2535
rect 6205 2485 6235 2515
rect 6205 2465 6210 2485
rect 6230 2465 6235 2485
rect 6205 2435 6235 2465
rect 6205 2415 6210 2435
rect 6230 2415 6235 2435
rect 6205 2405 6235 2415
rect 6295 2685 6325 2695
rect 6295 2665 6300 2685
rect 6320 2665 6325 2685
rect 6295 2635 6325 2665
rect 6295 2615 6300 2635
rect 6320 2615 6325 2635
rect 6295 2585 6325 2615
rect 6295 2565 6300 2585
rect 6320 2565 6325 2585
rect 6295 2535 6325 2565
rect 6295 2515 6300 2535
rect 6320 2515 6325 2535
rect 6295 2485 6325 2515
rect 6295 2465 6300 2485
rect 6320 2465 6325 2485
rect 6295 2435 6325 2465
rect 6295 2415 6300 2435
rect 6320 2415 6325 2435
rect 6295 2405 6325 2415
rect 6385 2685 6415 2695
rect 6385 2665 6390 2685
rect 6410 2665 6415 2685
rect 6385 2635 6415 2665
rect 6385 2615 6390 2635
rect 6410 2615 6415 2635
rect 6385 2585 6415 2615
rect 6385 2565 6390 2585
rect 6410 2565 6415 2585
rect 6385 2535 6415 2565
rect 6385 2515 6390 2535
rect 6410 2515 6415 2535
rect 6385 2485 6415 2515
rect 6385 2465 6390 2485
rect 6410 2465 6415 2485
rect 6385 2435 6415 2465
rect 6385 2415 6390 2435
rect 6410 2415 6415 2435
rect 6385 2405 6415 2415
rect 6475 2685 6505 2695
rect 6475 2665 6480 2685
rect 6500 2665 6505 2685
rect 6475 2635 6505 2665
rect 6475 2615 6480 2635
rect 6500 2615 6505 2635
rect 6475 2585 6505 2615
rect 6475 2565 6480 2585
rect 6500 2565 6505 2585
rect 6475 2535 6505 2565
rect 6475 2515 6480 2535
rect 6500 2515 6505 2535
rect 6475 2485 6505 2515
rect 6475 2465 6480 2485
rect 6500 2465 6505 2485
rect 6475 2435 6505 2465
rect 6475 2415 6480 2435
rect 6500 2415 6505 2435
rect 6475 2405 6505 2415
rect 6565 2685 6595 2695
rect 6565 2665 6570 2685
rect 6590 2665 6595 2685
rect 6565 2635 6595 2665
rect 6565 2615 6570 2635
rect 6590 2615 6595 2635
rect 6565 2585 6595 2615
rect 6565 2565 6570 2585
rect 6590 2565 6595 2585
rect 6565 2535 6595 2565
rect 6565 2515 6570 2535
rect 6590 2515 6595 2535
rect 6565 2485 6595 2515
rect 6565 2465 6570 2485
rect 6590 2465 6595 2485
rect 6565 2435 6595 2465
rect 6565 2415 6570 2435
rect 6590 2415 6595 2435
rect 6565 2405 6595 2415
rect 6655 2685 6685 2695
rect 6655 2665 6660 2685
rect 6680 2665 6685 2685
rect 6655 2635 6685 2665
rect 6655 2615 6660 2635
rect 6680 2615 6685 2635
rect 6655 2585 6685 2615
rect 6655 2565 6660 2585
rect 6680 2565 6685 2585
rect 6655 2535 6685 2565
rect 6655 2515 6660 2535
rect 6680 2515 6685 2535
rect 6655 2485 6685 2515
rect 6655 2465 6660 2485
rect 6680 2465 6685 2485
rect 6655 2435 6685 2465
rect 6655 2415 6660 2435
rect 6680 2415 6685 2435
rect 6655 2405 6685 2415
rect 6745 2685 6775 2695
rect 6745 2665 6750 2685
rect 6770 2665 6775 2685
rect 6745 2635 6775 2665
rect 6745 2615 6750 2635
rect 6770 2615 6775 2635
rect 6745 2585 6775 2615
rect 6745 2565 6750 2585
rect 6770 2565 6775 2585
rect 6745 2535 6775 2565
rect 6745 2515 6750 2535
rect 6770 2515 6775 2535
rect 6745 2485 6775 2515
rect 6745 2465 6750 2485
rect 6770 2465 6775 2485
rect 6745 2435 6775 2465
rect 6745 2415 6750 2435
rect 6770 2415 6775 2435
rect 6745 2405 6775 2415
rect 4410 2385 4430 2405
rect 4500 2385 4520 2405
rect 4680 2385 4700 2405
rect 4400 2375 4440 2385
rect 4400 2355 4410 2375
rect 4430 2355 4440 2375
rect 4400 2345 4440 2355
rect 4490 2375 4530 2385
rect 4490 2355 4500 2375
rect 4520 2355 4530 2375
rect 4490 2345 4530 2355
rect 4580 2370 4620 2380
rect 4580 2350 4590 2370
rect 4610 2350 4620 2370
rect 4215 2315 4245 2345
rect 4580 2340 4620 2350
rect 4670 2375 4710 2385
rect 4670 2355 4680 2375
rect 4700 2355 4710 2375
rect 4670 2345 4710 2355
rect 4860 2340 4880 2405
rect 5040 2385 5060 2405
rect 5030 2375 5070 2385
rect 5030 2355 5040 2375
rect 5060 2355 5070 2375
rect 5030 2345 5070 2355
rect 5220 2340 5240 2405
rect 5400 2385 5420 2405
rect 5580 2385 5600 2405
rect 5760 2385 5780 2405
rect 5335 2375 5375 2385
rect 5335 2355 5345 2375
rect 5365 2355 5375 2375
rect 5335 2345 5375 2355
rect 5400 2375 5440 2385
rect 5400 2355 5410 2375
rect 5430 2355 5440 2375
rect 5400 2345 5440 2355
rect 5570 2375 5610 2385
rect 5570 2355 5580 2375
rect 5600 2355 5610 2375
rect 5570 2345 5610 2355
rect 5740 2375 5780 2385
rect 5740 2355 5750 2375
rect 5770 2355 5780 2375
rect 5740 2345 5780 2355
rect 5940 2340 5960 2405
rect 6120 2385 6140 2405
rect 6110 2375 6150 2385
rect 6110 2355 6120 2375
rect 6140 2355 6150 2375
rect 6110 2345 6150 2355
rect 6300 2340 6320 2405
rect 6480 2385 6500 2405
rect 6660 2385 6680 2405
rect 6750 2385 6770 2405
rect 6470 2375 6510 2385
rect 6470 2355 6480 2375
rect 6500 2355 6510 2375
rect 6470 2345 6510 2355
rect 6650 2375 6690 2385
rect 6650 2355 6660 2375
rect 6680 2355 6690 2375
rect 6650 2345 6690 2355
rect 6740 2375 6780 2385
rect 6740 2355 6750 2375
rect 6770 2355 6780 2375
rect 6740 2345 6780 2355
rect 4850 2330 4890 2340
rect 4850 2310 4860 2330
rect 4880 2310 4890 2330
rect 4850 2300 4890 2310
rect 5210 2330 5250 2340
rect 5210 2310 5220 2330
rect 5240 2310 5250 2330
rect 5210 2300 5250 2310
rect 5930 2330 5970 2340
rect 5930 2310 5940 2330
rect 5960 2310 5970 2330
rect 5930 2300 5970 2310
rect 6290 2330 6330 2340
rect 6290 2310 6300 2330
rect 6320 2310 6330 2330
rect 6290 2300 6330 2310
rect 3835 2260 3865 2290
rect 5030 2285 5070 2295
rect 5030 2265 5040 2285
rect 5060 2265 5070 2285
rect 5030 2255 5070 2265
rect 6110 2285 6150 2295
rect 6110 2265 6120 2285
rect 6140 2265 6150 2285
rect 6110 2255 6150 2265
rect 6845 2260 6875 2290
rect 4060 2165 4090 2195
rect 4675 2165 4705 2195
rect 4010 2115 4040 2145
rect 4105 2070 4135 2100
rect 4855 2070 4885 2100
rect 5800 2065 5830 2095
rect 7040 2065 7070 2095
rect 125 2015 2135 2055
rect -45 1715 130 1725
rect -45 1695 -35 1715
rect -15 1695 15 1715
rect 35 1695 65 1715
rect 85 1695 130 1715
rect -45 1685 130 1695
rect 650 1375 775 2015
rect 2010 1375 2135 2015
rect 4455 2040 4495 2050
rect 4455 2020 4465 2040
rect 4485 2020 4495 2040
rect 4455 2010 4495 2020
rect 4575 2040 4615 2050
rect 4575 2020 4585 2040
rect 4605 2020 4615 2040
rect 4575 2010 4615 2020
rect 4695 2040 4735 2050
rect 4695 2020 4705 2040
rect 4725 2020 4735 2040
rect 4695 2010 4735 2020
rect 4815 2040 4855 2050
rect 4815 2020 4825 2040
rect 4845 2020 4855 2040
rect 4815 2010 4855 2020
rect 4935 2040 4975 2050
rect 4935 2020 4945 2040
rect 4965 2020 4975 2040
rect 4935 2010 4975 2020
rect 5055 2040 5095 2050
rect 5055 2020 5065 2040
rect 5085 2020 5095 2040
rect 5055 2010 5095 2020
rect 5175 2040 5215 2050
rect 5175 2020 5185 2040
rect 5205 2020 5215 2040
rect 5175 2010 5215 2020
rect 5295 2040 5335 2050
rect 5295 2020 5305 2040
rect 5325 2020 5335 2040
rect 5295 2010 5335 2020
rect 5415 2040 5455 2050
rect 5415 2020 5425 2040
rect 5445 2020 5455 2040
rect 5415 2010 5455 2020
rect 5725 2040 5765 2050
rect 5725 2020 5735 2040
rect 5755 2020 5765 2040
rect 5725 2010 5765 2020
rect 5845 2040 5885 2050
rect 5845 2020 5855 2040
rect 5875 2020 5885 2040
rect 5845 2010 5885 2020
rect 5965 2040 6005 2050
rect 5965 2020 5975 2040
rect 5995 2020 6005 2040
rect 5965 2010 6005 2020
rect 6085 2040 6125 2050
rect 6085 2020 6095 2040
rect 6115 2020 6125 2040
rect 6085 2010 6125 2020
rect 6205 2040 6245 2050
rect 6205 2020 6215 2040
rect 6235 2020 6245 2040
rect 6205 2010 6245 2020
rect 6325 2040 6365 2050
rect 6325 2020 6335 2040
rect 6355 2020 6365 2040
rect 6325 2010 6365 2020
rect 6445 2040 6485 2050
rect 6445 2020 6455 2040
rect 6475 2020 6485 2040
rect 6445 2010 6485 2020
rect 6565 2040 6605 2050
rect 6565 2020 6575 2040
rect 6595 2020 6605 2040
rect 6565 2010 6605 2020
rect 6685 2040 6725 2050
rect 6685 2020 6695 2040
rect 6715 2020 6725 2040
rect 6685 2010 6725 2020
rect 4210 1995 4250 2005
rect 4210 1975 4220 1995
rect 4240 1975 4250 1995
rect 4210 1965 4250 1975
rect 4335 1995 4375 2005
rect 4335 1975 4345 1995
rect 4365 1975 4375 1995
rect 4335 1965 4375 1975
rect 4395 1995 4435 2005
rect 4395 1975 4405 1995
rect 4425 1975 4435 1995
rect 4395 1965 4435 1975
rect 4220 1945 4240 1965
rect 4345 1945 4365 1965
rect 4405 1945 4425 1965
rect 4465 1945 4485 2010
rect 4585 1945 4605 2010
rect 4705 1945 4725 2010
rect 4755 1995 4795 2005
rect 4755 1975 4765 1995
rect 4785 1975 4795 1995
rect 4755 1965 4795 1975
rect 4765 1945 4785 1965
rect 4825 1945 4845 2010
rect 4945 1945 4965 2010
rect 5065 1945 5085 2010
rect 5115 1995 5155 2005
rect 5115 1975 5125 1995
rect 5145 1975 5155 1995
rect 5115 1965 5155 1975
rect 5125 1945 5145 1965
rect 5185 1945 5205 2010
rect 5305 1945 5325 2010
rect 5355 1995 5395 2005
rect 5355 1975 5365 1995
rect 5385 1975 5395 1995
rect 5355 1965 5395 1975
rect 5365 1945 5385 1965
rect 5425 1945 5445 2010
rect 5475 1995 5515 2005
rect 5475 1975 5485 1995
rect 5505 1975 5515 1995
rect 5475 1965 5515 1975
rect 5535 1995 5575 2005
rect 5535 1975 5545 1995
rect 5565 1975 5575 1995
rect 5535 1965 5575 1975
rect 5605 1995 5645 2005
rect 5605 1975 5615 1995
rect 5635 1975 5645 1995
rect 5605 1965 5645 1975
rect 5665 1995 5705 2005
rect 5665 1975 5675 1995
rect 5695 1975 5705 1995
rect 5665 1965 5705 1975
rect 5485 1945 5505 1965
rect 5545 1945 5565 1965
rect 5615 1945 5635 1965
rect 5675 1945 5695 1965
rect 5735 1945 5755 2010
rect 5785 1995 5825 2005
rect 5785 1975 5795 1995
rect 5815 1975 5825 1995
rect 5785 1965 5825 1975
rect 5795 1945 5815 1965
rect 5855 1945 5875 2010
rect 5975 1945 5995 2010
rect 6025 1995 6065 2005
rect 6025 1975 6035 1995
rect 6055 1975 6065 1995
rect 6025 1965 6065 1975
rect 6035 1945 6055 1965
rect 6095 1945 6115 2010
rect 6215 1945 6235 2010
rect 6335 1945 6355 2010
rect 6385 1995 6425 2005
rect 6385 1975 6395 1995
rect 6415 1975 6425 1995
rect 6385 1965 6425 1975
rect 6395 1945 6415 1965
rect 6455 1945 6475 2010
rect 6575 1945 6595 2010
rect 6695 1945 6715 2010
rect 6745 1995 6785 2005
rect 6745 1975 6755 1995
rect 6775 1975 6785 1995
rect 6745 1965 6785 1975
rect 6805 1995 6845 2005
rect 6805 1975 6815 1995
rect 6835 1975 6845 1995
rect 6805 1965 6845 1975
rect 6755 1945 6775 1965
rect 6815 1945 6835 1965
rect 4160 1935 4190 1945
rect 4160 1915 4165 1935
rect 4185 1915 4190 1935
rect 4160 1885 4190 1915
rect 4160 1865 4165 1885
rect 4185 1865 4190 1885
rect 4160 1855 4190 1865
rect 4215 1935 4245 1945
rect 4215 1915 4220 1935
rect 4240 1915 4245 1935
rect 4215 1885 4245 1915
rect 4215 1865 4220 1885
rect 4240 1865 4245 1885
rect 4215 1855 4245 1865
rect 4270 1935 4300 1945
rect 4270 1915 4275 1935
rect 4295 1915 4300 1935
rect 4270 1885 4300 1915
rect 4270 1865 4275 1885
rect 4295 1865 4300 1885
rect 4270 1855 4300 1865
rect 4340 1935 4370 1945
rect 4340 1915 4345 1935
rect 4365 1915 4370 1935
rect 4340 1885 4370 1915
rect 4340 1865 4345 1885
rect 4365 1865 4370 1885
rect 4340 1855 4370 1865
rect 4400 1935 4430 1945
rect 4400 1915 4405 1935
rect 4425 1915 4430 1935
rect 4400 1885 4430 1915
rect 4400 1865 4405 1885
rect 4425 1865 4430 1885
rect 4400 1855 4430 1865
rect 4460 1935 4490 1945
rect 4460 1915 4465 1935
rect 4485 1915 4490 1935
rect 4460 1885 4490 1915
rect 4460 1865 4465 1885
rect 4485 1865 4490 1885
rect 4460 1855 4490 1865
rect 4520 1935 4550 1945
rect 4520 1915 4525 1935
rect 4545 1915 4550 1935
rect 4520 1885 4550 1915
rect 4520 1865 4525 1885
rect 4545 1865 4550 1885
rect 4520 1855 4550 1865
rect 4580 1935 4610 1945
rect 4580 1915 4585 1935
rect 4605 1915 4610 1935
rect 4580 1885 4610 1915
rect 4580 1865 4585 1885
rect 4605 1865 4610 1885
rect 4580 1855 4610 1865
rect 4640 1935 4670 1945
rect 4640 1915 4645 1935
rect 4665 1915 4670 1935
rect 4640 1885 4670 1915
rect 4640 1865 4645 1885
rect 4665 1865 4670 1885
rect 4640 1855 4670 1865
rect 4700 1935 4730 1945
rect 4700 1915 4705 1935
rect 4725 1915 4730 1935
rect 4700 1885 4730 1915
rect 4700 1865 4705 1885
rect 4725 1865 4730 1885
rect 4700 1855 4730 1865
rect 4760 1935 4790 1945
rect 4760 1915 4765 1935
rect 4785 1915 4790 1935
rect 4760 1885 4790 1915
rect 4760 1865 4765 1885
rect 4785 1865 4790 1885
rect 4760 1855 4790 1865
rect 4820 1935 4850 1945
rect 4820 1915 4825 1935
rect 4845 1915 4850 1935
rect 4820 1885 4850 1915
rect 4820 1865 4825 1885
rect 4845 1865 4850 1885
rect 4820 1855 4850 1865
rect 4880 1935 4910 1945
rect 4880 1915 4885 1935
rect 4905 1915 4910 1935
rect 4880 1885 4910 1915
rect 4880 1865 4885 1885
rect 4905 1865 4910 1885
rect 4880 1855 4910 1865
rect 4940 1935 4970 1945
rect 4940 1915 4945 1935
rect 4965 1915 4970 1935
rect 4940 1885 4970 1915
rect 4940 1865 4945 1885
rect 4965 1865 4970 1885
rect 4940 1855 4970 1865
rect 5000 1935 5030 1945
rect 5000 1915 5005 1935
rect 5025 1915 5030 1935
rect 5000 1885 5030 1915
rect 5000 1865 5005 1885
rect 5025 1865 5030 1885
rect 5000 1855 5030 1865
rect 5060 1935 5090 1945
rect 5060 1915 5065 1935
rect 5085 1915 5090 1935
rect 5060 1885 5090 1915
rect 5060 1865 5065 1885
rect 5085 1865 5090 1885
rect 5060 1855 5090 1865
rect 5120 1935 5150 1945
rect 5120 1915 5125 1935
rect 5145 1915 5150 1935
rect 5120 1885 5150 1915
rect 5120 1865 5125 1885
rect 5145 1865 5150 1885
rect 5120 1855 5150 1865
rect 5180 1935 5210 1945
rect 5180 1915 5185 1935
rect 5205 1915 5210 1935
rect 5180 1885 5210 1915
rect 5180 1865 5185 1885
rect 5205 1865 5210 1885
rect 5180 1855 5210 1865
rect 5240 1935 5270 1945
rect 5240 1915 5245 1935
rect 5265 1915 5270 1935
rect 5240 1885 5270 1915
rect 5240 1865 5245 1885
rect 5265 1865 5270 1885
rect 5240 1855 5270 1865
rect 5300 1935 5330 1945
rect 5300 1915 5305 1935
rect 5325 1915 5330 1935
rect 5300 1885 5330 1915
rect 5300 1865 5305 1885
rect 5325 1865 5330 1885
rect 5300 1855 5330 1865
rect 5360 1935 5390 1945
rect 5360 1915 5365 1935
rect 5385 1915 5390 1935
rect 5360 1885 5390 1915
rect 5360 1865 5365 1885
rect 5385 1865 5390 1885
rect 5360 1855 5390 1865
rect 5420 1935 5450 1945
rect 5420 1915 5425 1935
rect 5445 1915 5450 1935
rect 5420 1885 5450 1915
rect 5420 1865 5425 1885
rect 5445 1865 5450 1885
rect 5420 1855 5450 1865
rect 5480 1935 5510 1945
rect 5480 1915 5485 1935
rect 5505 1915 5510 1935
rect 5480 1885 5510 1915
rect 5480 1865 5485 1885
rect 5505 1865 5510 1885
rect 5480 1855 5510 1865
rect 5540 1935 5570 1945
rect 5540 1915 5545 1935
rect 5565 1915 5570 1935
rect 5540 1885 5570 1915
rect 5540 1865 5545 1885
rect 5565 1865 5570 1885
rect 5540 1855 5570 1865
rect 5610 1935 5640 1945
rect 5610 1915 5615 1935
rect 5635 1915 5640 1935
rect 5610 1885 5640 1915
rect 5610 1865 5615 1885
rect 5635 1865 5640 1885
rect 5610 1855 5640 1865
rect 5670 1935 5700 1945
rect 5670 1915 5675 1935
rect 5695 1915 5700 1935
rect 5670 1885 5700 1915
rect 5670 1865 5675 1885
rect 5695 1865 5700 1885
rect 5670 1855 5700 1865
rect 5730 1935 5760 1945
rect 5730 1915 5735 1935
rect 5755 1915 5760 1935
rect 5730 1885 5760 1915
rect 5730 1865 5735 1885
rect 5755 1865 5760 1885
rect 5730 1855 5760 1865
rect 5790 1935 5820 1945
rect 5790 1915 5795 1935
rect 5815 1915 5820 1935
rect 5790 1885 5820 1915
rect 5790 1865 5795 1885
rect 5815 1865 5820 1885
rect 5790 1855 5820 1865
rect 5850 1935 5880 1945
rect 5850 1915 5855 1935
rect 5875 1915 5880 1935
rect 5850 1885 5880 1915
rect 5850 1865 5855 1885
rect 5875 1865 5880 1885
rect 5850 1855 5880 1865
rect 5910 1935 5940 1945
rect 5910 1915 5915 1935
rect 5935 1915 5940 1935
rect 5910 1885 5940 1915
rect 5910 1865 5915 1885
rect 5935 1865 5940 1885
rect 5910 1855 5940 1865
rect 5970 1935 6000 1945
rect 5970 1915 5975 1935
rect 5995 1915 6000 1935
rect 5970 1885 6000 1915
rect 5970 1865 5975 1885
rect 5995 1865 6000 1885
rect 5970 1855 6000 1865
rect 6030 1935 6060 1945
rect 6030 1915 6035 1935
rect 6055 1915 6060 1935
rect 6030 1885 6060 1915
rect 6030 1865 6035 1885
rect 6055 1865 6060 1885
rect 6030 1855 6060 1865
rect 6090 1935 6120 1945
rect 6090 1915 6095 1935
rect 6115 1915 6120 1935
rect 6090 1885 6120 1915
rect 6090 1865 6095 1885
rect 6115 1865 6120 1885
rect 6090 1855 6120 1865
rect 6150 1935 6180 1945
rect 6150 1915 6155 1935
rect 6175 1915 6180 1935
rect 6150 1885 6180 1915
rect 6150 1865 6155 1885
rect 6175 1865 6180 1885
rect 6150 1855 6180 1865
rect 6210 1935 6240 1945
rect 6210 1915 6215 1935
rect 6235 1915 6240 1935
rect 6210 1885 6240 1915
rect 6210 1865 6215 1885
rect 6235 1865 6240 1885
rect 6210 1855 6240 1865
rect 6270 1935 6300 1945
rect 6270 1915 6275 1935
rect 6295 1915 6300 1935
rect 6270 1885 6300 1915
rect 6270 1865 6275 1885
rect 6295 1865 6300 1885
rect 6270 1855 6300 1865
rect 6330 1935 6360 1945
rect 6330 1915 6335 1935
rect 6355 1915 6360 1935
rect 6330 1885 6360 1915
rect 6330 1865 6335 1885
rect 6355 1865 6360 1885
rect 6330 1855 6360 1865
rect 6390 1935 6420 1945
rect 6390 1915 6395 1935
rect 6415 1915 6420 1935
rect 6390 1885 6420 1915
rect 6390 1865 6395 1885
rect 6415 1865 6420 1885
rect 6390 1855 6420 1865
rect 6450 1935 6480 1945
rect 6450 1915 6455 1935
rect 6475 1915 6480 1935
rect 6450 1885 6480 1915
rect 6450 1865 6455 1885
rect 6475 1865 6480 1885
rect 6450 1855 6480 1865
rect 6510 1935 6540 1945
rect 6510 1915 6515 1935
rect 6535 1915 6540 1935
rect 6510 1885 6540 1915
rect 6510 1865 6515 1885
rect 6535 1865 6540 1885
rect 6510 1855 6540 1865
rect 6570 1935 6600 1945
rect 6570 1915 6575 1935
rect 6595 1915 6600 1935
rect 6570 1885 6600 1915
rect 6570 1865 6575 1885
rect 6595 1865 6600 1885
rect 6570 1855 6600 1865
rect 6630 1935 6660 1945
rect 6630 1915 6635 1935
rect 6655 1915 6660 1935
rect 6630 1885 6660 1915
rect 6630 1865 6635 1885
rect 6655 1865 6660 1885
rect 6630 1855 6660 1865
rect 6690 1935 6720 1945
rect 6690 1915 6695 1935
rect 6715 1915 6720 1935
rect 6690 1885 6720 1915
rect 6690 1865 6695 1885
rect 6715 1865 6720 1885
rect 6690 1855 6720 1865
rect 6750 1935 6780 1945
rect 6750 1915 6755 1935
rect 6775 1915 6780 1935
rect 6750 1885 6780 1915
rect 6750 1865 6755 1885
rect 6775 1865 6780 1885
rect 6750 1855 6780 1865
rect 6810 1935 6840 1945
rect 6810 1915 6815 1935
rect 6835 1915 6840 1935
rect 6810 1885 6840 1915
rect 6810 1865 6815 1885
rect 6835 1865 6840 1885
rect 6810 1855 6840 1865
rect 4165 1835 4185 1855
rect 4275 1835 4295 1855
rect 4525 1835 4545 1855
rect 4645 1835 4665 1855
rect 4885 1835 4905 1855
rect 5005 1835 5025 1855
rect 5245 1835 5265 1855
rect 5365 1835 5385 1855
rect 5795 1835 5815 1855
rect 5915 1835 5935 1855
rect 6155 1835 6175 1855
rect 6275 1835 6295 1855
rect 6515 1835 6535 1855
rect 6635 1835 6655 1855
rect 4010 1800 4040 1830
rect 4155 1825 4190 1835
rect 4155 1805 4165 1825
rect 4185 1805 4190 1825
rect 4155 1795 4190 1805
rect 4210 1825 4250 1835
rect 4210 1805 4220 1825
rect 4240 1805 4250 1825
rect 4210 1795 4250 1805
rect 4270 1825 4305 1835
rect 4270 1805 4275 1825
rect 4295 1805 4305 1825
rect 4270 1795 4305 1805
rect 4425 1825 4465 1835
rect 4425 1805 4435 1825
rect 4455 1805 4465 1825
rect 4425 1795 4465 1805
rect 4515 1825 4555 1835
rect 4515 1805 4525 1825
rect 4545 1805 4555 1825
rect 4515 1795 4555 1805
rect 4635 1825 4675 1835
rect 4635 1805 4645 1825
rect 4665 1805 4675 1825
rect 4635 1795 4675 1805
rect 4755 1825 4795 1835
rect 4755 1805 4765 1825
rect 4785 1805 4795 1825
rect 4755 1795 4795 1805
rect 4875 1825 4915 1835
rect 4875 1805 4885 1825
rect 4905 1805 4915 1825
rect 4875 1795 4915 1805
rect 4995 1825 5035 1835
rect 4995 1805 5005 1825
rect 5025 1805 5035 1825
rect 4995 1795 5035 1805
rect 5115 1825 5155 1835
rect 5115 1805 5125 1825
rect 5145 1805 5155 1825
rect 5115 1795 5155 1805
rect 5235 1825 5275 1835
rect 5235 1805 5245 1825
rect 5265 1805 5275 1825
rect 5235 1795 5275 1805
rect 5355 1825 5395 1835
rect 5355 1805 5365 1825
rect 5385 1805 5395 1825
rect 5355 1795 5395 1805
rect 5445 1825 5485 1835
rect 5445 1805 5455 1825
rect 5475 1805 5485 1825
rect 5445 1795 5485 1805
rect 5695 1825 5735 1835
rect 5695 1805 5705 1825
rect 5725 1805 5735 1825
rect 5695 1795 5735 1805
rect 5785 1825 5825 1835
rect 5785 1805 5795 1825
rect 5815 1805 5825 1825
rect 5785 1795 5825 1805
rect 5905 1825 5945 1835
rect 5905 1805 5915 1825
rect 5935 1805 5945 1825
rect 5905 1795 5945 1805
rect 6025 1825 6065 1835
rect 6025 1805 6035 1825
rect 6055 1805 6065 1825
rect 6025 1795 6065 1805
rect 6145 1825 6185 1835
rect 6145 1805 6155 1825
rect 6175 1805 6185 1825
rect 6145 1795 6185 1805
rect 6265 1825 6305 1835
rect 6265 1805 6275 1825
rect 6295 1805 6305 1825
rect 6265 1795 6305 1805
rect 6385 1825 6425 1835
rect 6385 1805 6395 1825
rect 6415 1805 6425 1825
rect 6385 1795 6425 1805
rect 6505 1825 6545 1835
rect 6505 1805 6515 1825
rect 6535 1805 6545 1825
rect 6505 1795 6545 1805
rect 6625 1825 6665 1835
rect 6625 1805 6635 1825
rect 6655 1805 6665 1825
rect 6625 1795 6665 1805
rect 6715 1825 6755 1835
rect 6715 1805 6725 1825
rect 6745 1805 6755 1825
rect 6715 1795 6755 1805
rect 4425 1735 4465 1775
rect 4635 1765 4675 1775
rect 4635 1745 4645 1765
rect 4665 1745 4675 1765
rect 4635 1735 4675 1745
rect 4755 1735 4795 1775
rect 4995 1765 5035 1775
rect 4995 1745 5005 1765
rect 5025 1745 5035 1765
rect 4995 1735 5035 1745
rect 5115 1735 5155 1775
rect 5355 1765 5395 1775
rect 5355 1745 5365 1765
rect 5385 1745 5395 1765
rect 5355 1735 5395 1745
rect 5445 1735 5485 1775
rect 5695 1735 5735 1775
rect 5785 1765 5825 1775
rect 5785 1745 5795 1765
rect 5815 1745 5825 1765
rect 5785 1735 5825 1745
rect 6025 1735 6065 1775
rect 6145 1765 6185 1775
rect 6145 1745 6155 1765
rect 6175 1745 6185 1765
rect 6145 1735 6185 1745
rect 6385 1735 6425 1775
rect 6505 1765 6545 1775
rect 6505 1745 6515 1765
rect 6535 1745 6545 1765
rect 6505 1735 6545 1745
rect 6715 1735 6755 1775
rect 3590 1680 3620 1710
rect 4105 1680 4135 1710
rect 4160 1680 4190 1710
rect 4270 1680 4300 1710
rect 4815 1705 4855 1715
rect 4815 1685 4825 1705
rect 4845 1685 4855 1705
rect 4815 1675 4855 1685
rect 4875 1705 4915 1715
rect 4875 1685 4885 1705
rect 4905 1685 4915 1705
rect 4875 1675 4915 1685
rect 5115 1705 5155 1715
rect 5115 1685 5125 1705
rect 5145 1685 5155 1705
rect 5115 1675 5155 1685
rect 5355 1705 5395 1715
rect 5355 1685 5365 1705
rect 5385 1685 5395 1705
rect 5355 1675 5395 1685
rect 5785 1705 5825 1715
rect 5785 1685 5795 1705
rect 5815 1685 5825 1705
rect 5785 1675 5825 1685
rect 6025 1705 6065 1715
rect 6025 1685 6035 1705
rect 6055 1685 6065 1705
rect 6025 1675 6065 1685
rect 6265 1705 6305 1715
rect 6265 1685 6275 1705
rect 6295 1685 6305 1705
rect 6265 1675 6305 1685
rect 6325 1705 6365 1715
rect 6325 1685 6335 1705
rect 6355 1685 6365 1705
rect 6325 1675 6365 1685
rect 6845 1680 6875 1710
rect 4755 1660 4795 1670
rect 4755 1640 4765 1660
rect 4785 1640 4795 1660
rect 4755 1630 4795 1640
rect 4765 1610 4785 1630
rect 4885 1610 4905 1675
rect 4995 1660 5035 1670
rect 4995 1640 5005 1660
rect 5025 1640 5035 1660
rect 4995 1630 5035 1640
rect 5005 1610 5025 1630
rect 5125 1610 5145 1675
rect 5235 1660 5275 1670
rect 5235 1640 5245 1660
rect 5265 1640 5275 1660
rect 5235 1630 5275 1640
rect 5245 1610 5265 1630
rect 5365 1610 5385 1675
rect 5795 1610 5815 1675
rect 5905 1660 5945 1670
rect 5905 1640 5915 1660
rect 5935 1640 5945 1660
rect 5905 1630 5945 1640
rect 5915 1610 5935 1630
rect 6035 1610 6055 1675
rect 6145 1660 6185 1670
rect 6145 1640 6155 1660
rect 6175 1640 6185 1660
rect 6145 1630 6185 1640
rect 6155 1610 6175 1630
rect 6275 1610 6295 1675
rect 6385 1660 6425 1670
rect 6385 1640 6395 1660
rect 6415 1640 6425 1660
rect 6385 1630 6425 1640
rect 6395 1610 6415 1630
rect 2345 1570 2385 1605
rect 3425 1600 3470 1605
rect 3425 1575 3435 1600
rect 3460 1575 3470 1600
rect 3590 1575 3620 1605
rect 4760 1600 4790 1610
rect 4760 1580 4765 1600
rect 4785 1580 4790 1600
rect 3425 1570 3470 1575
rect 4760 1570 4790 1580
rect 4820 1600 4850 1610
rect 4820 1580 4825 1600
rect 4845 1580 4850 1600
rect 4820 1570 4850 1580
rect 4880 1600 4910 1610
rect 4880 1580 4885 1600
rect 4905 1580 4910 1600
rect 4880 1570 4910 1580
rect 4940 1600 4970 1610
rect 4940 1580 4945 1600
rect 4965 1580 4970 1600
rect 4940 1570 4970 1580
rect 5000 1600 5030 1610
rect 5000 1580 5005 1600
rect 5025 1580 5030 1600
rect 5000 1570 5030 1580
rect 5060 1600 5090 1610
rect 5060 1580 5065 1600
rect 5085 1580 5090 1600
rect 5060 1570 5090 1580
rect 5120 1600 5150 1610
rect 5120 1580 5125 1600
rect 5145 1580 5150 1600
rect 5120 1570 5150 1580
rect 5180 1600 5210 1610
rect 5180 1580 5185 1600
rect 5205 1580 5210 1600
rect 5180 1570 5210 1580
rect 5240 1600 5270 1610
rect 5240 1580 5245 1600
rect 5265 1580 5270 1600
rect 5240 1570 5270 1580
rect 5300 1600 5330 1610
rect 5300 1580 5305 1600
rect 5325 1580 5330 1600
rect 5300 1570 5330 1580
rect 5360 1600 5390 1610
rect 5360 1580 5365 1600
rect 5385 1580 5390 1600
rect 5360 1570 5390 1580
rect 5790 1600 5820 1610
rect 5790 1580 5795 1600
rect 5815 1580 5820 1600
rect 5790 1570 5820 1580
rect 5850 1600 5880 1610
rect 5850 1580 5855 1600
rect 5875 1580 5880 1600
rect 5850 1570 5880 1580
rect 5910 1600 5940 1610
rect 5910 1580 5915 1600
rect 5935 1580 5940 1600
rect 5910 1570 5940 1580
rect 5970 1600 6000 1610
rect 5970 1580 5975 1600
rect 5995 1580 6000 1600
rect 5970 1570 6000 1580
rect 6030 1600 6060 1610
rect 6030 1580 6035 1600
rect 6055 1580 6060 1600
rect 6030 1570 6060 1580
rect 6090 1600 6120 1610
rect 6090 1580 6095 1600
rect 6115 1580 6120 1600
rect 6090 1570 6120 1580
rect 6150 1600 6180 1610
rect 6150 1580 6155 1600
rect 6175 1580 6180 1600
rect 6150 1570 6180 1580
rect 6210 1600 6240 1610
rect 6210 1580 6215 1600
rect 6235 1580 6240 1600
rect 6210 1570 6240 1580
rect 6270 1600 6300 1610
rect 6270 1580 6275 1600
rect 6295 1580 6300 1600
rect 6270 1570 6300 1580
rect 6330 1600 6360 1610
rect 6330 1580 6335 1600
rect 6355 1580 6360 1600
rect 6330 1570 6360 1580
rect 6390 1600 6420 1610
rect 6390 1580 6395 1600
rect 6415 1580 6420 1600
rect 6390 1570 6420 1580
rect 2345 1425 2365 1570
rect 3425 1540 3470 1545
rect 3425 1515 3435 1540
rect 3460 1515 3470 1540
rect 3590 1515 3620 1545
rect 4060 1515 4090 1545
rect 4755 1540 4795 1550
rect 4755 1520 4765 1540
rect 4785 1520 4795 1540
rect 3425 1510 3470 1515
rect 4755 1510 4795 1520
rect 2385 1485 2420 1510
rect 4825 1500 4845 1570
rect 4945 1500 4965 1570
rect 5065 1500 5085 1570
rect 5185 1500 5205 1570
rect 5305 1500 5325 1570
rect 5855 1500 5875 1570
rect 5975 1500 5995 1570
rect 6095 1500 6115 1570
rect 6215 1500 6235 1570
rect 6335 1500 6355 1570
rect 6385 1540 6425 1550
rect 6385 1520 6395 1540
rect 6415 1520 6425 1540
rect 6385 1510 6425 1520
rect 6845 1515 6875 1545
rect 4815 1490 4855 1500
rect 3425 1450 3465 1485
rect 4815 1470 4825 1490
rect 4845 1470 4855 1490
rect 4815 1460 4855 1470
rect 4935 1490 4975 1500
rect 4935 1470 4945 1490
rect 4965 1470 4975 1490
rect 4935 1460 4975 1470
rect 5055 1490 5095 1500
rect 5055 1470 5065 1490
rect 5085 1470 5095 1490
rect 5055 1460 5095 1470
rect 5175 1490 5215 1500
rect 5175 1470 5185 1490
rect 5205 1470 5215 1490
rect 5175 1460 5215 1470
rect 5295 1490 5335 1500
rect 5295 1470 5305 1490
rect 5325 1470 5335 1490
rect 5295 1460 5335 1470
rect 5845 1490 5885 1500
rect 5845 1470 5855 1490
rect 5875 1470 5885 1490
rect 5845 1460 5885 1470
rect 5965 1490 6005 1500
rect 5965 1470 5975 1490
rect 5995 1470 6005 1490
rect 5965 1460 6005 1470
rect 6085 1490 6125 1500
rect 6085 1470 6095 1490
rect 6115 1470 6125 1490
rect 6085 1460 6125 1470
rect 6205 1490 6245 1500
rect 6205 1470 6215 1490
rect 6235 1470 6245 1490
rect 6205 1460 6245 1470
rect 6325 1490 6365 1500
rect 6325 1470 6335 1490
rect 6355 1470 6365 1490
rect 6325 1460 6365 1470
rect 2345 1390 2385 1425
rect 125 1335 2135 1375
rect 3390 1365 3425 1390
rect 650 690 775 1335
rect 1330 690 1455 1335
rect 2010 695 2135 1335
rect 2340 1360 2385 1365
rect 2340 1335 2350 1360
rect 2375 1335 2385 1360
rect 2340 1330 2385 1335
rect 2340 1300 2385 1310
rect 3445 1305 3465 1450
rect 4425 1435 4465 1445
rect 4425 1415 4435 1435
rect 4455 1415 4465 1435
rect 4425 1405 4465 1415
rect 5505 1435 5545 1445
rect 5505 1415 5515 1435
rect 5535 1415 5545 1435
rect 5505 1405 5545 1415
rect 5635 1435 5675 1445
rect 5635 1415 5645 1435
rect 5665 1415 5675 1435
rect 5635 1405 5675 1415
rect 6715 1435 6755 1445
rect 6715 1415 6725 1435
rect 6745 1415 6755 1435
rect 6715 1405 6755 1415
rect 2340 1275 2350 1300
rect 2375 1275 2385 1300
rect 2340 1265 2385 1275
rect 3425 1270 3465 1305
rect 4430 1395 4460 1405
rect 4430 1375 4435 1395
rect 4455 1375 4460 1395
rect 4430 1345 4460 1375
rect 4430 1325 4435 1345
rect 4455 1325 4460 1345
rect 4430 1295 4460 1325
rect 4430 1275 4435 1295
rect 4455 1275 4460 1295
rect 4430 1245 4460 1275
rect 4430 1225 4435 1245
rect 4455 1225 4460 1245
rect 4430 1195 4460 1225
rect 4430 1175 4435 1195
rect 4455 1175 4460 1195
rect 4430 1165 4460 1175
rect 4970 1395 5000 1405
rect 4970 1375 4975 1395
rect 4995 1375 5000 1395
rect 4970 1345 5000 1375
rect 4970 1325 4975 1345
rect 4995 1325 5000 1345
rect 4970 1295 5000 1325
rect 4970 1275 4975 1295
rect 4995 1275 5000 1295
rect 4970 1245 5000 1275
rect 4970 1225 4975 1245
rect 4995 1225 5000 1245
rect 4970 1195 5000 1225
rect 4970 1175 4975 1195
rect 4995 1175 5000 1195
rect 4970 1165 5000 1175
rect 5510 1395 5540 1405
rect 5510 1375 5515 1395
rect 5535 1375 5540 1395
rect 5510 1345 5540 1375
rect 5510 1325 5515 1345
rect 5535 1325 5540 1345
rect 5510 1295 5540 1325
rect 5510 1275 5515 1295
rect 5535 1275 5540 1295
rect 5510 1245 5540 1275
rect 5510 1225 5515 1245
rect 5535 1225 5540 1245
rect 5510 1195 5540 1225
rect 5510 1175 5515 1195
rect 5535 1175 5540 1195
rect 5510 1165 5540 1175
rect 5640 1395 5670 1405
rect 5640 1375 5645 1395
rect 5665 1375 5670 1395
rect 5640 1345 5670 1375
rect 5640 1325 5645 1345
rect 5665 1325 5670 1345
rect 5640 1295 5670 1325
rect 5640 1275 5645 1295
rect 5665 1275 5670 1295
rect 5640 1245 5670 1275
rect 5640 1225 5645 1245
rect 5665 1225 5670 1245
rect 5640 1195 5670 1225
rect 5640 1175 5645 1195
rect 5665 1175 5670 1195
rect 5640 1165 5670 1175
rect 6180 1395 6210 1405
rect 6180 1375 6185 1395
rect 6205 1375 6210 1395
rect 6180 1345 6210 1375
rect 6180 1325 6185 1345
rect 6205 1325 6210 1345
rect 6180 1295 6210 1325
rect 6180 1275 6185 1295
rect 6205 1275 6210 1295
rect 6180 1245 6210 1275
rect 6180 1225 6185 1245
rect 6205 1225 6210 1245
rect 6180 1195 6210 1225
rect 6180 1175 6185 1195
rect 6205 1175 6210 1195
rect 6180 1165 6210 1175
rect 6720 1395 6750 1405
rect 6720 1375 6725 1395
rect 6745 1375 6750 1395
rect 6720 1345 6750 1375
rect 6720 1325 6725 1345
rect 6745 1325 6750 1345
rect 6720 1295 6750 1325
rect 6720 1275 6725 1295
rect 6745 1275 6750 1295
rect 6720 1245 6750 1275
rect 6720 1225 6725 1245
rect 6745 1225 6750 1245
rect 6720 1195 6750 1225
rect 6720 1175 6725 1195
rect 6745 1175 6750 1195
rect 6720 1165 6750 1175
rect 4530 1110 4570 1120
rect 4530 1090 4540 1110
rect 4560 1090 4570 1110
rect 4530 1080 4570 1090
rect 4610 1110 4650 1120
rect 4610 1090 4620 1110
rect 4640 1090 4650 1110
rect 4610 1080 4650 1090
rect 4690 1110 4730 1120
rect 4690 1090 4700 1110
rect 4720 1090 4730 1110
rect 4690 1080 4730 1090
rect 4770 1110 4810 1120
rect 4770 1090 4780 1110
rect 4800 1090 4810 1110
rect 4770 1080 4810 1090
rect 4850 1110 4890 1120
rect 4850 1090 4860 1110
rect 4880 1090 4890 1110
rect 4850 1080 4890 1090
rect 4930 1110 4970 1120
rect 4930 1090 4940 1110
rect 4960 1090 4970 1110
rect 4930 1080 4970 1090
rect 5010 1110 5050 1120
rect 5010 1090 5020 1110
rect 5040 1090 5050 1110
rect 5010 1080 5050 1090
rect 5090 1110 5130 1120
rect 5090 1090 5100 1110
rect 5120 1090 5130 1110
rect 5090 1080 5130 1090
rect 5170 1110 5210 1120
rect 5170 1090 5180 1110
rect 5200 1090 5210 1110
rect 5170 1080 5210 1090
rect 5250 1110 5290 1120
rect 5250 1090 5260 1110
rect 5280 1090 5290 1110
rect 5250 1080 5290 1090
rect 5330 1110 5370 1120
rect 5330 1090 5340 1110
rect 5360 1090 5370 1110
rect 5330 1080 5370 1090
rect 5410 1110 5450 1120
rect 5410 1090 5420 1110
rect 5440 1090 5450 1110
rect 5410 1080 5450 1090
rect 5490 1110 5530 1120
rect 5490 1090 5500 1110
rect 5520 1090 5530 1110
rect 5490 1080 5530 1090
rect 5570 1110 5610 1120
rect 5570 1090 5580 1110
rect 5600 1090 5610 1110
rect 5570 1080 5610 1090
rect 5650 1110 5690 1120
rect 5650 1090 5660 1110
rect 5680 1090 5690 1110
rect 5650 1080 5690 1090
rect 5730 1110 5770 1120
rect 5730 1090 5740 1110
rect 5760 1090 5770 1110
rect 5730 1080 5770 1090
rect 5810 1110 5850 1120
rect 5810 1090 5820 1110
rect 5840 1090 5850 1110
rect 5810 1080 5850 1090
rect 5890 1110 5930 1120
rect 5890 1090 5900 1110
rect 5920 1090 5930 1110
rect 5890 1080 5930 1090
rect 5970 1110 6010 1120
rect 5970 1090 5980 1110
rect 6000 1090 6010 1110
rect 5970 1080 6010 1090
rect 6050 1110 6090 1120
rect 6050 1090 6060 1110
rect 6080 1090 6090 1110
rect 6050 1080 6090 1090
rect 6130 1110 6170 1120
rect 6130 1090 6140 1110
rect 6160 1090 6170 1110
rect 6130 1080 6170 1090
rect 6210 1110 6250 1120
rect 6210 1090 6220 1110
rect 6240 1090 6250 1110
rect 6210 1080 6250 1090
rect 6290 1110 6330 1120
rect 6290 1090 6300 1110
rect 6320 1090 6330 1110
rect 6290 1080 6330 1090
rect 6370 1110 6410 1120
rect 6370 1090 6380 1110
rect 6400 1090 6410 1110
rect 6370 1080 6410 1090
rect 6450 1110 6490 1120
rect 6450 1090 6460 1110
rect 6480 1090 6490 1110
rect 6450 1080 6490 1090
rect 6530 1110 6570 1120
rect 6530 1090 6540 1110
rect 6560 1090 6570 1110
rect 6530 1080 6570 1090
rect 4540 1060 4560 1080
rect 5580 1060 5600 1080
rect 4535 1050 4565 1060
rect 4535 1035 4540 1050
rect 4520 1030 4540 1035
rect 4560 1030 4565 1050
rect 2345 1025 2390 1030
rect 2345 1000 2355 1025
rect 2380 1000 2390 1025
rect 2345 995 2390 1000
rect 3060 1025 3105 1030
rect 3060 1000 3070 1025
rect 3095 1000 3105 1025
rect 3590 1000 3620 1030
rect 4010 1000 4040 1030
rect 4495 1025 4565 1030
rect 4495 1005 4500 1025
rect 4520 1005 4565 1025
rect 4495 1000 4565 1005
rect 3060 995 3105 1000
rect 4520 995 4540 1000
rect 4535 980 4540 995
rect 4560 980 4565 1000
rect 4535 970 4565 980
rect 5575 1050 5605 1060
rect 5575 1030 5580 1050
rect 5600 1030 5605 1050
rect 5575 1000 5605 1030
rect 5575 980 5580 1000
rect 5600 980 5605 1000
rect 5575 970 5605 980
rect 6615 1050 6645 1060
rect 6615 1030 6620 1050
rect 6640 1030 6645 1050
rect 6615 1000 6645 1030
rect 6615 980 6620 1000
rect 6640 980 6645 1000
rect 6615 970 6645 980
rect 2460 965 2505 970
rect 2460 940 2470 965
rect 2495 940 2505 965
rect 2460 935 2505 940
rect 3530 910 3550 935
rect 2460 905 2505 910
rect 2460 880 2470 905
rect 2495 880 2505 905
rect 2460 875 2505 880
rect 4685 895 4715 905
rect 4685 875 4690 895
rect 4710 875 4715 895
rect 3835 840 3865 870
rect 4685 845 4715 875
rect 2460 825 2505 830
rect 2460 800 2470 825
rect 2495 800 2505 825
rect 2460 795 2505 800
rect 4685 825 4690 845
rect 4710 825 4715 845
rect 4685 815 4715 825
rect 4775 895 4805 905
rect 4775 875 4780 895
rect 4800 875 4805 895
rect 4775 845 4805 875
rect 4775 825 4780 845
rect 4800 825 4805 845
rect 4775 815 4805 825
rect 4845 895 4875 905
rect 4845 875 4850 895
rect 4870 875 4875 895
rect 4845 845 4875 875
rect 4845 825 4850 845
rect 4870 825 4875 845
rect 4845 815 4875 825
rect 4935 895 4965 905
rect 4935 875 4940 895
rect 4960 875 4965 895
rect 4935 845 4965 875
rect 4935 825 4940 845
rect 4960 825 4965 845
rect 4935 815 4965 825
rect 5025 895 5055 905
rect 5025 875 5030 895
rect 5050 875 5055 895
rect 5025 845 5055 875
rect 5025 825 5030 845
rect 5050 825 5055 845
rect 5025 815 5055 825
rect 5115 895 5145 905
rect 5115 875 5120 895
rect 5140 875 5145 895
rect 5115 845 5145 875
rect 5115 825 5120 845
rect 5140 825 5145 845
rect 5115 815 5145 825
rect 5205 895 5235 905
rect 5205 875 5210 895
rect 5230 875 5235 895
rect 5205 845 5235 875
rect 5205 825 5210 845
rect 5230 825 5235 845
rect 5205 815 5235 825
rect 5295 895 5325 905
rect 5295 875 5300 895
rect 5320 875 5325 895
rect 5295 845 5325 875
rect 5295 825 5300 845
rect 5320 825 5325 845
rect 5295 815 5325 825
rect 5385 895 5415 905
rect 5385 875 5390 895
rect 5410 875 5415 895
rect 5385 845 5415 875
rect 5385 825 5390 845
rect 5410 825 5415 845
rect 5385 815 5415 825
rect 5475 895 5505 905
rect 5475 875 5480 895
rect 5500 875 5505 895
rect 5475 845 5505 875
rect 5475 825 5480 845
rect 5500 825 5505 845
rect 5475 815 5505 825
rect 5565 895 5595 905
rect 5565 875 5570 895
rect 5590 875 5595 895
rect 5565 845 5595 875
rect 5565 825 5570 845
rect 5590 825 5595 845
rect 5565 815 5595 825
rect 5655 895 5685 905
rect 5655 875 5660 895
rect 5680 875 5685 895
rect 5655 845 5685 875
rect 5655 825 5660 845
rect 5680 825 5685 845
rect 5655 815 5685 825
rect 5745 895 5775 905
rect 5745 875 5750 895
rect 5770 875 5775 895
rect 5745 845 5775 875
rect 5745 825 5750 845
rect 5770 825 5775 845
rect 5745 815 5775 825
rect 5835 895 5865 905
rect 5835 875 5840 895
rect 5860 875 5865 895
rect 5835 845 5865 875
rect 5835 825 5840 845
rect 5860 825 5865 845
rect 5835 815 5865 825
rect 5925 895 5955 905
rect 5925 875 5930 895
rect 5950 875 5955 895
rect 5925 845 5955 875
rect 5925 825 5930 845
rect 5950 825 5955 845
rect 5925 815 5955 825
rect 6015 895 6045 905
rect 6015 875 6020 895
rect 6040 875 6045 895
rect 6015 845 6045 875
rect 6015 825 6020 845
rect 6040 825 6045 845
rect 6015 815 6045 825
rect 6105 895 6135 905
rect 6105 875 6110 895
rect 6130 875 6135 895
rect 6105 845 6135 875
rect 6105 825 6110 845
rect 6130 825 6135 845
rect 6105 815 6135 825
rect 6195 895 6225 905
rect 6195 875 6200 895
rect 6220 875 6225 895
rect 6195 845 6225 875
rect 6195 825 6200 845
rect 6220 825 6225 845
rect 6195 815 6225 825
rect 6285 895 6315 905
rect 6285 875 6290 895
rect 6310 875 6315 895
rect 6285 845 6315 875
rect 6285 825 6290 845
rect 6310 825 6315 845
rect 6285 815 6315 825
rect 6375 895 6405 905
rect 6375 875 6380 895
rect 6400 875 6405 895
rect 6375 845 6405 875
rect 6375 825 6380 845
rect 6400 825 6405 845
rect 6375 815 6405 825
rect 6465 895 6495 905
rect 6465 875 6470 895
rect 6490 875 6495 895
rect 6465 845 6495 875
rect 6465 825 6470 845
rect 6490 825 6495 845
rect 6465 815 6495 825
rect 6555 895 6585 905
rect 6555 875 6560 895
rect 6580 875 6585 895
rect 6555 845 6585 875
rect 6555 825 6560 845
rect 6580 825 6585 845
rect 6555 815 6585 825
rect 3525 770 3545 795
rect 2460 765 2505 770
rect 2460 740 2470 765
rect 2495 740 2505 765
rect 2460 735 2505 740
rect 6845 700 6875 730
rect -840 -405 -795 -400
rect -840 -430 -830 -405
rect -805 -430 -795 -405
rect -840 -435 -795 -430
rect 189 -435 269 -400
rect -840 -465 -795 -460
rect -840 -490 -830 -465
rect -805 -490 -795 -465
rect -840 -495 -795 -490
rect 189 -495 229 -460
rect -840 -525 -795 -520
rect -840 -550 -830 -525
rect -805 -550 -795 -525
rect -840 -555 -795 -550
rect 154 -580 189 -555
rect -875 -615 -795 -580
rect -875 -880 -855 -615
rect 209 -640 229 -495
rect -835 -675 -795 -640
rect 189 -675 229 -640
rect -835 -820 -815 -675
rect 249 -700 269 -435
rect 189 -735 269 -700
rect -795 -760 -760 -735
rect 189 -795 269 -760
rect -835 -855 -795 -820
rect 189 -855 229 -820
rect -875 -915 -795 -880
rect -975 -945 -935 -940
rect -975 -970 -970 -945
rect -945 -970 -935 -945
rect -975 -975 -935 -970
rect -840 -945 -795 -940
rect -840 -970 -830 -945
rect -805 -970 -795 -945
rect -840 -975 -795 -970
rect -21 -945 24 -940
rect -21 -970 -11 -945
rect 14 -970 24 -945
rect -21 -975 24 -970
rect 154 -1000 189 -915
rect -875 -1035 -795 -1000
rect -875 -1300 -855 -1035
rect 209 -1060 229 -855
rect -835 -1095 -795 -1060
rect 189 -1095 229 -1060
rect -835 -1240 -815 -1095
rect 249 -1120 269 -795
rect 189 -1155 269 -1120
rect -795 -1180 -760 -1155
rect 189 -1215 269 -1180
rect -835 -1275 -795 -1240
rect 189 -1275 229 -1240
rect -875 -1335 -795 -1300
rect 154 -1360 189 -1335
rect -840 -1365 -795 -1360
rect -840 -1390 -830 -1365
rect -805 -1390 -795 -1365
rect -840 -1395 -795 -1390
rect 209 -1420 229 -1275
rect -840 -1425 -795 -1420
rect -840 -1450 -830 -1425
rect -805 -1450 -795 -1425
rect -840 -1455 -795 -1450
rect 189 -1455 229 -1420
rect -840 -1485 -795 -1475
rect 249 -1480 269 -1215
rect -840 -1510 -830 -1485
rect -805 -1510 -795 -1485
rect -840 -1520 -795 -1510
rect 189 -1515 269 -1480
<< viali >>
rect 4555 2915 4575 2935
rect 4590 2725 4610 2745
rect 4770 2725 4790 2745
rect 4950 2725 4970 2745
rect 5130 2725 5150 2745
rect 5310 2725 5330 2745
rect 5490 2725 5510 2745
rect 5670 2725 5690 2745
rect 5850 2725 5870 2745
rect 6030 2725 6050 2745
rect 6210 2725 6230 2745
rect 6390 2725 6410 2745
rect 6570 2725 6590 2745
rect 4500 2355 4520 2375
rect 4590 2350 4610 2370
rect 4680 2355 4700 2375
rect 5040 2355 5060 2375
rect 5345 2355 5365 2375
rect 5410 2355 5430 2375
rect 5580 2355 5600 2375
rect 5750 2355 5770 2375
rect 6120 2355 6140 2375
rect 6480 2355 6500 2375
rect 6660 2355 6680 2375
rect 4860 2310 4880 2330
rect 5220 2310 5240 2330
rect 5940 2310 5960 2330
rect 6300 2310 6320 2330
rect 5040 2265 5060 2285
rect 6120 2265 6140 2285
rect -35 1695 -15 1715
rect 4465 2020 4485 2040
rect 4585 2020 4605 2040
rect 4705 2020 4725 2040
rect 4825 2020 4845 2040
rect 4945 2020 4965 2040
rect 5065 2020 5085 2040
rect 5185 2020 5205 2040
rect 5305 2020 5325 2040
rect 5425 2020 5445 2040
rect 5735 2020 5755 2040
rect 5855 2020 5875 2040
rect 5975 2020 5995 2040
rect 6095 2020 6115 2040
rect 6215 2020 6235 2040
rect 6335 2020 6355 2040
rect 6455 2020 6475 2040
rect 6575 2020 6595 2040
rect 6695 2020 6715 2040
rect 4220 1975 4240 1995
rect 4405 1975 4425 1995
rect 4765 1975 4785 1995
rect 5125 1975 5145 1995
rect 5365 1975 5385 1995
rect 5485 1975 5505 1995
rect 5675 1975 5695 1995
rect 5795 1975 5815 1995
rect 6035 1975 6055 1995
rect 6395 1975 6415 1995
rect 6755 1975 6775 1995
rect 4165 1805 4185 1825
rect 4220 1805 4240 1825
rect 4275 1805 4295 1825
rect 4435 1805 4455 1825
rect 4525 1805 4545 1825
rect 4645 1805 4665 1825
rect 4765 1805 4785 1825
rect 4885 1805 4905 1825
rect 5005 1805 5025 1825
rect 5125 1805 5145 1825
rect 5245 1805 5265 1825
rect 5365 1805 5385 1825
rect 5455 1805 5475 1825
rect 5705 1805 5725 1825
rect 5795 1805 5815 1825
rect 5915 1805 5935 1825
rect 6035 1805 6055 1825
rect 6155 1805 6175 1825
rect 6275 1805 6295 1825
rect 6395 1805 6415 1825
rect 6515 1805 6535 1825
rect 6635 1805 6655 1825
rect 6725 1805 6745 1825
rect 4645 1745 4665 1765
rect 5005 1745 5025 1765
rect 5365 1745 5385 1765
rect 5795 1745 5815 1765
rect 6155 1745 6175 1765
rect 6515 1745 6535 1765
rect 4825 1685 4845 1705
rect 4885 1685 4905 1705
rect 5125 1685 5145 1705
rect 5365 1685 5385 1705
rect 5795 1685 5815 1705
rect 6035 1685 6055 1705
rect 6275 1685 6295 1705
rect 6335 1685 6355 1705
rect 4765 1640 4785 1660
rect 5005 1640 5025 1660
rect 5245 1640 5265 1660
rect 5915 1640 5935 1660
rect 6155 1640 6175 1660
rect 6395 1640 6415 1660
rect 3435 1575 3460 1600
rect 3435 1515 3460 1540
rect 4765 1520 4785 1540
rect 6395 1520 6415 1540
rect 4825 1470 4845 1490
rect 4945 1470 4965 1490
rect 5065 1470 5085 1490
rect 5185 1470 5205 1490
rect 5305 1470 5325 1490
rect 5855 1470 5875 1490
rect 5975 1470 5995 1490
rect 6095 1470 6115 1490
rect 6215 1470 6235 1490
rect 6335 1470 6355 1490
rect 2350 1335 2375 1360
rect 4435 1415 4455 1435
rect 5515 1415 5535 1435
rect 5645 1415 5665 1435
rect 6725 1415 6745 1435
rect 2350 1275 2375 1300
rect 4540 1090 4560 1110
rect 4620 1090 4640 1110
rect 4700 1090 4720 1110
rect 4780 1090 4800 1110
rect 4860 1090 4880 1110
rect 4940 1090 4960 1110
rect 5020 1090 5040 1110
rect 5100 1090 5120 1110
rect 5180 1090 5200 1110
rect 5260 1090 5280 1110
rect 5340 1090 5360 1110
rect 5420 1090 5440 1110
rect 5500 1090 5520 1110
rect 5580 1090 5600 1110
rect 5660 1090 5680 1110
rect 5740 1090 5760 1110
rect 5820 1090 5840 1110
rect 5900 1090 5920 1110
rect 5980 1090 6000 1110
rect 6060 1090 6080 1110
rect 6140 1090 6160 1110
rect 6220 1090 6240 1110
rect 6300 1090 6320 1110
rect 6380 1090 6400 1110
rect 6460 1090 6480 1110
rect 6540 1090 6560 1110
rect 2355 1000 2380 1025
rect 3070 1000 3095 1025
rect 4500 1005 4520 1025
rect 2470 940 2495 965
rect 2470 880 2495 905
rect 2470 800 2495 825
rect 2470 740 2495 765
rect -830 -430 -805 -405
rect -830 -490 -805 -465
rect -830 -550 -805 -525
rect -970 -970 -945 -945
rect -830 -970 -805 -945
rect -11 -970 14 -945
rect -830 -1390 -805 -1365
rect -830 -1450 -805 -1425
rect -830 -1510 -805 -1485
<< metal1 >>
rect 3730 4360 3750 4675
rect 4545 3075 4585 3080
rect 4545 3045 4550 3075
rect 4580 3045 4585 3075
rect 4545 3040 4585 3045
rect 7035 3075 7075 3080
rect 7035 3045 7040 3075
rect 7070 3045 7075 3075
rect 7035 3040 7075 3045
rect 4555 2945 4575 3040
rect 4545 2935 4585 2945
rect 4545 2915 4555 2935
rect 4575 2915 4585 2935
rect 4545 2905 4585 2915
rect 4580 2750 4620 2755
rect 4580 2720 4585 2750
rect 4615 2720 4620 2750
rect 4580 2715 4620 2720
rect 4760 2750 4800 2755
rect 4760 2720 4765 2750
rect 4795 2720 4800 2750
rect 4760 2715 4800 2720
rect 4940 2750 4980 2755
rect 4940 2720 4945 2750
rect 4975 2720 4980 2750
rect 4940 2715 4980 2720
rect 5120 2750 5160 2755
rect 5120 2720 5125 2750
rect 5155 2720 5160 2750
rect 5120 2715 5160 2720
rect 5300 2750 5340 2755
rect 5300 2720 5305 2750
rect 5335 2720 5340 2750
rect 5300 2715 5340 2720
rect 5480 2750 5520 2755
rect 5480 2720 5485 2750
rect 5515 2720 5520 2750
rect 5480 2715 5520 2720
rect 5660 2750 5700 2755
rect 5660 2720 5665 2750
rect 5695 2720 5700 2750
rect 5660 2715 5700 2720
rect 5840 2750 5880 2755
rect 5840 2720 5845 2750
rect 5875 2720 5880 2750
rect 5840 2715 5880 2720
rect 6020 2750 6060 2755
rect 6020 2720 6025 2750
rect 6055 2720 6060 2750
rect 6020 2715 6060 2720
rect 6200 2750 6240 2755
rect 6200 2720 6205 2750
rect 6235 2720 6240 2750
rect 6200 2715 6240 2720
rect 6380 2750 6420 2755
rect 6380 2720 6385 2750
rect 6415 2720 6420 2750
rect 6380 2715 6420 2720
rect 6560 2750 6600 2755
rect 6560 2720 6565 2750
rect 6595 2720 6600 2750
rect 6560 2715 6600 2720
rect 275 2200 1985 2550
rect 4490 2375 4530 2385
rect 4670 2380 4710 2385
rect 4490 2355 4500 2375
rect 4520 2355 4530 2375
rect 4210 2345 4250 2350
rect 4490 2345 4530 2355
rect 4580 2375 4620 2380
rect 4580 2345 4585 2375
rect 4615 2345 4620 2375
rect 4670 2350 4675 2380
rect 4705 2350 4710 2380
rect 4670 2345 4710 2350
rect 5030 2375 5070 2385
rect 5030 2355 5040 2375
rect 5060 2355 5070 2375
rect 5030 2345 5070 2355
rect 5335 2375 5375 2385
rect 5335 2355 5345 2375
rect 5365 2355 5375 2375
rect 5335 2345 5375 2355
rect 5400 2380 5440 2385
rect 5400 2350 5405 2380
rect 5435 2350 5440 2380
rect 5400 2345 5440 2350
rect 5570 2375 5610 2385
rect 5570 2355 5580 2375
rect 5600 2355 5610 2375
rect 5570 2345 5610 2355
rect 5740 2380 5780 2385
rect 5740 2350 5745 2380
rect 5775 2350 5780 2380
rect 5740 2345 5780 2350
rect 6110 2375 6150 2385
rect 6110 2355 6120 2375
rect 6140 2355 6150 2375
rect 6110 2345 6150 2355
rect 6470 2380 6510 2385
rect 6470 2350 6475 2380
rect 6505 2350 6510 2380
rect 6470 2345 6510 2350
rect 6650 2375 6690 2385
rect 6650 2355 6660 2375
rect 6680 2355 6690 2375
rect 6650 2345 6690 2355
rect 4210 2315 4215 2345
rect 4245 2315 4250 2345
rect 4210 2310 4250 2315
rect 3830 2290 3870 2295
rect 3830 2260 3835 2290
rect 3865 2260 3870 2290
rect 3830 2255 3870 2260
rect -110 1720 -70 1725
rect -110 1690 -105 1720
rect -75 1715 -70 1720
rect -45 1720 -5 1725
rect -45 1715 -40 1720
rect -75 1695 -40 1715
rect -75 1690 -70 1695
rect -110 1685 -70 1690
rect -45 1690 -40 1695
rect -10 1690 -5 1720
rect -45 1685 -5 1690
rect 275 1190 625 2200
rect 955 1710 1305 1870
rect 955 1680 1270 1710
rect 1300 1680 1305 1710
rect 955 1520 1305 1680
rect 1635 1190 1985 2200
rect 3585 1710 3625 1715
rect 3585 1680 3590 1710
rect 3620 1680 3625 1710
rect 3585 1675 3625 1680
rect 3595 1610 3615 1675
rect 3585 1605 3625 1610
rect 3425 1570 3430 1605
rect 3465 1570 3470 1605
rect 3585 1575 3590 1605
rect 3620 1575 3625 1605
rect 3585 1570 3625 1575
rect 3585 1545 3625 1550
rect 3425 1510 3430 1545
rect 3465 1510 3470 1545
rect 3585 1515 3590 1545
rect 3620 1515 3625 1545
rect 3585 1510 3625 1515
rect 2340 1330 2345 1365
rect 2380 1330 2385 1365
rect 2340 1305 2385 1310
rect 2340 1270 2345 1305
rect 2380 1270 2385 1305
rect 2340 1265 2385 1270
rect 275 1035 2175 1190
rect 3595 1035 3615 1510
rect 275 1030 2215 1035
rect 3585 1030 3625 1035
rect 275 1000 2180 1030
rect 2210 1000 2215 1030
rect 275 995 2215 1000
rect 2345 995 2350 1030
rect 2385 995 2390 1030
rect 3060 995 3065 1030
rect 3100 995 3105 1030
rect 3585 1000 3590 1030
rect 3620 1000 3625 1030
rect 3585 995 3625 1000
rect 275 840 2175 995
rect 2320 970 2360 975
rect 2320 940 2325 970
rect 2355 940 2360 970
rect 2320 935 2360 940
rect 2460 935 2465 970
rect 2500 935 2505 970
rect 2330 835 2350 935
rect 2460 875 2465 910
rect 2500 875 2505 910
rect 3840 875 3860 2255
rect 4055 2195 4095 2200
rect 4055 2165 4060 2195
rect 4090 2165 4095 2195
rect 4055 2160 4095 2165
rect 4005 2145 4045 2150
rect 4005 2115 4010 2145
rect 4040 2115 4045 2145
rect 4005 2110 4045 2115
rect 4015 1835 4035 2110
rect 4005 1830 4045 1835
rect 4005 1800 4010 1830
rect 4040 1800 4045 1830
rect 4005 1795 4045 1800
rect 4015 1035 4035 1795
rect 4065 1550 4085 2160
rect 4100 2100 4140 2105
rect 4100 2070 4105 2100
rect 4135 2070 4140 2100
rect 4100 2065 4140 2070
rect 4110 1715 4130 2065
rect 4220 2005 4240 2310
rect 4500 2150 4520 2345
rect 4580 2340 4620 2345
rect 4680 2200 4700 2345
rect 4850 2335 4890 2340
rect 4850 2305 4855 2335
rect 4885 2305 4890 2335
rect 4850 2300 4890 2305
rect 4670 2195 4710 2200
rect 4670 2165 4675 2195
rect 4705 2165 4710 2195
rect 4670 2160 4710 2165
rect 4490 2145 4530 2150
rect 4490 2115 4495 2145
rect 4525 2115 4530 2145
rect 4490 2110 4530 2115
rect 4860 2105 4880 2300
rect 5040 2295 5060 2345
rect 5210 2335 5250 2340
rect 5210 2305 5215 2335
rect 5245 2305 5250 2335
rect 5210 2300 5250 2305
rect 5030 2290 5070 2295
rect 5030 2260 5035 2290
rect 5065 2260 5070 2290
rect 5030 2255 5070 2260
rect 4850 2100 4890 2105
rect 4850 2070 4855 2100
rect 4885 2070 4890 2100
rect 4850 2065 4890 2070
rect 4455 2045 4495 2050
rect 4455 2015 4460 2045
rect 4490 2015 4495 2045
rect 4455 2010 4495 2015
rect 4575 2045 4615 2050
rect 4575 2015 4580 2045
rect 4610 2015 4615 2045
rect 4575 2010 4615 2015
rect 4695 2045 4735 2050
rect 4695 2015 4700 2045
rect 4730 2015 4735 2045
rect 4695 2010 4735 2015
rect 4815 2045 4855 2050
rect 4815 2015 4820 2045
rect 4850 2015 4855 2045
rect 4815 2010 4855 2015
rect 4935 2045 4975 2050
rect 4935 2015 4940 2045
rect 4970 2015 4975 2045
rect 4935 2010 4975 2015
rect 5055 2045 5095 2050
rect 5055 2015 5060 2045
rect 5090 2015 5095 2045
rect 5055 2010 5095 2015
rect 5175 2045 5215 2050
rect 5175 2015 5180 2045
rect 5210 2015 5215 2045
rect 5175 2010 5215 2015
rect 5295 2045 5335 2050
rect 5295 2015 5300 2045
rect 5330 2015 5335 2045
rect 5295 2010 5335 2015
rect 5355 2005 5375 2345
rect 5580 2150 5600 2345
rect 5930 2335 5970 2340
rect 5930 2305 5935 2335
rect 5965 2305 5970 2335
rect 5930 2300 5970 2305
rect 6120 2295 6140 2345
rect 6290 2335 6330 2340
rect 6290 2305 6295 2335
rect 6325 2305 6330 2335
rect 6290 2300 6330 2305
rect 6110 2290 6150 2295
rect 6110 2260 6115 2290
rect 6145 2260 6150 2290
rect 6110 2255 6150 2260
rect 6660 2150 6680 2345
rect 6840 2290 6880 2295
rect 6840 2260 6845 2290
rect 6875 2260 6880 2290
rect 6840 2255 6880 2260
rect 5570 2145 5610 2150
rect 5570 2115 5575 2145
rect 5605 2115 5610 2145
rect 5570 2110 5610 2115
rect 6650 2145 6690 2150
rect 6650 2115 6655 2145
rect 6685 2115 6690 2145
rect 6650 2110 6690 2115
rect 5795 2095 5835 2100
rect 5795 2065 5800 2095
rect 5830 2065 5835 2095
rect 5795 2060 5835 2065
rect 5415 2045 5455 2050
rect 5415 2015 5420 2045
rect 5450 2015 5455 2045
rect 5415 2010 5455 2015
rect 5725 2045 5765 2050
rect 5725 2015 5730 2045
rect 5760 2015 5765 2045
rect 5725 2010 5765 2015
rect 5805 2005 5825 2060
rect 5845 2045 5885 2050
rect 5845 2015 5850 2045
rect 5880 2015 5885 2045
rect 5845 2010 5885 2015
rect 5965 2045 6005 2050
rect 5965 2015 5970 2045
rect 6000 2015 6005 2045
rect 5965 2010 6005 2015
rect 6085 2045 6125 2050
rect 6085 2015 6090 2045
rect 6120 2015 6125 2045
rect 6085 2010 6125 2015
rect 6205 2045 6245 2050
rect 6205 2015 6210 2045
rect 6240 2015 6245 2045
rect 6205 2010 6245 2015
rect 6325 2045 6365 2050
rect 6325 2015 6330 2045
rect 6360 2015 6365 2045
rect 6325 2010 6365 2015
rect 6445 2045 6485 2050
rect 6445 2015 6450 2045
rect 6480 2015 6485 2045
rect 6445 2010 6485 2015
rect 6565 2045 6605 2050
rect 6565 2015 6570 2045
rect 6600 2015 6605 2045
rect 6565 2010 6605 2015
rect 6685 2045 6725 2050
rect 6685 2015 6690 2045
rect 6720 2015 6725 2045
rect 6685 2010 6725 2015
rect 4210 2000 4250 2005
rect 4210 1970 4215 2000
rect 4245 1970 4250 2000
rect 4210 1965 4250 1970
rect 4395 2000 4435 2005
rect 4395 1970 4400 2000
rect 4430 1970 4435 2000
rect 4395 1965 4435 1970
rect 4755 2000 4795 2005
rect 4755 1970 4760 2000
rect 4790 1970 4795 2000
rect 4755 1965 4795 1970
rect 5115 2000 5155 2005
rect 5115 1970 5120 2000
rect 5150 1970 5155 2000
rect 5115 1965 5155 1970
rect 5355 1995 5395 2005
rect 5355 1975 5365 1995
rect 5385 1975 5395 1995
rect 5355 1965 5395 1975
rect 5475 2000 5535 2005
rect 5475 1970 5480 2000
rect 5510 1970 5535 2000
rect 5475 1965 5535 1970
rect 4155 1825 4190 1835
rect 4155 1805 4165 1825
rect 4185 1805 4190 1825
rect 4155 1795 4190 1805
rect 4210 1830 4250 1835
rect 4210 1800 4215 1830
rect 4245 1800 4250 1830
rect 4210 1795 4250 1800
rect 4270 1825 4305 1835
rect 4270 1805 4275 1825
rect 4295 1805 4305 1825
rect 4270 1795 4305 1805
rect 4425 1825 4465 1835
rect 4425 1805 4435 1825
rect 4455 1805 4465 1825
rect 4425 1795 4465 1805
rect 4515 1830 4555 1835
rect 4515 1800 4520 1830
rect 4550 1800 4555 1830
rect 4515 1795 4555 1800
rect 4635 1825 4675 1835
rect 4635 1805 4645 1825
rect 4665 1805 4675 1825
rect 4635 1795 4675 1805
rect 4755 1825 4795 1835
rect 4755 1805 4765 1825
rect 4785 1805 4795 1825
rect 4755 1795 4795 1805
rect 4875 1830 4915 1835
rect 4875 1800 4880 1830
rect 4910 1800 4915 1830
rect 4875 1795 4915 1800
rect 4995 1825 5035 1835
rect 4995 1805 5005 1825
rect 5025 1805 5035 1825
rect 4995 1795 5035 1805
rect 5115 1825 5155 1835
rect 5115 1805 5125 1825
rect 5145 1805 5155 1825
rect 5115 1795 5155 1805
rect 5235 1830 5275 1835
rect 5235 1800 5240 1830
rect 5270 1800 5275 1830
rect 5235 1795 5275 1800
rect 5355 1825 5395 1835
rect 5355 1805 5365 1825
rect 5385 1805 5395 1825
rect 5355 1795 5395 1805
rect 5445 1825 5485 1835
rect 5445 1805 5455 1825
rect 5475 1805 5485 1825
rect 5445 1795 5485 1805
rect 4165 1715 4185 1795
rect 4275 1715 4295 1795
rect 4435 1775 4455 1795
rect 4645 1775 4665 1795
rect 4765 1775 4785 1795
rect 4425 1770 4465 1775
rect 4425 1740 4430 1770
rect 4460 1740 4465 1770
rect 4425 1735 4465 1740
rect 4635 1770 4675 1775
rect 4635 1740 4640 1770
rect 4670 1740 4675 1770
rect 4635 1735 4675 1740
rect 4755 1770 4795 1775
rect 4755 1740 4760 1770
rect 4790 1740 4795 1770
rect 4755 1735 4795 1740
rect 4885 1715 4905 1795
rect 5005 1775 5025 1795
rect 5125 1775 5145 1795
rect 5365 1775 5385 1795
rect 5455 1775 5475 1795
rect 4995 1770 5035 1775
rect 4995 1740 5000 1770
rect 5030 1740 5035 1770
rect 4995 1735 5035 1740
rect 5115 1770 5155 1775
rect 5115 1740 5120 1770
rect 5150 1740 5155 1770
rect 5115 1735 5155 1740
rect 5355 1770 5395 1775
rect 5355 1740 5360 1770
rect 5390 1740 5395 1770
rect 5355 1735 5395 1740
rect 5445 1770 5485 1775
rect 5445 1740 5450 1770
rect 5480 1740 5485 1770
rect 5445 1735 5485 1740
rect 4100 1710 4140 1715
rect 4100 1680 4105 1710
rect 4135 1680 4140 1710
rect 4100 1675 4140 1680
rect 4155 1710 4195 1715
rect 4155 1680 4160 1710
rect 4190 1680 4195 1710
rect 4155 1675 4195 1680
rect 4265 1710 4305 1715
rect 4265 1680 4270 1710
rect 4300 1680 4305 1710
rect 4265 1675 4305 1680
rect 4815 1710 4855 1715
rect 4815 1680 4820 1710
rect 4850 1680 4855 1710
rect 4815 1675 4855 1680
rect 4875 1710 4915 1715
rect 4875 1680 4880 1710
rect 4910 1680 4915 1710
rect 4875 1675 4915 1680
rect 5005 1670 5025 1735
rect 5115 1710 5155 1715
rect 5115 1680 5120 1710
rect 5150 1680 5155 1710
rect 5115 1675 5155 1680
rect 5355 1710 5395 1715
rect 5355 1680 5360 1710
rect 5390 1680 5395 1710
rect 5355 1675 5395 1680
rect 4755 1665 4795 1670
rect 4755 1635 4760 1665
rect 4790 1635 4795 1665
rect 4755 1630 4795 1635
rect 4995 1665 5035 1670
rect 4995 1635 5000 1665
rect 5030 1635 5035 1665
rect 4995 1630 5035 1635
rect 5235 1665 5275 1670
rect 5235 1635 5240 1665
rect 5270 1635 5275 1665
rect 5235 1630 5275 1635
rect 4055 1545 4095 1550
rect 4055 1515 4060 1545
rect 4090 1515 4095 1545
rect 4055 1510 4095 1515
rect 4755 1545 4795 1550
rect 4755 1515 4760 1545
rect 4790 1515 4795 1545
rect 4755 1510 4795 1515
rect 4425 1495 4465 1500
rect 4425 1465 4430 1495
rect 4460 1465 4465 1495
rect 4425 1460 4465 1465
rect 4815 1495 4855 1500
rect 4815 1465 4820 1495
rect 4850 1465 4855 1495
rect 4815 1460 4855 1465
rect 4935 1495 4975 1500
rect 4935 1465 4940 1495
rect 4970 1465 4975 1495
rect 4935 1460 4975 1465
rect 5055 1495 5095 1500
rect 5055 1465 5060 1495
rect 5090 1465 5095 1495
rect 5055 1460 5095 1465
rect 5175 1495 5215 1500
rect 5175 1465 5180 1495
rect 5210 1465 5215 1495
rect 5175 1460 5215 1465
rect 5295 1495 5335 1500
rect 5295 1465 5300 1495
rect 5330 1465 5335 1495
rect 5295 1460 5335 1465
rect 4435 1445 4455 1460
rect 5515 1445 5535 1965
rect 5645 2000 5705 2005
rect 5645 1970 5670 2000
rect 5700 1970 5705 2000
rect 5645 1965 5705 1970
rect 5785 1995 5825 2005
rect 5785 1975 5795 1995
rect 5815 1975 5825 1995
rect 5785 1965 5825 1975
rect 6025 2000 6065 2005
rect 6025 1970 6030 2000
rect 6060 1970 6065 2000
rect 6025 1965 6065 1970
rect 6385 2000 6425 2005
rect 6385 1970 6390 2000
rect 6420 1970 6425 2000
rect 6385 1965 6425 1970
rect 6745 2000 6785 2005
rect 6745 1970 6750 2000
rect 6780 1970 6785 2000
rect 6745 1965 6785 1970
rect 5645 1445 5665 1965
rect 5695 1825 5735 1835
rect 5695 1805 5705 1825
rect 5725 1805 5735 1825
rect 5695 1795 5735 1805
rect 5785 1825 5825 1835
rect 5785 1805 5795 1825
rect 5815 1805 5825 1825
rect 5785 1795 5825 1805
rect 5905 1830 5945 1835
rect 5905 1800 5910 1830
rect 5940 1800 5945 1830
rect 5905 1795 5945 1800
rect 6025 1825 6065 1835
rect 6025 1805 6035 1825
rect 6055 1805 6065 1825
rect 6025 1795 6065 1805
rect 6145 1825 6185 1835
rect 6145 1805 6155 1825
rect 6175 1805 6185 1825
rect 6145 1795 6185 1805
rect 6265 1830 6305 1835
rect 6265 1800 6270 1830
rect 6300 1800 6305 1830
rect 6265 1795 6305 1800
rect 6385 1825 6425 1835
rect 6385 1805 6395 1825
rect 6415 1805 6425 1825
rect 6385 1795 6425 1805
rect 6505 1825 6545 1835
rect 6505 1805 6515 1825
rect 6535 1805 6545 1825
rect 6505 1795 6545 1805
rect 6625 1830 6665 1835
rect 6625 1800 6630 1830
rect 6660 1800 6665 1830
rect 6625 1795 6665 1800
rect 6715 1825 6755 1835
rect 6715 1805 6725 1825
rect 6745 1805 6755 1825
rect 6715 1795 6755 1805
rect 5705 1775 5725 1795
rect 5795 1775 5815 1795
rect 6035 1775 6055 1795
rect 6155 1775 6175 1795
rect 5695 1770 5735 1775
rect 5695 1740 5700 1770
rect 5730 1740 5735 1770
rect 5695 1735 5735 1740
rect 5785 1770 5825 1775
rect 5785 1740 5790 1770
rect 5820 1740 5825 1770
rect 5785 1735 5825 1740
rect 6025 1770 6065 1775
rect 6025 1740 6030 1770
rect 6060 1740 6065 1770
rect 6025 1735 6065 1740
rect 6145 1770 6185 1775
rect 6145 1740 6150 1770
rect 6180 1740 6185 1770
rect 6145 1735 6185 1740
rect 5785 1710 5825 1715
rect 5785 1680 5790 1710
rect 5820 1680 5825 1710
rect 5785 1675 5825 1680
rect 6025 1710 6065 1715
rect 6025 1680 6030 1710
rect 6060 1680 6065 1710
rect 6025 1675 6065 1680
rect 6155 1670 6175 1735
rect 6275 1715 6295 1795
rect 6395 1775 6415 1795
rect 6515 1775 6535 1795
rect 6725 1775 6745 1795
rect 6385 1770 6425 1775
rect 6385 1740 6390 1770
rect 6420 1740 6425 1770
rect 6385 1735 6425 1740
rect 6505 1770 6545 1775
rect 6505 1740 6510 1770
rect 6540 1740 6545 1770
rect 6505 1735 6545 1740
rect 6715 1770 6755 1775
rect 6715 1740 6720 1770
rect 6750 1740 6755 1770
rect 6715 1735 6755 1740
rect 6850 1715 6870 2255
rect 7045 2100 7065 3040
rect 7035 2095 7075 2100
rect 7035 2065 7040 2095
rect 7070 2065 7075 2095
rect 7035 2060 7075 2065
rect 6265 1710 6305 1715
rect 6265 1680 6270 1710
rect 6300 1680 6305 1710
rect 6265 1675 6305 1680
rect 6325 1710 6365 1715
rect 6325 1680 6330 1710
rect 6360 1680 6365 1710
rect 6325 1675 6365 1680
rect 6840 1710 6880 1715
rect 6840 1680 6845 1710
rect 6875 1680 6880 1710
rect 6840 1675 6880 1680
rect 5905 1665 5945 1670
rect 5905 1635 5910 1665
rect 5940 1635 5945 1665
rect 5905 1630 5945 1635
rect 6145 1665 6185 1670
rect 6145 1635 6150 1665
rect 6180 1635 6185 1665
rect 6145 1630 6185 1635
rect 6385 1665 6425 1670
rect 6385 1635 6390 1665
rect 6420 1635 6425 1665
rect 6385 1630 6425 1635
rect 6385 1545 6425 1550
rect 6385 1515 6390 1545
rect 6420 1515 6425 1545
rect 6385 1510 6425 1515
rect 6840 1545 6880 1550
rect 6840 1515 6845 1545
rect 6875 1515 6880 1545
rect 6840 1510 6880 1515
rect 5845 1495 5885 1500
rect 5845 1465 5850 1495
rect 5880 1465 5885 1495
rect 5845 1460 5885 1465
rect 5965 1495 6005 1500
rect 5965 1465 5970 1495
rect 6000 1465 6005 1495
rect 5965 1460 6005 1465
rect 6085 1495 6125 1500
rect 6085 1465 6090 1495
rect 6120 1465 6125 1495
rect 6085 1460 6125 1465
rect 6205 1495 6245 1500
rect 6205 1465 6210 1495
rect 6240 1465 6245 1495
rect 6205 1460 6245 1465
rect 6325 1495 6365 1500
rect 6325 1465 6330 1495
rect 6360 1465 6365 1495
rect 6325 1460 6365 1465
rect 6715 1495 6755 1500
rect 6715 1465 6720 1495
rect 6750 1465 6755 1495
rect 6715 1460 6755 1465
rect 6725 1445 6745 1460
rect 4425 1435 4465 1445
rect 4425 1415 4435 1435
rect 4455 1415 4465 1435
rect 4425 1405 4465 1415
rect 5505 1435 5545 1445
rect 5505 1415 5515 1435
rect 5535 1415 5545 1435
rect 5505 1405 5545 1415
rect 5635 1435 5675 1445
rect 5635 1415 5645 1435
rect 5665 1415 5675 1435
rect 5635 1405 5675 1415
rect 6715 1435 6755 1445
rect 6715 1415 6725 1435
rect 6745 1415 6755 1435
rect 6715 1405 6755 1415
rect 4530 1115 4570 1120
rect 4530 1085 4535 1115
rect 4565 1085 4570 1115
rect 4530 1080 4570 1085
rect 4610 1115 4650 1120
rect 4610 1085 4615 1115
rect 4645 1085 4650 1115
rect 4610 1080 4650 1085
rect 4690 1115 4730 1120
rect 4690 1085 4695 1115
rect 4725 1085 4730 1115
rect 4690 1080 4730 1085
rect 4770 1115 4810 1120
rect 4770 1085 4775 1115
rect 4805 1085 4810 1115
rect 4770 1080 4810 1085
rect 4850 1115 4890 1120
rect 4850 1085 4855 1115
rect 4885 1085 4890 1115
rect 4850 1080 4890 1085
rect 4930 1115 4970 1120
rect 4930 1085 4935 1115
rect 4965 1085 4970 1115
rect 4930 1080 4970 1085
rect 5010 1115 5050 1120
rect 5010 1085 5015 1115
rect 5045 1085 5050 1115
rect 5010 1080 5050 1085
rect 5090 1115 5130 1120
rect 5090 1085 5095 1115
rect 5125 1085 5130 1115
rect 5090 1080 5130 1085
rect 5170 1115 5210 1120
rect 5170 1085 5175 1115
rect 5205 1085 5210 1115
rect 5170 1080 5210 1085
rect 5250 1115 5290 1120
rect 5250 1085 5255 1115
rect 5285 1085 5290 1115
rect 5250 1080 5290 1085
rect 5330 1115 5370 1120
rect 5330 1085 5335 1115
rect 5365 1085 5370 1115
rect 5330 1080 5370 1085
rect 5410 1115 5450 1120
rect 5410 1085 5415 1115
rect 5445 1085 5450 1115
rect 5410 1080 5450 1085
rect 5490 1115 5530 1120
rect 5490 1085 5495 1115
rect 5525 1085 5530 1115
rect 5490 1080 5530 1085
rect 5570 1115 5610 1120
rect 5570 1085 5575 1115
rect 5605 1085 5610 1115
rect 5570 1080 5610 1085
rect 5650 1115 5690 1120
rect 5650 1085 5655 1115
rect 5685 1085 5690 1115
rect 5650 1080 5690 1085
rect 5730 1115 5770 1120
rect 5730 1085 5735 1115
rect 5765 1085 5770 1115
rect 5730 1080 5770 1085
rect 5810 1115 5850 1120
rect 5810 1085 5815 1115
rect 5845 1085 5850 1115
rect 5810 1080 5850 1085
rect 5890 1115 5930 1120
rect 5890 1085 5895 1115
rect 5925 1085 5930 1115
rect 5890 1080 5930 1085
rect 5970 1115 6010 1120
rect 5970 1085 5975 1115
rect 6005 1085 6010 1115
rect 5970 1080 6010 1085
rect 6050 1115 6090 1120
rect 6050 1085 6055 1115
rect 6085 1085 6090 1115
rect 6050 1080 6090 1085
rect 6130 1115 6170 1120
rect 6130 1085 6135 1115
rect 6165 1085 6170 1115
rect 6130 1080 6170 1085
rect 6210 1115 6250 1120
rect 6210 1085 6215 1115
rect 6245 1085 6250 1115
rect 6210 1080 6250 1085
rect 6290 1115 6330 1120
rect 6290 1085 6295 1115
rect 6325 1085 6330 1115
rect 6290 1080 6330 1085
rect 6370 1115 6410 1120
rect 6370 1085 6375 1115
rect 6405 1085 6410 1115
rect 6370 1080 6410 1085
rect 6450 1115 6490 1120
rect 6450 1085 6455 1115
rect 6485 1085 6490 1115
rect 6450 1080 6490 1085
rect 6530 1115 6570 1120
rect 6530 1085 6535 1115
rect 6565 1085 6570 1115
rect 6530 1080 6570 1085
rect 4005 1030 4045 1035
rect 4005 1000 4010 1030
rect 4040 1000 4045 1030
rect 4005 995 4045 1000
rect 4490 1030 4530 1035
rect 4490 1000 4495 1030
rect 4525 1000 4530 1030
rect 4490 995 4530 1000
rect 3830 870 3870 875
rect 3830 840 3835 870
rect 3865 840 3870 870
rect 3830 835 3870 840
rect 2320 830 2360 835
rect 2320 800 2325 830
rect 2355 800 2360 830
rect 2320 795 2360 800
rect 2460 795 2465 830
rect 2500 795 2505 830
rect 2330 650 2350 795
rect 2460 735 2465 770
rect 2500 735 2505 770
rect 6850 735 6870 1510
rect 6840 730 6880 735
rect 6840 700 6845 730
rect 6875 700 6880 730
rect 6840 695 6880 700
rect 3115 640 3135 645
rect 3100 630 3150 640
rect 3100 600 3110 630
rect 3140 600 3150 630
rect 3100 590 3150 600
rect -930 -520 -910 -395
rect -880 -460 -860 -395
rect -830 -400 -810 -395
rect -840 -435 -835 -400
rect -800 -435 -795 -400
rect -890 -465 -855 -460
rect -890 -495 -885 -465
rect -840 -495 -835 -460
rect -800 -495 -795 -460
rect -890 -500 -855 -495
rect -940 -525 -900 -520
rect -940 -555 -935 -525
rect -905 -555 -900 -525
rect -840 -555 -835 -520
rect -800 -555 -795 -520
rect -940 -560 -900 -555
rect -940 -975 -935 -940
rect -840 -975 -835 -940
rect -800 -975 -795 -940
rect -21 -975 -16 -940
rect 19 -975 24 -940
rect -950 -1365 -910 -1360
rect -950 -1395 -945 -1365
rect -915 -1395 -910 -1365
rect -840 -1395 -835 -1360
rect -800 -1395 -795 -1360
rect -950 -1400 -910 -1395
rect -940 -1600 -920 -1400
rect -895 -1425 -855 -1420
rect -895 -1455 -890 -1425
rect -860 -1455 -855 -1425
rect -840 -1455 -835 -1420
rect -800 -1455 -795 -1420
rect -895 -1460 -855 -1455
rect -885 -1555 -865 -1460
rect -840 -1480 -795 -1475
rect -840 -1515 -835 -1480
rect -800 -1515 -795 -1480
rect -840 -1520 -795 -1515
rect -895 -1560 -855 -1555
rect -895 -1590 -890 -1560
rect -860 -1590 -855 -1560
rect -895 -1595 -855 -1590
<< via1 >>
rect 4550 3045 4580 3075
rect 7040 3045 7070 3075
rect 4585 2745 4615 2750
rect 4585 2725 4590 2745
rect 4590 2725 4610 2745
rect 4610 2725 4615 2745
rect 4585 2720 4615 2725
rect 4765 2745 4795 2750
rect 4765 2725 4770 2745
rect 4770 2725 4790 2745
rect 4790 2725 4795 2745
rect 4765 2720 4795 2725
rect 4945 2745 4975 2750
rect 4945 2725 4950 2745
rect 4950 2725 4970 2745
rect 4970 2725 4975 2745
rect 4945 2720 4975 2725
rect 5125 2745 5155 2750
rect 5125 2725 5130 2745
rect 5130 2725 5150 2745
rect 5150 2725 5155 2745
rect 5125 2720 5155 2725
rect 5305 2745 5335 2750
rect 5305 2725 5310 2745
rect 5310 2725 5330 2745
rect 5330 2725 5335 2745
rect 5305 2720 5335 2725
rect 5485 2745 5515 2750
rect 5485 2725 5490 2745
rect 5490 2725 5510 2745
rect 5510 2725 5515 2745
rect 5485 2720 5515 2725
rect 5665 2745 5695 2750
rect 5665 2725 5670 2745
rect 5670 2725 5690 2745
rect 5690 2725 5695 2745
rect 5665 2720 5695 2725
rect 5845 2745 5875 2750
rect 5845 2725 5850 2745
rect 5850 2725 5870 2745
rect 5870 2725 5875 2745
rect 5845 2720 5875 2725
rect 6025 2745 6055 2750
rect 6025 2725 6030 2745
rect 6030 2725 6050 2745
rect 6050 2725 6055 2745
rect 6025 2720 6055 2725
rect 6205 2745 6235 2750
rect 6205 2725 6210 2745
rect 6210 2725 6230 2745
rect 6230 2725 6235 2745
rect 6205 2720 6235 2725
rect 6385 2745 6415 2750
rect 6385 2725 6390 2745
rect 6390 2725 6410 2745
rect 6410 2725 6415 2745
rect 6385 2720 6415 2725
rect 6565 2745 6595 2750
rect 6565 2725 6570 2745
rect 6570 2725 6590 2745
rect 6590 2725 6595 2745
rect 6565 2720 6595 2725
rect 4585 2370 4615 2375
rect 4585 2350 4590 2370
rect 4590 2350 4610 2370
rect 4610 2350 4615 2370
rect 4585 2345 4615 2350
rect 4675 2375 4705 2380
rect 4675 2355 4680 2375
rect 4680 2355 4700 2375
rect 4700 2355 4705 2375
rect 4675 2350 4705 2355
rect 5405 2375 5435 2380
rect 5405 2355 5410 2375
rect 5410 2355 5430 2375
rect 5430 2355 5435 2375
rect 5405 2350 5435 2355
rect 5745 2375 5775 2380
rect 5745 2355 5750 2375
rect 5750 2355 5770 2375
rect 5770 2355 5775 2375
rect 5745 2350 5775 2355
rect 6475 2375 6505 2380
rect 6475 2355 6480 2375
rect 6480 2355 6500 2375
rect 6500 2355 6505 2375
rect 6475 2350 6505 2355
rect 4215 2315 4245 2345
rect 3835 2260 3865 2290
rect -105 1690 -75 1720
rect -40 1715 -10 1720
rect -40 1695 -35 1715
rect -35 1695 -15 1715
rect -15 1695 -10 1715
rect -40 1690 -10 1695
rect 1270 1680 1300 1710
rect 3590 1680 3620 1710
rect 3430 1600 3465 1605
rect 3430 1575 3435 1600
rect 3435 1575 3460 1600
rect 3460 1575 3465 1600
rect 3430 1570 3465 1575
rect 3590 1575 3620 1605
rect 3430 1540 3465 1545
rect 3430 1515 3435 1540
rect 3435 1515 3460 1540
rect 3460 1515 3465 1540
rect 3430 1510 3465 1515
rect 3590 1515 3620 1545
rect 2345 1360 2380 1365
rect 2345 1335 2350 1360
rect 2350 1335 2375 1360
rect 2375 1335 2380 1360
rect 2345 1330 2380 1335
rect 2345 1300 2380 1305
rect 2345 1275 2350 1300
rect 2350 1275 2375 1300
rect 2375 1275 2380 1300
rect 2345 1270 2380 1275
rect 2180 1000 2210 1030
rect 2350 1025 2385 1030
rect 2350 1000 2355 1025
rect 2355 1000 2380 1025
rect 2380 1000 2385 1025
rect 2350 995 2385 1000
rect 3065 1025 3100 1030
rect 3065 1000 3070 1025
rect 3070 1000 3095 1025
rect 3095 1000 3100 1025
rect 3065 995 3100 1000
rect 3590 1000 3620 1030
rect 2325 940 2355 970
rect 2465 965 2500 970
rect 2465 940 2470 965
rect 2470 940 2495 965
rect 2495 940 2500 965
rect 2465 935 2500 940
rect 2465 905 2500 910
rect 2465 880 2470 905
rect 2470 880 2495 905
rect 2495 880 2500 905
rect 2465 875 2500 880
rect 4060 2165 4090 2195
rect 4010 2115 4040 2145
rect 4010 1800 4040 1830
rect 4105 2070 4135 2100
rect 4855 2330 4885 2335
rect 4855 2310 4860 2330
rect 4860 2310 4880 2330
rect 4880 2310 4885 2330
rect 4855 2305 4885 2310
rect 4675 2165 4705 2195
rect 4495 2115 4525 2145
rect 5215 2330 5245 2335
rect 5215 2310 5220 2330
rect 5220 2310 5240 2330
rect 5240 2310 5245 2330
rect 5215 2305 5245 2310
rect 5035 2285 5065 2290
rect 5035 2265 5040 2285
rect 5040 2265 5060 2285
rect 5060 2265 5065 2285
rect 5035 2260 5065 2265
rect 4855 2070 4885 2100
rect 4460 2040 4490 2045
rect 4460 2020 4465 2040
rect 4465 2020 4485 2040
rect 4485 2020 4490 2040
rect 4460 2015 4490 2020
rect 4580 2040 4610 2045
rect 4580 2020 4585 2040
rect 4585 2020 4605 2040
rect 4605 2020 4610 2040
rect 4580 2015 4610 2020
rect 4700 2040 4730 2045
rect 4700 2020 4705 2040
rect 4705 2020 4725 2040
rect 4725 2020 4730 2040
rect 4700 2015 4730 2020
rect 4820 2040 4850 2045
rect 4820 2020 4825 2040
rect 4825 2020 4845 2040
rect 4845 2020 4850 2040
rect 4820 2015 4850 2020
rect 4940 2040 4970 2045
rect 4940 2020 4945 2040
rect 4945 2020 4965 2040
rect 4965 2020 4970 2040
rect 4940 2015 4970 2020
rect 5060 2040 5090 2045
rect 5060 2020 5065 2040
rect 5065 2020 5085 2040
rect 5085 2020 5090 2040
rect 5060 2015 5090 2020
rect 5180 2040 5210 2045
rect 5180 2020 5185 2040
rect 5185 2020 5205 2040
rect 5205 2020 5210 2040
rect 5180 2015 5210 2020
rect 5300 2040 5330 2045
rect 5300 2020 5305 2040
rect 5305 2020 5325 2040
rect 5325 2020 5330 2040
rect 5300 2015 5330 2020
rect 5935 2330 5965 2335
rect 5935 2310 5940 2330
rect 5940 2310 5960 2330
rect 5960 2310 5965 2330
rect 5935 2305 5965 2310
rect 6295 2330 6325 2335
rect 6295 2310 6300 2330
rect 6300 2310 6320 2330
rect 6320 2310 6325 2330
rect 6295 2305 6325 2310
rect 6115 2285 6145 2290
rect 6115 2265 6120 2285
rect 6120 2265 6140 2285
rect 6140 2265 6145 2285
rect 6115 2260 6145 2265
rect 6845 2260 6875 2290
rect 5575 2115 5605 2145
rect 6655 2115 6685 2145
rect 5800 2065 5830 2095
rect 5420 2040 5450 2045
rect 5420 2020 5425 2040
rect 5425 2020 5445 2040
rect 5445 2020 5450 2040
rect 5420 2015 5450 2020
rect 5730 2040 5760 2045
rect 5730 2020 5735 2040
rect 5735 2020 5755 2040
rect 5755 2020 5760 2040
rect 5730 2015 5760 2020
rect 5850 2040 5880 2045
rect 5850 2020 5855 2040
rect 5855 2020 5875 2040
rect 5875 2020 5880 2040
rect 5850 2015 5880 2020
rect 5970 2040 6000 2045
rect 5970 2020 5975 2040
rect 5975 2020 5995 2040
rect 5995 2020 6000 2040
rect 5970 2015 6000 2020
rect 6090 2040 6120 2045
rect 6090 2020 6095 2040
rect 6095 2020 6115 2040
rect 6115 2020 6120 2040
rect 6090 2015 6120 2020
rect 6210 2040 6240 2045
rect 6210 2020 6215 2040
rect 6215 2020 6235 2040
rect 6235 2020 6240 2040
rect 6210 2015 6240 2020
rect 6330 2040 6360 2045
rect 6330 2020 6335 2040
rect 6335 2020 6355 2040
rect 6355 2020 6360 2040
rect 6330 2015 6360 2020
rect 6450 2040 6480 2045
rect 6450 2020 6455 2040
rect 6455 2020 6475 2040
rect 6475 2020 6480 2040
rect 6450 2015 6480 2020
rect 6570 2040 6600 2045
rect 6570 2020 6575 2040
rect 6575 2020 6595 2040
rect 6595 2020 6600 2040
rect 6570 2015 6600 2020
rect 6690 2040 6720 2045
rect 6690 2020 6695 2040
rect 6695 2020 6715 2040
rect 6715 2020 6720 2040
rect 6690 2015 6720 2020
rect 4215 1995 4245 2000
rect 4215 1975 4220 1995
rect 4220 1975 4240 1995
rect 4240 1975 4245 1995
rect 4215 1970 4245 1975
rect 4400 1995 4430 2000
rect 4400 1975 4405 1995
rect 4405 1975 4425 1995
rect 4425 1975 4430 1995
rect 4400 1970 4430 1975
rect 4760 1995 4790 2000
rect 4760 1975 4765 1995
rect 4765 1975 4785 1995
rect 4785 1975 4790 1995
rect 4760 1970 4790 1975
rect 5120 1995 5150 2000
rect 5120 1975 5125 1995
rect 5125 1975 5145 1995
rect 5145 1975 5150 1995
rect 5120 1970 5150 1975
rect 5480 1995 5510 2000
rect 5480 1975 5485 1995
rect 5485 1975 5505 1995
rect 5505 1975 5510 1995
rect 5480 1970 5510 1975
rect 4215 1825 4245 1830
rect 4215 1805 4220 1825
rect 4220 1805 4240 1825
rect 4240 1805 4245 1825
rect 4215 1800 4245 1805
rect 4520 1825 4550 1830
rect 4520 1805 4525 1825
rect 4525 1805 4545 1825
rect 4545 1805 4550 1825
rect 4520 1800 4550 1805
rect 4880 1825 4910 1830
rect 4880 1805 4885 1825
rect 4885 1805 4905 1825
rect 4905 1805 4910 1825
rect 4880 1800 4910 1805
rect 5240 1825 5270 1830
rect 5240 1805 5245 1825
rect 5245 1805 5265 1825
rect 5265 1805 5270 1825
rect 5240 1800 5270 1805
rect 4430 1740 4460 1770
rect 4640 1765 4670 1770
rect 4640 1745 4645 1765
rect 4645 1745 4665 1765
rect 4665 1745 4670 1765
rect 4640 1740 4670 1745
rect 4760 1740 4790 1770
rect 5000 1765 5030 1770
rect 5000 1745 5005 1765
rect 5005 1745 5025 1765
rect 5025 1745 5030 1765
rect 5000 1740 5030 1745
rect 5120 1740 5150 1770
rect 5360 1765 5390 1770
rect 5360 1745 5365 1765
rect 5365 1745 5385 1765
rect 5385 1745 5390 1765
rect 5360 1740 5390 1745
rect 5450 1740 5480 1770
rect 4105 1680 4135 1710
rect 4160 1680 4190 1710
rect 4270 1680 4300 1710
rect 4820 1705 4850 1710
rect 4820 1685 4825 1705
rect 4825 1685 4845 1705
rect 4845 1685 4850 1705
rect 4820 1680 4850 1685
rect 4880 1705 4910 1710
rect 4880 1685 4885 1705
rect 4885 1685 4905 1705
rect 4905 1685 4910 1705
rect 4880 1680 4910 1685
rect 5120 1705 5150 1710
rect 5120 1685 5125 1705
rect 5125 1685 5145 1705
rect 5145 1685 5150 1705
rect 5120 1680 5150 1685
rect 5360 1705 5390 1710
rect 5360 1685 5365 1705
rect 5365 1685 5385 1705
rect 5385 1685 5390 1705
rect 5360 1680 5390 1685
rect 4760 1660 4790 1665
rect 4760 1640 4765 1660
rect 4765 1640 4785 1660
rect 4785 1640 4790 1660
rect 4760 1635 4790 1640
rect 5000 1660 5030 1665
rect 5000 1640 5005 1660
rect 5005 1640 5025 1660
rect 5025 1640 5030 1660
rect 5000 1635 5030 1640
rect 5240 1660 5270 1665
rect 5240 1640 5245 1660
rect 5245 1640 5265 1660
rect 5265 1640 5270 1660
rect 5240 1635 5270 1640
rect 4060 1515 4090 1545
rect 4760 1540 4790 1545
rect 4760 1520 4765 1540
rect 4765 1520 4785 1540
rect 4785 1520 4790 1540
rect 4760 1515 4790 1520
rect 4430 1465 4460 1495
rect 4820 1490 4850 1495
rect 4820 1470 4825 1490
rect 4825 1470 4845 1490
rect 4845 1470 4850 1490
rect 4820 1465 4850 1470
rect 4940 1490 4970 1495
rect 4940 1470 4945 1490
rect 4945 1470 4965 1490
rect 4965 1470 4970 1490
rect 4940 1465 4970 1470
rect 5060 1490 5090 1495
rect 5060 1470 5065 1490
rect 5065 1470 5085 1490
rect 5085 1470 5090 1490
rect 5060 1465 5090 1470
rect 5180 1490 5210 1495
rect 5180 1470 5185 1490
rect 5185 1470 5205 1490
rect 5205 1470 5210 1490
rect 5180 1465 5210 1470
rect 5300 1490 5330 1495
rect 5300 1470 5305 1490
rect 5305 1470 5325 1490
rect 5325 1470 5330 1490
rect 5300 1465 5330 1470
rect 5670 1995 5700 2000
rect 5670 1975 5675 1995
rect 5675 1975 5695 1995
rect 5695 1975 5700 1995
rect 5670 1970 5700 1975
rect 6030 1995 6060 2000
rect 6030 1975 6035 1995
rect 6035 1975 6055 1995
rect 6055 1975 6060 1995
rect 6030 1970 6060 1975
rect 6390 1995 6420 2000
rect 6390 1975 6395 1995
rect 6395 1975 6415 1995
rect 6415 1975 6420 1995
rect 6390 1970 6420 1975
rect 6750 1995 6780 2000
rect 6750 1975 6755 1995
rect 6755 1975 6775 1995
rect 6775 1975 6780 1995
rect 6750 1970 6780 1975
rect 5910 1825 5940 1830
rect 5910 1805 5915 1825
rect 5915 1805 5935 1825
rect 5935 1805 5940 1825
rect 5910 1800 5940 1805
rect 6270 1825 6300 1830
rect 6270 1805 6275 1825
rect 6275 1805 6295 1825
rect 6295 1805 6300 1825
rect 6270 1800 6300 1805
rect 6630 1825 6660 1830
rect 6630 1805 6635 1825
rect 6635 1805 6655 1825
rect 6655 1805 6660 1825
rect 6630 1800 6660 1805
rect 5700 1740 5730 1770
rect 5790 1765 5820 1770
rect 5790 1745 5795 1765
rect 5795 1745 5815 1765
rect 5815 1745 5820 1765
rect 5790 1740 5820 1745
rect 6030 1740 6060 1770
rect 6150 1765 6180 1770
rect 6150 1745 6155 1765
rect 6155 1745 6175 1765
rect 6175 1745 6180 1765
rect 6150 1740 6180 1745
rect 5790 1705 5820 1710
rect 5790 1685 5795 1705
rect 5795 1685 5815 1705
rect 5815 1685 5820 1705
rect 5790 1680 5820 1685
rect 6030 1705 6060 1710
rect 6030 1685 6035 1705
rect 6035 1685 6055 1705
rect 6055 1685 6060 1705
rect 6030 1680 6060 1685
rect 6390 1740 6420 1770
rect 6510 1765 6540 1770
rect 6510 1745 6515 1765
rect 6515 1745 6535 1765
rect 6535 1745 6540 1765
rect 6510 1740 6540 1745
rect 6720 1740 6750 1770
rect 7040 2065 7070 2095
rect 6270 1705 6300 1710
rect 6270 1685 6275 1705
rect 6275 1685 6295 1705
rect 6295 1685 6300 1705
rect 6270 1680 6300 1685
rect 6330 1705 6360 1710
rect 6330 1685 6335 1705
rect 6335 1685 6355 1705
rect 6355 1685 6360 1705
rect 6330 1680 6360 1685
rect 6845 1680 6875 1710
rect 5910 1660 5940 1665
rect 5910 1640 5915 1660
rect 5915 1640 5935 1660
rect 5935 1640 5940 1660
rect 5910 1635 5940 1640
rect 6150 1660 6180 1665
rect 6150 1640 6155 1660
rect 6155 1640 6175 1660
rect 6175 1640 6180 1660
rect 6150 1635 6180 1640
rect 6390 1660 6420 1665
rect 6390 1640 6395 1660
rect 6395 1640 6415 1660
rect 6415 1640 6420 1660
rect 6390 1635 6420 1640
rect 6390 1540 6420 1545
rect 6390 1520 6395 1540
rect 6395 1520 6415 1540
rect 6415 1520 6420 1540
rect 6390 1515 6420 1520
rect 6845 1515 6875 1545
rect 5850 1490 5880 1495
rect 5850 1470 5855 1490
rect 5855 1470 5875 1490
rect 5875 1470 5880 1490
rect 5850 1465 5880 1470
rect 5970 1490 6000 1495
rect 5970 1470 5975 1490
rect 5975 1470 5995 1490
rect 5995 1470 6000 1490
rect 5970 1465 6000 1470
rect 6090 1490 6120 1495
rect 6090 1470 6095 1490
rect 6095 1470 6115 1490
rect 6115 1470 6120 1490
rect 6090 1465 6120 1470
rect 6210 1490 6240 1495
rect 6210 1470 6215 1490
rect 6215 1470 6235 1490
rect 6235 1470 6240 1490
rect 6210 1465 6240 1470
rect 6330 1490 6360 1495
rect 6330 1470 6335 1490
rect 6335 1470 6355 1490
rect 6355 1470 6360 1490
rect 6330 1465 6360 1470
rect 6720 1465 6750 1495
rect 4535 1110 4565 1115
rect 4535 1090 4540 1110
rect 4540 1090 4560 1110
rect 4560 1090 4565 1110
rect 4535 1085 4565 1090
rect 4615 1110 4645 1115
rect 4615 1090 4620 1110
rect 4620 1090 4640 1110
rect 4640 1090 4645 1110
rect 4615 1085 4645 1090
rect 4695 1110 4725 1115
rect 4695 1090 4700 1110
rect 4700 1090 4720 1110
rect 4720 1090 4725 1110
rect 4695 1085 4725 1090
rect 4775 1110 4805 1115
rect 4775 1090 4780 1110
rect 4780 1090 4800 1110
rect 4800 1090 4805 1110
rect 4775 1085 4805 1090
rect 4855 1110 4885 1115
rect 4855 1090 4860 1110
rect 4860 1090 4880 1110
rect 4880 1090 4885 1110
rect 4855 1085 4885 1090
rect 4935 1110 4965 1115
rect 4935 1090 4940 1110
rect 4940 1090 4960 1110
rect 4960 1090 4965 1110
rect 4935 1085 4965 1090
rect 5015 1110 5045 1115
rect 5015 1090 5020 1110
rect 5020 1090 5040 1110
rect 5040 1090 5045 1110
rect 5015 1085 5045 1090
rect 5095 1110 5125 1115
rect 5095 1090 5100 1110
rect 5100 1090 5120 1110
rect 5120 1090 5125 1110
rect 5095 1085 5125 1090
rect 5175 1110 5205 1115
rect 5175 1090 5180 1110
rect 5180 1090 5200 1110
rect 5200 1090 5205 1110
rect 5175 1085 5205 1090
rect 5255 1110 5285 1115
rect 5255 1090 5260 1110
rect 5260 1090 5280 1110
rect 5280 1090 5285 1110
rect 5255 1085 5285 1090
rect 5335 1110 5365 1115
rect 5335 1090 5340 1110
rect 5340 1090 5360 1110
rect 5360 1090 5365 1110
rect 5335 1085 5365 1090
rect 5415 1110 5445 1115
rect 5415 1090 5420 1110
rect 5420 1090 5440 1110
rect 5440 1090 5445 1110
rect 5415 1085 5445 1090
rect 5495 1110 5525 1115
rect 5495 1090 5500 1110
rect 5500 1090 5520 1110
rect 5520 1090 5525 1110
rect 5495 1085 5525 1090
rect 5575 1110 5605 1115
rect 5575 1090 5580 1110
rect 5580 1090 5600 1110
rect 5600 1090 5605 1110
rect 5575 1085 5605 1090
rect 5655 1110 5685 1115
rect 5655 1090 5660 1110
rect 5660 1090 5680 1110
rect 5680 1090 5685 1110
rect 5655 1085 5685 1090
rect 5735 1110 5765 1115
rect 5735 1090 5740 1110
rect 5740 1090 5760 1110
rect 5760 1090 5765 1110
rect 5735 1085 5765 1090
rect 5815 1110 5845 1115
rect 5815 1090 5820 1110
rect 5820 1090 5840 1110
rect 5840 1090 5845 1110
rect 5815 1085 5845 1090
rect 5895 1110 5925 1115
rect 5895 1090 5900 1110
rect 5900 1090 5920 1110
rect 5920 1090 5925 1110
rect 5895 1085 5925 1090
rect 5975 1110 6005 1115
rect 5975 1090 5980 1110
rect 5980 1090 6000 1110
rect 6000 1090 6005 1110
rect 5975 1085 6005 1090
rect 6055 1110 6085 1115
rect 6055 1090 6060 1110
rect 6060 1090 6080 1110
rect 6080 1090 6085 1110
rect 6055 1085 6085 1090
rect 6135 1110 6165 1115
rect 6135 1090 6140 1110
rect 6140 1090 6160 1110
rect 6160 1090 6165 1110
rect 6135 1085 6165 1090
rect 6215 1110 6245 1115
rect 6215 1090 6220 1110
rect 6220 1090 6240 1110
rect 6240 1090 6245 1110
rect 6215 1085 6245 1090
rect 6295 1110 6325 1115
rect 6295 1090 6300 1110
rect 6300 1090 6320 1110
rect 6320 1090 6325 1110
rect 6295 1085 6325 1090
rect 6375 1110 6405 1115
rect 6375 1090 6380 1110
rect 6380 1090 6400 1110
rect 6400 1090 6405 1110
rect 6375 1085 6405 1090
rect 6455 1110 6485 1115
rect 6455 1090 6460 1110
rect 6460 1090 6480 1110
rect 6480 1090 6485 1110
rect 6455 1085 6485 1090
rect 6535 1110 6565 1115
rect 6535 1090 6540 1110
rect 6540 1090 6560 1110
rect 6560 1090 6565 1110
rect 6535 1085 6565 1090
rect 4010 1000 4040 1030
rect 4495 1025 4525 1030
rect 4495 1005 4500 1025
rect 4500 1005 4520 1025
rect 4520 1005 4525 1025
rect 4495 1000 4525 1005
rect 3835 840 3865 870
rect 2325 800 2355 830
rect 2465 825 2500 830
rect 2465 800 2470 825
rect 2470 800 2495 825
rect 2495 800 2500 825
rect 2465 795 2500 800
rect 2465 765 2500 770
rect 2465 740 2470 765
rect 2470 740 2495 765
rect 2495 740 2500 765
rect 2465 735 2500 740
rect 6845 700 6875 730
rect 3110 600 3140 630
rect -835 -405 -800 -400
rect -835 -430 -830 -405
rect -830 -430 -805 -405
rect -805 -430 -800 -405
rect -835 -435 -800 -430
rect -885 -495 -855 -465
rect -835 -465 -800 -460
rect -835 -490 -830 -465
rect -830 -490 -805 -465
rect -805 -490 -800 -465
rect -835 -495 -800 -490
rect -935 -555 -905 -525
rect -835 -525 -800 -520
rect -835 -550 -830 -525
rect -830 -550 -805 -525
rect -805 -550 -800 -525
rect -835 -555 -800 -550
rect -975 -945 -940 -940
rect -975 -970 -970 -945
rect -970 -970 -945 -945
rect -945 -970 -940 -945
rect -975 -975 -940 -970
rect -835 -945 -800 -940
rect -835 -970 -830 -945
rect -830 -970 -805 -945
rect -805 -970 -800 -945
rect -835 -975 -800 -970
rect -16 -945 19 -940
rect -16 -970 -11 -945
rect -11 -970 14 -945
rect 14 -970 19 -945
rect -16 -975 19 -970
rect -945 -1395 -915 -1365
rect -835 -1365 -800 -1360
rect -835 -1390 -830 -1365
rect -830 -1390 -805 -1365
rect -805 -1390 -800 -1365
rect -835 -1395 -800 -1390
rect -890 -1455 -860 -1425
rect -835 -1425 -800 -1420
rect -835 -1450 -830 -1425
rect -830 -1450 -805 -1425
rect -805 -1450 -800 -1425
rect -835 -1455 -800 -1450
rect -835 -1485 -800 -1480
rect -835 -1510 -830 -1485
rect -830 -1510 -805 -1485
rect -805 -1510 -800 -1485
rect -835 -1515 -800 -1510
rect -890 -1590 -860 -1560
<< metal2 >>
rect -195 4485 -155 4490
rect -195 4455 -190 4485
rect -160 4455 -155 4485
rect -195 4450 -155 4455
rect 7375 4485 7415 4490
rect 7375 4455 7380 4485
rect 7410 4455 7415 4485
rect 7375 4450 7415 4455
rect -195 4350 -155 4355
rect -195 4320 -190 4350
rect -160 4345 -155 4350
rect 7375 4350 7415 4355
rect 7375 4345 7380 4350
rect -160 4325 2755 4345
rect 7290 4325 7380 4345
rect -160 4320 -155 4325
rect -195 4315 -155 4320
rect 7375 4320 7380 4325
rect 7410 4320 7415 4350
rect 7375 4315 7415 4320
rect 4545 3075 4585 3080
rect 4545 3045 4550 3075
rect 4580 3070 4585 3075
rect 7035 3075 7075 3080
rect 7035 3070 7040 3075
rect 4580 3050 7040 3070
rect 4580 3045 4585 3050
rect 4545 3040 4585 3045
rect 7035 3045 7040 3050
rect 7070 3045 7075 3075
rect 7035 3040 7075 3045
rect 4545 2905 4585 2945
rect 4580 2750 4620 2755
rect 4580 2720 4585 2750
rect 4615 2745 4620 2750
rect 4760 2750 4800 2755
rect 4760 2745 4765 2750
rect 4615 2725 4765 2745
rect 4615 2720 4620 2725
rect 4580 2715 4620 2720
rect 4760 2720 4765 2725
rect 4795 2745 4800 2750
rect 4940 2750 4980 2755
rect 4940 2745 4945 2750
rect 4795 2725 4945 2745
rect 4795 2720 4800 2725
rect 4760 2715 4800 2720
rect 4940 2720 4945 2725
rect 4975 2745 4980 2750
rect 5120 2750 5160 2755
rect 5120 2745 5125 2750
rect 4975 2725 5125 2745
rect 4975 2720 4980 2725
rect 4940 2715 4980 2720
rect 5120 2720 5125 2725
rect 5155 2745 5160 2750
rect 5300 2750 5340 2755
rect 5300 2745 5305 2750
rect 5155 2725 5305 2745
rect 5155 2720 5160 2725
rect 5120 2715 5160 2720
rect 5300 2720 5305 2725
rect 5335 2745 5340 2750
rect 5480 2750 5520 2755
rect 5480 2745 5485 2750
rect 5335 2725 5485 2745
rect 5335 2720 5340 2725
rect 5300 2715 5340 2720
rect 5480 2720 5485 2725
rect 5515 2745 5520 2750
rect 5660 2750 5700 2755
rect 5660 2745 5665 2750
rect 5515 2725 5665 2745
rect 5515 2720 5520 2725
rect 5480 2715 5520 2720
rect 5660 2720 5665 2725
rect 5695 2745 5700 2750
rect 5840 2750 5880 2755
rect 5840 2745 5845 2750
rect 5695 2725 5845 2745
rect 5695 2720 5700 2725
rect 5660 2715 5700 2720
rect 5840 2720 5845 2725
rect 5875 2745 5880 2750
rect 6020 2750 6060 2755
rect 6020 2745 6025 2750
rect 5875 2725 6025 2745
rect 5875 2720 5880 2725
rect 5840 2715 5880 2720
rect 6020 2720 6025 2725
rect 6055 2745 6060 2750
rect 6200 2750 6240 2755
rect 6200 2745 6205 2750
rect 6055 2725 6205 2745
rect 6055 2720 6060 2725
rect 6020 2715 6060 2720
rect 6200 2720 6205 2725
rect 6235 2745 6240 2750
rect 6380 2750 6420 2755
rect 6380 2745 6385 2750
rect 6235 2725 6385 2745
rect 6235 2720 6240 2725
rect 6200 2715 6240 2720
rect 6380 2720 6385 2725
rect 6415 2745 6420 2750
rect 6560 2750 6600 2755
rect 6560 2745 6565 2750
rect 6415 2725 6565 2745
rect 6415 2720 6420 2725
rect 6380 2715 6420 2720
rect 6560 2720 6565 2725
rect 6595 2720 6600 2750
rect 6560 2715 6600 2720
rect 4670 2380 4710 2385
rect 4580 2375 4620 2380
rect 4210 2345 4250 2350
rect 4210 2315 4215 2345
rect 4245 2340 4250 2345
rect 4580 2345 4585 2375
rect 4615 2345 4620 2375
rect 4670 2350 4675 2380
rect 4705 2375 4710 2380
rect 5400 2380 5440 2385
rect 5400 2375 5405 2380
rect 4705 2355 5405 2375
rect 4705 2350 4710 2355
rect 4670 2345 4710 2350
rect 5400 2350 5405 2355
rect 5435 2375 5440 2380
rect 5740 2380 5780 2385
rect 5740 2375 5745 2380
rect 5435 2355 5745 2375
rect 5435 2350 5440 2355
rect 5400 2345 5440 2350
rect 5740 2350 5745 2355
rect 5775 2375 5780 2380
rect 6470 2380 6510 2385
rect 6470 2375 6475 2380
rect 5775 2355 6475 2375
rect 5775 2350 5780 2355
rect 5740 2345 5780 2350
rect 6470 2350 6475 2355
rect 6505 2350 6510 2380
rect 6470 2345 6510 2350
rect 4580 2340 4620 2345
rect 4245 2320 4620 2340
rect 4850 2335 4890 2340
rect 4245 2315 4250 2320
rect 4210 2310 4250 2315
rect 4850 2305 4855 2335
rect 4885 2330 4890 2335
rect 5210 2335 5250 2340
rect 5210 2330 5215 2335
rect 4885 2310 5215 2330
rect 4885 2305 4890 2310
rect 4850 2300 4890 2305
rect 5210 2305 5215 2310
rect 5245 2330 5250 2335
rect 5930 2335 5970 2340
rect 5930 2330 5935 2335
rect 5245 2310 5935 2330
rect 5245 2305 5250 2310
rect 5210 2300 5250 2305
rect 5930 2305 5935 2310
rect 5965 2330 5970 2335
rect 6290 2335 6330 2340
rect 6290 2330 6295 2335
rect 5965 2310 6295 2330
rect 5965 2305 5970 2310
rect 5930 2300 5970 2305
rect 6290 2305 6295 2310
rect 6325 2305 6330 2335
rect 6290 2300 6330 2305
rect 3830 2290 3870 2295
rect 3830 2260 3835 2290
rect 3865 2285 3870 2290
rect 5030 2290 5070 2295
rect 5030 2285 5035 2290
rect 3865 2265 5035 2285
rect 3865 2260 3870 2265
rect 3830 2255 3870 2260
rect 5030 2260 5035 2265
rect 5065 2285 5070 2290
rect 6110 2290 6150 2295
rect 6110 2285 6115 2290
rect 5065 2265 6115 2285
rect 5065 2260 5070 2265
rect 5030 2255 5070 2260
rect 6110 2260 6115 2265
rect 6145 2285 6150 2290
rect 6840 2290 6880 2295
rect 6840 2285 6845 2290
rect 6145 2265 6845 2285
rect 6145 2260 6150 2265
rect 6110 2255 6150 2260
rect 6840 2260 6845 2265
rect 6875 2260 6880 2290
rect 6840 2255 6880 2260
rect 7375 2230 7415 2235
rect 7375 2225 7380 2230
rect 7290 2205 7380 2225
rect 7375 2200 7380 2205
rect 7410 2200 7415 2230
rect 4055 2195 4095 2200
rect 4055 2165 4060 2195
rect 4090 2190 4095 2195
rect 4670 2195 4710 2200
rect 7375 2195 7415 2200
rect 4670 2190 4675 2195
rect 4090 2170 4675 2190
rect 4090 2165 4095 2170
rect 4055 2160 4095 2165
rect 4670 2165 4675 2170
rect 4705 2165 4710 2195
rect 4670 2160 4710 2165
rect 4005 2145 4045 2150
rect 4005 2115 4010 2145
rect 4040 2140 4045 2145
rect 4490 2145 4530 2150
rect 4490 2140 4495 2145
rect 4040 2120 4495 2140
rect 4040 2115 4045 2120
rect 4005 2110 4045 2115
rect 4490 2115 4495 2120
rect 4525 2140 4530 2145
rect 5570 2145 5610 2150
rect 5570 2140 5575 2145
rect 4525 2120 5575 2140
rect 4525 2115 4530 2120
rect 4490 2110 4530 2115
rect 5570 2115 5575 2120
rect 5605 2140 5610 2145
rect 6650 2145 6690 2150
rect 6650 2140 6655 2145
rect 5605 2120 6655 2140
rect 5605 2115 5610 2120
rect 5570 2110 5610 2115
rect 6650 2115 6655 2120
rect 6685 2115 6690 2145
rect 6650 2110 6690 2115
rect 4100 2100 4140 2105
rect 4100 2070 4105 2100
rect 4135 2095 4140 2100
rect 4850 2100 4890 2105
rect 4850 2095 4855 2100
rect 4135 2075 4855 2095
rect 4135 2070 4140 2075
rect 4100 2065 4140 2070
rect 4850 2070 4855 2075
rect 4885 2070 4890 2100
rect 4850 2065 4890 2070
rect 5795 2095 5835 2100
rect 5795 2065 5800 2095
rect 5830 2090 5835 2095
rect 7035 2095 7075 2100
rect 7035 2090 7040 2095
rect 5830 2070 7040 2090
rect 5830 2065 5835 2070
rect 5795 2060 5835 2065
rect 7035 2065 7040 2070
rect 7070 2065 7075 2095
rect 7035 2060 7075 2065
rect 4455 2045 4495 2050
rect 4455 2015 4460 2045
rect 4490 2040 4495 2045
rect 4575 2045 4615 2050
rect 4575 2040 4580 2045
rect 4490 2020 4580 2040
rect 4490 2015 4495 2020
rect 4455 2010 4495 2015
rect 4575 2015 4580 2020
rect 4610 2040 4615 2045
rect 4695 2045 4735 2050
rect 4695 2040 4700 2045
rect 4610 2020 4700 2040
rect 4610 2015 4615 2020
rect 4575 2010 4615 2015
rect 4695 2015 4700 2020
rect 4730 2040 4735 2045
rect 4815 2045 4855 2050
rect 4815 2040 4820 2045
rect 4730 2020 4820 2040
rect 4730 2015 4735 2020
rect 4695 2010 4735 2015
rect 4815 2015 4820 2020
rect 4850 2040 4855 2045
rect 4935 2045 4975 2050
rect 4935 2040 4940 2045
rect 4850 2020 4940 2040
rect 4850 2015 4855 2020
rect 4815 2010 4855 2015
rect 4935 2015 4940 2020
rect 4970 2040 4975 2045
rect 5055 2045 5095 2050
rect 5055 2040 5060 2045
rect 4970 2020 5060 2040
rect 4970 2015 4975 2020
rect 4935 2010 4975 2015
rect 5055 2015 5060 2020
rect 5090 2040 5095 2045
rect 5175 2045 5215 2050
rect 5175 2040 5180 2045
rect 5090 2020 5180 2040
rect 5090 2015 5095 2020
rect 5055 2010 5095 2015
rect 5175 2015 5180 2020
rect 5210 2040 5215 2045
rect 5295 2045 5335 2050
rect 5295 2040 5300 2045
rect 5210 2020 5300 2040
rect 5210 2015 5215 2020
rect 5175 2010 5215 2015
rect 5295 2015 5300 2020
rect 5330 2040 5335 2045
rect 5415 2045 5455 2050
rect 5415 2040 5420 2045
rect 5330 2020 5420 2040
rect 5330 2015 5335 2020
rect 5295 2010 5335 2015
rect 5415 2015 5420 2020
rect 5450 2015 5455 2045
rect 5415 2010 5455 2015
rect 5725 2045 5765 2050
rect 5725 2015 5730 2045
rect 5760 2040 5765 2045
rect 5845 2045 5885 2050
rect 5845 2040 5850 2045
rect 5760 2020 5850 2040
rect 5760 2015 5765 2020
rect 5725 2010 5765 2015
rect 5845 2015 5850 2020
rect 5880 2040 5885 2045
rect 5965 2045 6005 2050
rect 5965 2040 5970 2045
rect 5880 2020 5970 2040
rect 5880 2015 5885 2020
rect 5845 2010 5885 2015
rect 5965 2015 5970 2020
rect 6000 2040 6005 2045
rect 6085 2045 6125 2050
rect 6085 2040 6090 2045
rect 6000 2020 6090 2040
rect 6000 2015 6005 2020
rect 5965 2010 6005 2015
rect 6085 2015 6090 2020
rect 6120 2040 6125 2045
rect 6205 2045 6245 2050
rect 6205 2040 6210 2045
rect 6120 2020 6210 2040
rect 6120 2015 6125 2020
rect 6085 2010 6125 2015
rect 6205 2015 6210 2020
rect 6240 2040 6245 2045
rect 6325 2045 6365 2050
rect 6325 2040 6330 2045
rect 6240 2020 6330 2040
rect 6240 2015 6245 2020
rect 6205 2010 6245 2015
rect 6325 2015 6330 2020
rect 6360 2040 6365 2045
rect 6445 2045 6485 2050
rect 6445 2040 6450 2045
rect 6360 2020 6450 2040
rect 6360 2015 6365 2020
rect 6325 2010 6365 2015
rect 6445 2015 6450 2020
rect 6480 2040 6485 2045
rect 6565 2045 6605 2050
rect 6565 2040 6570 2045
rect 6480 2020 6570 2040
rect 6480 2015 6485 2020
rect 6445 2010 6485 2015
rect 6565 2015 6570 2020
rect 6600 2040 6605 2045
rect 6685 2045 6725 2050
rect 6685 2040 6690 2045
rect 6600 2020 6690 2040
rect 6600 2015 6605 2020
rect 6565 2010 6605 2015
rect 6685 2015 6690 2020
rect 6720 2015 6725 2045
rect 6685 2010 6725 2015
rect 4210 2000 4250 2005
rect 4210 1970 4215 2000
rect 4245 1970 4250 2000
rect 4210 1965 4250 1970
rect 4395 2000 4435 2005
rect 4395 1970 4400 2000
rect 4430 1995 4435 2000
rect 4755 2000 4795 2005
rect 4755 1995 4760 2000
rect 4430 1975 4760 1995
rect 4430 1970 4435 1975
rect 4395 1965 4435 1970
rect 4755 1970 4760 1975
rect 4790 1995 4795 2000
rect 5115 2000 5155 2005
rect 5115 1995 5120 2000
rect 4790 1975 5120 1995
rect 4790 1970 4795 1975
rect 4755 1965 4795 1970
rect 5115 1970 5120 1975
rect 5150 1995 5155 2000
rect 5475 2000 5515 2005
rect 5475 1995 5480 2000
rect 5150 1975 5480 1995
rect 5150 1970 5155 1975
rect 5115 1965 5155 1970
rect 5475 1970 5480 1975
rect 5510 1970 5515 2000
rect 5475 1965 5515 1970
rect 5665 2000 5705 2005
rect 5665 1970 5670 2000
rect 5700 1995 5705 2000
rect 6025 2000 6065 2005
rect 6025 1995 6030 2000
rect 5700 1975 6030 1995
rect 5700 1970 5705 1975
rect 5665 1965 5705 1970
rect 6025 1970 6030 1975
rect 6060 1995 6065 2000
rect 6385 2000 6425 2005
rect 6385 1995 6390 2000
rect 6060 1975 6390 1995
rect 6060 1970 6065 1975
rect 6025 1965 6065 1970
rect 6385 1970 6390 1975
rect 6420 1995 6425 2000
rect 6745 2000 6785 2005
rect 6745 1995 6750 2000
rect 6420 1975 6750 1995
rect 6420 1970 6425 1975
rect 6385 1965 6425 1970
rect 6745 1970 6750 1975
rect 6780 1970 6785 2000
rect 6745 1965 6785 1970
rect 4005 1830 4045 1835
rect 4005 1800 4010 1830
rect 4040 1825 4045 1830
rect 4210 1830 4250 1835
rect 4210 1825 4215 1830
rect 4040 1805 4215 1825
rect 4040 1800 4045 1805
rect 4005 1795 4045 1800
rect 4210 1800 4215 1805
rect 4245 1800 4250 1830
rect 4210 1795 4250 1800
rect 4515 1830 4555 1835
rect 4515 1800 4520 1830
rect 4550 1825 4555 1830
rect 4635 1825 4675 1835
rect 4875 1830 4915 1835
rect 4875 1825 4880 1830
rect 4550 1805 4880 1825
rect 4550 1800 4555 1805
rect 4515 1795 4555 1800
rect 4635 1795 4675 1805
rect 4875 1800 4880 1805
rect 4910 1825 4915 1830
rect 4995 1825 5035 1835
rect 5235 1830 5275 1835
rect 5235 1825 5240 1830
rect 4910 1805 5240 1825
rect 4910 1800 4915 1805
rect 4875 1795 4915 1800
rect 4995 1795 5035 1805
rect 5235 1800 5240 1805
rect 5270 1800 5275 1830
rect 5235 1795 5275 1800
rect 5355 1795 5395 1835
rect 5785 1795 5825 1835
rect 5905 1830 5945 1835
rect 5905 1800 5910 1830
rect 5940 1825 5945 1830
rect 6145 1825 6185 1835
rect 6265 1830 6305 1835
rect 6265 1825 6270 1830
rect 5940 1805 6270 1825
rect 5940 1800 5945 1805
rect 5905 1795 5945 1800
rect 6145 1795 6185 1805
rect 6265 1800 6270 1805
rect 6300 1825 6305 1830
rect 6505 1825 6545 1835
rect 6625 1830 6665 1835
rect 6625 1825 6630 1830
rect 6300 1805 6630 1825
rect 6300 1800 6305 1805
rect 6265 1795 6305 1800
rect 6505 1795 6545 1805
rect 6625 1800 6630 1805
rect 6660 1800 6665 1830
rect 6625 1795 6665 1800
rect 4425 1770 4465 1775
rect 4425 1740 4430 1770
rect 4460 1765 4465 1770
rect 4635 1770 4675 1775
rect 4635 1765 4640 1770
rect 4460 1745 4640 1765
rect 4460 1740 4465 1745
rect 4425 1735 4465 1740
rect 4635 1740 4640 1745
rect 4670 1765 4675 1770
rect 4755 1770 4795 1775
rect 4755 1765 4760 1770
rect 4670 1745 4760 1765
rect 4670 1740 4675 1745
rect 4635 1735 4675 1740
rect 4755 1740 4760 1745
rect 4790 1765 4795 1770
rect 4995 1770 5035 1775
rect 4995 1765 5000 1770
rect 4790 1745 5000 1765
rect 4790 1740 4795 1745
rect 4755 1735 4795 1740
rect 4995 1740 5000 1745
rect 5030 1765 5035 1770
rect 5115 1770 5155 1775
rect 5115 1765 5120 1770
rect 5030 1745 5120 1765
rect 5030 1740 5035 1745
rect 4995 1735 5035 1740
rect 5115 1740 5120 1745
rect 5150 1765 5155 1770
rect 5355 1770 5395 1775
rect 5355 1765 5360 1770
rect 5150 1745 5360 1765
rect 5150 1740 5155 1745
rect 5115 1735 5155 1740
rect 5355 1740 5360 1745
rect 5390 1765 5395 1770
rect 5445 1770 5485 1775
rect 5445 1765 5450 1770
rect 5390 1745 5450 1765
rect 5390 1740 5395 1745
rect 5355 1735 5395 1740
rect 5445 1740 5450 1745
rect 5480 1740 5485 1770
rect 5445 1735 5485 1740
rect 5695 1770 5735 1775
rect 5695 1740 5700 1770
rect 5730 1765 5735 1770
rect 5785 1770 5825 1775
rect 5785 1765 5790 1770
rect 5730 1745 5790 1765
rect 5730 1740 5735 1745
rect 5695 1735 5735 1740
rect 5785 1740 5790 1745
rect 5820 1765 5825 1770
rect 6025 1770 6065 1775
rect 6025 1765 6030 1770
rect 5820 1745 6030 1765
rect 5820 1740 5825 1745
rect 5785 1735 5825 1740
rect 6025 1740 6030 1745
rect 6060 1765 6065 1770
rect 6145 1770 6185 1775
rect 6145 1765 6150 1770
rect 6060 1745 6150 1765
rect 6060 1740 6065 1745
rect 6025 1735 6065 1740
rect 6145 1740 6150 1745
rect 6180 1765 6185 1770
rect 6385 1770 6425 1775
rect 6385 1765 6390 1770
rect 6180 1745 6390 1765
rect 6180 1740 6185 1745
rect 6145 1735 6185 1740
rect 6385 1740 6390 1745
rect 6420 1765 6425 1770
rect 6505 1770 6545 1775
rect 6505 1765 6510 1770
rect 6420 1745 6510 1765
rect 6420 1740 6425 1745
rect 6385 1735 6425 1740
rect 6505 1740 6510 1745
rect 6540 1765 6545 1770
rect 6715 1770 6755 1775
rect 6715 1765 6720 1770
rect 6540 1745 6720 1765
rect 6540 1740 6545 1745
rect 6505 1735 6545 1740
rect 6715 1740 6720 1745
rect 6750 1740 6755 1770
rect 6715 1735 6755 1740
rect -110 1720 -70 1725
rect -110 1690 -105 1720
rect -75 1690 -70 1720
rect -110 1685 -70 1690
rect -45 1720 -5 1725
rect -45 1690 -40 1720
rect -10 1690 -5 1720
rect -45 1685 -5 1690
rect 1265 1710 1305 1715
rect 1265 1680 1270 1710
rect 1300 1705 1305 1710
rect 3585 1710 3625 1715
rect 3585 1705 3590 1710
rect 1300 1685 3590 1705
rect 1300 1680 1305 1685
rect 1265 1675 1305 1680
rect 3585 1680 3590 1685
rect 3620 1705 3625 1710
rect 4100 1710 4140 1715
rect 4100 1705 4105 1710
rect 3620 1685 4105 1705
rect 3620 1680 3625 1685
rect 3585 1675 3625 1680
rect 4100 1680 4105 1685
rect 4135 1705 4140 1710
rect 4155 1710 4195 1715
rect 4155 1705 4160 1710
rect 4135 1685 4160 1705
rect 4135 1680 4140 1685
rect 4100 1675 4140 1680
rect 4155 1680 4160 1685
rect 4190 1705 4195 1710
rect 4265 1710 4305 1715
rect 4265 1705 4270 1710
rect 4190 1685 4270 1705
rect 4190 1680 4195 1685
rect 4155 1675 4195 1680
rect 4265 1680 4270 1685
rect 4300 1705 4305 1710
rect 4815 1710 4855 1715
rect 4815 1705 4820 1710
rect 4300 1685 4820 1705
rect 4300 1680 4305 1685
rect 4265 1675 4305 1680
rect 4815 1680 4820 1685
rect 4850 1680 4855 1710
rect 4815 1675 4855 1680
rect 4875 1710 4915 1715
rect 4875 1680 4880 1710
rect 4910 1705 4915 1710
rect 5115 1710 5155 1715
rect 5115 1705 5120 1710
rect 4910 1685 5120 1705
rect 4910 1680 4915 1685
rect 4875 1675 4915 1680
rect 5115 1680 5120 1685
rect 5150 1705 5155 1710
rect 5355 1710 5395 1715
rect 5355 1705 5360 1710
rect 5150 1685 5360 1705
rect 5150 1680 5155 1685
rect 5115 1675 5155 1680
rect 5355 1680 5360 1685
rect 5390 1680 5395 1710
rect 5355 1675 5395 1680
rect 5785 1710 5825 1715
rect 5785 1680 5790 1710
rect 5820 1705 5825 1710
rect 6025 1710 6065 1715
rect 6025 1705 6030 1710
rect 5820 1685 6030 1705
rect 5820 1680 5825 1685
rect 5785 1675 5825 1680
rect 6025 1680 6030 1685
rect 6060 1705 6065 1710
rect 6265 1710 6305 1715
rect 6265 1705 6270 1710
rect 6060 1685 6270 1705
rect 6060 1680 6065 1685
rect 6025 1675 6065 1680
rect 6265 1680 6270 1685
rect 6300 1680 6305 1710
rect 6265 1675 6305 1680
rect 6325 1710 6365 1715
rect 6325 1680 6330 1710
rect 6360 1705 6365 1710
rect 6840 1710 6880 1715
rect 6840 1705 6845 1710
rect 6360 1685 6845 1705
rect 6360 1680 6365 1685
rect 6325 1675 6365 1680
rect 6840 1680 6845 1685
rect 6875 1680 6880 1710
rect 6840 1675 6880 1680
rect 4755 1665 4795 1670
rect 4755 1635 4760 1665
rect 4790 1660 4795 1665
rect 4995 1665 5035 1670
rect 4995 1660 5000 1665
rect 4790 1640 5000 1660
rect 4790 1635 4795 1640
rect 4755 1630 4795 1635
rect 4995 1635 5000 1640
rect 5030 1660 5035 1665
rect 5235 1665 5275 1670
rect 5235 1660 5240 1665
rect 5030 1640 5240 1660
rect 5030 1635 5035 1640
rect 4995 1630 5035 1635
rect 5235 1635 5240 1640
rect 5270 1635 5275 1665
rect 5235 1630 5275 1635
rect 5905 1665 5945 1670
rect 5905 1635 5910 1665
rect 5940 1660 5945 1665
rect 6145 1665 6185 1670
rect 6145 1660 6150 1665
rect 5940 1640 6150 1660
rect 5940 1635 5945 1640
rect 5905 1630 5945 1635
rect 6145 1635 6150 1640
rect 6180 1660 6185 1665
rect 6385 1665 6425 1670
rect 6385 1660 6390 1665
rect 6180 1640 6390 1660
rect 6180 1635 6185 1640
rect 6145 1630 6185 1635
rect 6385 1635 6390 1640
rect 6420 1635 6425 1665
rect 6385 1630 6425 1635
rect 3585 1605 3625 1610
rect 3425 1570 3430 1605
rect 3465 1600 3470 1605
rect 3585 1600 3590 1605
rect 3465 1580 3590 1600
rect 3465 1570 3470 1580
rect 3585 1575 3590 1580
rect 3620 1575 3625 1605
rect 3585 1570 3625 1575
rect 3585 1545 3625 1550
rect 3425 1510 3430 1545
rect 3465 1540 3470 1545
rect 3585 1540 3590 1545
rect 3465 1520 3590 1540
rect 3465 1510 3470 1520
rect 3585 1515 3590 1520
rect 3620 1540 3625 1545
rect 4055 1545 4095 1550
rect 4055 1540 4060 1545
rect 3620 1520 4060 1540
rect 3620 1515 3625 1520
rect 3585 1510 3625 1515
rect 4055 1515 4060 1520
rect 4090 1540 4095 1545
rect 4755 1545 4795 1550
rect 4755 1540 4760 1545
rect 4090 1520 4760 1540
rect 4090 1515 4095 1520
rect 4055 1510 4095 1515
rect 4755 1515 4760 1520
rect 4790 1515 4795 1545
rect 4755 1510 4795 1515
rect 6385 1545 6425 1550
rect 6385 1515 6390 1545
rect 6420 1540 6425 1545
rect 6840 1545 6880 1550
rect 6840 1540 6845 1545
rect 6420 1520 6845 1540
rect 6420 1515 6425 1520
rect 6385 1510 6425 1515
rect 6840 1515 6845 1520
rect 6875 1515 6880 1545
rect 6840 1510 6880 1515
rect 7290 1545 7330 1550
rect 7290 1515 7295 1545
rect 7325 1515 7330 1545
rect 7290 1510 7330 1515
rect 4425 1495 4465 1500
rect 4425 1465 4430 1495
rect 4460 1490 4465 1495
rect 4815 1495 4855 1500
rect 4815 1490 4820 1495
rect 4460 1470 4820 1490
rect 4460 1465 4465 1470
rect 4425 1460 4465 1465
rect 4815 1465 4820 1470
rect 4850 1490 4855 1495
rect 4935 1495 4975 1500
rect 4935 1490 4940 1495
rect 4850 1470 4940 1490
rect 4850 1465 4855 1470
rect 4815 1460 4855 1465
rect 4935 1465 4940 1470
rect 4970 1490 4975 1495
rect 5055 1495 5095 1500
rect 5055 1490 5060 1495
rect 4970 1470 5060 1490
rect 4970 1465 4975 1470
rect 4935 1460 4975 1465
rect 5055 1465 5060 1470
rect 5090 1490 5095 1495
rect 5175 1495 5215 1500
rect 5175 1490 5180 1495
rect 5090 1470 5180 1490
rect 5090 1465 5095 1470
rect 5055 1460 5095 1465
rect 5175 1465 5180 1470
rect 5210 1490 5215 1495
rect 5295 1495 5335 1500
rect 5295 1490 5300 1495
rect 5210 1470 5300 1490
rect 5210 1465 5215 1470
rect 5175 1460 5215 1465
rect 5295 1465 5300 1470
rect 5330 1465 5335 1495
rect 5295 1460 5335 1465
rect 5845 1495 5885 1500
rect 5845 1465 5850 1495
rect 5880 1490 5885 1495
rect 5965 1495 6005 1500
rect 5965 1490 5970 1495
rect 5880 1470 5970 1490
rect 5880 1465 5885 1470
rect 5845 1460 5885 1465
rect 5965 1465 5970 1470
rect 6000 1490 6005 1495
rect 6085 1495 6125 1500
rect 6085 1490 6090 1495
rect 6000 1470 6090 1490
rect 6000 1465 6005 1470
rect 5965 1460 6005 1465
rect 6085 1465 6090 1470
rect 6120 1490 6125 1495
rect 6205 1495 6245 1500
rect 6205 1490 6210 1495
rect 6120 1470 6210 1490
rect 6120 1465 6125 1470
rect 6085 1460 6125 1465
rect 6205 1465 6210 1470
rect 6240 1490 6245 1495
rect 6325 1495 6365 1500
rect 6325 1490 6330 1495
rect 6240 1470 6330 1490
rect 6240 1465 6245 1470
rect 6205 1460 6245 1465
rect 6325 1465 6330 1470
rect 6360 1490 6365 1495
rect 6715 1495 6755 1500
rect 6715 1490 6720 1495
rect 6360 1470 6720 1490
rect 6360 1465 6365 1470
rect 6325 1460 6365 1465
rect 6715 1465 6720 1470
rect 6750 1465 6755 1495
rect 6715 1460 6755 1465
rect 2340 1330 2345 1365
rect 2380 1330 2385 1365
rect 2340 1305 2385 1310
rect 2340 1270 2345 1305
rect 2380 1270 2385 1305
rect 2340 1265 2385 1270
rect 4530 1115 4570 1120
rect 4530 1085 4535 1115
rect 4565 1110 4570 1115
rect 4610 1115 4650 1120
rect 4610 1110 4615 1115
rect 4565 1090 4615 1110
rect 4565 1085 4570 1090
rect 4530 1080 4570 1085
rect 4610 1085 4615 1090
rect 4645 1110 4650 1115
rect 4690 1115 4730 1120
rect 4690 1110 4695 1115
rect 4645 1090 4695 1110
rect 4645 1085 4650 1090
rect 4610 1080 4650 1085
rect 4690 1085 4695 1090
rect 4725 1110 4730 1115
rect 4770 1115 4810 1120
rect 4770 1110 4775 1115
rect 4725 1090 4775 1110
rect 4725 1085 4730 1090
rect 4690 1080 4730 1085
rect 4770 1085 4775 1090
rect 4805 1110 4810 1115
rect 4850 1115 4890 1120
rect 4850 1110 4855 1115
rect 4805 1090 4855 1110
rect 4805 1085 4810 1090
rect 4770 1080 4810 1085
rect 4850 1085 4855 1090
rect 4885 1110 4890 1115
rect 4930 1115 4970 1120
rect 4930 1110 4935 1115
rect 4885 1090 4935 1110
rect 4885 1085 4890 1090
rect 4850 1080 4890 1085
rect 4930 1085 4935 1090
rect 4965 1110 4970 1115
rect 5010 1115 5050 1120
rect 5010 1110 5015 1115
rect 4965 1090 5015 1110
rect 4965 1085 4970 1090
rect 4930 1080 4970 1085
rect 5010 1085 5015 1090
rect 5045 1110 5050 1115
rect 5090 1115 5130 1120
rect 5090 1110 5095 1115
rect 5045 1090 5095 1110
rect 5045 1085 5050 1090
rect 5010 1080 5050 1085
rect 5090 1085 5095 1090
rect 5125 1110 5130 1115
rect 5170 1115 5210 1120
rect 5170 1110 5175 1115
rect 5125 1090 5175 1110
rect 5125 1085 5130 1090
rect 5090 1080 5130 1085
rect 5170 1085 5175 1090
rect 5205 1110 5210 1115
rect 5250 1115 5290 1120
rect 5250 1110 5255 1115
rect 5205 1090 5255 1110
rect 5205 1085 5210 1090
rect 5170 1080 5210 1085
rect 5250 1085 5255 1090
rect 5285 1110 5290 1115
rect 5330 1115 5370 1120
rect 5330 1110 5335 1115
rect 5285 1090 5335 1110
rect 5285 1085 5290 1090
rect 5250 1080 5290 1085
rect 5330 1085 5335 1090
rect 5365 1110 5370 1115
rect 5410 1115 5450 1120
rect 5410 1110 5415 1115
rect 5365 1090 5415 1110
rect 5365 1085 5370 1090
rect 5330 1080 5370 1085
rect 5410 1085 5415 1090
rect 5445 1110 5450 1115
rect 5490 1115 5530 1120
rect 5490 1110 5495 1115
rect 5445 1090 5495 1110
rect 5445 1085 5450 1090
rect 5410 1080 5450 1085
rect 5490 1085 5495 1090
rect 5525 1085 5530 1115
rect 5490 1080 5530 1085
rect 5570 1115 5610 1120
rect 5570 1085 5575 1115
rect 5605 1110 5610 1115
rect 5650 1115 5690 1120
rect 5650 1110 5655 1115
rect 5605 1090 5655 1110
rect 5605 1085 5610 1090
rect 5570 1080 5610 1085
rect 5650 1085 5655 1090
rect 5685 1110 5690 1115
rect 5730 1115 5770 1120
rect 5730 1110 5735 1115
rect 5685 1090 5735 1110
rect 5685 1085 5690 1090
rect 5650 1080 5690 1085
rect 5730 1085 5735 1090
rect 5765 1110 5770 1115
rect 5810 1115 5850 1120
rect 5810 1110 5815 1115
rect 5765 1090 5815 1110
rect 5765 1085 5770 1090
rect 5730 1080 5770 1085
rect 5810 1085 5815 1090
rect 5845 1110 5850 1115
rect 5890 1115 5930 1120
rect 5890 1110 5895 1115
rect 5845 1090 5895 1110
rect 5845 1085 5850 1090
rect 5810 1080 5850 1085
rect 5890 1085 5895 1090
rect 5925 1110 5930 1115
rect 5970 1115 6010 1120
rect 5970 1110 5975 1115
rect 5925 1090 5975 1110
rect 5925 1085 5930 1090
rect 5890 1080 5930 1085
rect 5970 1085 5975 1090
rect 6005 1110 6010 1115
rect 6050 1115 6090 1120
rect 6050 1110 6055 1115
rect 6005 1090 6055 1110
rect 6005 1085 6010 1090
rect 5970 1080 6010 1085
rect 6050 1085 6055 1090
rect 6085 1110 6090 1115
rect 6130 1115 6170 1120
rect 6130 1110 6135 1115
rect 6085 1090 6135 1110
rect 6085 1085 6090 1090
rect 6050 1080 6090 1085
rect 6130 1085 6135 1090
rect 6165 1110 6170 1115
rect 6210 1115 6250 1120
rect 6210 1110 6215 1115
rect 6165 1090 6215 1110
rect 6165 1085 6170 1090
rect 6130 1080 6170 1085
rect 6210 1085 6215 1090
rect 6245 1110 6250 1115
rect 6290 1115 6330 1120
rect 6290 1110 6295 1115
rect 6245 1090 6295 1110
rect 6245 1085 6250 1090
rect 6210 1080 6250 1085
rect 6290 1085 6295 1090
rect 6325 1110 6330 1115
rect 6370 1115 6410 1120
rect 6370 1110 6375 1115
rect 6325 1090 6375 1110
rect 6325 1085 6330 1090
rect 6290 1080 6330 1085
rect 6370 1085 6375 1090
rect 6405 1110 6410 1115
rect 6450 1115 6490 1120
rect 6450 1110 6455 1115
rect 6405 1090 6455 1110
rect 6405 1085 6410 1090
rect 6370 1080 6410 1085
rect 6450 1085 6455 1090
rect 6485 1110 6490 1115
rect 6530 1115 6570 1120
rect 6530 1110 6535 1115
rect 6485 1090 6535 1110
rect 6485 1085 6490 1090
rect 6450 1080 6490 1085
rect 6530 1085 6535 1090
rect 6565 1085 6570 1115
rect 6530 1080 6570 1085
rect 2175 1030 2215 1035
rect 3585 1030 3625 1035
rect 2175 1000 2180 1030
rect 2210 1025 2215 1030
rect 2345 1025 2350 1030
rect 2210 1005 2350 1025
rect 2210 1000 2215 1005
rect 2175 995 2215 1000
rect 2345 995 2350 1005
rect 2385 995 2390 1030
rect 3060 995 3065 1030
rect 3100 1025 3105 1030
rect 3585 1025 3590 1030
rect 3100 1005 3590 1025
rect 3100 995 3105 1005
rect 3585 1000 3590 1005
rect 3620 1000 3625 1030
rect 3585 995 3625 1000
rect 4005 1030 4045 1035
rect 4005 1000 4010 1030
rect 4040 1025 4045 1030
rect 4490 1030 4530 1035
rect 4490 1025 4495 1030
rect 4040 1005 4495 1025
rect 4040 1000 4045 1005
rect 4005 995 4045 1000
rect 4490 1000 4495 1005
rect 4525 1000 4530 1030
rect 4490 995 4530 1000
rect 2320 970 2360 975
rect 2320 940 2325 970
rect 2355 965 2360 970
rect 2460 965 2465 970
rect 2355 945 2465 965
rect 2355 940 2360 945
rect 2320 935 2360 940
rect 2460 935 2465 945
rect 2500 935 2505 970
rect 7290 965 7330 970
rect 7290 935 7295 965
rect 7325 935 7330 965
rect 7290 930 7330 935
rect 2460 875 2465 910
rect 2500 875 2505 910
rect 2460 865 2505 875
rect 3830 870 3870 875
rect 3830 865 3835 870
rect 2460 845 3835 865
rect 3830 840 3835 845
rect 3865 840 3870 870
rect 3830 835 3870 840
rect 2320 830 2360 835
rect 2320 800 2325 830
rect 2355 825 2360 830
rect 2460 825 2465 830
rect 2355 805 2465 825
rect 2355 800 2360 805
rect 2320 795 2360 800
rect 2460 795 2465 805
rect 2500 795 2505 830
rect 7290 820 7330 825
rect 7290 790 7295 820
rect 7325 790 7330 820
rect 7290 785 7330 790
rect 2460 735 2465 770
rect 2500 735 2505 770
rect 2460 725 2505 735
rect 6840 730 6880 735
rect 6840 725 6845 730
rect 2460 705 6845 725
rect 6840 700 6845 705
rect 6875 700 6880 730
rect 6840 695 6880 700
rect 3100 630 3150 640
rect 3100 600 3110 630
rect 3140 600 3150 630
rect 3100 590 3150 600
rect -195 550 -155 555
rect -195 520 -190 550
rect -160 520 -155 550
rect -195 515 -155 520
rect -840 -435 -835 -400
rect -800 -435 -795 -400
rect -890 -465 -855 -460
rect -840 -465 -835 -460
rect -890 -495 -885 -465
rect -855 -490 -835 -465
rect -840 -495 -835 -490
rect -800 -495 -795 -460
rect -890 -500 -855 -495
rect -940 -525 -900 -520
rect -840 -525 -835 -520
rect -940 -555 -935 -525
rect -905 -550 -835 -525
rect -905 -555 -900 -550
rect -840 -555 -835 -550
rect -800 -555 -795 -520
rect -940 -560 -900 -555
rect -940 -945 -935 -940
rect -840 -945 -835 -940
rect -940 -970 -835 -945
rect -940 -975 -935 -970
rect -840 -975 -835 -970
rect -800 -975 -795 -940
rect -21 -975 -16 -940
rect 19 -945 24 -940
rect 19 -970 285 -945
rect 19 -975 24 -970
rect -950 -1365 -910 -1360
rect -840 -1365 -835 -1360
rect -950 -1395 -945 -1365
rect -915 -1390 -835 -1365
rect -915 -1395 -910 -1390
rect -840 -1395 -835 -1390
rect -800 -1395 -795 -1360
rect -950 -1400 -910 -1395
rect -895 -1425 -855 -1420
rect -840 -1425 -835 -1420
rect -895 -1455 -890 -1425
rect -860 -1450 -835 -1425
rect -860 -1455 -855 -1450
rect -840 -1455 -835 -1450
rect -800 -1455 -795 -1420
rect -895 -1460 -855 -1455
rect -840 -1480 -795 -1475
rect -840 -1515 -835 -1480
rect -800 -1515 -795 -1480
rect -840 -1520 -795 -1515
rect -840 -1540 285 -1520
rect -895 -1560 -855 -1555
rect -895 -1590 -890 -1560
rect -860 -1565 -855 -1560
rect -860 -1585 285 -1565
rect -860 -1590 -855 -1585
rect -895 -1595 -855 -1590
<< via2 >>
rect -190 4455 -160 4485
rect 7380 4455 7410 4485
rect -190 4320 -160 4350
rect 7380 4320 7410 4350
rect 7380 2200 7410 2230
rect -105 1690 -75 1720
rect 7295 1515 7325 1545
rect 7295 935 7325 965
rect 7295 790 7325 820
rect 3110 600 3140 630
rect -190 520 -160 550
<< metal3 >>
rect -200 4490 -150 4495
rect -200 4450 -195 4490
rect -155 4450 -150 4490
rect -200 4445 -150 4450
rect 7370 4490 7420 4495
rect 7370 4450 7375 4490
rect 7415 4450 7420 4490
rect 7370 4445 7420 4450
rect -195 4350 -155 4445
rect -115 4405 -65 4410
rect -115 4365 -110 4405
rect -70 4365 -65 4405
rect -115 4360 -65 4365
rect 7285 4405 7335 4410
rect 7285 4365 7290 4405
rect 7330 4365 7335 4405
rect 7285 4360 7335 4365
rect -195 4320 -190 4350
rect -160 4320 -155 4350
rect -195 560 -155 4320
rect -110 1720 -70 4360
rect -110 1690 -105 1720
rect -75 1690 -70 1720
rect -110 640 -70 1690
rect 7290 1545 7330 4360
rect 7290 1515 7295 1545
rect 7325 1515 7330 1545
rect 7290 965 7330 1515
rect 7290 935 7295 965
rect 7325 935 7330 965
rect 7290 820 7330 935
rect 7290 790 7295 820
rect 7325 790 7330 820
rect 7290 640 7330 790
rect 7375 4350 7415 4445
rect 7375 4320 7380 4350
rect 7410 4320 7415 4350
rect 7375 2230 7415 4320
rect 7375 2200 7380 2230
rect 7410 2200 7415 2230
rect -115 635 -65 640
rect -115 595 -110 635
rect -70 595 -65 635
rect -115 590 -65 595
rect 3100 635 3150 640
rect 3100 595 3105 635
rect 3145 595 3150 635
rect 3100 590 3150 595
rect 7285 635 7335 640
rect 7285 595 7290 635
rect 7330 595 7335 635
rect 7285 590 7335 595
rect 7375 560 7415 2200
rect -200 555 -150 560
rect -200 515 -195 555
rect -155 515 -150 555
rect -200 510 -150 515
rect 7370 555 7420 560
rect 7370 515 7375 555
rect 7415 515 7420 555
rect 7370 510 7420 515
<< via3 >>
rect -195 4485 -155 4490
rect -195 4455 -190 4485
rect -190 4455 -160 4485
rect -160 4455 -155 4485
rect -195 4450 -155 4455
rect 7375 4485 7415 4490
rect 7375 4455 7380 4485
rect 7380 4455 7410 4485
rect 7410 4455 7415 4485
rect 7375 4450 7415 4455
rect -110 4365 -70 4405
rect 7290 4365 7330 4405
rect -110 595 -70 635
rect 3105 630 3145 635
rect 3105 600 3110 630
rect 3110 600 3140 630
rect 3140 600 3145 630
rect 3105 595 3145 600
rect 7290 595 7330 635
rect -195 550 -155 555
rect -195 520 -190 550
rect -190 520 -160 550
rect -160 520 -155 550
rect -195 515 -155 520
rect 7375 515 7415 555
<< metal4 >>
rect -200 4490 7420 4495
rect -200 4450 -195 4490
rect -155 4450 7375 4490
rect 7415 4450 7420 4490
rect -200 4445 7420 4450
rect -115 4405 7335 4410
rect -115 4365 -110 4405
rect -70 4365 7290 4405
rect 7330 4365 7335 4405
rect -115 4360 7335 4365
rect -115 635 7335 640
rect -115 595 -110 635
rect -70 595 3105 635
rect 3145 595 7290 635
rect 7330 595 7335 635
rect -115 590 7335 595
rect -200 555 7420 560
rect -200 515 -195 555
rect -155 515 7375 555
rect 7415 515 7420 555
rect -200 510 7420 515
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0 $PDKPATH/libs.ref/sky130_fd_pr/mag
timestamp 1723858470
transform 1 0 795 0 1 1360
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_1
timestamp 1723858470
transform 1 0 795 0 1 2040
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_2
timestamp 1723858470
transform 1 0 795 0 1 680
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_3
timestamp 1723858470
transform 1 0 115 0 1 2040
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_4
timestamp 1723858470
transform 1 0 115 0 1 1360
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5
timestamp 1723858470
transform 1 0 115 0 1 680
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_6
timestamp 1723858470
transform 1 0 1475 0 1 2040
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_7
timestamp 1723858470
transform 1 0 1475 0 1 680
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8
timestamp 1723858470
transform 1 0 1475 0 1 1360
box 0 0 670 670
<< labels >>
flabel metal3 7330 1175 7330 1175 3 FreeSans 800 0 80 0 GNDA
port 6 e
flabel metal3 7415 1400 7415 1400 3 FreeSans 800 0 80 0 VDDA
port 1 e
flabel metal1 3740 4675 3740 4675 1 FreeSans 800 0 0 400 V_OUT
port 2 n
<< end >>
