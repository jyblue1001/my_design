magic
tech sky130A
timestamp 1740153552
<< nwell >>
rect 2345 650 2870 940
rect 2910 920 4470 1880
<< poly >>
rect -130 960 -90 975
rect 2180 945 2220 955
rect 2180 930 2190 945
rect 2090 925 2190 930
rect 2210 925 2220 945
rect 2090 915 2220 925
rect 3090 680 3130 690
rect 3090 660 3100 680
rect 3120 660 3130 680
rect 3090 650 3130 660
rect 3850 680 3890 690
rect 3850 660 3860 680
rect 3880 660 3890 680
rect 3850 650 3890 660
rect 4070 490 4110 500
rect 4070 470 4080 490
rect 4100 470 4110 490
rect 4070 460 4110 470
rect -130 260 -90 270
rect -130 240 -120 260
rect -100 240 -90 260
rect -130 230 -90 240
rect 2075 85 2115 95
rect 2075 65 2085 85
rect 2105 65 2115 85
rect 2075 55 2115 65
<< polycont >>
rect 2190 925 2210 945
rect 3100 660 3120 680
rect 3860 660 3880 680
rect 4080 470 4100 490
rect -120 240 -100 260
rect 2085 65 2105 85
<< locali >>
rect 2775 2815 2825 2830
rect 2775 2795 2790 2815
rect 2810 2795 2825 2815
rect 2775 2780 2825 2795
rect 4820 2540 4860 2550
rect 4820 2520 4830 2540
rect 4850 2520 4860 2540
rect 4820 2510 4860 2520
rect 2775 2220 2825 2235
rect 2775 2200 2790 2220
rect 2810 2200 2825 2220
rect 2775 2185 2825 2200
rect 2380 1220 2430 1230
rect 2380 1210 2390 1220
rect 2355 1190 2390 1210
rect 2420 1190 2430 1220
rect 2380 1180 2430 1190
rect 2040 1155 2080 1165
rect 2040 1135 2050 1155
rect 2070 1135 2080 1155
rect 2040 1125 2080 1135
rect 2040 1105 2060 1125
rect 2735 1015 2785 1030
rect 2735 995 2750 1015
rect 2770 995 2785 1015
rect 2735 980 2785 995
rect 2180 945 2220 955
rect 2180 925 2190 945
rect 2210 925 2220 945
rect 2180 915 2220 925
rect 2300 945 2340 955
rect 2300 925 2310 945
rect 2330 925 2340 945
rect 2300 915 2340 925
rect 3090 680 3130 690
rect 3090 660 3100 680
rect 3120 660 3130 680
rect 3850 680 3890 690
rect 3090 650 3130 660
rect 3155 645 3195 665
rect 3850 660 3860 680
rect 3880 660 3890 680
rect 3850 650 3890 660
rect -190 625 -140 635
rect -190 595 -180 625
rect -150 620 -140 625
rect 2460 625 2510 640
rect 2460 620 2475 625
rect -150 600 -130 620
rect 2370 600 2400 620
rect 2420 605 2475 620
rect 2495 605 2510 625
rect 3155 625 3165 645
rect 3185 625 3195 645
rect 3155 615 3195 625
rect 2420 600 2510 605
rect -150 595 -140 600
rect -190 585 -140 595
rect 2460 590 2510 600
rect 4450 595 4490 605
rect 4450 575 4460 595
rect 4480 575 4490 595
rect 4450 565 4490 575
rect 2040 550 2220 560
rect 2040 540 2190 550
rect 2040 505 2060 540
rect 2180 530 2190 540
rect 2210 530 2220 550
rect 2180 520 2220 530
rect 4070 490 4110 500
rect 4070 470 4080 490
rect 4100 470 4110 490
rect 4070 460 4110 470
rect 2305 275 2345 285
rect -130 260 -90 270
rect -130 240 -120 260
rect -100 240 -90 260
rect 2305 255 2315 275
rect 2335 255 2345 275
rect 2305 245 2345 255
rect -130 230 -90 240
rect 2735 165 2785 180
rect 2735 145 2750 165
rect 2770 145 2785 165
rect 2735 130 2785 145
rect 2075 85 2115 95
rect 2075 65 2085 85
rect 2105 65 2115 85
rect 2075 55 2115 65
rect 2380 30 2430 40
rect 2355 10 2390 30
rect 2380 0 2390 10
rect 2420 0 2430 30
rect 2380 -10 2430 0
rect 2380 -225 2430 -215
rect 2380 -255 2390 -225
rect 2420 -235 2430 -225
rect 6950 -235 6970 -135
rect 2420 -255 2460 -235
rect 2480 -255 2510 -235
rect 2530 -255 2560 -235
rect 2580 -255 2610 -235
rect 2630 -255 2660 -235
rect 2680 -255 2710 -235
rect 2730 -255 2760 -235
rect 2780 -255 2810 -235
rect 2830 -255 2860 -235
rect 2880 -255 2910 -235
rect 2930 -255 2960 -235
rect 2980 -255 3010 -235
rect 3030 -255 3060 -235
rect 3080 -255 3110 -235
rect 3130 -255 3160 -235
rect 3180 -255 3210 -235
rect 3230 -255 3260 -235
rect 3280 -255 3310 -235
rect 3330 -255 3360 -235
rect 3380 -255 3410 -235
rect 3430 -255 3460 -235
rect 3480 -255 3510 -235
rect 3530 -255 3560 -235
rect 3580 -255 3610 -235
rect 3630 -255 3660 -235
rect 3680 -255 3710 -235
rect 3730 -255 3760 -235
rect 3780 -255 3810 -235
rect 3830 -255 3860 -235
rect 3880 -255 3910 -235
rect 3930 -255 3960 -235
rect 3980 -255 4010 -235
rect 4030 -255 4060 -235
rect 4080 -255 4110 -235
rect 4130 -255 4160 -235
rect 4180 -255 4210 -235
rect 4230 -255 4260 -235
rect 4280 -255 4310 -235
rect 4330 -255 4360 -235
rect 4380 -255 4410 -235
rect 4430 -255 4460 -235
rect 4480 -255 4510 -235
rect 4530 -255 4560 -235
rect 4580 -255 4610 -235
rect 4630 -255 4660 -235
rect 4680 -255 4710 -235
rect 4730 -255 4760 -235
rect 4780 -255 4810 -235
rect 4830 -255 4860 -235
rect 4880 -255 4910 -235
rect 4930 -255 4960 -235
rect 4980 -255 5010 -235
rect 5030 -255 5060 -235
rect 5080 -255 5110 -235
rect 5130 -255 5160 -235
rect 5180 -255 5210 -235
rect 5230 -255 5260 -235
rect 5280 -255 5310 -235
rect 5330 -255 5360 -235
rect 5380 -255 5410 -235
rect 5430 -255 5460 -235
rect 5480 -255 5510 -235
rect 5530 -255 5560 -235
rect 5580 -255 5610 -235
rect 5630 -255 5660 -235
rect 5680 -255 5710 -235
rect 5730 -255 5760 -235
rect 5780 -255 5810 -235
rect 5830 -255 5860 -235
rect 5880 -255 5910 -235
rect 5930 -255 5960 -235
rect 5980 -255 6010 -235
rect 6030 -255 6060 -235
rect 6080 -255 6110 -235
rect 6130 -255 6160 -235
rect 6180 -255 6210 -235
rect 6230 -255 6260 -235
rect 6280 -255 6310 -235
rect 6330 -255 6360 -235
rect 6380 -255 6410 -235
rect 6430 -255 6460 -235
rect 6480 -255 6510 -235
rect 6530 -255 6560 -235
rect 6580 -255 6610 -235
rect 6630 -255 6660 -235
rect 6680 -255 6710 -235
rect 6730 -255 6760 -235
rect 6780 -255 6810 -235
rect 6830 -255 6860 -235
rect 6880 -255 6910 -235
rect 6930 -255 6970 -235
rect 2380 -265 2430 -255
<< viali >>
rect 2790 2795 2810 2815
rect 4830 2520 4850 2540
rect 2790 2200 2810 2220
rect 2390 1190 2420 1220
rect 2050 1135 2070 1155
rect 2750 995 2770 1015
rect 2190 925 2210 945
rect 2310 925 2330 945
rect 3100 660 3120 680
rect 3860 660 3880 680
rect -180 595 -150 625
rect 2350 600 2370 620
rect 2400 600 2420 620
rect 2475 605 2495 625
rect 3165 625 3185 645
rect 4460 575 4480 595
rect 2190 530 2210 550
rect 3065 520 3085 540
rect 4080 470 4100 490
rect -120 240 -100 260
rect 2315 255 2335 275
rect 2750 145 2770 165
rect 2085 65 2105 85
rect 2390 0 2420 30
rect 2390 -255 2420 -225
rect 2460 -255 2480 -235
rect 2510 -255 2530 -235
rect 2560 -255 2580 -235
rect 2610 -255 2630 -235
rect 2660 -255 2680 -235
rect 2710 -255 2730 -235
rect 2760 -255 2780 -235
rect 2810 -255 2830 -235
rect 2860 -255 2880 -235
rect 2910 -255 2930 -235
rect 2960 -255 2980 -235
rect 3010 -255 3030 -235
rect 3060 -255 3080 -235
rect 3110 -255 3130 -235
rect 3160 -255 3180 -235
rect 3210 -255 3230 -235
rect 3260 -255 3280 -235
rect 3310 -255 3330 -235
rect 3360 -255 3380 -235
rect 3410 -255 3430 -235
rect 3460 -255 3480 -235
rect 3510 -255 3530 -235
rect 3560 -255 3580 -235
rect 3610 -255 3630 -235
rect 3660 -255 3680 -235
rect 3710 -255 3730 -235
rect 3760 -255 3780 -235
rect 3810 -255 3830 -235
rect 3860 -255 3880 -235
rect 3910 -255 3930 -235
rect 3960 -255 3980 -235
rect 4010 -255 4030 -235
rect 4060 -255 4080 -235
rect 4110 -255 4130 -235
rect 4160 -255 4180 -235
rect 4210 -255 4230 -235
rect 4260 -255 4280 -235
rect 4310 -255 4330 -235
rect 4360 -255 4380 -235
rect 4410 -255 4430 -235
rect 4460 -255 4480 -235
rect 4510 -255 4530 -235
rect 4560 -255 4580 -235
rect 4610 -255 4630 -235
rect 4660 -255 4680 -235
rect 4710 -255 4730 -235
rect 4760 -255 4780 -235
rect 4810 -255 4830 -235
rect 4860 -255 4880 -235
rect 4910 -255 4930 -235
rect 4960 -255 4980 -235
rect 5010 -255 5030 -235
rect 5060 -255 5080 -235
rect 5110 -255 5130 -235
rect 5160 -255 5180 -235
rect 5210 -255 5230 -235
rect 5260 -255 5280 -235
rect 5310 -255 5330 -235
rect 5360 -255 5380 -235
rect 5410 -255 5430 -235
rect 5460 -255 5480 -235
rect 5510 -255 5530 -235
rect 5560 -255 5580 -235
rect 5610 -255 5630 -235
rect 5660 -255 5680 -235
rect 5710 -255 5730 -235
rect 5760 -255 5780 -235
rect 5810 -255 5830 -235
rect 5860 -255 5880 -235
rect 5910 -255 5930 -235
rect 5960 -255 5980 -235
rect 6010 -255 6030 -235
rect 6060 -255 6080 -235
rect 6110 -255 6130 -235
rect 6160 -255 6180 -235
rect 6210 -255 6230 -235
rect 6260 -255 6280 -235
rect 6310 -255 6330 -235
rect 6360 -255 6380 -235
rect 6410 -255 6430 -235
rect 6460 -255 6480 -235
rect 6510 -255 6530 -235
rect 6560 -255 6580 -235
rect 6610 -255 6630 -235
rect 6660 -255 6680 -235
rect 6710 -255 6730 -235
rect 6760 -255 6780 -235
rect 6810 -255 6830 -235
rect 6860 -255 6880 -235
rect 6910 -255 6930 -235
<< metal1 >>
rect 2775 2820 2825 2830
rect 2775 2790 2785 2820
rect 2815 2790 2825 2820
rect 2775 2780 2825 2790
rect 2635 2595 2675 2600
rect 2635 2565 2640 2595
rect 2670 2580 2675 2595
rect 2670 2565 3005 2580
rect 2635 2560 2675 2565
rect 4820 2540 4860 2550
rect 5975 2545 6015 2550
rect 5975 2540 5980 2545
rect 4820 2520 4830 2540
rect 4850 2525 5980 2540
rect 4850 2520 4860 2525
rect 2580 2510 2620 2515
rect 4820 2510 4860 2520
rect 5975 2515 5980 2525
rect 6010 2515 6015 2545
rect 5975 2510 6015 2515
rect 2580 2480 2585 2510
rect 2615 2500 2620 2510
rect 2615 2485 3005 2500
rect 2615 2480 2620 2485
rect 2580 2475 2620 2480
rect 2775 2225 2825 2235
rect 2775 2195 2785 2225
rect 2815 2195 2825 2225
rect 2775 2185 2825 2195
rect 2690 1390 2730 1395
rect 2690 1360 2695 1390
rect 2725 1380 2730 1390
rect 5975 1385 6015 1390
rect 5975 1380 5980 1385
rect 2725 1365 5980 1380
rect 2725 1360 2730 1365
rect 2690 1355 2730 1360
rect 5975 1355 5980 1365
rect 6010 1355 6015 1385
rect 5975 1350 6015 1355
rect 2580 1335 2620 1340
rect 2580 1305 2585 1335
rect 2615 1325 2620 1335
rect 2615 1310 5480 1325
rect 2615 1305 2620 1310
rect 2580 1300 2620 1305
rect 2540 1280 2580 1285
rect 2540 1250 2545 1280
rect 2575 1275 2580 1280
rect 2575 1260 2805 1275
rect 2575 1250 2580 1260
rect 2540 1245 2580 1250
rect 2380 1220 2430 1230
rect 2355 1190 2390 1220
rect 2420 1190 2430 1220
rect 2355 1180 2430 1190
rect 2040 1155 2080 1165
rect 2040 1135 2050 1155
rect 2070 1150 2080 1155
rect 2580 1160 2620 1165
rect 2580 1150 2585 1160
rect 2070 1135 2585 1150
rect 2040 1125 2080 1135
rect 2580 1130 2585 1135
rect 2615 1130 2620 1160
rect 2580 1125 2620 1130
rect 2180 1095 2220 1100
rect 2180 1065 2185 1095
rect 2215 1085 2220 1095
rect 2535 1095 2575 1100
rect 2535 1085 2540 1095
rect 2215 1070 2540 1085
rect 2215 1065 2220 1070
rect 2180 1060 2220 1065
rect 2535 1065 2540 1070
rect 2570 1065 2575 1095
rect 2535 1060 2575 1065
rect 2735 1020 2785 1030
rect 2735 990 2745 1020
rect 2775 990 2785 1020
rect 2735 980 2785 990
rect 2180 950 2220 955
rect 2180 920 2185 950
rect 2215 920 2220 950
rect 2180 915 2220 920
rect 2300 945 2340 955
rect 2300 925 2310 945
rect 2330 940 2340 945
rect 2535 950 2575 955
rect 2535 940 2540 950
rect 2330 925 2540 940
rect 2300 915 2340 925
rect 2535 920 2540 925
rect 2570 920 2575 950
rect 2535 915 2575 920
rect 2580 695 2620 700
rect 2580 665 2585 695
rect 2615 685 2620 695
rect 2690 695 2730 700
rect 2690 685 2695 695
rect 2615 670 2695 685
rect 2615 665 2620 670
rect 2580 660 2620 665
rect 2690 665 2695 670
rect 2725 675 2730 695
rect 3090 680 3130 690
rect 3090 675 3100 680
rect 2725 665 3100 675
rect 2690 660 3100 665
rect 3120 660 3130 680
rect 2635 650 2675 655
rect 3090 650 3130 660
rect 3850 685 3890 690
rect 3850 655 3855 685
rect 3885 655 3890 685
rect -190 630 -140 635
rect 2460 630 2510 640
rect -190 625 -115 630
rect -190 595 -180 625
rect -150 595 -115 625
rect 2355 620 2470 630
rect 2370 600 2400 620
rect 2420 600 2470 620
rect 2500 600 2510 630
rect 2635 620 2640 650
rect 2670 635 2675 650
rect 3155 645 3195 655
rect 3850 650 3890 655
rect 3155 635 3165 645
rect 2670 625 3165 635
rect 3185 625 3195 645
rect 2670 620 3195 625
rect 2635 615 2675 620
rect 3155 615 3195 620
rect 3850 615 3890 620
rect -190 590 -115 595
rect 2355 590 2510 600
rect 2535 610 2575 615
rect -190 585 -140 590
rect 2535 580 2540 610
rect 2570 600 2575 610
rect 3850 600 3855 615
rect 2570 585 3855 600
rect 3885 585 3890 615
rect 2570 580 2575 585
rect 3850 580 3890 585
rect 4450 595 4490 605
rect 2535 575 2575 580
rect 4450 575 4460 595
rect 4480 590 4490 595
rect 5465 590 5480 1310
rect 4480 575 5480 590
rect 4450 565 4490 575
rect 2180 550 2220 560
rect 2180 530 2190 550
rect 2210 535 2220 550
rect 3055 540 3095 550
rect 3055 535 3065 540
rect 2210 530 3065 535
rect 2180 520 3065 530
rect 3085 520 3095 540
rect 3055 510 3095 520
rect 2535 495 2575 500
rect 2535 465 2540 495
rect 2570 490 2575 495
rect 4070 490 4110 500
rect 2570 475 4080 490
rect 2570 465 2575 475
rect 2535 460 2575 465
rect 4070 470 4080 475
rect 4100 470 4110 490
rect 4070 460 4110 470
rect 2305 275 2345 285
rect -130 260 -90 270
rect -130 240 -120 260
rect -100 240 -90 260
rect 2305 255 2315 275
rect 2335 270 2345 275
rect 2535 280 2575 285
rect 2535 270 2540 280
rect 2335 255 2540 270
rect 2305 245 2345 255
rect 2535 250 2540 255
rect 2570 250 2575 280
rect 2535 245 2575 250
rect -130 230 -90 240
rect 2735 170 2785 180
rect 2735 140 2745 170
rect 2775 140 2785 170
rect 2735 130 2785 140
rect 2075 85 2115 95
rect 2075 65 2085 85
rect 2105 70 2740 85
rect 2105 65 2115 70
rect 2075 55 2115 65
rect 2355 30 2430 40
rect 2355 0 2390 30
rect 2420 0 2430 30
rect 2380 -10 2430 0
rect 5465 -15 5480 575
rect 5465 -30 6610 -15
rect 2380 -225 2430 -215
rect 2380 -255 2390 -225
rect 2420 -235 6970 -225
rect 2420 -255 2460 -235
rect 2480 -255 2510 -235
rect 2530 -255 2560 -235
rect 2580 -255 2610 -235
rect 2630 -255 2660 -235
rect 2680 -255 2710 -235
rect 2730 -255 2760 -235
rect 2780 -255 2810 -235
rect 2830 -255 2860 -235
rect 2880 -255 2910 -235
rect 2930 -255 2960 -235
rect 2980 -255 3010 -235
rect 3030 -255 3060 -235
rect 3080 -255 3110 -235
rect 3130 -255 3160 -235
rect 3180 -255 3210 -235
rect 3230 -255 3260 -235
rect 3280 -255 3310 -235
rect 3330 -255 3360 -235
rect 3380 -255 3410 -235
rect 3430 -255 3460 -235
rect 3480 -255 3510 -235
rect 3530 -255 3560 -235
rect 3580 -255 3610 -235
rect 3630 -255 3660 -235
rect 3680 -255 3710 -235
rect 3730 -255 3760 -235
rect 3780 -255 3810 -235
rect 3830 -255 3860 -235
rect 3880 -255 3910 -235
rect 3930 -255 3960 -235
rect 3980 -255 4010 -235
rect 4030 -255 4060 -235
rect 4080 -255 4110 -235
rect 4130 -255 4160 -235
rect 4180 -255 4210 -235
rect 4230 -255 4260 -235
rect 4280 -255 4310 -235
rect 4330 -255 4360 -235
rect 4380 -255 4410 -235
rect 4430 -255 4460 -235
rect 4480 -255 4510 -235
rect 4530 -255 4560 -235
rect 4580 -255 4610 -235
rect 4630 -255 4660 -235
rect 4680 -255 4710 -235
rect 4730 -255 4760 -235
rect 4780 -255 4810 -235
rect 4830 -255 4860 -235
rect 4880 -255 4910 -235
rect 4930 -255 4960 -235
rect 4980 -255 5010 -235
rect 5030 -255 5060 -235
rect 5080 -255 5110 -235
rect 5130 -255 5160 -235
rect 5180 -255 5210 -235
rect 5230 -255 5260 -235
rect 5280 -255 5310 -235
rect 5330 -255 5360 -235
rect 5380 -255 5410 -235
rect 5430 -255 5460 -235
rect 5480 -255 5510 -235
rect 5530 -255 5560 -235
rect 5580 -255 5610 -235
rect 5630 -255 5660 -235
rect 5680 -255 5710 -235
rect 5730 -255 5760 -235
rect 5780 -255 5810 -235
rect 5830 -255 5860 -235
rect 5880 -255 5910 -235
rect 5930 -255 5960 -235
rect 5980 -255 6010 -235
rect 6030 -255 6060 -235
rect 6080 -255 6110 -235
rect 6130 -255 6160 -235
rect 6180 -255 6210 -235
rect 6230 -255 6260 -235
rect 6280 -255 6310 -235
rect 6330 -255 6360 -235
rect 6380 -255 6410 -235
rect 6430 -255 6460 -235
rect 6480 -255 6510 -235
rect 6530 -255 6560 -235
rect 6580 -255 6610 -235
rect 6630 -255 6660 -235
rect 6680 -255 6710 -235
rect 6730 -255 6760 -235
rect 6780 -255 6810 -235
rect 6830 -255 6860 -235
rect 6880 -255 6910 -235
rect 6930 -255 6970 -235
rect 2380 -265 6970 -255
<< via1 >>
rect 2785 2815 2815 2820
rect 2785 2795 2790 2815
rect 2790 2795 2810 2815
rect 2810 2795 2815 2815
rect 2785 2790 2815 2795
rect 2640 2565 2670 2595
rect 5980 2515 6010 2545
rect 2585 2480 2615 2510
rect 2785 2220 2815 2225
rect 2785 2200 2790 2220
rect 2790 2200 2810 2220
rect 2810 2200 2815 2220
rect 2785 2195 2815 2200
rect 2695 1360 2725 1390
rect 5980 1355 6010 1385
rect 2585 1305 2615 1335
rect 2545 1250 2575 1280
rect 2390 1190 2420 1220
rect 2585 1130 2615 1160
rect 2185 1065 2215 1095
rect 2540 1065 2570 1095
rect 2745 1015 2775 1020
rect 2745 995 2750 1015
rect 2750 995 2770 1015
rect 2770 995 2775 1015
rect 2745 990 2775 995
rect 2185 945 2215 950
rect 2185 925 2190 945
rect 2190 925 2210 945
rect 2210 925 2215 945
rect 2185 920 2215 925
rect 2540 920 2570 950
rect 2585 665 2615 695
rect 2695 665 2725 695
rect 3855 680 3885 685
rect 3855 660 3860 680
rect 3860 660 3880 680
rect 3880 660 3885 680
rect 3855 655 3885 660
rect -180 595 -150 625
rect 2470 625 2500 630
rect 2470 605 2475 625
rect 2475 605 2495 625
rect 2495 605 2500 625
rect 2470 600 2500 605
rect 2640 620 2670 650
rect 2540 580 2570 610
rect 3855 585 3885 615
rect 2540 465 2570 495
rect 2540 250 2570 280
rect 2745 165 2775 170
rect 2745 145 2750 165
rect 2750 145 2770 165
rect 2770 145 2775 165
rect 2745 140 2775 145
rect 2390 0 2420 30
rect 2390 -255 2420 -225
<< metal2 >>
rect 2775 2820 2825 2830
rect 2775 2790 2785 2820
rect 2815 2790 2825 2820
rect 2775 2780 2825 2790
rect 2635 2595 2675 2600
rect 2635 2565 2640 2595
rect 2670 2565 2675 2595
rect 2635 2560 2675 2565
rect 2580 2510 2620 2515
rect 2580 2480 2585 2510
rect 2615 2480 2620 2510
rect 2580 2475 2620 2480
rect 2590 1340 2605 2475
rect 2580 1335 2620 1340
rect 2580 1305 2585 1335
rect 2615 1305 2620 1335
rect 2580 1300 2620 1305
rect 2540 1280 2580 1285
rect 2540 1250 2545 1280
rect 2575 1250 2580 1280
rect 2540 1245 2580 1250
rect 2380 1220 2430 1230
rect 2380 1190 2390 1220
rect 2420 1190 2430 1220
rect 2380 1180 2430 1190
rect 2550 1100 2565 1245
rect 2580 1160 2620 1165
rect 2580 1130 2585 1160
rect 2615 1130 2620 1160
rect 2580 1125 2620 1130
rect 2180 1095 2220 1100
rect 2180 1065 2185 1095
rect 2215 1065 2220 1095
rect 2180 1060 2220 1065
rect 2535 1095 2575 1100
rect 2535 1065 2540 1095
rect 2570 1065 2575 1095
rect 2535 1060 2575 1065
rect 2195 955 2210 1060
rect 2180 950 2220 955
rect 2180 920 2185 950
rect 2215 920 2220 950
rect 2180 915 2220 920
rect 2535 950 2575 955
rect 2535 920 2540 950
rect 2570 920 2575 950
rect 2535 915 2575 920
rect -190 625 -140 635
rect -190 595 -180 625
rect -150 595 -140 625
rect -190 585 -140 595
rect 2460 630 2510 640
rect 2460 600 2470 630
rect 2500 600 2510 630
rect 2550 615 2565 915
rect 2590 700 2605 1125
rect 2580 695 2620 700
rect 2580 665 2585 695
rect 2615 665 2620 695
rect 2580 660 2620 665
rect 2650 655 2665 2560
rect 5975 2545 6015 2550
rect 5975 2515 5980 2545
rect 6010 2515 6015 2545
rect 5975 2510 6015 2515
rect 2775 2225 2825 2235
rect 2775 2195 2785 2225
rect 2815 2195 2825 2225
rect 2775 2185 2825 2195
rect 2690 1390 2730 1395
rect 5985 1390 6000 2510
rect 2690 1360 2695 1390
rect 2725 1360 2730 1390
rect 2690 1355 2730 1360
rect 5975 1385 6015 1390
rect 5975 1355 5980 1385
rect 6010 1355 6015 1385
rect 2705 700 2720 1355
rect 5975 1350 6015 1355
rect 2735 1020 2785 1030
rect 2735 990 2745 1020
rect 2775 990 2785 1020
rect 2735 980 2785 990
rect 2690 695 2730 700
rect 2690 665 2695 695
rect 2725 665 2730 695
rect 2690 660 2730 665
rect 3850 685 3890 690
rect 3850 655 3855 685
rect 3885 655 3890 685
rect 2635 650 2675 655
rect 3850 650 3890 655
rect 2635 620 2640 650
rect 2670 620 2675 650
rect 3860 620 3875 650
rect 2635 615 2675 620
rect 3850 615 3890 620
rect 2460 590 2510 600
rect 2535 610 2575 615
rect 2535 580 2540 610
rect 2570 580 2575 610
rect 3850 585 3855 615
rect 3885 585 3890 615
rect 3850 580 3890 585
rect 2535 575 2575 580
rect 2535 495 2575 500
rect 2535 465 2540 495
rect 2570 465 2575 495
rect 2535 460 2575 465
rect 2550 285 2565 460
rect 2535 280 2575 285
rect 2535 250 2540 280
rect 2570 250 2575 280
rect 2535 245 2575 250
rect 2735 170 2785 180
rect 2735 140 2745 170
rect 2775 140 2785 170
rect 2735 130 2785 140
rect 2380 30 2430 40
rect 2380 0 2390 30
rect 2420 0 2430 30
rect 2380 -10 2430 0
rect 2380 -225 2430 -215
rect 2380 -255 2390 -225
rect 2420 -255 2430 -225
rect 2380 -265 2430 -255
<< via2 >>
rect 2785 2790 2815 2820
rect 2390 1190 2420 1220
rect -180 595 -150 625
rect 2470 600 2500 630
rect 2785 2195 2815 2225
rect 2745 990 2775 1020
rect 2745 140 2775 170
rect 2390 0 2420 30
rect 2390 -255 2420 -225
<< metal3 >>
rect 2380 2825 2825 2830
rect 2380 2785 2385 2825
rect 2425 2820 2825 2825
rect 2425 2790 2785 2820
rect 2815 2790 2825 2820
rect 2425 2785 2825 2790
rect 2380 2780 2825 2785
rect 2460 2230 2825 2235
rect 2460 2190 2465 2230
rect 2505 2225 2825 2230
rect 2505 2195 2785 2225
rect 2815 2195 2825 2225
rect 2505 2190 2825 2195
rect 2460 2185 2825 2190
rect 2380 1225 2430 1230
rect 2380 1185 2385 1225
rect 2425 1185 2430 1225
rect 2380 1180 2430 1185
rect 2460 1025 2785 1030
rect 2460 985 2465 1025
rect 2505 1020 2785 1025
rect 2505 990 2745 1020
rect 2775 990 2785 1020
rect 2505 985 2785 990
rect 2460 980 2785 985
rect 2460 635 2510 640
rect -280 625 -140 635
rect -280 595 -180 625
rect -150 595 -140 625
rect -280 585 -140 595
rect 2460 595 2465 635
rect 2505 595 2510 635
rect 2460 590 2510 595
rect 2380 175 2785 180
rect 2380 135 2385 175
rect 2425 170 2785 175
rect 2425 140 2745 170
rect 2775 140 2785 170
rect 2425 135 2785 140
rect 2380 130 2785 135
rect 2380 35 2430 40
rect 2380 -5 2385 35
rect 2425 -5 2430 35
rect 2380 -10 2430 -5
rect 2380 -220 2430 -215
rect 2380 -260 2385 -220
rect 2425 -260 2430 -220
rect 2380 -265 2430 -260
<< via3 >>
rect 2385 2785 2425 2825
rect 2465 2190 2505 2230
rect 2385 1220 2425 1225
rect 2385 1190 2390 1220
rect 2390 1190 2420 1220
rect 2420 1190 2425 1220
rect 2385 1185 2425 1190
rect 2465 985 2505 1025
rect 2465 630 2505 635
rect 2465 600 2470 630
rect 2470 600 2500 630
rect 2500 600 2505 630
rect 2465 595 2505 600
rect 2385 135 2425 175
rect 2385 30 2425 35
rect 2385 0 2390 30
rect 2390 0 2420 30
rect 2420 0 2425 30
rect 2385 -5 2425 0
rect 2385 -225 2425 -220
rect 2385 -255 2390 -225
rect 2390 -255 2420 -225
rect 2420 -255 2425 -225
rect 2385 -260 2425 -255
<< metal4 >>
rect 2380 2825 2430 2830
rect 2380 2785 2385 2825
rect 2425 2785 2430 2825
rect 2380 1225 2430 2785
rect 2380 1185 2385 1225
rect 2425 1185 2430 1225
rect 2380 175 2430 1185
rect 2460 2230 2510 2235
rect 2460 2190 2465 2230
rect 2505 2190 2510 2230
rect 2460 1025 2510 2190
rect 2460 985 2465 1025
rect 2505 985 2510 1025
rect 2460 635 2510 985
rect 2460 595 2465 635
rect 2505 595 2510 635
rect 2460 590 2510 595
rect -280 105 -230 155
rect 2380 135 2385 175
rect 2425 135 2430 175
rect 2380 35 2430 135
rect 2380 -5 2385 35
rect 2425 -5 2430 35
rect 2380 -220 2430 -5
rect 2380 -260 2385 -220
rect 2425 -260 2430 -220
rect 2380 -265 2430 -260
use charge_pump_cell_6  charge_pump_cell_6_0
timestamp 1740147043
transform 1 0 -6370 0 1 -1565
box 9105 1615 11810 2860
use loop_filter_2  loop_filter_2_0
timestamp 1740116583
transform 1 0 4330 0 1 -345
box 1135 -5975 9720 330
use opamp_cell_4  opamp_cell_4_0
timestamp 1740145811
transform 1 0 -425 0 -1 4625
box 3110 897 6365 3205
use pfd_8  pfd_8_0
timestamp 1739770731
transform 1 0 -930 0 1 4655
box 650 -4655 3290 -3435
<< labels >>
flabel metal1 -140 610 -140 610 7 FreeSans 400 0 -200 0 VDDA
port 2 w
flabel poly -130 250 -130 250 7 FreeSans 400 0 -200 0 F_VCO
port 5 w
flabel poly -130 965 -130 965 7 FreeSans 400 0 -200 0 F_REF
port 4 w
flabel metal1 5480 585 5480 585 3 FreeSans 400 0 200 0 V_OUT
port 1 e
flabel metal4 -280 130 -280 130 7 FreeSans 400 0 -200 0 GNDA
port 3 w
flabel metal1 2800 535 2800 535 1 FreeSans 400 0 0 200 I_IN
port 6 n
<< end >>
