magic
tech sky130A
timestamp 1737896025
<< nmos >>
rect 1070 445 1120 695
rect 1170 445 1220 695
rect 1270 445 1320 695
rect 1370 445 1420 695
rect 1470 445 1520 695
rect 1570 445 1620 695
rect 1670 445 1720 695
rect 1770 445 1820 695
rect 1055 245 1070 345
rect 1120 245 1135 345
rect 1185 245 1200 345
rect 1250 245 1265 345
rect 1410 245 1425 345
rect 1475 245 1490 345
rect 1540 245 1555 345
rect 1605 245 1620 345
rect 1790 245 1805 345
rect 1855 245 1870 345
rect 1920 245 1935 345
rect 1985 245 2000 345
rect 1055 90 1070 140
rect 1120 90 1135 140
rect 1185 90 1200 140
rect 1250 90 1265 140
rect 1410 90 1425 140
rect 1475 90 1490 140
rect 1540 90 1555 140
rect 1605 90 1620 140
rect 1790 90 1805 140
rect 1855 90 1870 140
rect 1920 90 1935 140
rect 1985 90 2000 140
rect 1615 -260 1665 -10
rect 1715 -260 1765 -10
rect 1815 -260 1865 -10
rect 1915 -260 1965 -10
<< ndiff >>
rect 1020 680 1070 695
rect 1020 460 1035 680
rect 1055 460 1070 680
rect 1020 445 1070 460
rect 1120 680 1170 695
rect 1120 460 1135 680
rect 1155 460 1170 680
rect 1120 445 1170 460
rect 1220 680 1270 695
rect 1220 460 1235 680
rect 1255 460 1270 680
rect 1220 445 1270 460
rect 1320 680 1370 695
rect 1320 460 1335 680
rect 1355 460 1370 680
rect 1320 445 1370 460
rect 1420 680 1470 695
rect 1420 460 1435 680
rect 1455 460 1470 680
rect 1420 445 1470 460
rect 1520 680 1570 695
rect 1520 460 1535 680
rect 1555 460 1570 680
rect 1520 445 1570 460
rect 1620 680 1670 695
rect 1620 460 1635 680
rect 1655 460 1670 680
rect 1620 445 1670 460
rect 1720 680 1770 695
rect 1720 460 1735 680
rect 1755 460 1770 680
rect 1720 445 1770 460
rect 1820 680 1870 695
rect 1820 460 1835 680
rect 1855 460 1870 680
rect 1820 445 1870 460
rect 1005 330 1055 345
rect 1005 260 1020 330
rect 1040 260 1055 330
rect 1005 245 1055 260
rect 1070 330 1120 345
rect 1070 260 1085 330
rect 1105 260 1120 330
rect 1070 245 1120 260
rect 1135 330 1185 345
rect 1135 260 1150 330
rect 1170 260 1185 330
rect 1135 245 1185 260
rect 1200 330 1250 345
rect 1200 260 1215 330
rect 1235 260 1250 330
rect 1200 245 1250 260
rect 1265 330 1315 345
rect 1265 260 1280 330
rect 1300 260 1315 330
rect 1265 245 1315 260
rect 1360 330 1410 345
rect 1360 260 1375 330
rect 1395 260 1410 330
rect 1360 245 1410 260
rect 1425 330 1475 345
rect 1425 260 1440 330
rect 1460 260 1475 330
rect 1425 245 1475 260
rect 1490 330 1540 345
rect 1490 260 1505 330
rect 1525 260 1540 330
rect 1490 245 1540 260
rect 1555 330 1605 345
rect 1555 260 1570 330
rect 1590 260 1605 330
rect 1555 245 1605 260
rect 1620 330 1670 345
rect 1620 260 1635 330
rect 1655 260 1670 330
rect 1620 245 1670 260
rect 1740 330 1790 345
rect 1740 260 1755 330
rect 1775 260 1790 330
rect 1740 245 1790 260
rect 1805 330 1855 345
rect 1805 260 1820 330
rect 1840 260 1855 330
rect 1805 245 1855 260
rect 1870 330 1920 345
rect 1870 260 1885 330
rect 1905 260 1920 330
rect 1870 245 1920 260
rect 1935 330 1985 345
rect 1935 260 1950 330
rect 1970 260 1985 330
rect 1935 245 1985 260
rect 2000 330 2050 345
rect 2000 260 2015 330
rect 2035 260 2050 330
rect 2000 245 2050 260
rect 1005 125 1055 140
rect 1005 105 1020 125
rect 1040 105 1055 125
rect 1005 90 1055 105
rect 1070 125 1120 140
rect 1070 105 1085 125
rect 1105 105 1120 125
rect 1070 90 1120 105
rect 1135 125 1185 140
rect 1135 105 1150 125
rect 1170 105 1185 125
rect 1135 90 1185 105
rect 1200 125 1250 140
rect 1200 105 1215 125
rect 1235 105 1250 125
rect 1200 90 1250 105
rect 1265 125 1315 140
rect 1265 105 1280 125
rect 1300 105 1315 125
rect 1265 90 1315 105
rect 1360 125 1410 140
rect 1360 105 1375 125
rect 1395 105 1410 125
rect 1360 90 1410 105
rect 1425 125 1475 140
rect 1425 105 1440 125
rect 1460 105 1475 125
rect 1425 90 1475 105
rect 1490 125 1540 140
rect 1490 105 1505 125
rect 1525 105 1540 125
rect 1490 90 1540 105
rect 1555 125 1605 140
rect 1555 105 1570 125
rect 1590 105 1605 125
rect 1555 90 1605 105
rect 1620 125 1670 140
rect 1620 105 1635 125
rect 1655 105 1670 125
rect 1620 90 1670 105
rect 1740 125 1790 140
rect 1740 105 1755 125
rect 1775 105 1790 125
rect 1740 90 1790 105
rect 1805 125 1855 140
rect 1805 105 1820 125
rect 1840 105 1855 125
rect 1805 90 1855 105
rect 1870 125 1920 140
rect 1870 105 1885 125
rect 1905 105 1920 125
rect 1870 90 1920 105
rect 1935 125 1985 140
rect 1935 105 1950 125
rect 1970 105 1985 125
rect 1935 90 1985 105
rect 2000 125 2050 140
rect 2000 105 2015 125
rect 2035 105 2050 125
rect 2000 90 2050 105
rect 1565 -25 1615 -10
rect 1565 -245 1580 -25
rect 1600 -245 1615 -25
rect 1565 -260 1615 -245
rect 1665 -25 1715 -10
rect 1665 -245 1680 -25
rect 1700 -245 1715 -25
rect 1665 -260 1715 -245
rect 1765 -25 1815 -10
rect 1765 -245 1780 -25
rect 1800 -245 1815 -25
rect 1765 -260 1815 -245
rect 1865 -25 1915 -10
rect 1865 -245 1880 -25
rect 1900 -245 1915 -25
rect 1865 -260 1915 -245
rect 1965 -25 2015 -10
rect 1965 -245 1980 -25
rect 2000 -245 2015 -25
rect 1965 -260 2015 -245
<< ndiffc >>
rect 1035 460 1055 680
rect 1135 460 1155 680
rect 1235 460 1255 680
rect 1335 460 1355 680
rect 1435 460 1455 680
rect 1535 460 1555 680
rect 1635 460 1655 680
rect 1735 460 1755 680
rect 1835 460 1855 680
rect 1020 260 1040 330
rect 1085 260 1105 330
rect 1150 260 1170 330
rect 1215 260 1235 330
rect 1280 260 1300 330
rect 1375 260 1395 330
rect 1440 260 1460 330
rect 1505 260 1525 330
rect 1570 260 1590 330
rect 1635 260 1655 330
rect 1755 260 1775 330
rect 1820 260 1840 330
rect 1885 260 1905 330
rect 1950 260 1970 330
rect 2015 260 2035 330
rect 1020 105 1040 125
rect 1085 105 1105 125
rect 1150 105 1170 125
rect 1215 105 1235 125
rect 1280 105 1300 125
rect 1375 105 1395 125
rect 1440 105 1460 125
rect 1505 105 1525 125
rect 1570 105 1590 125
rect 1635 105 1655 125
rect 1755 105 1775 125
rect 1820 105 1840 125
rect 1885 105 1905 125
rect 1950 105 1970 125
rect 2015 105 2035 125
rect 1580 -245 1600 -25
rect 1680 -245 1700 -25
rect 1780 -245 1800 -25
rect 1880 -245 1900 -25
rect 1980 -245 2000 -25
<< poly >>
rect 1125 740 1165 750
rect 1125 725 1135 740
rect 1070 720 1135 725
rect 1155 725 1165 740
rect 1525 740 1565 750
rect 1525 725 1535 740
rect 1155 720 1535 725
rect 1555 725 1565 740
rect 1555 720 1820 725
rect 1070 710 1820 720
rect 1070 695 1120 710
rect 1170 695 1220 710
rect 1270 695 1320 710
rect 1370 695 1420 710
rect 1470 695 1520 710
rect 1570 695 1620 710
rect 1670 695 1720 710
rect 1770 695 1820 710
rect 1070 430 1120 445
rect 1170 430 1220 445
rect 1270 430 1320 445
rect 1370 430 1420 445
rect 1470 430 1520 445
rect 1570 430 1620 445
rect 1670 430 1720 445
rect 1770 430 1820 445
rect 860 385 1200 400
rect 1055 345 1070 360
rect 1120 345 1135 360
rect 1185 345 1200 385
rect 1250 345 1265 360
rect 1410 345 1425 360
rect 1475 345 1490 360
rect 1540 345 1555 360
rect 1605 345 1620 360
rect 1790 345 1805 360
rect 1855 345 1870 360
rect 1920 345 1935 360
rect 1985 345 2000 360
rect 1055 235 1070 245
rect 1120 235 1135 245
rect 980 220 1135 235
rect 1185 235 1200 245
rect 1250 235 1265 245
rect 1410 235 1425 245
rect 1475 235 1490 245
rect 1540 235 1555 245
rect 1605 235 1620 245
rect 1185 220 1350 235
rect 980 50 995 220
rect 1075 185 1115 195
rect 1075 165 1085 185
rect 1105 165 1115 185
rect 1335 165 1350 220
rect 1410 220 1620 235
rect 1410 215 1440 220
rect 1430 200 1440 215
rect 1460 215 1620 220
rect 1685 240 1725 250
rect 2065 250 2105 260
rect 1685 220 1695 240
rect 1715 235 1725 240
rect 1790 235 1805 245
rect 1855 235 1870 245
rect 1920 235 1935 245
rect 1985 235 2000 245
rect 2065 235 2075 250
rect 1715 230 2075 235
rect 2095 230 2105 250
rect 1715 220 2105 230
rect 1460 200 1470 215
rect 1685 210 1725 220
rect 1430 190 1470 200
rect 1685 175 1725 185
rect 1055 150 1265 165
rect 1335 150 1490 165
rect 1685 155 1695 175
rect 1715 165 1725 175
rect 1715 155 2105 165
rect 1055 140 1070 150
rect 1120 140 1135 150
rect 1185 140 1200 150
rect 1250 140 1265 150
rect 1410 140 1425 150
rect 1475 140 1490 150
rect 1540 140 1555 155
rect 1605 140 1620 155
rect 1685 150 2075 155
rect 1685 145 1725 150
rect 1790 140 1805 150
rect 1855 140 1870 150
rect 1920 140 1935 150
rect 1985 140 2000 150
rect 2065 135 2075 150
rect 2095 135 2105 155
rect 2065 125 2105 135
rect 1055 75 1070 90
rect 1120 75 1135 90
rect 1185 75 1200 90
rect 1250 75 1265 90
rect 1410 75 1425 90
rect 1475 75 1490 90
rect 1540 80 1555 90
rect 1605 80 1620 90
rect 1540 65 1620 80
rect 1790 75 1805 90
rect 1855 75 1870 90
rect 1920 75 1935 90
rect 1985 75 2000 90
rect 1540 50 1555 65
rect 865 35 1555 50
rect 1615 -10 1665 5
rect 1715 -10 1765 5
rect 1815 -10 1865 5
rect 1915 -10 1965 5
rect 1615 -275 1665 -260
rect 1715 -275 1765 -260
rect 1815 -275 1865 -260
rect 1915 -275 1965 -260
rect 1615 -285 1965 -275
rect 1615 -290 1680 -285
rect 1670 -305 1680 -290
rect 1700 -290 1965 -285
rect 1700 -305 1710 -290
rect 1670 -315 1710 -305
<< polycont >>
rect 1135 720 1155 740
rect 1535 720 1555 740
rect 1085 165 1105 185
rect 1440 200 1460 220
rect 1695 220 1715 240
rect 2075 230 2095 250
rect 1695 155 1715 175
rect 2075 135 2095 155
rect 1680 -305 1700 -285
<< xpolycontact >>
rect 2070 745 2105 965
rect 2070 410 2105 630
rect 1020 -305 1240 -20
rect 1290 -305 1510 -20
rect 2070 -190 2105 30
rect 2070 -495 2105 -275
<< xpolyres >>
rect 2070 630 2105 745
rect 1240 -305 1290 -20
rect 2070 -275 2105 -190
<< locali >>
rect 2125 1070 2165 1080
rect 2085 1050 2165 1070
rect 2085 965 2105 1050
rect 2125 1040 2165 1050
rect 1085 740 1165 750
rect 1085 730 1135 740
rect 1025 680 1065 690
rect 1025 460 1035 680
rect 1055 460 1065 680
rect 1025 450 1065 460
rect 1085 430 1105 730
rect 1125 720 1135 730
rect 1155 720 1165 740
rect 1125 710 1165 720
rect 1525 740 1565 750
rect 1525 720 1535 740
rect 1555 720 1565 740
rect 1525 710 1565 720
rect 1135 690 1155 710
rect 1535 690 1555 710
rect 1125 680 1165 690
rect 1125 460 1135 680
rect 1155 460 1165 680
rect 1125 450 1165 460
rect 1225 680 1265 690
rect 1225 460 1235 680
rect 1255 460 1265 680
rect 1225 450 1265 460
rect 1325 680 1365 690
rect 1325 460 1335 680
rect 1355 460 1365 680
rect 1325 450 1365 460
rect 1425 680 1465 690
rect 1425 460 1435 680
rect 1455 460 1465 680
rect 1425 450 1465 460
rect 1525 680 1565 690
rect 1525 460 1535 680
rect 1555 460 1565 680
rect 1525 450 1565 460
rect 1625 680 1665 690
rect 1625 460 1635 680
rect 1655 460 1665 680
rect 1625 450 1665 460
rect 1725 680 1765 690
rect 1725 460 1735 680
rect 1755 460 1765 680
rect 1725 450 1765 460
rect 1825 680 1865 690
rect 1825 460 1835 680
rect 1855 460 1865 680
rect 1825 450 1865 460
rect 970 410 1105 430
rect 1335 420 1355 450
rect 1735 420 1755 450
rect 970 -20 990 410
rect 1335 400 1755 420
rect 1280 380 1300 400
rect 2085 380 2105 410
rect 1020 360 1300 380
rect 1020 340 1040 360
rect 1150 340 1170 360
rect 1280 340 1300 360
rect 1820 360 2105 380
rect 1820 340 1840 360
rect 1950 340 1970 360
rect 1010 330 1050 340
rect 1010 260 1020 330
rect 1040 260 1050 330
rect 1010 250 1050 260
rect 1075 330 1115 340
rect 1075 260 1085 330
rect 1105 260 1115 330
rect 1075 250 1115 260
rect 1140 330 1180 340
rect 1140 260 1150 330
rect 1170 260 1180 330
rect 1140 250 1180 260
rect 1205 330 1245 340
rect 1205 260 1215 330
rect 1235 260 1245 330
rect 1205 250 1245 260
rect 1270 330 1310 340
rect 1270 260 1280 330
rect 1300 260 1310 330
rect 1270 250 1310 260
rect 1365 330 1405 340
rect 1365 260 1375 330
rect 1395 260 1405 330
rect 1365 250 1405 260
rect 1430 330 1470 340
rect 1430 260 1440 330
rect 1460 260 1470 330
rect 1430 250 1470 260
rect 1495 330 1535 340
rect 1495 260 1505 330
rect 1525 260 1535 330
rect 1495 250 1535 260
rect 1560 330 1600 340
rect 1560 260 1570 330
rect 1590 260 1600 330
rect 1560 250 1600 260
rect 1625 330 1665 340
rect 1625 260 1635 330
rect 1655 260 1665 330
rect 1625 250 1665 260
rect 1745 330 1785 340
rect 1745 260 1755 330
rect 1775 260 1785 330
rect 1745 250 1785 260
rect 1810 330 1850 340
rect 1810 260 1820 330
rect 1840 260 1850 330
rect 1810 250 1850 260
rect 1875 330 1915 340
rect 1875 260 1885 330
rect 1905 260 1915 330
rect 1875 250 1915 260
rect 1940 330 1980 340
rect 1940 260 1950 330
rect 1970 260 1980 330
rect 1940 250 1980 260
rect 2005 330 2045 340
rect 2005 260 2015 330
rect 2035 260 2045 330
rect 2085 260 2105 360
rect 2005 250 2045 260
rect 2065 250 2105 260
rect 1085 195 1105 250
rect 1215 205 1235 250
rect 1440 230 1460 250
rect 1570 230 1590 250
rect 1685 240 1725 250
rect 1685 230 1695 240
rect 1430 220 1470 230
rect 1215 195 1255 205
rect 1075 185 1115 195
rect 1075 165 1085 185
rect 1105 165 1115 185
rect 1075 155 1115 165
rect 1215 175 1225 195
rect 1245 175 1255 195
rect 1430 200 1440 220
rect 1460 200 1470 220
rect 1430 190 1470 200
rect 1570 220 1695 230
rect 1715 220 1725 240
rect 2065 230 2075 250
rect 2095 240 2105 250
rect 2125 275 2165 315
rect 2125 240 2145 275
rect 2095 230 3210 240
rect 2065 220 3210 230
rect 1570 210 1725 220
rect 1215 165 1255 175
rect 1085 135 1105 155
rect 1215 135 1235 165
rect 1440 135 1460 190
rect 1570 135 1590 210
rect 1685 175 1725 185
rect 1685 155 1695 175
rect 1715 155 1725 175
rect 1685 145 1725 155
rect 2065 155 3210 165
rect 2065 135 2075 155
rect 2095 145 3210 155
rect 2095 135 2105 145
rect 1010 125 1050 135
rect 1010 105 1020 125
rect 1040 105 1050 125
rect 1010 95 1050 105
rect 1075 125 1115 135
rect 1075 105 1085 125
rect 1105 105 1115 125
rect 1075 95 1115 105
rect 1140 125 1180 135
rect 1140 105 1150 125
rect 1170 105 1180 125
rect 1140 95 1180 105
rect 1205 125 1245 135
rect 1205 105 1215 125
rect 1235 105 1245 125
rect 1205 95 1245 105
rect 1270 125 1310 135
rect 1270 105 1280 125
rect 1300 105 1310 125
rect 1270 95 1310 105
rect 1365 125 1405 135
rect 1365 105 1375 125
rect 1395 105 1405 125
rect 1365 95 1405 105
rect 1430 125 1470 135
rect 1430 105 1440 125
rect 1460 105 1470 125
rect 1430 95 1470 105
rect 1495 125 1535 135
rect 1495 105 1505 125
rect 1525 105 1535 125
rect 1495 95 1535 105
rect 1560 125 1600 135
rect 1560 105 1570 125
rect 1590 105 1600 125
rect 1560 95 1600 105
rect 1625 125 1665 135
rect 1625 105 1635 125
rect 1655 105 1665 125
rect 1625 95 1665 105
rect 1745 125 1785 135
rect 1745 105 1755 125
rect 1775 105 1785 125
rect 1745 95 1785 105
rect 1810 125 1850 135
rect 1810 105 1820 125
rect 1840 105 1850 125
rect 1810 95 1850 105
rect 1875 125 1915 135
rect 1875 105 1885 125
rect 1905 105 1915 125
rect 1875 95 1915 105
rect 1940 125 1980 135
rect 1940 105 1950 125
rect 1970 105 1980 125
rect 1940 95 1980 105
rect 2005 125 2045 135
rect 2065 125 2105 135
rect 2005 105 2015 125
rect 2035 105 2045 125
rect 2005 95 2045 105
rect 1020 75 1040 95
rect 1150 75 1170 95
rect 1280 75 1300 95
rect 1020 55 1300 75
rect 1375 75 1395 95
rect 1505 75 1525 95
rect 1635 75 1655 95
rect 1820 75 1840 95
rect 1950 75 1970 95
rect 2085 75 2105 125
rect 1375 55 1700 75
rect 1820 55 2105 75
rect 2125 110 2145 145
rect 2125 70 2165 110
rect 1680 35 1700 55
rect 1680 15 1900 35
rect 2085 30 2105 55
rect 1880 -15 1900 15
rect 970 -40 1020 -20
rect 1570 -25 1610 -15
rect 1570 -245 1580 -25
rect 1600 -245 1610 -25
rect 1570 -255 1610 -245
rect 1670 -25 1710 -15
rect 1670 -245 1680 -25
rect 1700 -245 1710 -25
rect 1670 -255 1710 -245
rect 1770 -25 1810 -15
rect 1770 -245 1780 -25
rect 1800 -245 1810 -25
rect 1770 -255 1810 -245
rect 1870 -25 1910 -15
rect 1870 -245 1880 -25
rect 1900 -245 1910 -25
rect 1870 -255 1910 -245
rect 1970 -25 2010 -15
rect 1970 -245 1980 -25
rect 2000 -245 2010 -25
rect 1970 -255 2010 -245
rect 1680 -275 1700 -255
rect 1670 -285 1710 -275
rect 1510 -305 1680 -285
rect 1700 -305 1710 -285
rect 1670 -315 1710 -305
rect 2085 -665 2105 -495
rect 2125 -665 2165 -655
rect 2085 -685 2165 -665
rect 2125 -695 2165 -685
<< viali >>
rect 1225 175 1245 195
rect 1695 155 1715 175
<< metal1 >>
rect 1215 195 1255 205
rect 1215 175 1225 195
rect 1245 185 1255 195
rect 1245 175 1725 185
rect 1215 165 1695 175
rect 1685 155 1695 165
rect 1715 155 1725 175
rect 1685 145 1725 155
<< metal3 >>
rect 2125 1040 3010 1085
rect 2180 255 3010 1040
rect 2180 -655 3010 130
rect 2125 -700 3010 -655
<< mimcap >>
rect 2195 315 2995 1070
rect 2195 280 2205 315
rect 2240 280 2995 315
rect 2195 270 2995 280
rect 2195 105 2995 115
rect 2195 70 2205 105
rect 2240 70 2995 105
rect 2195 -685 2995 70
<< mimcapcontact >>
rect 2205 280 2240 315
rect 2205 70 2240 105
<< metal4 >>
rect 2125 315 2245 320
rect 2125 280 2205 315
rect 2240 280 2245 315
rect 2125 275 2245 280
rect 2125 105 2245 110
rect 2125 70 2205 105
rect 2240 70 2245 105
rect 2125 65 2245 70
<< end >>
