magic
tech sky130A
timestamp 1756257297
<< nwell >>
rect 9230 2215 10840 2505
<< nmos >>
rect 9250 1795 9310 1995
rect 9360 1795 9420 1995
rect 9470 1795 9530 1995
rect 9580 1795 9640 1995
rect 9790 1795 9850 1995
rect 9900 1795 9960 1995
rect 10010 1795 10070 1995
rect 10120 1795 10180 1995
rect 10330 1795 10390 1995
rect 10440 1795 10500 1995
rect 10550 1795 10610 1995
rect 10660 1795 10720 1995
<< pmos >>
rect 9350 2285 9410 2485
rect 9460 2285 9520 2485
rect 9570 2285 9630 2485
rect 9680 2285 9740 2485
rect 9790 2285 9850 2485
rect 9900 2285 9960 2485
rect 10110 2285 10170 2485
rect 10220 2285 10280 2485
rect 10330 2285 10390 2485
rect 10440 2285 10500 2485
rect 10550 2285 10610 2485
rect 10660 2285 10720 2485
<< ndiff >>
rect 9200 1980 9250 1995
rect 9200 1960 9215 1980
rect 9235 1960 9250 1980
rect 9200 1930 9250 1960
rect 9200 1910 9215 1930
rect 9235 1910 9250 1930
rect 9200 1880 9250 1910
rect 9200 1860 9215 1880
rect 9235 1860 9250 1880
rect 9200 1830 9250 1860
rect 9200 1810 9215 1830
rect 9235 1810 9250 1830
rect 9200 1795 9250 1810
rect 9310 1980 9360 1995
rect 9310 1960 9325 1980
rect 9345 1960 9360 1980
rect 9310 1930 9360 1960
rect 9310 1910 9325 1930
rect 9345 1910 9360 1930
rect 9310 1880 9360 1910
rect 9310 1860 9325 1880
rect 9345 1860 9360 1880
rect 9310 1830 9360 1860
rect 9310 1810 9325 1830
rect 9345 1810 9360 1830
rect 9310 1795 9360 1810
rect 9420 1980 9470 1995
rect 9420 1960 9435 1980
rect 9455 1960 9470 1980
rect 9420 1930 9470 1960
rect 9420 1910 9435 1930
rect 9455 1910 9470 1930
rect 9420 1880 9470 1910
rect 9420 1860 9435 1880
rect 9455 1860 9470 1880
rect 9420 1830 9470 1860
rect 9420 1810 9435 1830
rect 9455 1810 9470 1830
rect 9420 1795 9470 1810
rect 9530 1980 9580 1995
rect 9530 1960 9545 1980
rect 9565 1960 9580 1980
rect 9530 1930 9580 1960
rect 9530 1910 9545 1930
rect 9565 1910 9580 1930
rect 9530 1880 9580 1910
rect 9530 1860 9545 1880
rect 9565 1860 9580 1880
rect 9530 1830 9580 1860
rect 9530 1810 9545 1830
rect 9565 1810 9580 1830
rect 9530 1795 9580 1810
rect 9640 1980 9690 1995
rect 9740 1980 9790 1995
rect 9640 1960 9655 1980
rect 9675 1960 9690 1980
rect 9740 1960 9755 1980
rect 9775 1960 9790 1980
rect 9640 1930 9690 1960
rect 9740 1930 9790 1960
rect 9640 1910 9655 1930
rect 9675 1910 9690 1930
rect 9740 1910 9755 1930
rect 9775 1910 9790 1930
rect 9640 1880 9690 1910
rect 9740 1880 9790 1910
rect 9640 1860 9655 1880
rect 9675 1860 9690 1880
rect 9740 1860 9755 1880
rect 9775 1860 9790 1880
rect 9640 1830 9690 1860
rect 9740 1830 9790 1860
rect 9640 1810 9655 1830
rect 9675 1810 9690 1830
rect 9740 1810 9755 1830
rect 9775 1810 9790 1830
rect 9640 1795 9690 1810
rect 9740 1795 9790 1810
rect 9850 1980 9900 1995
rect 9850 1960 9865 1980
rect 9885 1960 9900 1980
rect 9850 1930 9900 1960
rect 9850 1910 9865 1930
rect 9885 1910 9900 1930
rect 9850 1880 9900 1910
rect 9850 1860 9865 1880
rect 9885 1860 9900 1880
rect 9850 1830 9900 1860
rect 9850 1810 9865 1830
rect 9885 1810 9900 1830
rect 9850 1795 9900 1810
rect 9960 1980 10010 1995
rect 9960 1960 9975 1980
rect 9995 1960 10010 1980
rect 9960 1930 10010 1960
rect 9960 1910 9975 1930
rect 9995 1910 10010 1930
rect 9960 1880 10010 1910
rect 9960 1860 9975 1880
rect 9995 1860 10010 1880
rect 9960 1830 10010 1860
rect 9960 1810 9975 1830
rect 9995 1810 10010 1830
rect 9960 1795 10010 1810
rect 10070 1980 10120 1995
rect 10070 1960 10085 1980
rect 10105 1960 10120 1980
rect 10070 1930 10120 1960
rect 10070 1910 10085 1930
rect 10105 1910 10120 1930
rect 10070 1880 10120 1910
rect 10070 1860 10085 1880
rect 10105 1860 10120 1880
rect 10070 1830 10120 1860
rect 10070 1810 10085 1830
rect 10105 1810 10120 1830
rect 10070 1795 10120 1810
rect 10180 1980 10230 1995
rect 10280 1980 10330 1995
rect 10180 1960 10195 1980
rect 10215 1960 10230 1980
rect 10280 1960 10295 1980
rect 10315 1960 10330 1980
rect 10180 1930 10230 1960
rect 10280 1930 10330 1960
rect 10180 1910 10195 1930
rect 10215 1910 10230 1930
rect 10280 1910 10295 1930
rect 10315 1910 10330 1930
rect 10180 1880 10230 1910
rect 10280 1880 10330 1910
rect 10180 1860 10195 1880
rect 10215 1860 10230 1880
rect 10280 1860 10295 1880
rect 10315 1860 10330 1880
rect 10180 1830 10230 1860
rect 10280 1830 10330 1860
rect 10180 1810 10195 1830
rect 10215 1810 10230 1830
rect 10280 1810 10295 1830
rect 10315 1810 10330 1830
rect 10180 1795 10230 1810
rect 10280 1795 10330 1810
rect 10390 1980 10440 1995
rect 10390 1960 10405 1980
rect 10425 1960 10440 1980
rect 10390 1930 10440 1960
rect 10390 1910 10405 1930
rect 10425 1910 10440 1930
rect 10390 1880 10440 1910
rect 10390 1860 10405 1880
rect 10425 1860 10440 1880
rect 10390 1830 10440 1860
rect 10390 1810 10405 1830
rect 10425 1810 10440 1830
rect 10390 1795 10440 1810
rect 10500 1980 10550 1995
rect 10500 1960 10515 1980
rect 10535 1960 10550 1980
rect 10500 1930 10550 1960
rect 10500 1910 10515 1930
rect 10535 1910 10550 1930
rect 10500 1880 10550 1910
rect 10500 1860 10515 1880
rect 10535 1860 10550 1880
rect 10500 1830 10550 1860
rect 10500 1810 10515 1830
rect 10535 1810 10550 1830
rect 10500 1795 10550 1810
rect 10610 1980 10660 1995
rect 10610 1960 10625 1980
rect 10645 1960 10660 1980
rect 10610 1930 10660 1960
rect 10610 1910 10625 1930
rect 10645 1910 10660 1930
rect 10610 1880 10660 1910
rect 10610 1860 10625 1880
rect 10645 1860 10660 1880
rect 10610 1830 10660 1860
rect 10610 1810 10625 1830
rect 10645 1810 10660 1830
rect 10610 1795 10660 1810
rect 10720 1980 10770 1995
rect 10720 1960 10735 1980
rect 10755 1960 10770 1980
rect 10720 1930 10770 1960
rect 10720 1910 10735 1930
rect 10755 1910 10770 1930
rect 10720 1880 10770 1910
rect 10720 1860 10735 1880
rect 10755 1860 10770 1880
rect 10720 1830 10770 1860
rect 10720 1810 10735 1830
rect 10755 1810 10770 1830
rect 10720 1795 10770 1810
<< pdiff >>
rect 9300 2470 9350 2485
rect 9300 2450 9315 2470
rect 9335 2450 9350 2470
rect 9300 2420 9350 2450
rect 9300 2400 9315 2420
rect 9335 2400 9350 2420
rect 9300 2370 9350 2400
rect 9300 2350 9315 2370
rect 9335 2350 9350 2370
rect 9300 2320 9350 2350
rect 9300 2300 9315 2320
rect 9335 2300 9350 2320
rect 9300 2285 9350 2300
rect 9410 2470 9460 2485
rect 9410 2450 9425 2470
rect 9445 2450 9460 2470
rect 9410 2420 9460 2450
rect 9410 2400 9425 2420
rect 9445 2400 9460 2420
rect 9410 2370 9460 2400
rect 9410 2350 9425 2370
rect 9445 2350 9460 2370
rect 9410 2320 9460 2350
rect 9410 2300 9425 2320
rect 9445 2300 9460 2320
rect 9410 2285 9460 2300
rect 9520 2470 9570 2485
rect 9520 2450 9535 2470
rect 9555 2450 9570 2470
rect 9520 2420 9570 2450
rect 9520 2400 9535 2420
rect 9555 2400 9570 2420
rect 9520 2370 9570 2400
rect 9520 2350 9535 2370
rect 9555 2350 9570 2370
rect 9520 2320 9570 2350
rect 9520 2300 9535 2320
rect 9555 2300 9570 2320
rect 9520 2285 9570 2300
rect 9630 2470 9680 2485
rect 9630 2450 9645 2470
rect 9665 2450 9680 2470
rect 9630 2420 9680 2450
rect 9630 2400 9645 2420
rect 9665 2400 9680 2420
rect 9630 2370 9680 2400
rect 9630 2350 9645 2370
rect 9665 2350 9680 2370
rect 9630 2320 9680 2350
rect 9630 2300 9645 2320
rect 9665 2300 9680 2320
rect 9630 2285 9680 2300
rect 9740 2470 9790 2485
rect 9740 2450 9755 2470
rect 9775 2450 9790 2470
rect 9740 2420 9790 2450
rect 9740 2400 9755 2420
rect 9775 2400 9790 2420
rect 9740 2370 9790 2400
rect 9740 2350 9755 2370
rect 9775 2350 9790 2370
rect 9740 2320 9790 2350
rect 9740 2300 9755 2320
rect 9775 2300 9790 2320
rect 9740 2285 9790 2300
rect 9850 2470 9900 2485
rect 9850 2450 9865 2470
rect 9885 2450 9900 2470
rect 9850 2420 9900 2450
rect 9850 2400 9865 2420
rect 9885 2400 9900 2420
rect 9850 2370 9900 2400
rect 9850 2350 9865 2370
rect 9885 2350 9900 2370
rect 9850 2320 9900 2350
rect 9850 2300 9865 2320
rect 9885 2300 9900 2320
rect 9850 2285 9900 2300
rect 9960 2470 10010 2485
rect 10060 2470 10110 2485
rect 9960 2450 9975 2470
rect 9995 2450 10010 2470
rect 10060 2450 10075 2470
rect 10095 2450 10110 2470
rect 9960 2420 10010 2450
rect 10060 2420 10110 2450
rect 9960 2400 9975 2420
rect 9995 2400 10010 2420
rect 10060 2400 10075 2420
rect 10095 2400 10110 2420
rect 9960 2370 10010 2400
rect 10060 2370 10110 2400
rect 9960 2350 9975 2370
rect 9995 2350 10010 2370
rect 10060 2350 10075 2370
rect 10095 2350 10110 2370
rect 9960 2320 10010 2350
rect 10060 2320 10110 2350
rect 9960 2300 9975 2320
rect 9995 2300 10010 2320
rect 10060 2300 10075 2320
rect 10095 2300 10110 2320
rect 9960 2285 10010 2300
rect 10060 2285 10110 2300
rect 10170 2470 10220 2485
rect 10170 2450 10185 2470
rect 10205 2450 10220 2470
rect 10170 2420 10220 2450
rect 10170 2400 10185 2420
rect 10205 2400 10220 2420
rect 10170 2370 10220 2400
rect 10170 2350 10185 2370
rect 10205 2350 10220 2370
rect 10170 2320 10220 2350
rect 10170 2300 10185 2320
rect 10205 2300 10220 2320
rect 10170 2285 10220 2300
rect 10280 2470 10330 2485
rect 10280 2450 10295 2470
rect 10315 2450 10330 2470
rect 10280 2420 10330 2450
rect 10280 2400 10295 2420
rect 10315 2400 10330 2420
rect 10280 2370 10330 2400
rect 10280 2350 10295 2370
rect 10315 2350 10330 2370
rect 10280 2320 10330 2350
rect 10280 2300 10295 2320
rect 10315 2300 10330 2320
rect 10280 2285 10330 2300
rect 10390 2470 10440 2485
rect 10390 2450 10405 2470
rect 10425 2450 10440 2470
rect 10390 2420 10440 2450
rect 10390 2400 10405 2420
rect 10425 2400 10440 2420
rect 10390 2370 10440 2400
rect 10390 2350 10405 2370
rect 10425 2350 10440 2370
rect 10390 2320 10440 2350
rect 10390 2300 10405 2320
rect 10425 2300 10440 2320
rect 10390 2285 10440 2300
rect 10500 2470 10550 2485
rect 10500 2450 10515 2470
rect 10535 2450 10550 2470
rect 10500 2420 10550 2450
rect 10500 2400 10515 2420
rect 10535 2400 10550 2420
rect 10500 2370 10550 2400
rect 10500 2350 10515 2370
rect 10535 2350 10550 2370
rect 10500 2320 10550 2350
rect 10500 2300 10515 2320
rect 10535 2300 10550 2320
rect 10500 2285 10550 2300
rect 10610 2470 10660 2485
rect 10610 2450 10625 2470
rect 10645 2450 10660 2470
rect 10610 2420 10660 2450
rect 10610 2400 10625 2420
rect 10645 2400 10660 2420
rect 10610 2370 10660 2400
rect 10610 2350 10625 2370
rect 10645 2350 10660 2370
rect 10610 2320 10660 2350
rect 10610 2300 10625 2320
rect 10645 2300 10660 2320
rect 10610 2285 10660 2300
rect 10720 2470 10770 2485
rect 10720 2450 10735 2470
rect 10755 2450 10770 2470
rect 10720 2420 10770 2450
rect 10720 2400 10735 2420
rect 10755 2400 10770 2420
rect 10720 2370 10770 2400
rect 10720 2350 10735 2370
rect 10755 2350 10770 2370
rect 10720 2320 10770 2350
rect 10720 2300 10735 2320
rect 10755 2300 10770 2320
rect 10720 2285 10770 2300
<< ndiffc >>
rect 9215 1960 9235 1980
rect 9215 1910 9235 1930
rect 9215 1860 9235 1880
rect 9215 1810 9235 1830
rect 9325 1960 9345 1980
rect 9325 1910 9345 1930
rect 9325 1860 9345 1880
rect 9325 1810 9345 1830
rect 9435 1960 9455 1980
rect 9435 1910 9455 1930
rect 9435 1860 9455 1880
rect 9435 1810 9455 1830
rect 9545 1960 9565 1980
rect 9545 1910 9565 1930
rect 9545 1860 9565 1880
rect 9545 1810 9565 1830
rect 9655 1960 9675 1980
rect 9755 1960 9775 1980
rect 9655 1910 9675 1930
rect 9755 1910 9775 1930
rect 9655 1860 9675 1880
rect 9755 1860 9775 1880
rect 9655 1810 9675 1830
rect 9755 1810 9775 1830
rect 9865 1960 9885 1980
rect 9865 1910 9885 1930
rect 9865 1860 9885 1880
rect 9865 1810 9885 1830
rect 9975 1960 9995 1980
rect 9975 1910 9995 1930
rect 9975 1860 9995 1880
rect 9975 1810 9995 1830
rect 10085 1960 10105 1980
rect 10085 1910 10105 1930
rect 10085 1860 10105 1880
rect 10085 1810 10105 1830
rect 10195 1960 10215 1980
rect 10295 1960 10315 1980
rect 10195 1910 10215 1930
rect 10295 1910 10315 1930
rect 10195 1860 10215 1880
rect 10295 1860 10315 1880
rect 10195 1810 10215 1830
rect 10295 1810 10315 1830
rect 10405 1960 10425 1980
rect 10405 1910 10425 1930
rect 10405 1860 10425 1880
rect 10405 1810 10425 1830
rect 10515 1960 10535 1980
rect 10515 1910 10535 1930
rect 10515 1860 10535 1880
rect 10515 1810 10535 1830
rect 10625 1960 10645 1980
rect 10625 1910 10645 1930
rect 10625 1860 10645 1880
rect 10625 1810 10645 1830
rect 10735 1960 10755 1980
rect 10735 1910 10755 1930
rect 10735 1860 10755 1880
rect 10735 1810 10755 1830
<< pdiffc >>
rect 9315 2450 9335 2470
rect 9315 2400 9335 2420
rect 9315 2350 9335 2370
rect 9315 2300 9335 2320
rect 9425 2450 9445 2470
rect 9425 2400 9445 2420
rect 9425 2350 9445 2370
rect 9425 2300 9445 2320
rect 9535 2450 9555 2470
rect 9535 2400 9555 2420
rect 9535 2350 9555 2370
rect 9535 2300 9555 2320
rect 9645 2450 9665 2470
rect 9645 2400 9665 2420
rect 9645 2350 9665 2370
rect 9645 2300 9665 2320
rect 9755 2450 9775 2470
rect 9755 2400 9775 2420
rect 9755 2350 9775 2370
rect 9755 2300 9775 2320
rect 9865 2450 9885 2470
rect 9865 2400 9885 2420
rect 9865 2350 9885 2370
rect 9865 2300 9885 2320
rect 9975 2450 9995 2470
rect 10075 2450 10095 2470
rect 9975 2400 9995 2420
rect 10075 2400 10095 2420
rect 9975 2350 9995 2370
rect 10075 2350 10095 2370
rect 9975 2300 9995 2320
rect 10075 2300 10095 2320
rect 10185 2450 10205 2470
rect 10185 2400 10205 2420
rect 10185 2350 10205 2370
rect 10185 2300 10205 2320
rect 10295 2450 10315 2470
rect 10295 2400 10315 2420
rect 10295 2350 10315 2370
rect 10295 2300 10315 2320
rect 10405 2450 10425 2470
rect 10405 2400 10425 2420
rect 10405 2350 10425 2370
rect 10405 2300 10425 2320
rect 10515 2450 10535 2470
rect 10515 2400 10535 2420
rect 10515 2350 10535 2370
rect 10515 2300 10535 2320
rect 10625 2450 10645 2470
rect 10625 2400 10645 2420
rect 10625 2350 10645 2370
rect 10625 2300 10645 2320
rect 10735 2450 10755 2470
rect 10735 2400 10755 2420
rect 10735 2350 10755 2370
rect 10735 2300 10755 2320
<< psubdiff >>
rect 9150 1980 9200 1995
rect 9150 1960 9165 1980
rect 9185 1960 9200 1980
rect 9150 1930 9200 1960
rect 9150 1910 9165 1930
rect 9185 1910 9200 1930
rect 9150 1880 9200 1910
rect 9150 1860 9165 1880
rect 9185 1860 9200 1880
rect 9150 1830 9200 1860
rect 9150 1810 9165 1830
rect 9185 1810 9200 1830
rect 9150 1795 9200 1810
rect 9690 1980 9740 1995
rect 9690 1960 9705 1980
rect 9725 1960 9740 1980
rect 9690 1930 9740 1960
rect 9690 1910 9705 1930
rect 9725 1910 9740 1930
rect 9690 1880 9740 1910
rect 9690 1860 9705 1880
rect 9725 1860 9740 1880
rect 9690 1830 9740 1860
rect 9690 1810 9705 1830
rect 9725 1810 9740 1830
rect 9690 1795 9740 1810
rect 10230 1980 10280 1995
rect 10230 1960 10245 1980
rect 10265 1960 10280 1980
rect 10230 1930 10280 1960
rect 10230 1910 10245 1930
rect 10265 1910 10280 1930
rect 10230 1880 10280 1910
rect 10230 1860 10245 1880
rect 10265 1860 10280 1880
rect 10230 1830 10280 1860
rect 10230 1810 10245 1830
rect 10265 1810 10280 1830
rect 10230 1795 10280 1810
rect 10770 1980 10820 1995
rect 10770 1960 10785 1980
rect 10805 1960 10820 1980
rect 10770 1930 10820 1960
rect 10770 1910 10785 1930
rect 10805 1910 10820 1930
rect 10770 1880 10820 1910
rect 10770 1860 10785 1880
rect 10805 1860 10820 1880
rect 10770 1830 10820 1860
rect 10770 1810 10785 1830
rect 10805 1810 10820 1830
rect 10770 1795 10820 1810
<< nsubdiff >>
rect 9250 2470 9300 2485
rect 9250 2450 9265 2470
rect 9285 2450 9300 2470
rect 9250 2420 9300 2450
rect 9250 2400 9265 2420
rect 9285 2400 9300 2420
rect 9250 2370 9300 2400
rect 9250 2350 9265 2370
rect 9285 2350 9300 2370
rect 9250 2320 9300 2350
rect 9250 2300 9265 2320
rect 9285 2300 9300 2320
rect 9250 2285 9300 2300
rect 10010 2470 10060 2485
rect 10010 2450 10025 2470
rect 10045 2450 10060 2470
rect 10010 2420 10060 2450
rect 10010 2400 10025 2420
rect 10045 2400 10060 2420
rect 10010 2370 10060 2400
rect 10010 2350 10025 2370
rect 10045 2350 10060 2370
rect 10010 2320 10060 2350
rect 10010 2300 10025 2320
rect 10045 2300 10060 2320
rect 10010 2285 10060 2300
rect 10770 2470 10820 2485
rect 10770 2450 10785 2470
rect 10805 2450 10820 2470
rect 10770 2420 10820 2450
rect 10770 2400 10785 2420
rect 10805 2400 10820 2420
rect 10770 2370 10820 2400
rect 10770 2350 10785 2370
rect 10805 2350 10820 2370
rect 10770 2320 10820 2350
rect 10770 2300 10785 2320
rect 10805 2300 10820 2320
rect 10770 2285 10820 2300
<< psubdiffcont >>
rect 9165 1960 9185 1980
rect 9165 1910 9185 1930
rect 9165 1860 9185 1880
rect 9165 1810 9185 1830
rect 9705 1960 9725 1980
rect 9705 1910 9725 1930
rect 9705 1860 9725 1880
rect 9705 1810 9725 1830
rect 10245 1960 10265 1980
rect 10245 1910 10265 1930
rect 10245 1860 10265 1880
rect 10245 1810 10265 1830
rect 10785 1960 10805 1980
rect 10785 1910 10805 1930
rect 10785 1860 10805 1880
rect 10785 1810 10805 1830
<< nsubdiffcont >>
rect 9265 2450 9285 2470
rect 9265 2400 9285 2420
rect 9265 2350 9285 2370
rect 9265 2300 9285 2320
rect 10025 2450 10045 2470
rect 10025 2400 10045 2420
rect 10025 2350 10045 2370
rect 10025 2300 10045 2320
rect 10785 2450 10805 2470
rect 10785 2400 10805 2420
rect 10785 2350 10805 2370
rect 10785 2300 10805 2320
<< poly >>
rect 9305 2530 9345 2540
rect 9305 2510 9315 2530
rect 9335 2515 9345 2530
rect 10725 2530 10765 2540
rect 10725 2515 10735 2530
rect 9335 2510 9410 2515
rect 9305 2500 9410 2510
rect 9350 2485 9410 2500
rect 9460 2495 9850 2515
rect 9460 2485 9520 2495
rect 9570 2485 9630 2495
rect 9680 2485 9740 2495
rect 9790 2485 9850 2495
rect 9900 2485 9960 2500
rect 10110 2485 10170 2500
rect 10220 2495 10610 2515
rect 10220 2485 10280 2495
rect 10330 2485 10390 2495
rect 10440 2485 10500 2495
rect 10550 2485 10610 2495
rect 10660 2510 10735 2515
rect 10755 2510 10765 2530
rect 10660 2500 10765 2510
rect 10660 2485 10720 2500
rect 9350 2270 9410 2285
rect 9460 2275 9520 2285
rect 9570 2275 9630 2285
rect 9680 2275 9740 2285
rect 9790 2275 9850 2285
rect 9460 2255 9850 2275
rect 9900 2275 9960 2285
rect 10110 2275 10170 2285
rect 9900 2260 10170 2275
rect 10220 2270 10280 2285
rect 10330 2270 10390 2285
rect 10440 2270 10500 2285
rect 10550 2270 10610 2285
rect 10660 2270 10720 2285
rect 10015 2240 10025 2260
rect 10045 2240 10055 2260
rect 10220 2255 10610 2270
rect 10015 2230 10055 2240
rect 10570 2245 10610 2255
rect 10570 2225 10580 2245
rect 10600 2225 10610 2245
rect 10570 2215 10610 2225
rect 9425 2105 9465 2115
rect 9425 2085 9435 2105
rect 9455 2085 9465 2105
rect 9425 2025 9465 2085
rect 10570 2055 10610 2065
rect 9695 2040 9735 2050
rect 9250 1995 9310 2010
rect 9360 2005 9530 2025
rect 9695 2020 9705 2040
rect 9725 2020 9735 2040
rect 10235 2040 10275 2050
rect 10235 2020 10245 2040
rect 10265 2020 10275 2040
rect 10570 2035 10580 2055
rect 10600 2035 10610 2055
rect 10570 2025 10610 2035
rect 9360 1995 9420 2005
rect 9470 1995 9530 2005
rect 9580 2005 9850 2020
rect 9580 1995 9640 2005
rect 9790 1995 9850 2005
rect 9900 2005 10070 2020
rect 9900 1995 9960 2005
rect 10010 1995 10070 2005
rect 10120 2005 10390 2020
rect 10120 1995 10180 2005
rect 10330 1995 10390 2005
rect 10440 2010 10610 2025
rect 10440 1995 10500 2010
rect 10550 1995 10610 2010
rect 10660 1995 10720 2010
rect 9250 1780 9310 1795
rect 9205 1770 9310 1780
rect 9205 1750 9215 1770
rect 9235 1765 9310 1770
rect 9360 1785 9420 1795
rect 9470 1785 9530 1795
rect 9360 1765 9530 1785
rect 9580 1780 9640 1795
rect 9790 1780 9850 1795
rect 9900 1785 9960 1795
rect 10010 1785 10070 1795
rect 9235 1750 9245 1765
rect 9205 1740 9245 1750
rect 9470 1755 9530 1765
rect 9900 1765 10070 1785
rect 10120 1780 10180 1795
rect 10330 1780 10390 1795
rect 10440 1785 10500 1795
rect 10550 1785 10610 1795
rect 10440 1765 10610 1785
rect 10660 1780 10720 1795
rect 10660 1770 10765 1780
rect 10660 1765 10735 1770
rect 9900 1755 9960 1765
rect 9470 1740 9960 1755
rect 10725 1750 10735 1765
rect 10755 1750 10765 1770
rect 10725 1740 10765 1750
<< polycont >>
rect 9315 2510 9335 2530
rect 10735 2510 10755 2530
rect 10025 2240 10045 2260
rect 10580 2225 10600 2245
rect 9435 2085 9455 2105
rect 9705 2020 9725 2040
rect 10245 2020 10265 2040
rect 10580 2035 10600 2055
rect 9215 1750 9235 1770
rect 10735 1750 10755 1770
<< locali >>
rect 11025 2850 11080 2860
rect 11025 2815 11035 2850
rect 11070 2815 11080 2850
rect 11025 2805 11080 2815
rect 9150 2565 9180 2585
rect 9200 2565 9230 2585
rect 9250 2565 9280 2585
rect 9300 2565 9330 2585
rect 9350 2565 9380 2585
rect 9400 2565 9430 2585
rect 9450 2565 9480 2585
rect 9500 2565 9530 2585
rect 9550 2565 9580 2585
rect 9600 2565 9630 2585
rect 9650 2565 9680 2585
rect 9700 2565 9730 2585
rect 9750 2565 9780 2585
rect 9800 2565 9830 2585
rect 9850 2565 9880 2585
rect 9900 2565 9930 2585
rect 9950 2565 9980 2585
rect 10000 2565 10030 2585
rect 10050 2565 10080 2585
rect 10100 2565 10130 2585
rect 10150 2565 10180 2585
rect 10200 2565 10230 2585
rect 10250 2565 10280 2585
rect 10300 2565 10330 2585
rect 10350 2565 10380 2585
rect 10400 2565 10430 2585
rect 10450 2565 10480 2585
rect 10500 2565 10530 2585
rect 10550 2565 10580 2585
rect 10600 2565 10630 2585
rect 10650 2565 10680 2585
rect 10700 2565 10730 2585
rect 10750 2565 10765 2585
rect 9305 2530 9345 2565
rect 9305 2510 9315 2530
rect 9335 2510 9345 2530
rect 9305 2480 9345 2510
rect 9255 2470 9345 2480
rect 9255 2450 9265 2470
rect 9285 2450 9315 2470
rect 9335 2450 9345 2470
rect 9255 2420 9345 2450
rect 9255 2400 9265 2420
rect 9285 2400 9315 2420
rect 9335 2400 9345 2420
rect 9255 2370 9345 2400
rect 9255 2350 9265 2370
rect 9285 2350 9315 2370
rect 9335 2350 9345 2370
rect 9255 2320 9345 2350
rect 9255 2300 9265 2320
rect 9285 2300 9315 2320
rect 9335 2300 9345 2320
rect 9255 2290 9345 2300
rect 9415 2470 9455 2565
rect 9415 2450 9425 2470
rect 9445 2450 9455 2470
rect 9415 2420 9455 2450
rect 9415 2400 9425 2420
rect 9445 2400 9455 2420
rect 9415 2370 9455 2400
rect 9415 2350 9425 2370
rect 9445 2350 9455 2370
rect 9415 2320 9455 2350
rect 9415 2300 9425 2320
rect 9445 2300 9455 2320
rect 9415 2290 9455 2300
rect 9525 2470 9565 2480
rect 9525 2450 9535 2470
rect 9555 2450 9565 2470
rect 9525 2420 9565 2450
rect 9525 2400 9535 2420
rect 9555 2400 9565 2420
rect 9525 2370 9565 2400
rect 9525 2350 9535 2370
rect 9555 2350 9565 2370
rect 9525 2320 9565 2350
rect 9525 2300 9535 2320
rect 9555 2300 9565 2320
rect 9525 2270 9565 2300
rect 9635 2470 9675 2565
rect 9635 2450 9645 2470
rect 9665 2450 9675 2470
rect 9635 2420 9675 2450
rect 9635 2400 9645 2420
rect 9665 2400 9675 2420
rect 9635 2370 9675 2400
rect 9635 2350 9645 2370
rect 9665 2350 9675 2370
rect 9635 2320 9675 2350
rect 9635 2300 9645 2320
rect 9665 2300 9675 2320
rect 9635 2290 9675 2300
rect 9745 2470 9785 2480
rect 9745 2450 9755 2470
rect 9775 2450 9785 2470
rect 9745 2420 9785 2450
rect 9745 2400 9755 2420
rect 9775 2400 9785 2420
rect 9745 2370 9785 2400
rect 9745 2350 9755 2370
rect 9775 2350 9785 2370
rect 9745 2320 9785 2350
rect 9745 2300 9755 2320
rect 9775 2300 9785 2320
rect 9745 2270 9785 2300
rect 9855 2470 9895 2565
rect 10015 2480 10055 2565
rect 9855 2450 9865 2470
rect 9885 2450 9895 2470
rect 9855 2420 9895 2450
rect 9855 2400 9865 2420
rect 9885 2400 9895 2420
rect 9855 2370 9895 2400
rect 9855 2350 9865 2370
rect 9885 2350 9895 2370
rect 9855 2320 9895 2350
rect 9855 2300 9865 2320
rect 9885 2300 9895 2320
rect 9855 2290 9895 2300
rect 9965 2470 10105 2480
rect 9965 2450 9975 2470
rect 9995 2450 10025 2470
rect 10045 2450 10075 2470
rect 10095 2450 10105 2470
rect 9965 2420 10105 2450
rect 9965 2400 9975 2420
rect 9995 2400 10025 2420
rect 10045 2400 10075 2420
rect 10095 2400 10105 2420
rect 9965 2370 10105 2400
rect 9965 2350 9975 2370
rect 9995 2350 10025 2370
rect 10045 2350 10075 2370
rect 10095 2350 10105 2370
rect 9965 2320 10105 2350
rect 9965 2300 9975 2320
rect 9995 2300 10025 2320
rect 10045 2300 10075 2320
rect 10095 2300 10105 2320
rect 9965 2290 10105 2300
rect 10175 2470 10215 2565
rect 10175 2450 10185 2470
rect 10205 2450 10215 2470
rect 10175 2420 10215 2450
rect 10175 2400 10185 2420
rect 10205 2400 10215 2420
rect 10175 2370 10215 2400
rect 10175 2350 10185 2370
rect 10205 2350 10215 2370
rect 10175 2320 10215 2350
rect 10175 2300 10185 2320
rect 10205 2300 10215 2320
rect 10175 2290 10215 2300
rect 10285 2470 10325 2480
rect 10285 2450 10295 2470
rect 10315 2450 10325 2470
rect 10285 2420 10325 2450
rect 10285 2400 10295 2420
rect 10315 2400 10325 2420
rect 10285 2370 10325 2400
rect 10285 2350 10295 2370
rect 10315 2350 10325 2370
rect 10285 2320 10325 2350
rect 10285 2300 10295 2320
rect 10315 2300 10325 2320
rect 9525 2230 9785 2270
rect 10015 2260 10055 2290
rect 10015 2240 10025 2260
rect 10045 2240 10055 2260
rect 10015 2230 10055 2240
rect 10285 2270 10325 2300
rect 10395 2470 10435 2565
rect 10395 2450 10405 2470
rect 10425 2450 10435 2470
rect 10395 2420 10435 2450
rect 10395 2400 10405 2420
rect 10425 2400 10435 2420
rect 10395 2370 10435 2400
rect 10395 2350 10405 2370
rect 10425 2350 10435 2370
rect 10395 2320 10435 2350
rect 10395 2300 10405 2320
rect 10425 2300 10435 2320
rect 10395 2290 10435 2300
rect 10505 2470 10545 2480
rect 10505 2450 10515 2470
rect 10535 2450 10545 2470
rect 10505 2420 10545 2450
rect 10505 2400 10515 2420
rect 10535 2400 10545 2420
rect 10505 2370 10545 2400
rect 10505 2350 10515 2370
rect 10535 2350 10545 2370
rect 10505 2320 10545 2350
rect 10505 2300 10515 2320
rect 10535 2300 10545 2320
rect 10505 2270 10545 2300
rect 10615 2470 10655 2565
rect 10615 2450 10625 2470
rect 10645 2450 10655 2470
rect 10615 2420 10655 2450
rect 10615 2400 10625 2420
rect 10645 2400 10655 2420
rect 10615 2370 10655 2400
rect 10615 2350 10625 2370
rect 10645 2350 10655 2370
rect 10615 2320 10655 2350
rect 10615 2300 10625 2320
rect 10645 2300 10655 2320
rect 10615 2290 10655 2300
rect 10725 2530 10765 2565
rect 10725 2510 10735 2530
rect 10755 2510 10765 2530
rect 10725 2480 10765 2510
rect 10725 2470 10815 2480
rect 10725 2450 10735 2470
rect 10755 2450 10785 2470
rect 10805 2450 10815 2470
rect 10725 2420 10815 2450
rect 10725 2400 10735 2420
rect 10755 2400 10785 2420
rect 10805 2400 10815 2420
rect 10725 2370 10815 2400
rect 10725 2350 10735 2370
rect 10755 2350 10785 2370
rect 10805 2350 10815 2370
rect 10725 2320 10815 2350
rect 10725 2300 10735 2320
rect 10755 2300 10785 2320
rect 10805 2300 10815 2320
rect 10725 2290 10815 2300
rect 10285 2230 10545 2270
rect 10905 2260 10960 2270
rect 10905 2255 10915 2260
rect 9745 2155 9785 2230
rect 10505 2160 10545 2230
rect 10570 2245 10915 2255
rect 10570 2225 10580 2245
rect 10600 2225 10915 2245
rect 10950 2225 10960 2260
rect 10570 2215 10960 2225
rect 9745 2115 10005 2155
rect 9425 2105 9465 2115
rect 9425 2085 9435 2105
rect 9455 2085 9465 2105
rect 9155 1980 9245 1990
rect 9155 1960 9165 1980
rect 9185 1960 9215 1980
rect 9235 1960 9245 1980
rect 9155 1930 9245 1960
rect 9155 1910 9165 1930
rect 9185 1910 9215 1930
rect 9235 1910 9245 1930
rect 9155 1880 9245 1910
rect 9155 1860 9165 1880
rect 9185 1860 9215 1880
rect 9235 1860 9245 1880
rect 9155 1830 9245 1860
rect 9155 1810 9165 1830
rect 9185 1810 9215 1830
rect 9235 1810 9245 1830
rect 9155 1800 9245 1810
rect 9205 1770 9245 1800
rect 9205 1750 9215 1770
rect 9235 1750 9245 1770
rect 9205 1725 9245 1750
rect 9315 1980 9355 1990
rect 9315 1960 9325 1980
rect 9345 1960 9355 1980
rect 9315 1930 9355 1960
rect 9315 1910 9325 1930
rect 9345 1910 9355 1930
rect 9315 1880 9355 1910
rect 9315 1860 9325 1880
rect 9345 1860 9355 1880
rect 9315 1830 9355 1860
rect 9315 1810 9325 1830
rect 9345 1810 9355 1830
rect 9315 1725 9355 1810
rect 9425 1980 9465 2085
rect 9695 2040 9735 2050
rect 9695 2020 9705 2040
rect 9725 2020 9735 2040
rect 9695 1990 9735 2020
rect 9425 1960 9435 1980
rect 9455 1960 9465 1980
rect 9425 1930 9465 1960
rect 9425 1910 9435 1930
rect 9455 1910 9465 1930
rect 9425 1880 9465 1910
rect 9425 1860 9435 1880
rect 9455 1860 9465 1880
rect 9425 1830 9465 1860
rect 9425 1810 9435 1830
rect 9455 1810 9465 1830
rect 9425 1800 9465 1810
rect 9535 1980 9575 1990
rect 9535 1960 9545 1980
rect 9565 1960 9575 1980
rect 9535 1930 9575 1960
rect 9535 1910 9545 1930
rect 9565 1910 9575 1930
rect 9535 1880 9575 1910
rect 9535 1860 9545 1880
rect 9565 1860 9575 1880
rect 9535 1830 9575 1860
rect 9535 1810 9545 1830
rect 9565 1810 9575 1830
rect 9535 1725 9575 1810
rect 9645 1980 9785 1990
rect 9645 1960 9655 1980
rect 9675 1960 9705 1980
rect 9725 1960 9755 1980
rect 9775 1960 9785 1980
rect 9645 1930 9785 1960
rect 9645 1910 9655 1930
rect 9675 1910 9705 1930
rect 9725 1910 9755 1930
rect 9775 1910 9785 1930
rect 9645 1880 9785 1910
rect 9645 1860 9655 1880
rect 9675 1860 9705 1880
rect 9725 1860 9755 1880
rect 9775 1860 9785 1880
rect 9645 1830 9785 1860
rect 9645 1810 9655 1830
rect 9675 1810 9705 1830
rect 9725 1810 9755 1830
rect 9775 1810 9785 1830
rect 9645 1800 9785 1810
rect 9855 1980 9895 1990
rect 9855 1960 9865 1980
rect 9885 1960 9895 1980
rect 9855 1930 9895 1960
rect 9855 1910 9865 1930
rect 9885 1910 9895 1930
rect 9855 1880 9895 1910
rect 9855 1860 9865 1880
rect 9885 1860 9895 1880
rect 9855 1830 9895 1860
rect 9855 1810 9865 1830
rect 9885 1810 9895 1830
rect 9695 1725 9735 1800
rect 9855 1725 9895 1810
rect 9965 1980 10005 2115
rect 10505 2120 10860 2160
rect 10235 2040 10275 2050
rect 10235 2020 10245 2040
rect 10265 2020 10275 2040
rect 10235 1990 10275 2020
rect 9965 1960 9975 1980
rect 9995 1960 10005 1980
rect 9965 1930 10005 1960
rect 9965 1910 9975 1930
rect 9995 1910 10005 1930
rect 9965 1880 10005 1910
rect 9965 1860 9975 1880
rect 9995 1860 10005 1880
rect 9965 1830 10005 1860
rect 9965 1810 9975 1830
rect 9995 1810 10005 1830
rect 9965 1800 10005 1810
rect 10075 1980 10115 1990
rect 10075 1960 10085 1980
rect 10105 1960 10115 1980
rect 10075 1930 10115 1960
rect 10075 1910 10085 1930
rect 10105 1910 10115 1930
rect 10075 1880 10115 1910
rect 10075 1860 10085 1880
rect 10105 1860 10115 1880
rect 10075 1830 10115 1860
rect 10075 1810 10085 1830
rect 10105 1810 10115 1830
rect 10075 1725 10115 1810
rect 10185 1980 10325 1990
rect 10185 1960 10195 1980
rect 10215 1960 10245 1980
rect 10265 1960 10295 1980
rect 10315 1960 10325 1980
rect 10185 1930 10325 1960
rect 10185 1910 10195 1930
rect 10215 1910 10245 1930
rect 10265 1910 10295 1930
rect 10315 1910 10325 1930
rect 10185 1880 10325 1910
rect 10185 1860 10195 1880
rect 10215 1860 10245 1880
rect 10265 1860 10295 1880
rect 10315 1860 10325 1880
rect 10185 1830 10325 1860
rect 10185 1810 10195 1830
rect 10215 1810 10245 1830
rect 10265 1810 10295 1830
rect 10315 1810 10325 1830
rect 10185 1800 10325 1810
rect 10395 1980 10435 1990
rect 10395 1960 10405 1980
rect 10425 1960 10435 1980
rect 10395 1930 10435 1960
rect 10395 1910 10405 1930
rect 10425 1910 10435 1930
rect 10395 1880 10435 1910
rect 10395 1860 10405 1880
rect 10425 1860 10435 1880
rect 10395 1830 10435 1860
rect 10395 1810 10405 1830
rect 10425 1810 10435 1830
rect 10235 1725 10275 1800
rect 10395 1725 10435 1810
rect 10505 1980 10545 2120
rect 10570 2055 10960 2065
rect 10570 2035 10580 2055
rect 10600 2035 10915 2055
rect 10570 2025 10915 2035
rect 10905 2020 10915 2025
rect 10950 2020 10960 2055
rect 10905 2010 10960 2020
rect 10505 1960 10515 1980
rect 10535 1960 10545 1980
rect 10505 1930 10545 1960
rect 10505 1910 10515 1930
rect 10535 1910 10545 1930
rect 10505 1880 10545 1910
rect 10505 1860 10515 1880
rect 10535 1860 10545 1880
rect 10505 1830 10545 1860
rect 10505 1810 10515 1830
rect 10535 1810 10545 1830
rect 10505 1800 10545 1810
rect 10615 1980 10655 1990
rect 10615 1960 10625 1980
rect 10645 1960 10655 1980
rect 10615 1930 10655 1960
rect 10615 1910 10625 1930
rect 10645 1910 10655 1930
rect 10615 1880 10655 1910
rect 10615 1860 10625 1880
rect 10645 1860 10655 1880
rect 10615 1830 10655 1860
rect 10615 1810 10625 1830
rect 10645 1810 10655 1830
rect 10615 1725 10655 1810
rect 10725 1980 10815 1990
rect 10725 1960 10735 1980
rect 10755 1960 10785 1980
rect 10805 1960 10815 1980
rect 10725 1930 10815 1960
rect 10725 1910 10735 1930
rect 10755 1910 10785 1930
rect 10805 1910 10815 1930
rect 10725 1880 10815 1910
rect 10725 1860 10735 1880
rect 10755 1860 10785 1880
rect 10805 1860 10815 1880
rect 10725 1830 10815 1860
rect 10725 1810 10735 1830
rect 10755 1810 10785 1830
rect 10805 1810 10815 1830
rect 10725 1800 10815 1810
rect 10725 1770 10765 1800
rect 10725 1750 10735 1770
rect 10755 1750 10765 1770
rect 10725 1725 10765 1750
rect 9155 1705 9185 1725
rect 9205 1705 9235 1725
rect 9255 1705 9285 1725
rect 9305 1705 9335 1725
rect 9355 1705 9385 1725
rect 9405 1705 9435 1725
rect 9455 1705 9485 1725
rect 9505 1705 9535 1725
rect 9555 1705 9585 1725
rect 9605 1705 9635 1725
rect 9655 1705 9685 1725
rect 9705 1705 9735 1725
rect 9755 1705 9785 1725
rect 9805 1705 9835 1725
rect 9855 1705 9885 1725
rect 9905 1705 9935 1725
rect 9955 1705 9985 1725
rect 10005 1705 10035 1725
rect 10055 1705 10085 1725
rect 10105 1705 10135 1725
rect 10155 1705 10185 1725
rect 10205 1705 10235 1725
rect 10255 1705 10285 1725
rect 10305 1705 10335 1725
rect 10355 1705 10385 1725
rect 10405 1705 10435 1725
rect 10455 1705 10485 1725
rect 10505 1705 10535 1725
rect 10555 1705 10585 1725
rect 10605 1705 10635 1725
rect 10655 1705 10685 1725
rect 10705 1705 10735 1725
rect 10755 1705 10765 1725
rect 11080 1660 11135 1670
rect 11080 1625 11090 1660
rect 11125 1625 11135 1660
rect 11080 1615 11135 1625
<< viali >>
rect 11035 2815 11070 2850
rect 9180 2565 9200 2585
rect 9230 2565 9250 2585
rect 9280 2565 9300 2585
rect 9330 2565 9350 2585
rect 9380 2565 9400 2585
rect 9430 2565 9450 2585
rect 9480 2565 9500 2585
rect 9530 2565 9550 2585
rect 9580 2565 9600 2585
rect 9630 2565 9650 2585
rect 9680 2565 9700 2585
rect 9730 2565 9750 2585
rect 9780 2565 9800 2585
rect 9830 2565 9850 2585
rect 9880 2565 9900 2585
rect 9930 2565 9950 2585
rect 9980 2565 10000 2585
rect 10030 2565 10050 2585
rect 10080 2565 10100 2585
rect 10130 2565 10150 2585
rect 10180 2565 10200 2585
rect 10230 2565 10250 2585
rect 10280 2565 10300 2585
rect 10330 2565 10350 2585
rect 10380 2565 10400 2585
rect 10430 2565 10450 2585
rect 10480 2565 10500 2585
rect 10530 2565 10550 2585
rect 10580 2565 10600 2585
rect 10630 2565 10650 2585
rect 10680 2565 10700 2585
rect 10730 2565 10750 2585
rect 10915 2225 10950 2260
rect 10915 2020 10950 2055
rect 9185 1705 9205 1725
rect 9235 1705 9255 1725
rect 9285 1705 9305 1725
rect 9335 1705 9355 1725
rect 9385 1705 9405 1725
rect 9435 1705 9455 1725
rect 9485 1705 9505 1725
rect 9535 1705 9555 1725
rect 9585 1705 9605 1725
rect 9635 1705 9655 1725
rect 9685 1705 9705 1725
rect 9735 1705 9755 1725
rect 9785 1705 9805 1725
rect 9835 1705 9855 1725
rect 9885 1705 9905 1725
rect 9935 1705 9955 1725
rect 9985 1705 10005 1725
rect 10035 1705 10055 1725
rect 10085 1705 10105 1725
rect 10135 1705 10155 1725
rect 10185 1705 10205 1725
rect 10235 1705 10255 1725
rect 10285 1705 10305 1725
rect 10335 1705 10355 1725
rect 10385 1705 10405 1725
rect 10435 1705 10455 1725
rect 10485 1705 10505 1725
rect 10535 1705 10555 1725
rect 10585 1705 10605 1725
rect 10635 1705 10655 1725
rect 10685 1705 10705 1725
rect 10735 1705 10755 1725
rect 11090 1625 11125 1660
<< metal1 >>
rect 11025 2850 11080 2860
rect 11025 2815 11035 2850
rect 11070 2815 11080 2850
rect 11025 2805 11080 2815
rect 9150 2585 10765 2595
rect 9150 2565 9180 2585
rect 9200 2565 9230 2585
rect 9250 2565 9280 2585
rect 9300 2565 9330 2585
rect 9350 2565 9380 2585
rect 9400 2565 9430 2585
rect 9450 2565 9480 2585
rect 9500 2565 9530 2585
rect 9550 2565 9580 2585
rect 9600 2565 9630 2585
rect 9650 2565 9680 2585
rect 9700 2565 9730 2585
rect 9750 2565 9780 2585
rect 9800 2565 9830 2585
rect 9850 2565 9880 2585
rect 9900 2565 9930 2585
rect 9950 2565 9980 2585
rect 10000 2565 10030 2585
rect 10050 2565 10080 2585
rect 10100 2565 10130 2585
rect 10150 2565 10180 2585
rect 10200 2565 10230 2585
rect 10250 2565 10280 2585
rect 10300 2565 10330 2585
rect 10350 2565 10380 2585
rect 10400 2565 10430 2585
rect 10450 2565 10480 2585
rect 10500 2565 10530 2585
rect 10550 2565 10580 2585
rect 10600 2565 10630 2585
rect 10650 2565 10680 2585
rect 10700 2565 10730 2585
rect 10750 2565 10765 2585
rect 9150 2555 10765 2565
rect 10905 2260 10960 2270
rect 10905 2225 10915 2260
rect 10950 2225 10960 2260
rect 10905 2215 10960 2225
rect 10905 2055 10960 2065
rect 10905 2020 10915 2055
rect 10950 2020 10960 2055
rect 10905 2010 10960 2020
rect 9155 1725 10765 1735
rect 9155 1705 9185 1725
rect 9205 1705 9235 1725
rect 9255 1705 9285 1725
rect 9305 1705 9335 1725
rect 9355 1705 9385 1725
rect 9405 1705 9435 1725
rect 9455 1705 9485 1725
rect 9505 1705 9535 1725
rect 9555 1705 9585 1725
rect 9605 1705 9635 1725
rect 9655 1705 9685 1725
rect 9705 1705 9735 1725
rect 9755 1705 9785 1725
rect 9805 1705 9835 1725
rect 9855 1705 9885 1725
rect 9905 1705 9935 1725
rect 9955 1705 9985 1725
rect 10005 1705 10035 1725
rect 10055 1705 10085 1725
rect 10105 1705 10135 1725
rect 10155 1705 10185 1725
rect 10205 1705 10235 1725
rect 10255 1705 10285 1725
rect 10305 1705 10335 1725
rect 10355 1705 10385 1725
rect 10405 1705 10435 1725
rect 10455 1705 10485 1725
rect 10505 1705 10535 1725
rect 10555 1705 10585 1725
rect 10605 1705 10635 1725
rect 10655 1705 10685 1725
rect 10705 1705 10735 1725
rect 10755 1705 10765 1725
rect 9155 1695 10765 1705
rect 11080 1660 11135 1670
rect 11080 1625 11090 1660
rect 11125 1625 11135 1660
rect 11080 1615 11135 1625
<< via1 >>
rect 11035 2815 11070 2850
rect 10915 2225 10950 2260
rect 10915 2020 10950 2055
rect 11090 1625 11125 1660
<< metal2 >>
rect 11025 2850 11080 2860
rect 11025 2840 11035 2850
rect 9105 2825 11035 2840
rect 11025 2815 11035 2825
rect 11070 2815 11080 2850
rect 11025 2805 11080 2815
rect 10905 2260 10960 2270
rect 10905 2225 10915 2260
rect 10950 2225 10960 2260
rect 10905 2215 10960 2225
rect 10905 2055 10960 2065
rect 10905 2020 10915 2055
rect 10950 2020 10960 2055
rect 10905 2010 10960 2020
rect 11080 1660 11135 1670
rect 11080 1650 11090 1660
rect 9105 1635 11090 1650
rect 11080 1625 11090 1635
rect 11125 1625 11135 1660
rect 11080 1615 11135 1625
<< via2 >>
rect 11035 2815 11070 2850
rect 10915 2225 10950 2260
rect 10915 2020 10950 2055
rect 11090 1625 11125 1660
<< metal3 >>
rect 11025 2850 11630 2860
rect 11025 2815 11035 2850
rect 11070 2815 11630 2850
rect 11025 2805 11630 2815
rect 10905 2260 10960 2270
rect 10905 2225 10915 2260
rect 10950 2225 10960 2260
rect 10905 2215 10960 2225
rect 11080 2200 11630 2805
rect 10905 2055 10960 2065
rect 10905 2020 10915 2055
rect 10950 2020 10960 2055
rect 10905 2010 10960 2020
rect 11080 1670 11380 2080
rect 11080 1660 11135 1670
rect 11080 1625 11090 1660
rect 11125 1625 11135 1660
rect 11080 1615 11135 1625
<< via3 >>
rect 10915 2225 10950 2260
rect 10915 2020 10950 2055
<< mimcap >>
rect 11095 2260 11615 2845
rect 11095 2225 11105 2260
rect 11140 2225 11615 2260
rect 11095 2215 11615 2225
rect 11095 2055 11365 2065
rect 11095 2020 11105 2055
rect 11140 2020 11365 2055
rect 11095 1685 11365 2020
<< mimcapcontact >>
rect 11105 2225 11140 2260
rect 11105 2020 11140 2055
<< metal4 >>
rect 10905 2260 11150 2270
rect 10905 2225 10915 2260
rect 10950 2225 11105 2260
rect 11140 2225 11150 2260
rect 10905 2215 11150 2225
rect 10905 2055 11150 2065
rect 10905 2020 10915 2055
rect 10950 2020 11105 2055
rect 11140 2020 11150 2055
rect 10905 2010 11150 2020
<< labels >>
flabel metal1 9150 2575 9150 2575 7 FreeSans 400 0 -200 0 VDDA
port 1 w
flabel poly 10610 2270 10610 2270 3 FreeSans 400 0 200 0 UP_input
port 8 e
flabel poly 9510 2255 9510 2255 5 FreeSans 400 0 0 -200 opamp_out
port 10 s
flabel locali 9425 2105 9425 2105 7 FreeSans 400 0 -200 0 I_IN
port 7 w
flabel locali 10005 2140 10005 2140 3 FreeSans 400 0 200 0 x
port 3 e
flabel poly 10610 2010 10610 2010 3 FreeSans 400 0 200 0 DOWN_input
port 9 e
flabel metal1 9155 1715 9155 1715 7 FreeSans 400 0 -200 0 GNDA
port 2 w
flabel locali 10545 2095 10545 2095 3 FreeSans 400 0 160 0 vout
port 4 e
flabel metal2 9105 2830 9105 2830 7 FreeSans 400 0 -200 0 UP_b
port 5 w
flabel metal2 9105 1640 9105 1640 7 FreeSans 400 0 -200 0 DOWN
port 6 w
<< end >>
