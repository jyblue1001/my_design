** sch_path: /foss/designs/my_design/projects/opamp/xschem_ngspice/vds_vgs_sweep_pfet_2.sch
**.subckt vds_vgs_sweep_pfet_2
VGS GND VGS 1.05
VDS GND VDS 1.8
XM1 VDS VGS GND GND sky130_fd_pr__pfet_01v8 L=0.15 W=30 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 VDS VGS GND GND sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=4 m=4
**** begin user architecture code
.lib /foss/pdks/sky130A/libs.tech/combined/sky130.lib.spice tt



.option method=gear
.option wnflag=1
.option savecurrents
*.temp = 120

.save
+@m.xm1.msky130_fd_pr__pfet_01v8[gm]
+@m.xm1.msky130_fd_pr__pfet_01v8[vth]
+@m.xm2.msky130_fd_pr__pfet_01v8[gm]
+@m.xm2.msky130_fd_pr__pfet_01v8[vth]
+@m.xm3.msky130_fd_pr__pfet_01v8[gm]
+@m.xm4.msky130_fd_pr__pfet_01v8[gm]
+@m.xm5.msky130_fd_pr__pfet_01v8[gm]
+@m.xm6.msky130_fd_pr__pfet_01v8[gm]
+@m.xm7.msky130_fd_pr__pfet_01v8[gm]
+@m.xm8.msky130_fd_pr__pfet_01v8[gm]
+@m.xm9.msky130_fd_pr__pfet_01v8[gm]
+@m.xm10.msky130_fd_pr__pfet_01v8[gm]


.control
  save all
  * dc VGS 0 1.8 0.1 VDS 0 1.8 0.1
  * dc VDS 0 1.0 0.001 VGS 0.6 1.3 0.01
  dc VDS 0.1 0.9 0.001 VGS 0.3 1.6 0.01
  remzerovec
  write vds_vgs_sweep_pfet_2.raw
  set appendwrite
  let rout = deriv(vds)/deriv(@m.xm10.msky130_fd_pr__pfet_01v8[id])
  save rout
  show
.endc



**** end user architecture code
**.ends
.GLOBAL GND
.end
