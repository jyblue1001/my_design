* PEX produced on Mon Feb  3 03:58:52 AM CET 2025 using /foss/tools/osic-multitool/iic-pex.sh with m=3 and s=1
* NGSPICE file created from TSPC_FF_ratioed_divide120_magic.ext - technology: sky130A

.subckt TSPC_FF_ratioed_divide120_magic VOUT VIN VDDA GNDA
X0 VDDA.t66 div2.t2 div2_3_1.A.t1 VDDA.t65 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X1 div5_0.A.t2 div5_0.Q2_b.t2 VDDA.t60 VDDA.t59 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X2 div2_3_0.C.t2 div2_3_0.CLK.t3 GNDA.t30 GNDA.t29 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X3 div2.t1 div2_3_1.C.t4 GNDA.t23 GNDA.t22 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X4 div5_0.H.t1 div24.t3 div5_0.G.t2 GNDA.t40 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X5 div2_3_0.A.t0 div2_3_0.CLK.t4 div2_3_0.B.t0 GNDA.t28 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X6 GNDA.t27 div2_3_0.CLK.t5 div2_3_0.C.t1 GNDA.t26 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X7 VDDA.t64 div2.t3 div2_3_2.CLK.t2 VDDA.t63 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X8 GNDA.t3 div3_2_0.I.t2 div3_2_0.G.t1 GNDA.t2 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X9 VDDA.t18 div3_2_0.I.t3 div24.t0 VDDA.t17 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X10 div5_0.G.t0 VOUT.t2 div5_0.F.t1 VDDA.t12 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X11 div2_3_0.CLK.t0 div4.t2 VDDA.t14 VDDA.t13 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X12 div2_3_0.B.t1 div8.t2 GNDA.t36 GNDA.t35 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X13 div3_2_0.G.t0 div3_2_0.D.t2 div3_2_0.F.t1 GNDA.t10 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X14 VDDA.t38 div3_2_0.E.t3 div3_2_0.H.t3 VDDA.t37 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X15 VDDA.t1 div5_0.Q2_b.t3 div5_0.G.t1 VDDA.t0 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X16 GNDA.t58 div2_3_1.CLK.t3 div2_3_1.C.t1 GNDA.t57 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X17 GNDA.t71 div4.t3 div2_3_0.CLK.t1 GNDA.t70 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X18 div3_2_0.D.t1 div3_2_0.C.t4 GNDA.t42 GNDA.t41 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X19 div24.t2 div3_2_0.I.t4 GNDA.t44 GNDA.t43 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X20 div5_0.D.t0 div5_0.B.t2 VDDA.t20 VDDA.t19 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X21 div3_2_0.F.t0 div3_2_0.CLK.t3 div3_2_0.E.t0 GNDA.t21 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X22 div2_3_1.C.t3 div2_3_1.CLK.t4 GNDA.t93 GNDA.t92 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X23 VDDA.t72 div8.t3 div2_3_0.A.t1 VDDA.t71 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X24 GNDA.t54 div3_2_0.CLK.t4 div3_2_0.C.t2 GNDA.t53 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X25 div5_0.M.t0 div5_0.K.t2 VDDA.t24 VDDA.t23 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X26 VDDA.t34 div8.t4 div3_2_0.CLK.t2 VDDA.t33 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X27 div2_3_2.C.t0 div2_3_2.A.t2 VDDA.t36 VDDA.t35 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X28 div3_2_0.C.t0 div3_2_0.A.t2 VDDA.t9 VDDA.t8 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X29 GNDA.t56 div2_3_1.CLK.t5 div2_3_1.C.t0 GNDA.t55 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X30 div5_0.K.t0 div5_0.Q2_b.t4 div5_0.L.t0 GNDA.t89 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X31 VDDA.t70 VIN.t0 div2_3_1.CLK.t2 VDDA.t69 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X32 div2_3_1.C.t2 div2_3_1.A.t2 VDDA.t68 VDDA.t67 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X33 GNDA.t95 div2_3_2.CLK.t3 div2_3_2.C.t3 GNDA.t94 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X34 div3_2_0.C.t1 div3_2_0.CLK.t5 GNDA.t48 GNDA.t47 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X35 div3_2_0.D.t0 div3_2_0.CLK.t6 VDDA.t42 VDDA.t41 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X36 VDDA.t54 div3_2_0.D.t3 div3_2_0.E.t1 VDDA.t53 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X37 div4.t0 div2_3_2.C.t4 GNDA.t12 GNDA.t11 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X38 div5_0.J.t3 div24.t4 GNDA.t1 GNDA.t0 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X39 div4.t1 div2_3_2.CLK.t4 VDDA.t16 VDDA.t15 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X40 VDDA.t48 div5_0.G.t3 div5_0.J.t0 VDDA.t47 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X41 div5_0.L.t1 VOUT.t3 GNDA.t69 GNDA.t68 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X42 GNDA.t50 div2_3_2.CLK.t5 div2_3_2.C.t2 GNDA.t49 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X43 GNDA.t61 div3_2_0.CLK.t7 div3_2_0.C.t3 GNDA.t60 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X44 div5_0.A.t0 div5_0.Q2_b.t5 GNDA.t88 GNDA.t87 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X45 div5_0.Q2_b.t0 div5_0.J.t4 GNDA.t16 GNDA.t15 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X46 div3_2_0.CLK.t1 div8.t5 VDDA.t58 VDDA.t57 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X47 VDDA.t52 div5_0.Q2_b.t6 div5_0.A.t1 VDDA.t51 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X48 div5_0.B.t1 div24.t5 div5_0.C.t1 GNDA.t39 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X49 GNDA.t34 div24.t6 div5_0.J.t2 GNDA.t33 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X50 div2_3_1.A.t0 div2_3_1.CLK.t6 div2_3_1.B.t0 GNDA.t6 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X51 div2_3_2.C.t1 div2_3_2.CLK.t6 GNDA.t9 GNDA.t8 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X52 GNDA.t99 div24.t7 div5_0.J.t1 GNDA.t98 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X53 div2_3_2.A.t1 div2_3_2.CLK.t7 div2_3_2.B.t1 GNDA.t7 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X54 GNDA.t63 div8.t6 div3_2_0.CLK.t0 GNDA.t62 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X55 VOUT.t1 div5_0.Q2_b.t7 VDDA.t50 VDDA.t49 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X56 div5_0.C.t0 div5_0.A.t3 GNDA.t91 GNDA.t90 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X57 VDDA.t32 div24.t8 div3_2_0.A.t1 VDDA.t31 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X58 div2_3_1.B.t1 div2.t4 GNDA.t79 GNDA.t78 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X59 GNDA.t73 div3_2_0.CLK.t8 div3_2_0.H.t2 GNDA.t72 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X60 div5_0.E.t0 div5_0.D.t4 GNDA.t46 GNDA.t45 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X61 div5_0.M.t3 div5_0.Q2_b.t8 GNDA.t86 GNDA.t85 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X62 div24.t1 div3_2_0.I.t5 VDDA.t40 VDDA.t39 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X63 div5_0.F.t0 div5_0.E.t2 VDDA.t3 VDDA.t2 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X64 VDDA.t74 div4.t4 div2_3_0.CLK.t2 VDDA.t73 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X65 div2_3_2.B.t0 div4.t5 GNDA.t14 GNDA.t13 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X66 div3_2_0.A.t0 div3_2_0.CLK.t9 div3_2_0.B.t0 GNDA.t59 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X67 GNDA.t97 div24.t9 div5_0.D.t3 GNDA.t96 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X68 GNDA.t84 div5_0.Q2_b.t9 div5_0.M.t2 GNDA.t83 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X69 div2.t0 div2_3_1.CLK.t7 VDDA.t28 VDDA.t27 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X70 div2_3_0.C.t3 div2_3_0.A.t2 VDDA.t76 VDDA.t75 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X71 GNDA.t67 VIN.t1 div2_3_1.CLK.t1 GNDA.t66 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X72 div3_2_0.H.t0 div3_2_0.CLK.t10 GNDA.t20 GNDA.t19 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X73 div5_0.I.t2 VOUT.t4 GNDA.t65 GNDA.t64 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X74 VDDA.t5 div5_0.A.t4 div5_0.B.t0 VDDA.t4 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X75 div5_0.E.t1 div24.t10 VDDA.t44 VDDA.t43 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X76 div2_3_2.CLK.t1 div2.t5 VDDA.t62 VDDA.t61 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X77 div8.t0 div2_3_0.CLK.t6 VDDA.t11 VDDA.t10 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X78 GNDA.t77 div2.t6 div2_3_2.CLK.t0 GNDA.t76 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X79 div8.t1 div2_3_0.C.t4 GNDA.t32 GNDA.t31 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X80 div3_2_0.B.t1 div24.t11 GNDA.t75 GNDA.t74 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X81 div5_0.D.t2 div24.t12 GNDA.t103 GNDA.t102 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X82 div2_3_1.CLK.t0 VIN.t2 VDDA.t30 VDDA.t29 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X83 div3_2_0.I.t1 div3_2_0.H.t4 GNDA.t38 GNDA.t37 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X84 GNDA.t5 div5_0.E.t3 div5_0.I.t0 GNDA.t4 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X85 VOUT.t0 div5_0.M.t4 GNDA.t18 GNDA.t17 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X86 GNDA.t52 div3_2_0.CLK.t11 div3_2_0.H.t1 GNDA.t51 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X87 VDDA.t26 VOUT.t5 div5_0.K.t1 VDDA.t25 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X88 GNDA.t101 div24.t13 div5_0.D.t1 GNDA.t100 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X89 div3_2_0.E.t2 div3_2_0.I.t6 VDDA.t56 VDDA.t55 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X90 GNDA.t25 div2_3_0.CLK.t7 div2_3_0.C.t0 GNDA.t24 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X91 div5_0.Q2_b.t1 div24.t14 VDDA.t46 VDDA.t45 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X92 div5_0.I.t1 div5_0.Q2_b.t10 div5_0.H.t0 GNDA.t82 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X93 GNDA.t81 div5_0.Q2_b.t11 div5_0.M.t1 GNDA.t80 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X94 VDDA.t7 div4.t6 div2_3_2.A.t0 VDDA.t6 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X95 div3_2_0.I.t0 div3_2_0.CLK.t12 VDDA.t22 VDDA.t21 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
R0 div2.t2 div2.t4 819.4
R1 div2.n0 div2.t0 663.801
R2 div2.n0 div2.t2 489.168
R3 div2.t3 div2.t5 401.668
R4 div2.n1 div2.t1 270.12
R5 div2.n2 div2.t3 257.067
R6 div2_3_2.VIN div2.n2 216.9
R7 div2.n2 div2.t6 208.868
R8 div2.n3 div2_3_2.VIN 192.167
R9 div2.n1 div2.n0 67.2005
R10 div2.n3 div2.n1 25.6005
R11 div2_3_1.VOUT div2.n3 4.8005
R12 div2_3_1.A.n0 div2_3_1.A.t1 713.933
R13 div2_3_1.A.n0 div2_3_1.A.t2 314.233
R14 div2_3_1.A.t0 div2_3_1.A.n0 308.2
R15 VDDA.t43 VDDA.t0 2804.76
R16 VDDA.t45 VDDA.t25 2533.33
R17 VDDA.t53 VDDA.t41 2307.14
R18 VDDA.t39 VDDA.t21 2126.19
R19 VDDA.t10 VDDA.t33 2080.95
R20 VDDA.t73 VDDA.t15 2080.95
R21 VDDA.t27 VDDA.t63 2080.95
R22 VDDA.t4 VDDA.t59 1538.1
R23 VDDA.t12 VDDA.t47 1492.86
R24 VDDA.t37 VDDA.t55 1492.86
R25 VDDA.t23 VDDA.n15 1289.29
R26 VDDA.n16 VDDA.t19 1289.29
R27 VDDA.t51 VDDA.t17 1130.95
R28 VDDA.t57 VDDA.t31 1130.95
R29 VDDA.t71 VDDA.t13 1130.95
R30 VDDA.t61 VDDA.t6 1130.95
R31 VDDA.t65 VDDA.t29 1130.95
R32 VDDA.t8 VDDA.n36 927.381
R33 VDDA.n37 VDDA.t75 927.381
R34 VDDA.t35 VDDA.n51 927.381
R35 VDDA.n52 VDDA.t67 927.381
R36 VDDA.n24 VDDA.t40 673.101
R37 VDDA.n23 VDDA.t18 673.101
R38 VDDA.n14 VDDA.t50 667.62
R39 VDDA.n1 VDDA.t28 663.801
R40 VDDA.n2 VDDA.t16 663.801
R41 VDDA.n4 VDDA.t11 663.801
R42 VDDA.n5 VDDA.t42 663.801
R43 VDDA.n7 VDDA.t44 663.801
R44 VDDA.n15 VDDA.t49 610.715
R45 VDDA.n16 VDDA.t43 610.715
R46 VDDA.n36 VDDA.t41 610.715
R47 VDDA.n37 VDDA.t10 610.715
R48 VDDA.n51 VDDA.t15 610.715
R49 VDDA.n52 VDDA.t27 610.715
R50 VDDA.n58 VDDA.n57 594.301
R51 VDDA.n56 VDDA.n55 594.301
R52 VDDA.n46 VDDA.n45 594.301
R53 VDDA.n48 VDDA.n47 594.301
R54 VDDA.n43 VDDA.n42 594.301
R55 VDDA.n41 VDDA.n40 594.301
R56 VDDA.n31 VDDA.n30 594.301
R57 VDDA.n33 VDDA.n32 594.301
R58 VDDA.n28 VDDA.n27 594.301
R59 VDDA.n26 VDDA.n25 594.301
R60 VDDA.n22 VDDA.n21 594.301
R61 VDDA.n20 VDDA.n19 594.301
R62 VDDA.n9 VDDA.n8 594.301
R63 VDDA.n11 VDDA.n10 594.301
R64 VDDA.n13 VDDA.n12 594.301
R65 VDDA.t25 VDDA.t23 497.62
R66 VDDA.t47 VDDA.t45 497.62
R67 VDDA.t2 VDDA.t12 497.62
R68 VDDA.t0 VDDA.t2 497.62
R69 VDDA.t19 VDDA.t4 497.62
R70 VDDA.t59 VDDA.t51 497.62
R71 VDDA.t17 VDDA.t39 497.62
R72 VDDA.t21 VDDA.t37 497.62
R73 VDDA.t55 VDDA.t53 497.62
R74 VDDA.t31 VDDA.t8 497.62
R75 VDDA.t33 VDDA.t57 497.62
R76 VDDA.t75 VDDA.t71 497.62
R77 VDDA.t13 VDDA.t73 497.62
R78 VDDA.t6 VDDA.t35 497.62
R79 VDDA.t63 VDDA.t61 497.62
R80 VDDA.t67 VDDA.t65 497.62
R81 VDDA.t29 VDDA.t69 497.62
R82 VDDA.n15 VDDA.n14 373.781
R83 VDDA.n17 VDDA.n16 370
R84 VDDA.n36 VDDA.n35 370
R85 VDDA.n38 VDDA.n37 370
R86 VDDA.n51 VDDA.n50 370
R87 VDDA.n53 VDDA.n52 370
R88 VDDA.n57 VDDA.t30 78.8005
R89 VDDA.n57 VDDA.t70 78.8005
R90 VDDA.n55 VDDA.t68 78.8005
R91 VDDA.n55 VDDA.t66 78.8005
R92 VDDA.n45 VDDA.t62 78.8005
R93 VDDA.n45 VDDA.t64 78.8005
R94 VDDA.n47 VDDA.t36 78.8005
R95 VDDA.n47 VDDA.t7 78.8005
R96 VDDA.n42 VDDA.t14 78.8005
R97 VDDA.n42 VDDA.t74 78.8005
R98 VDDA.n40 VDDA.t76 78.8005
R99 VDDA.n40 VDDA.t72 78.8005
R100 VDDA.n30 VDDA.t58 78.8005
R101 VDDA.n30 VDDA.t34 78.8005
R102 VDDA.n32 VDDA.t9 78.8005
R103 VDDA.n32 VDDA.t32 78.8005
R104 VDDA.n27 VDDA.t56 78.8005
R105 VDDA.n27 VDDA.t54 78.8005
R106 VDDA.n25 VDDA.t22 78.8005
R107 VDDA.n25 VDDA.t38 78.8005
R108 VDDA.n21 VDDA.t60 78.8005
R109 VDDA.n21 VDDA.t52 78.8005
R110 VDDA.n19 VDDA.t20 78.8005
R111 VDDA.n19 VDDA.t5 78.8005
R112 VDDA.n8 VDDA.t3 78.8005
R113 VDDA.n8 VDDA.t1 78.8005
R114 VDDA.n10 VDDA.t46 78.8005
R115 VDDA.n10 VDDA.t48 78.8005
R116 VDDA.n12 VDDA.t24 78.8005
R117 VDDA.n12 VDDA.t26 78.8005
R118 VDDA.n53 VDDA.n1 12.8005
R119 VDDA.n50 VDDA.n2 12.8005
R120 VDDA.n38 VDDA.n4 12.8005
R121 VDDA.n35 VDDA.n5 12.8005
R122 VDDA.n17 VDDA.n7 12.8005
R123 VDDA.n7 VDDA.n6 9.3005
R124 VDDA.n18 VDDA.n17 9.3005
R125 VDDA.n29 VDDA.n5 9.3005
R126 VDDA.n35 VDDA.n34 9.3005
R127 VDDA.n4 VDDA.n3 9.3005
R128 VDDA.n39 VDDA.n38 9.3005
R129 VDDA.n44 VDDA.n2 9.3005
R130 VDDA.n50 VDDA.n49 9.3005
R131 VDDA.n1 VDDA.n0 9.3005
R132 VDDA.n54 VDDA.n53 9.3005
R133 VDDA.n14 VDDA.n13 3.20124
R134 VDDA.n9 VDDA.n6 0.913
R135 VDDA.n13 VDDA.n11 0.838
R136 VDDA.n29 VDDA.n28 0.7755
R137 VDDA.n11 VDDA.n9 0.688
R138 VDDA.n26 VDDA.n24 0.588
R139 VDDA.n22 VDDA.n20 0.563
R140 VDDA.n28 VDDA.n26 0.5505
R141 VDDA VDDA.n3 0.4755
R142 VDDA.n44 VDDA 0.4755
R143 VDDA VDDA.n0 0.4755
R144 VDDA.n33 VDDA.n31 0.4505
R145 VDDA.n43 VDDA.n41 0.4505
R146 VDDA.n48 VDDA.n46 0.4505
R147 VDDA.n58 VDDA.n56 0.4505
R148 VDDA.n20 VDDA.n18 0.4255
R149 VDDA.n34 VDDA.n33 0.3255
R150 VDDA.n41 VDDA.n39 0.3255
R151 VDDA.n49 VDDA.n48 0.3255
R152 VDDA.n56 VDDA.n54 0.3255
R153 VDDA.n24 VDDA.n23 0.2755
R154 VDDA VDDA.n22 0.238
R155 VDDA.n31 VDDA 0.238
R156 VDDA VDDA.n43 0.238
R157 VDDA.n46 VDDA 0.238
R158 VDDA VDDA.n58 0.238
R159 VDDA.n18 VDDA.n6 0.1005
R160 VDDA.n34 VDDA.n29 0.1005
R161 VDDA.n39 VDDA.n3 0.1005
R162 VDDA.n49 VDDA.n44 0.1005
R163 VDDA.n54 VDDA.n0 0.1005
R164 VDDA.n23 VDDA 0.0755
R165 div5_0.Q2_b.n6 div5_0.Q2_b.t5 2779.53
R166 div5_0.Q2_b.n7 div5_0.Q2_b.n6 1206
R167 div5_0.Q2_b.n4 div5_0.Q2_b.t1 777.4
R168 div5_0.Q2_b.t10 div5_0.Q2_b.t3 514.134
R169 div5_0.Q2_b.n3 div5_0.Q2_b.n2 364.178
R170 div5_0.Q2_b.n0 div5_0.Q2_b.t7 353.467
R171 div5_0.Q2_b.t5 div5_0.Q2_b.n5 353.467
R172 div5_0.Q2_b.n5 div5_0.Q2_b.t2 289.2
R173 div5_0.Q2_b.n4 div5_0.Q2_b.n3 257.079
R174 div5_0.Q2_b.t0 div5_0.Q2_b.n7 233
R175 div5_0.Q2_b.n6 div5_0.Q2_b.t10 208.868
R176 div5_0.Q2_b.n0 div5_0.Q2_b.t11 192.8
R177 div5_0.Q2_b.n2 div5_0.Q2_b.n1 176.733
R178 div5_0.Q2_b.n2 div5_0.Q2_b.t9 112.468
R179 div5_0.Q2_b.n1 div5_0.Q2_b.t8 112.468
R180 div5_0.Q2_b.n3 div5_0.Q2_b.t4 112.468
R181 div5_0.Q2_b.n5 div5_0.Q2_b.t6 112.468
R182 div5_0.Q2_b.n1 div5_0.Q2_b.n0 96.4005
R183 div5_0.Q2_b.n7 div5_0.Q2_b.n4 21.3338
R184 div5_0.A.n2 div5_0.A.t1 755.534
R185 div5_0.A.t2 div5_0.A.n2 685.134
R186 div5_0.A.n1 div5_0.A.n0 389.733
R187 div5_0.A.n1 div5_0.A.t0 340.2
R188 div5_0.A.n0 div5_0.A.t3 321.334
R189 div5_0.A.n0 div5_0.A.t4 144.601
R190 div5_0.A.n2 div5_0.A.n1 19.2005
R191 div2_3_0.CLK.n5 div2_3_0.CLK.t2 723.534
R192 div2_3_0.CLK.n4 div2_3_0.CLK.t0 723.534
R193 div2_3_0.CLK.n0 div2_3_0.CLK.t6 369.534
R194 div2_3_0.CLK.n3 div2_3_0.CLK.n2 366.856
R195 div2_3_0.CLK.t1 div2_3_0.CLK.n5 254.333
R196 div2_3_0.CLK.n3 div2_3_0.CLK.t4 190.123
R197 div2_3_0.CLK.n4 div2_3_0.CLK.n3 187.201
R198 div2_3_0.CLK.n1 div2_3_0.CLK.n0 176.733
R199 div2_3_0.CLK.n2 div2_3_0.CLK.n1 176.733
R200 div2_3_0.CLK.n0 div2_3_0.CLK.t7 112.468
R201 div2_3_0.CLK.n2 div2_3_0.CLK.t5 112.468
R202 div2_3_0.CLK.n1 div2_3_0.CLK.t3 112.468
R203 div2_3_0.CLK.n5 div2_3_0.CLK.n4 70.4005
R204 GNDA.t66 GNDA.t17 1.00944e+06
R205 GNDA.t43 GNDA.t87 3600
R206 GNDA.t40 GNDA.t45 3500
R207 GNDA.t68 GNDA.t15 3400
R208 GNDA.t33 GNDA.t64 3300
R209 GNDA.t21 GNDA.t41 3300
R210 GNDA.t60 GNDA.t59 3300
R211 GNDA.t28 GNDA.t26 3300
R212 GNDA.t94 GNDA.t7 3300
R213 GNDA.t55 GNDA.t6 3300
R214 GNDA.n51 GNDA.t87 3150
R215 GNDA.t83 GNDA.t89 2500
R216 GNDA.t100 GNDA.t39 2500
R217 GNDA.t37 GNDA.t43 2500
R218 GNDA.n40 GNDA.t51 1950
R219 GNDA.t62 GNDA.n39 1950
R220 GNDA.n39 GNDA.t31 1950
R221 GNDA.n30 GNDA.t70 1950
R222 GNDA.n30 GNDA.t11 1950
R223 GNDA.n52 GNDA.t76 1950
R224 GNDA.n52 GNDA.t22 1950
R225 GNDA.t90 GNDA.n51 1350
R226 GNDA.n40 GNDA.t2 1350
R227 GNDA.n39 GNDA.n38 1179.3
R228 GNDA.n31 GNDA.n30 1179.3
R229 GNDA.n53 GNDA.n52 1179.3
R230 GNDA.n41 GNDA.n40 1170
R231 GNDA.n51 GNDA.n50 1170
R232 GNDA.t17 GNDA.t80 1100
R233 GNDA.t80 GNDA.t85 1100
R234 GNDA.t85 GNDA.t83 1100
R235 GNDA.t89 GNDA.t68 1100
R236 GNDA.t15 GNDA.t98 1100
R237 GNDA.t98 GNDA.t0 1100
R238 GNDA.t0 GNDA.t33 1100
R239 GNDA.t64 GNDA.t4 1100
R240 GNDA.t4 GNDA.t82 1100
R241 GNDA.t82 GNDA.t40 1100
R242 GNDA.t45 GNDA.t96 1100
R243 GNDA.t96 GNDA.t102 1100
R244 GNDA.t102 GNDA.t100 1100
R245 GNDA.t39 GNDA.t90 1100
R246 GNDA.t72 GNDA.t37 1100
R247 GNDA.t19 GNDA.t72 1100
R248 GNDA.t51 GNDA.t19 1100
R249 GNDA.t2 GNDA.t10 1100
R250 GNDA.t10 GNDA.t21 1100
R251 GNDA.t41 GNDA.t53 1100
R252 GNDA.t53 GNDA.t47 1100
R253 GNDA.t47 GNDA.t60 1100
R254 GNDA.t59 GNDA.t74 1100
R255 GNDA.t74 GNDA.t62 1100
R256 GNDA.t24 GNDA.t31 1100
R257 GNDA.t29 GNDA.t24 1100
R258 GNDA.t26 GNDA.t29 1100
R259 GNDA.t35 GNDA.t28 1100
R260 GNDA.t70 GNDA.t35 1100
R261 GNDA.t11 GNDA.t49 1100
R262 GNDA.t49 GNDA.t8 1100
R263 GNDA.t8 GNDA.t94 1100
R264 GNDA.t7 GNDA.t13 1100
R265 GNDA.t13 GNDA.t76 1100
R266 GNDA.t22 GNDA.t57 1100
R267 GNDA.t57 GNDA.t92 1100
R268 GNDA.t92 GNDA.t55 1100
R269 GNDA.t6 GNDA.t78 1100
R270 GNDA.t78 GNDA.t66 1100
R271 GNDA.n47 GNDA.t44 242.3
R272 GNDA.n48 GNDA.t88 242.3
R273 GNDA.n4 GNDA.t69 242.3
R274 GNDA.n17 GNDA.t3 233
R275 GNDA.n0 GNDA.t91 233
R276 GNDA.n3 GNDA.n1 194.576
R277 GNDA.n59 GNDA.n58 194.3
R278 GNDA.n57 GNDA.n56 194.3
R279 GNDA.n55 GNDA.n54 194.3
R280 GNDA.n25 GNDA.n24 194.3
R281 GNDA.n27 GNDA.n26 194.3
R282 GNDA.n29 GNDA.n28 194.3
R283 GNDA.n33 GNDA.n32 194.3
R284 GNDA.n35 GNDA.n34 194.3
R285 GNDA.n37 GNDA.n36 194.3
R286 GNDA.n23 GNDA.n22 194.3
R287 GNDA.n21 GNDA.n20 194.3
R288 GNDA.n19 GNDA.n18 194.3
R289 GNDA.n44 GNDA.n43 194.3
R290 GNDA.n46 GNDA.n45 194.3
R291 GNDA.n14 GNDA.n13 194.3
R292 GNDA.n12 GNDA.n11 194.3
R293 GNDA.n10 GNDA.n9 194.3
R294 GNDA.n8 GNDA.n7 194.3
R295 GNDA.n6 GNDA.n5 194.3
R296 GNDA.n3 GNDA.n2 194.3
R297 GNDA.n58 GNDA.t79 48.0005
R298 GNDA.n58 GNDA.t67 48.0005
R299 GNDA.n56 GNDA.t93 48.0005
R300 GNDA.n56 GNDA.t56 48.0005
R301 GNDA.n54 GNDA.t23 48.0005
R302 GNDA.n54 GNDA.t58 48.0005
R303 GNDA.n24 GNDA.t14 48.0005
R304 GNDA.n24 GNDA.t77 48.0005
R305 GNDA.n26 GNDA.t9 48.0005
R306 GNDA.n26 GNDA.t95 48.0005
R307 GNDA.n28 GNDA.t12 48.0005
R308 GNDA.n28 GNDA.t50 48.0005
R309 GNDA.n32 GNDA.t36 48.0005
R310 GNDA.n32 GNDA.t71 48.0005
R311 GNDA.n34 GNDA.t30 48.0005
R312 GNDA.n34 GNDA.t27 48.0005
R313 GNDA.n36 GNDA.t32 48.0005
R314 GNDA.n36 GNDA.t25 48.0005
R315 GNDA.n22 GNDA.t75 48.0005
R316 GNDA.n22 GNDA.t63 48.0005
R317 GNDA.n20 GNDA.t48 48.0005
R318 GNDA.n20 GNDA.t61 48.0005
R319 GNDA.n18 GNDA.t42 48.0005
R320 GNDA.n18 GNDA.t54 48.0005
R321 GNDA.n43 GNDA.t20 48.0005
R322 GNDA.n43 GNDA.t52 48.0005
R323 GNDA.n45 GNDA.t38 48.0005
R324 GNDA.n45 GNDA.t73 48.0005
R325 GNDA.n13 GNDA.t103 48.0005
R326 GNDA.n13 GNDA.t101 48.0005
R327 GNDA.n11 GNDA.t46 48.0005
R328 GNDA.n11 GNDA.t97 48.0005
R329 GNDA.n9 GNDA.t65 48.0005
R330 GNDA.n9 GNDA.t5 48.0005
R331 GNDA.n7 GNDA.t1 48.0005
R332 GNDA.n7 GNDA.t34 48.0005
R333 GNDA.n5 GNDA.t16 48.0005
R334 GNDA.n5 GNDA.t99 48.0005
R335 GNDA.n2 GNDA.t86 48.0005
R336 GNDA.n2 GNDA.t84 48.0005
R337 GNDA.n1 GNDA.t18 48.0005
R338 GNDA.n1 GNDA.t81 48.0005
R339 GNDA.n41 GNDA.n17 12.8005
R340 GNDA.n50 GNDA.n0 12.8005
R341 GNDA.n15 GNDA.n0 9.3005
R342 GNDA.n50 GNDA.n49 9.3005
R343 GNDA.n42 GNDA.n41 9.3005
R344 GNDA.n17 GNDA.n16 9.3005
R345 GNDA.n12 GNDA.n10 0.8505
R346 GNDA.n19 GNDA.n16 0.8255
R347 GNDA.n23 GNDA.n21 0.688
R348 GNDA.n35 GNDA.n33 0.688
R349 GNDA.n27 GNDA.n25 0.688
R350 GNDA.n59 GNDA.n57 0.688
R351 GNDA.n4 GNDA.n3 0.588
R352 GNDA.n15 GNDA.n14 0.588
R353 GNDA.n10 GNDA.n8 0.5505
R354 GNDA.n49 GNDA.n48 0.463
R355 GNDA.n6 GNDA.n4 0.4255
R356 GNDA GNDA.n47 0.3505
R357 GNDA.n47 GNDA.n46 0.313
R358 GNDA.n44 GNDA.n42 0.313
R359 GNDA.n38 GNDA.n37 0.313
R360 GNDA.n31 GNDA.n29 0.313
R361 GNDA.n55 GNDA.n53 0.313
R362 GNDA.n8 GNDA.n6 0.2755
R363 GNDA.n14 GNDA.n12 0.2755
R364 GNDA.n46 GNDA.n44 0.2755
R365 GNDA.n21 GNDA.n19 0.2755
R366 GNDA.n37 GNDA.n35 0.2755
R367 GNDA.n29 GNDA.n27 0.2755
R368 GNDA.n57 GNDA.n55 0.2755
R369 GNDA GNDA.n23 0.238
R370 GNDA.n33 GNDA 0.238
R371 GNDA.n25 GNDA 0.238
R372 GNDA GNDA.n59 0.238
R373 GNDA.n49 GNDA.n15 0.1005
R374 GNDA.n48 GNDA 0.1005
R375 GNDA.n42 GNDA.n16 0.1005
R376 GNDA.n38 GNDA 0.0755
R377 GNDA GNDA.n31 0.0755
R378 GNDA.n53 GNDA 0.0755
R379 div2_3_0.C.n0 div2_3_0.C.t3 721.4
R380 div2_3_0.C.n1 div2_3_0.C.t4 349.433
R381 div2_3_0.C.n0 div2_3_0.C.t1 276.733
R382 div2_3_0.C.n2 div2_3_0.C.n1 206.333
R383 div2_3_0.C.n1 div2_3_0.C.n0 48.0005
R384 div2_3_0.C.n2 div2_3_0.C.t0 48.0005
R385 div2_3_0.C.t2 div2_3_0.C.n2 48.0005
R386 div2_3_1.C.n2 div2_3_1.C.t2 721.4
R387 div2_3_1.C.n1 div2_3_1.C.t4 349.433
R388 div2_3_1.C.t0 div2_3_1.C.n2 276.733
R389 div2_3_1.C.n1 div2_3_1.C.n0 206.333
R390 div2_3_1.C.n0 div2_3_1.C.t1 48.0005
R391 div2_3_1.C.n0 div2_3_1.C.t3 48.0005
R392 div2_3_1.C.n2 div2_3_1.C.n1 48.0005
R393 div24.n10 div24.t11 4546.23
R394 div24.n3 div24.n2 919.244
R395 div3_2_0.VOUT div24.n7 886.702
R396 div24.t11 div24.t8 819.4
R397 div24.n2 div24.n1 758.606
R398 div24.n9 div24.n8 628.734
R399 div24.n7 div24.n6 364.178
R400 div24.n0 div24.t14 337.401
R401 div24.n0 div24.t7 305.267
R402 div24.n9 div24.t2 257.534
R403 div24.n4 div24.t9 192.8
R404 div24.n1 div24.n0 176.733
R405 div24.n6 div24.n5 176.733
R406 div24.n4 div24.n3 160.667
R407 div24.n3 div24.t10 144.601
R408 div24.n2 div24.t3 131.976
R409 div24.n0 div24.t4 128.534
R410 div24.n1 div24.t6 128.534
R411 div24.n6 div24.t13 112.468
R412 div24.n5 div24.t12 112.468
R413 div24.n7 div24.t5 112.468
R414 div24.n5 div24.n4 96.4005
R415 div24.n8 div24.t0 78.8005
R416 div24.n8 div24.t1 78.8005
R417 div5_0.VIN div24.n10 28.8005
R418 div24.n10 div24.n9 9.6005
R419 div5_0.VIN div3_2_0.VOUT 6.4005
R420 div5_0.G.n0 div5_0.G.t0 685.134
R421 div5_0.G.n1 div5_0.G.t1 685.134
R422 div5_0.G.n0 div5_0.G.t3 534.268
R423 div5_0.G.t2 div5_0.G.n1 340.521
R424 div5_0.G.n1 div5_0.G.n0 105.6
R425 div5_0.H.t0 div5_0.H.t1 96.0005
R426 div2_3_0.B.t0 div2_3_0.B.t1 96.0005
R427 div2_3_0.A.n0 div2_3_0.A.t1 713.933
R428 div2_3_0.A.n0 div2_3_0.A.t2 314.233
R429 div2_3_0.A.t0 div2_3_0.A.n0 308.2
R430 div2_3_2.CLK.n4 div2_3_2.CLK.t1 723.534
R431 div2_3_2.CLK.t2 div2_3_2.CLK.n5 723.534
R432 div2_3_2.CLK.n0 div2_3_2.CLK.t4 369.534
R433 div2_3_2.CLK.n3 div2_3_2.CLK.n2 366.856
R434 div2_3_2.CLK.n5 div2_3_2.CLK.t0 254.333
R435 div2_3_2.CLK.n3 div2_3_2.CLK.t7 190.123
R436 div2_3_2.CLK.n4 div2_3_2.CLK.n3 187.201
R437 div2_3_2.CLK.n1 div2_3_2.CLK.n0 176.733
R438 div2_3_2.CLK.n2 div2_3_2.CLK.n1 176.733
R439 div2_3_2.CLK.n0 div2_3_2.CLK.t5 112.468
R440 div2_3_2.CLK.n2 div2_3_2.CLK.t3 112.468
R441 div2_3_2.CLK.n1 div2_3_2.CLK.t6 112.468
R442 div2_3_2.CLK.n5 div2_3_2.CLK.n4 70.4005
R443 div3_2_0.I.n0 div3_2_0.I.t0 663.801
R444 div3_2_0.I.n0 div3_2_0.I.t6 568.067
R445 div3_2_0.I.t6 div3_2_0.I.t2 514.134
R446 div3_2_0.I.n3 div3_2_0.I.n2 344.8
R447 div3_2_0.I.n1 div3_2_0.I.t3 289.2
R448 div3_2_0.I.t1 div3_2_0.I.n3 275.454
R449 div3_2_0.I.n2 div3_2_0.I.t4 241
R450 div3_2_0.I.n1 div3_2_0.I.t5 112.468
R451 div3_2_0.I.n3 div3_2_0.I.n0 97.9205
R452 div3_2_0.I.n2 div3_2_0.I.n1 64.2672
R453 div3_2_0.G.t0 div3_2_0.G.t1 96.0005
R454 VOUT.n2 VOUT.n1 2120.39
R455 VOUT.n1 VOUT.t2 1992.27
R456 VOUT.n3 VOUT.t1 751.801
R457 VOUT.t2 VOUT.t4 514.134
R458 VOUT.n0 VOUT.t3 289.2
R459 VOUT.n2 VOUT.t0 233
R460 VOUT.n1 VOUT.n0 208.868
R461 VOUT.n0 VOUT.t5 176.733
R462 VOUT.n3 VOUT.n2 40.3205
R463 VOUT VOUT.n3 32.0005
R464 div5_0.F.t0 div5_0.F.t1 157.601
R465 div4.t6 div4.t5 819.4
R466 div4.n0 div4.t1 663.801
R467 div4.n0 div4.t6 489.168
R468 div4.t4 div4.t2 401.668
R469 div4.n1 div4.t0 270.12
R470 div4.n2 div4.t4 257.067
R471 div2_3_0.VIN div4.n2 216.9
R472 div4.n2 div4.t3 208.868
R473 div4.n3 div2_3_0.VIN 192.167
R474 div4.n1 div4.n0 67.2005
R475 div4.n3 div4.n1 25.6005
R476 div2_3_2.VOUT div4.n3 4.8005
R477 div8.t3 div8.t2 819.4
R478 div8.n0 div8.t0 663.801
R479 div8.n0 div8.t3 489.168
R480 div8.t4 div8.t5 401.668
R481 div8.n1 div8.t1 270.12
R482 div8.n2 div8.t4 257.067
R483 div3_2_0.VIN div8.n2 216.9
R484 div8.n2 div8.t6 208.868
R485 div8.n3 div3_2_0.VIN 192.167
R486 div8.n1 div8.n0 67.2005
R487 div8.n3 div8.n1 25.6005
R488 div2_3_0.VOUT div8.n3 4.8005
R489 div3_2_0.D.n1 div3_2_0.D.n0 701.467
R490 div3_2_0.D.n1 div3_2_0.D.t0 694.201
R491 div3_2_0.D.n0 div3_2_0.D.t2 321.334
R492 div3_2_0.D.t1 div3_2_0.D.n1 314.921
R493 div3_2_0.D.n0 div3_2_0.D.t3 144.601
R494 div3_2_0.F.t0 div3_2_0.F.t1 96.0005
R495 div3_2_0.E.n0 div3_2_0.E.t2 685.134
R496 div3_2_0.E.n1 div3_2_0.E.t1 663.801
R497 div3_2_0.E.n0 div3_2_0.E.t3 534.268
R498 div3_2_0.E.t0 div3_2_0.E.n1 362.921
R499 div3_2_0.E.n1 div3_2_0.E.n0 91.7338
R500 div3_2_0.H.n0 div3_2_0.H.t3 723.534
R501 div3_2_0.H.n1 div3_2_0.H.t4 553.534
R502 div3_2_0.H.n0 div3_2_0.H.t1 254.333
R503 div3_2_0.H.n2 div3_2_0.H.n1 206.333
R504 div3_2_0.H.n1 div3_2_0.H.n0 70.4005
R505 div3_2_0.H.n2 div3_2_0.H.t2 48.0005
R506 div3_2_0.H.t0 div3_2_0.H.n2 48.0005
R507 div2_3_1.CLK.n5 div2_3_1.CLK.t2 723.534
R508 div2_3_1.CLK.n4 div2_3_1.CLK.t0 723.534
R509 div2_3_1.CLK.n0 div2_3_1.CLK.t7 369.534
R510 div2_3_1.CLK.n3 div2_3_1.CLK.n2 366.856
R511 div2_3_1.CLK.t1 div2_3_1.CLK.n5 254.333
R512 div2_3_1.CLK.n3 div2_3_1.CLK.t6 190.123
R513 div2_3_1.CLK.n4 div2_3_1.CLK.n3 187.201
R514 div2_3_1.CLK.n1 div2_3_1.CLK.n0 176.733
R515 div2_3_1.CLK.n2 div2_3_1.CLK.n1 176.733
R516 div2_3_1.CLK.n0 div2_3_1.CLK.t3 112.468
R517 div2_3_1.CLK.n2 div2_3_1.CLK.t5 112.468
R518 div2_3_1.CLK.n1 div2_3_1.CLK.t4 112.468
R519 div2_3_1.CLK.n5 div2_3_1.CLK.n4 70.4005
R520 div3_2_0.C.n0 div3_2_0.C.t0 721.4
R521 div3_2_0.C.n1 div3_2_0.C.t4 350.349
R522 div3_2_0.C.n0 div3_2_0.C.t3 276.733
R523 div3_2_0.C.n2 div3_2_0.C.n1 206.333
R524 div3_2_0.C.n1 div3_2_0.C.n0 48.0005
R525 div3_2_0.C.n2 div3_2_0.C.t2 48.0005
R526 div3_2_0.C.t1 div3_2_0.C.n2 48.0005
R527 div5_0.B.n0 div5_0.B.t0 663.801
R528 div5_0.B.n0 div5_0.B.t2 380.368
R529 div5_0.B div5_0.B.t1 282.921
R530 div5_0.B div5_0.B.n0 114.133
R531 div5_0.D.n0 div5_0.D.t0 761.4
R532 div5_0.D.n1 div5_0.D.t4 350.349
R533 div5_0.D.n0 div5_0.D.t1 254.333
R534 div5_0.D.n2 div5_0.D.n1 206.333
R535 div5_0.D.n1 div5_0.D.n0 70.4005
R536 div5_0.D.t3 div5_0.D.n2 48.0005
R537 div5_0.D.n2 div5_0.D.t2 48.0005
R538 div3_2_0.CLK.n3 div3_2_0.CLK.n2 742.51
R539 div3_2_0.CLK.n8 div3_2_0.CLK.t1 723.534
R540 div3_2_0.CLK.t2 div3_2_0.CLK.n9 723.534
R541 div3_2_0.CLK.n2 div3_2_0.CLK.n1 684.806
R542 div3_2_0.CLK.n7 div3_2_0.CLK.n6 366.856
R543 div3_2_0.CLK.n0 div3_2_0.CLK.t12 337.401
R544 div3_2_0.CLK.n0 div3_2_0.CLK.t8 305.267
R545 div3_2_0.CLK.n9 div3_2_0.CLK.t0 254.333
R546 div3_2_0.CLK.n4 div3_2_0.CLK.n3 224.934
R547 div3_2_0.CLK.n7 div3_2_0.CLK.t9 190.123
R548 div3_2_0.CLK.n8 div3_2_0.CLK.n7 187.201
R549 div3_2_0.CLK.n1 div3_2_0.CLK.n0 176.733
R550 div3_2_0.CLK.n5 div3_2_0.CLK.n4 176.733
R551 div3_2_0.CLK.n6 div3_2_0.CLK.n5 176.733
R552 div3_2_0.CLK.n3 div3_2_0.CLK.t6 144.601
R553 div3_2_0.CLK.n2 div3_2_0.CLK.t3 131.976
R554 div3_2_0.CLK.n0 div3_2_0.CLK.t10 128.534
R555 div3_2_0.CLK.n1 div3_2_0.CLK.t11 128.534
R556 div3_2_0.CLK.n4 div3_2_0.CLK.t4 112.468
R557 div3_2_0.CLK.n6 div3_2_0.CLK.t7 112.468
R558 div3_2_0.CLK.n5 div3_2_0.CLK.t5 112.468
R559 div3_2_0.CLK.n9 div3_2_0.CLK.n8 70.4005
R560 div5_0.K.n0 div5_0.K.t1 663.801
R561 div5_0.K.t0 div5_0.K.n0 397.053
R562 div5_0.K.n0 div5_0.K.t2 380.368
R563 div5_0.M.n0 div5_0.M.t0 761.4
R564 div5_0.M.n1 div5_0.M.t4 349.433
R565 div5_0.M.n0 div5_0.M.t2 254.333
R566 div5_0.M.n2 div5_0.M.n1 206.333
R567 div5_0.M.n1 div5_0.M.n0 70.4005
R568 div5_0.M.n2 div5_0.M.t1 48.0005
R569 div5_0.M.t3 div5_0.M.n2 48.0005
R570 div2_3_2.A.n0 div2_3_2.A.t0 713.933
R571 div2_3_2.A.n0 div2_3_2.A.t2 314.233
R572 div2_3_2.A.t1 div2_3_2.A.n0 308.2
R573 div2_3_2.C.n2 div2_3_2.C.t0 721.4
R574 div2_3_2.C.n1 div2_3_2.C.t4 349.433
R575 div2_3_2.C.t3 div2_3_2.C.n2 276.733
R576 div2_3_2.C.n1 div2_3_2.C.n0 206.333
R577 div2_3_2.C.n0 div2_3_2.C.t2 48.0005
R578 div2_3_2.C.n0 div2_3_2.C.t1 48.0005
R579 div2_3_2.C.n2 div2_3_2.C.n1 48.0005
R580 div3_2_0.A.n0 div3_2_0.A.t1 713.933
R581 div3_2_0.A.n0 div3_2_0.A.t2 314.233
R582 div3_2_0.A.t0 div3_2_0.A.n0 308.2
R583 div5_0.L.t0 div5_0.L.t1 96.0005
R584 VIN.t0 VIN.t2 401.668
R585 VIN.n0 VIN.t0 257.067
R586 VIN VIN.n0 216.9
R587 VIN.n0 VIN.t1 208.868
R588 div5_0.J.n0 div5_0.J.t0 723.534
R589 div5_0.J.n1 div5_0.J.t4 553.534
R590 div5_0.J.n0 div5_0.J.t2 254.333
R591 div5_0.J.n2 div5_0.J.n1 206.333
R592 div5_0.J.n1 div5_0.J.n0 70.4005
R593 div5_0.J.n2 div5_0.J.t1 48.0005
R594 div5_0.J.t3 div5_0.J.n2 48.0005
R595 div5_0.C.t0 div5_0.C.t1 96.0005
R596 div2_3_1.B.t0 div2_3_1.B.t1 96.0005
R597 div2_3_2.B.t0 div2_3_2.B.t1 96.0005
R598 div5_0.E.n0 div5_0.E.t2 1207.57
R599 div5_0.E.n0 div5_0.E.t1 723
R600 div5_0.E.t2 div5_0.E.t3 514.134
R601 div5_0.E.t0 div5_0.E.n0 314.921
R602 div3_2_0.B.t0 div3_2_0.B.t1 96.0005
R603 div5_0.I.n0 div5_0.I.t2 531.067
R604 div5_0.I.t0 div5_0.I.n0 48.0005
R605 div5_0.I.n0 div5_0.I.t1 48.0005
C0 VDDA VIN 0.125773f
C1 div5_0.B VDDA 0.308332f
C2 VOUT VDDA 0.659192f
C3 VOUT GNDA 1.87185f
C4 VIN GNDA 0.304628f
C5 VDDA GNDA 10.4898f
C6 div5_0.B GNDA 0.250854f
.ends

