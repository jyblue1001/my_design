* PEX produced on Sun Aug 24 11:20:01 PM CEST 2025 using /foss/tools/osic-multitool/iic-pex.sh with m=3 and s=1
* NGSPICE file created from bgr_opamp_dummy_magic_19.ext - technology: sky130A

.subckt bgr_opamp_dummy_magic_19 VDDA GNDA VOUT+ VOUT- VIN+ VIN- GNDA_2 VDDA_2
X0 VDDA.t217 bgr_11_0.1st_Vout_2.t7 bgr_11_0.PFET_GATE_10uA.t5 VDDA.t216 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X1 VOUT+.t19 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t143 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2 VOUT+.t20 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t142 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3 VOUT+.t21 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t141 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4 VOUT+.t22 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t140 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5 GNDA_2.t163 GNDA_2.t161 two_stage_opamp_dummy_magic_29_0.Vb2.t3 GNDA_2.t162 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X6 VDDA.t20 two_stage_opamp_dummy_magic_29_0.Y.t25 VOUT+.t0 VDDA.t19 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X7 VDDA.t111 two_stage_opamp_dummy_magic_29_0.Y.t26 VOUT+.t5 VDDA.t110 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X8 GNDA_2.t278 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.t2 VOUT-.t9 GNDA_2.t277 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X9 two_stage_opamp_dummy_magic_29_0.Vb2_2.t9 two_stage_opamp_dummy_magic_29_0.Vb2.t8 two_stage_opamp_dummy_magic_29_0.Vb2.t9 two_stage_opamp_dummy_magic_29_0.Vb2_2.t8 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X10 VOUT+.t23 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t139 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X11 VDDA.t368 bgr_11_0.V_TOP.t14 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref.t3 VDDA.t367 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X12 VOUT-.t19 two_stage_opamp_dummy_magic_29_0.cap_res_X.t142 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X13 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.t10 two_stage_opamp_dummy_magic_29_0.X.t25 GNDA_2.t180 VDDA.t75 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X14 bgr_11_0.1st_Vout_1.t7 bgr_11_0.cap_res1.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X15 VOUT+.t24 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t138 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X16 VOUT-.t20 two_stage_opamp_dummy_magic_29_0.cap_res_X.t141 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X17 two_stage_opamp_dummy_magic_29_0.Vb2.t5 bgr_11_0.NFET_GATE_10uA.t5 GNDA_2.t232 GNDA_2.t231 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X18 VOUT-.t21 two_stage_opamp_dummy_magic_29_0.cap_res_X.t140 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X19 bgr_11_0.V_TOP.t15 VDDA.t369 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X20 GNDA_2.t36 bgr_11_0.NFET_GATE_10uA.t6 two_stage_opamp_dummy_magic_29_0.Vb2.t1 GNDA_2.t35 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X21 two_stage_opamp_dummy_magic_29_0.Y.t17 two_stage_opamp_dummy_magic_29_0.Vb2.t11 two_stage_opamp_dummy_magic_29_0.VD4.t31 two_stage_opamp_dummy_magic_29_0.VD4.t30 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X22 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.t13 two_stage_opamp_dummy_magic_29_0.X.t26 VDDA.t73 GNDA_2.t178 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X23 VOUT+.t25 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t137 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X24 VOUT+.t26 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t136 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X25 VOUT+.t27 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t135 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X26 bgr_11_0.START_UP_NFET1.t0 bgr_11_0.START_UP_NFET1 GNDA_2.t49 GNDA_2.t48 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X27 bgr_11_0.1st_Vout_1.t0 bgr_11_0.V_mir1.t13 VDDA.t8 VDDA.t7 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X28 VOUT-.t22 two_stage_opamp_dummy_magic_29_0.cap_res_X.t139 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X29 VOUT+.t28 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t134 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X30 VOUT-.t23 two_stage_opamp_dummy_magic_29_0.cap_res_X.t138 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X31 VOUT+.t29 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t133 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X32 two_stage_opamp_dummy_magic_29_0.Vb1_2.t3 two_stage_opamp_dummy_magic_29_0.Vb1.t9 two_stage_opamp_dummy_magic_29_0.Vb1.t10 GNDA_2.t106 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X33 two_stage_opamp_dummy_magic_29_0.VD2.t15 two_stage_opamp_dummy_magic_29_0.Vb1.t12 two_stage_opamp_dummy_magic_29_0.Y.t7 GNDA_2.t229 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X34 VOUT+.t30 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t132 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X35 two_stage_opamp_dummy_magic_29_0.VD3.t36 two_stage_opamp_dummy_magic_29_0.Vb2.t12 two_stage_opamp_dummy_magic_29_0.X.t17 two_stage_opamp_dummy_magic_29_0.VD3.t35 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X36 VOUT-.t24 two_stage_opamp_dummy_magic_29_0.cap_res_X.t137 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X37 two_stage_opamp_dummy_magic_29_0.VD4.t5 two_stage_opamp_dummy_magic_29_0.Vb3.t8 VDDA.t117 VDDA.t116 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X38 bgr_11_0.V_TOP.t16 VDDA.t87 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X39 VOUT-.t25 two_stage_opamp_dummy_magic_29_0.cap_res_X.t136 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X40 VDDA.t45 two_stage_opamp_dummy_magic_29_0.X.t27 VOUT-.t1 VDDA.t44 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X41 VOUT+.t31 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t131 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X42 VOUT-.t26 two_stage_opamp_dummy_magic_29_0.cap_res_X.t135 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X43 VOUT+.t32 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t130 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X44 a_6350_30238.t0 bgr_11_0.Vin+.t4 GNDA_2.t16 sky130_fd_pr__res_xhigh_po_0p35 l=6
X45 VDDA.t36 two_stage_opamp_dummy_magic_29_0.Vb3.t9 two_stage_opamp_dummy_magic_29_0.VD3.t1 VDDA.t35 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X46 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.t16 two_stage_opamp_dummy_magic_29_0.Y.t27 GNDA_2.t236 VDDA.t165 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X47 VOUT-.t27 two_stage_opamp_dummy_magic_29_0.cap_res_X.t134 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X48 VOUT-.t28 two_stage_opamp_dummy_magic_29_0.cap_res_X.t133 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X49 VOUT+.t33 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t129 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X50 bgr_11_0.V_TOP.t17 VDDA.t88 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X51 two_stage_opamp_dummy_magic_29_0.V_err_gate.t2 bgr_11_0.NFET_GATE_10uA.t7 GNDA_2.t291 GNDA_2.t290 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X52 VDDA.t377 a_6540_22450.t11 a_6540_22450.t12 VDDA.t376 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X53 VOUT-.t29 two_stage_opamp_dummy_magic_29_0.cap_res_X.t132 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X54 VDDA.t197 bgr_11_0.V_mir1.t11 bgr_11_0.V_mir1.t12 VDDA.t196 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X55 VOUT+.t34 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t128 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X56 VOUT+.t35 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t127 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X57 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.t14 two_stage_opamp_dummy_magic_29_0.Y.t28 VDDA.t153 GNDA_2.t228 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X58 two_stage_opamp_dummy_magic_29_0.VD2.t0 VIN+.t0 two_stage_opamp_dummy_magic_29_0.V_source.t37 GNDA_2.t25 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X59 VOUT+.t36 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t126 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X60 VOUT+.t37 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t125 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X61 VOUT+.t38 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t124 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X62 VOUT+.t39 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t123 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X63 VOUT-.t30 two_stage_opamp_dummy_magic_29_0.cap_res_X.t131 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X64 two_stage_opamp_dummy_magic_29_0.V_source.t12 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t12 GNDA_2.t63 GNDA_2.t6 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X65 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.t4 bgr_11_0.PFET_GATE_10uA.t10 VDDA.t253 VDDA.t252 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X66 VOUT-.t31 two_stage_opamp_dummy_magic_29_0.cap_res_X.t130 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X67 VDDA.t251 bgr_11_0.PFET_GATE_10uA.t11 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.t3 VDDA.t250 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X68 bgr_11_0.V_TOP.t18 VDDA.t81 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X69 bgr_11_0.cap_res1.t20 bgr_11_0.V_TOP.t13 GNDA_2.t284 sky130_fd_pr__res_high_po_0p35 l=2.05
X70 two_stage_opamp_dummy_magic_29_0.VD3.t34 two_stage_opamp_dummy_magic_29_0.Vb2.t13 two_stage_opamp_dummy_magic_29_0.X.t15 two_stage_opamp_dummy_magic_29_0.VD3.t33 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X71 VOUT-.t32 two_stage_opamp_dummy_magic_29_0.cap_res_X.t129 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X72 VOUT+.t40 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t122 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X73 a_14420_3878.t1 two_stage_opamp_dummy_magic_29_0.V_tot.t3 GNDA_2.t289 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X74 VOUT+.t41 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t121 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X75 VDDA.t390 two_stage_opamp_dummy_magic_29_0.Y.t29 VOUT+.t15 VDDA.t389 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X76 VOUT-.t33 two_stage_opamp_dummy_magic_29_0.cap_res_X.t128 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X77 VOUT+.t42 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t120 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X78 VOUT-.t34 two_stage_opamp_dummy_magic_29_0.cap_res_X.t127 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X79 bgr_11_0.V_TOP.t19 VDDA.t82 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X80 VDDA.t363 VDDA.t361 two_stage_opamp_dummy_magic_29_0.VD3.t16 VDDA.t362 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X81 bgr_11_0.1st_Vout_2.t8 bgr_11_0.cap_res2.t20 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X82 GNDA_2.t73 GNDA_2.t160 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t7 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X83 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.t9 two_stage_opamp_dummy_magic_29_0.X.t28 GNDA_2.t211 VDDA.t113 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X84 VOUT+.t43 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t119 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X85 VOUT+.t44 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t118 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X86 VOUT-.t35 two_stage_opamp_dummy_magic_29_0.cap_res_X.t126 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X87 VDDA.t411 two_stage_opamp_dummy_magic_29_0.Y.t30 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.t13 GNDA_2.t288 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X88 VOUT+.t45 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t117 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X89 GNDA_2.t64 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t13 two_stage_opamp_dummy_magic_29_0.V_source.t13 GNDA_2.t6 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X90 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.t12 two_stage_opamp_dummy_magic_29_0.X.t29 VDDA.t131 GNDA_2.t220 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X91 GNDA_2.t57 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t14 two_stage_opamp_dummy_magic_29_0.V_source.t11 GNDA_2.t6 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X92 VDDA.t215 bgr_11_0.1st_Vout_2.t9 bgr_11_0.PFET_GATE_10uA.t3 VDDA.t214 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X93 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t0 two_stage_opamp_dummy_magic_29_0.Y.t2 GNDA_2.t54 sky130_fd_pr__res_high_po_1p41 l=1.41
X94 bgr_11_0.1st_Vout_2.t10 bgr_11_0.cap_res2.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X95 two_stage_opamp_dummy_magic_29_0.Vb1.t4 two_stage_opamp_dummy_magic_29_0.Vb1.t3 two_stage_opamp_dummy_magic_29_0.Vb1_2.t2 GNDA_2.t106 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X96 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t11 bgr_11_0.PFET_GATE_10uA.t12 VDDA.t249 VDDA.t248 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X97 two_stage_opamp_dummy_magic_29_0.VD2.t14 two_stage_opamp_dummy_magic_29_0.Vb1.t13 two_stage_opamp_dummy_magic_29_0.Y.t1 GNDA_2.t43 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X98 VOUT-.t36 two_stage_opamp_dummy_magic_29_0.cap_res_X.t125 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X99 VOUT+.t46 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t116 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X100 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t8 bgr_11_0.Vin+.t5 GNDA_2.t276 sky130_fd_pr__res_xhigh_po_0p35 l=2.3
X101 VOUT+.t47 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t115 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X102 bgr_11_0.1st_Vout_1.t8 bgr_11_0.cap_res1.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X103 VDDA.t49 two_stage_opamp_dummy_magic_29_0.X.t30 VOUT-.t2 VDDA.t48 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X104 bgr_11_0.1st_Vout_2.t11 bgr_11_0.cap_res2.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X105 VOUT+.t48 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t114 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X106 bgr_11_0.V_TOP.t20 VDDA.t395 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X107 VOUT+.t49 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t113 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X108 VOUT+.t50 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t112 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X109 VDDA.t247 bgr_11_0.PFET_GATE_10uA.t13 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.t14 VDDA.t246 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X110 VOUT+.t51 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t111 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X111 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.t16 VDDA.t358 VDDA.t360 VDDA.t359 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X112 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.t15 two_stage_opamp_dummy_magic_29_0.Y.t31 GNDA_2.t58 VDDA.t52 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X113 GNDA_2.t159 GNDA_2.t157 VOUT+.t14 GNDA_2.t158 sky130_fd_pr__nfet_01v8 ad=2.8 pd=14.8 as=1.4 ps=7.4 w=7 l=0.6
X114 VOUT+.t52 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t110 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X115 VOUT+.t53 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t109 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X116 VDDA.t127 a_6540_22450.t13 bgr_11_0.1st_Vout_2.t3 VDDA.t126 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X117 VDDA.t397 bgr_11_0.V_TOP.t21 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref.t2 VDDA.t396 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X118 a_3230_3878.t0 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.t0 GNDA_2.t169 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X119 VOUT-.t37 two_stage_opamp_dummy_magic_29_0.cap_res_X.t124 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X120 two_stage_opamp_dummy_magic_29_0.VD2.t5 VIN+.t1 two_stage_opamp_dummy_magic_29_0.V_source.t36 GNDA_2.t183 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X121 VOUT-.t38 two_stage_opamp_dummy_magic_29_0.cap_res_X.t123 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X122 VOUT-.t8 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.t3 GNDA_2.t283 GNDA_2.t282 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X123 two_stage_opamp_dummy_magic_29_0.V_source.t25 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t15 GNDA_2.t239 GNDA_2.t238 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X124 VOUT-.t39 two_stage_opamp_dummy_magic_29_0.cap_res_X.t122 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X125 VOUT+.t54 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t108 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X126 two_stage_opamp_dummy_magic_29_0.Vb2_2.t5 two_stage_opamp_dummy_magic_29_0.Vb2_2.t3 two_stage_opamp_dummy_magic_29_0.Vb2_2.t5 two_stage_opamp_dummy_magic_29_0.Vb2_2.t4 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0 ps=0 w=3.5 l=0.2
X127 VOUT-.t40 two_stage_opamp_dummy_magic_29_0.cap_res_X.t121 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X128 VOUT+.t55 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t107 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X129 bgr_11_0.1st_Vout_2.t12 bgr_11_0.cap_res2.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X130 VOUT-.t41 two_stage_opamp_dummy_magic_29_0.cap_res_X.t120 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X131 VDDA.t124 two_stage_opamp_dummy_magic_29_0.Y.t32 VOUT+.t6 VDDA.t123 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X132 VOUT+.t56 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t106 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X133 bgr_11_0.V_TOP.t22 VDDA.t379 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X134 VOUT-.t42 two_stage_opamp_dummy_magic_29_0.cap_res_X.t119 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X135 two_stage_opamp_dummy_magic_29_0.err_amp_out.t3 two_stage_opamp_dummy_magic_29_0.err_amp_mir.t5 GNDA_2.t187 GNDA_2.t52 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X136 VOUT+.t57 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t105 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X137 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref.t6 VDDA.t355 VDDA.t357 VDDA.t356 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=1.2 ps=6.8 w=3 l=0.5
X138 GNDA_2.t210 two_stage_opamp_dummy_magic_29_0.Y.t33 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.t14 VDDA.t112 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X139 two_stage_opamp_dummy_magic_29_0.VD4.t37 two_stage_opamp_dummy_magic_29_0.VD4.t35 two_stage_opamp_dummy_magic_29_0.Y.t24 two_stage_opamp_dummy_magic_29_0.VD4.t36 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X140 VOUT-.t43 two_stage_opamp_dummy_magic_29_0.cap_res_X.t118 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X141 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.t8 two_stage_opamp_dummy_magic_29_0.X.t31 GNDA_2.t33 VDDA.t32 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X142 VOUT+.t4 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.t4 GNDA_2.t186 GNDA_2.t185 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X143 GNDA_2.t222 bgr_11_0.NFET_GATE_10uA.t8 two_stage_opamp_dummy_magic_29_0.Vb3.t5 GNDA_2.t221 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X144 two_stage_opamp_dummy_magic_29_0.VD1.t19 two_stage_opamp_dummy_magic_29_0.Vb1.t14 two_stage_opamp_dummy_magic_29_0.X.t11 GNDA_2.t235 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X145 VDDA.t78 a_6540_22450.t9 a_6540_22450.t10 VDDA.t77 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X146 VOUT-.t44 two_stage_opamp_dummy_magic_29_0.cap_res_X.t117 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X147 GNDA_2.t212 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t16 two_stage_opamp_dummy_magic_29_0.V_source.t21 GNDA_2.t6 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X148 bgr_11_0.START_UP.t3 bgr_11_0.V_TOP.t23 VDDA.t381 VDDA.t380 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X149 VOUT+.t58 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t104 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X150 VDDA.t354 VDDA.t352 two_stage_opamp_dummy_magic_29_0.VD4.t11 VDDA.t353 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X151 two_stage_opamp_dummy_magic_29_0.X.t16 two_stage_opamp_dummy_magic_29_0.Vb2.t14 two_stage_opamp_dummy_magic_29_0.VD3.t32 two_stage_opamp_dummy_magic_29_0.VD3.t31 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X152 VOUT-.t45 two_stage_opamp_dummy_magic_29_0.cap_res_X.t116 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X153 a_11420_30238.t1 bgr_11_0.Vin-.t5 GNDA_2.t196 sky130_fd_pr__res_xhigh_po_0p35 l=6
X154 bgr_11_0.V_TOP.t12 VDDA.t349 VDDA.t351 VDDA.t350 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.45 ps=2.9 w=1 l=0.15
X155 VOUT-.t46 two_stage_opamp_dummy_magic_29_0.cap_res_X.t115 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X156 VOUT-.t47 two_stage_opamp_dummy_magic_29_0.cap_res_X.t114 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X157 GNDA_2.t191 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.t5 VOUT-.t7 GNDA_2.t190 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X158 GNDA_2.t195 a_11950_28880.t0 GNDA_2.t194 sky130_fd_pr__res_xhigh_po_0p35 l=4
X159 VOUT+.t59 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t103 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X160 two_stage_opamp_dummy_magic_29_0.VD2.t13 two_stage_opamp_dummy_magic_29_0.Vb1.t15 two_stage_opamp_dummy_magic_29_0.Y.t5 GNDA_2.t50 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X161 bgr_11_0.V_TOP.t24 VDDA.t101 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X162 VOUT+.t16 two_stage_opamp_dummy_magic_29_0.Y.t34 VDDA.t392 VDDA.t391 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X163 two_stage_opamp_dummy_magic_29_0.err_amp_out.t0 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref.t7 two_stage_opamp_dummy_magic_29_0.V_err_p.t0 VDDA.t378 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X164 two_stage_opamp_dummy_magic_29_0.VD1.t18 two_stage_opamp_dummy_magic_29_0.Vb1.t16 two_stage_opamp_dummy_magic_29_0.X.t4 GNDA_2.t61 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X165 bgr_11_0.Vin+.t3 bgr_11_0.V_TOP.t25 VDDA.t103 VDDA.t102 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X166 two_stage_opamp_dummy_magic_29_0.VD3.t9 two_stage_opamp_dummy_magic_29_0.Vb3.t10 VDDA.t84 VDDA.t83 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X167 VDDA.t130 two_stage_opamp_dummy_magic_29_0.X.t32 VOUT-.t11 VDDA.t129 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X168 VOUT-.t48 two_stage_opamp_dummy_magic_29_0.cap_res_X.t113 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X169 VDDA.t191 bgr_11_0.V_mir1.t14 bgr_11_0.1st_Vout_1.t6 VDDA.t190 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X170 two_stage_opamp_dummy_magic_29_0.VD1.t0 VIN-.t0 two_stage_opamp_dummy_magic_29_0.V_source.t3 GNDA_2.t15 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X171 VOUT+.t60 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t102 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X172 bgr_11_0.1st_Vout_2.t13 bgr_11_0.cap_res2.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X173 VDDA_2.t6 VDDA_2.t3 VDDA_2.t5 VDDA_2.t4 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0 ps=0 w=2 l=0.15
X174 VDDA.t348 VDDA.t345 VDDA.t347 VDDA.t346 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0 ps=0 w=1 l=0.15
X175 VDDA.t245 bgr_11_0.PFET_GATE_10uA.t14 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t10 VDDA.t244 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X176 two_stage_opamp_dummy_magic_29_0.VD2.t3 GNDA_2.t155 GNDA_2.t156 GNDA_2.t96 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X177 VOUT-.t49 two_stage_opamp_dummy_magic_29_0.cap_res_X.t112 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X178 VOUT-.t50 two_stage_opamp_dummy_magic_29_0.cap_res_X.t111 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X179 VOUT-.t51 two_stage_opamp_dummy_magic_29_0.cap_res_X.t110 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X180 VOUT+.t61 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t101 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X181 two_stage_opamp_dummy_magic_29_0.X.t20 two_stage_opamp_dummy_magic_29_0.Vb2.t15 two_stage_opamp_dummy_magic_29_0.VD3.t30 two_stage_opamp_dummy_magic_29_0.VD3.t29 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X182 VOUT+.t62 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t100 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X183 VOUT+.t63 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t99 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X184 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.t4 bgr_11_0.NFET_GATE_10uA.t9 GNDA_2.t56 GNDA_2.t55 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X185 GNDA_2.t154 GNDA_2.t153 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t2 GNDA_2.t24 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X186 two_stage_opamp_dummy_magic_29_0.VD1.t1 VIN-.t1 two_stage_opamp_dummy_magic_29_0.V_source.t4 GNDA_2.t24 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X187 VOUT-.t52 two_stage_opamp_dummy_magic_29_0.cap_res_X.t109 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X188 VOUT-.t53 two_stage_opamp_dummy_magic_29_0.cap_res_X.t108 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X189 two_stage_opamp_dummy_magic_29_0.Vb2.t6 bgr_11_0.NFET_GATE_10uA.t10 GNDA_2.t242 GNDA_2.t241 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X190 VDDA.t406 bgr_11_0.V_TOP.t26 bgr_11_0.Vin-.t3 VDDA.t405 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X191 VDDA.t344 VDDA.t342 bgr_11_0.V_TOP.t11 VDDA.t343 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.2
X192 VOUT+.t64 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t98 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X193 GNDA_2.t73 GNDA_2.t72 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t6 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X194 VOUT+.t65 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t97 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X195 bgr_11_0.1st_Vout_1.t9 bgr_11_0.cap_res1.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X196 GNDA_2.t76 GNDA_2.t75 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t5 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X197 VDDA.t69 bgr_11_0.1st_Vout_1.t10 bgr_11_0.V_TOP.t3 VDDA.t68 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X198 bgr_11_0.START_UP.t5 bgr_11_0.START_UP.t4 bgr_11_0.START_UP_NFET1.t0 GNDA_2.t29 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X199 VDDA.t136 two_stage_opamp_dummy_magic_29_0.Y.t35 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.t12 GNDA_2.t225 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X200 VOUT-.t54 two_stage_opamp_dummy_magic_29_0.cap_res_X.t107 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X201 VOUT-.t55 two_stage_opamp_dummy_magic_29_0.cap_res_X.t106 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X202 VOUT+.t66 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t96 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X203 VOUT+.t67 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t95 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X204 two_stage_opamp_dummy_magic_29_0.VD1.t17 two_stage_opamp_dummy_magic_29_0.Vb1.t17 two_stage_opamp_dummy_magic_29_0.X.t24 GNDA_2.t164 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X205 VOUT-.t56 two_stage_opamp_dummy_magic_29_0.cap_res_X.t105 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X206 VOUT+.t68 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t94 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X207 GNDA_2.t32 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t17 two_stage_opamp_dummy_magic_29_0.V_source.t5 GNDA_2.t6 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X208 bgr_11_0.NFET_GATE_10uA.t2 bgr_11_0.NFET_GATE_10uA.t1 GNDA_2.t38 GNDA_2.t37 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X209 VDDA.t408 bgr_11_0.V_TOP.t27 bgr_11_0.Vin+.t2 VDDA.t407 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X210 VOUT-.t57 two_stage_opamp_dummy_magic_29_0.cap_res_X.t104 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X211 bgr_11_0.1st_Vout_1.t11 bgr_11_0.cap_res1.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X212 VOUT+.t69 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t93 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X213 two_stage_opamp_dummy_magic_29_0.V_err_mir_p.t0 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref.t8 two_stage_opamp_dummy_magic_29_0.V_err_gate.t0 VDDA.t72 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X214 two_stage_opamp_dummy_magic_29_0.VD2.t12 two_stage_opamp_dummy_magic_29_0.Vb1.t18 two_stage_opamp_dummy_magic_29_0.Y.t10 GNDA_2.t3 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X215 bgr_11_0.V_TOP.t28 VDDA.t382 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X216 VDDA.t59 two_stage_opamp_dummy_magic_29_0.V_err_gate.t6 two_stage_opamp_dummy_magic_29_0.V_err_p.t3 VDDA.t58 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X217 two_stage_opamp_dummy_magic_29_0.VD1.t16 two_stage_opamp_dummy_magic_29_0.Vb1.t19 two_stage_opamp_dummy_magic_29_0.X.t1 GNDA_2.t3 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X218 GNDA_2.t73 GNDA_2.t152 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t4 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X219 GNDA_2.t151 GNDA_2.t149 GNDA_2.t151 GNDA_2.t150 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0 ps=0 w=2.5 l=0.15
X220 VDDA.t40 bgr_11_0.V_mir1.t9 bgr_11_0.V_mir1.t10 VDDA.t39 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X221 VOUT-.t58 two_stage_opamp_dummy_magic_29_0.cap_res_X.t103 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X222 GNDA_2.t148 GNDA_2.t145 GNDA_2.t147 GNDA_2.t146 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0 ps=0 w=1 l=0.15
X223 VDDA.t341 VDDA.t339 bgr_11_0.NFET_GATE_10uA.t4 VDDA.t340 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X224 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.t7 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.t4 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.t6 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.t5 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0 ps=0 w=3.5 l=0.2
X225 VOUT-.t59 two_stage_opamp_dummy_magic_29_0.cap_res_X.t102 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X226 bgr_11_0.1st_Vout_1.t12 bgr_11_0.cap_res1.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X227 a_3110_3878.t0 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.t1 GNDA_2.t168 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X228 VOUT+.t70 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t92 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X229 two_stage_opamp_dummy_magic_29_0.VD1.t4 VIN-.t2 two_stage_opamp_dummy_magic_29_0.V_source.t10 GNDA_2.t41 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X230 VOUT-.t60 two_stage_opamp_dummy_magic_29_0.cap_res_X.t101 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X231 VOUT+.t71 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t91 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X232 VDDA.t155 bgr_11_0.1st_Vout_1.t13 bgr_11_0.V_TOP.t6 VDDA.t154 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X233 VOUT-.t61 two_stage_opamp_dummy_magic_29_0.cap_res_X.t100 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X234 VOUT+.t72 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t90 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X235 VOUT-.t62 two_stage_opamp_dummy_magic_29_0.cap_res_X.t99 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X236 VOUT+.t73 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t89 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X237 VOUT+.t74 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t88 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X238 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.t1 a_13940_76.t1 GNDA_2.t215 sky130_fd_pr__res_xhigh_po_0p35 l=2.63
X239 VOUT-.t63 two_stage_opamp_dummy_magic_29_0.cap_res_X.t98 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X240 VOUT+.t75 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t87 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X241 VOUT+.t76 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t86 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X242 bgr_11_0.Vin+.t1 bgr_11_0.V_TOP.t29 VDDA.t384 VDDA.t383 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X243 VDDA.t93 two_stage_opamp_dummy_magic_29_0.X.t33 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.t11 GNDA_2.t199 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X244 two_stage_opamp_dummy_magic_29_0.VD1.t21 VIN-.t3 two_stage_opamp_dummy_magic_29_0.V_source.t39 GNDA_2.t24 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X245 VOUT-.t64 two_stage_opamp_dummy_magic_29_0.cap_res_X.t97 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X246 bgr_11_0.V_TOP.t30 VDDA.t143 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X247 two_stage_opamp_dummy_magic_29_0.Vb1.t1 GNDA_2.t143 GNDA_2.t144 GNDA_2.t106 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X248 bgr_11_0.PFET_GATE_10uA.t2 bgr_11_0.1st_Vout_2.t14 VDDA.t213 VDDA.t212 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X249 two_stage_opamp_dummy_magic_29_0.Vb2.t7 bgr_11_0.NFET_GATE_10uA.t11 GNDA_2.t253 GNDA_2.t252 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X250 VOUT+.t77 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t85 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X251 VOUT-.t65 two_stage_opamp_dummy_magic_29_0.cap_res_X.t96 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X252 bgr_11_0.1st_Vout_1.t14 bgr_11_0.cap_res1.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X253 GNDA_2.t275 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.t6 VOUT+.t13 GNDA_2.t274 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X254 VDDA.t366 bgr_11_0.V_mir1.t7 bgr_11_0.V_mir1.t8 VDDA.t365 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X255 two_stage_opamp_dummy_magic_29_0.VD4.t1 two_stage_opamp_dummy_magic_29_0.Vb3.t11 VDDA.t10 VDDA.t9 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X256 VOUT-.t66 two_stage_opamp_dummy_magic_29_0.cap_res_X.t95 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X257 VOUT-.t67 two_stage_opamp_dummy_magic_29_0.cap_res_X.t94 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X258 bgr_11_0.V_TOP.t31 VDDA.t144 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X259 GNDA_2.t0 two_stage_opamp_dummy_magic_29_0.Y.t36 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.t13 VDDA.t0 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X260 GNDA_2.t142 GNDA_2.t141 two_stage_opamp_dummy_magic_29_0.VD1.t6 GNDA_2.t87 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X261 VDDA.t211 bgr_11_0.1st_Vout_2.t15 bgr_11_0.PFET_GATE_10uA.t4 VDDA.t210 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X262 VOUT-.t68 two_stage_opamp_dummy_magic_29_0.cap_res_X.t93 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X263 VOUT+.t78 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t84 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X264 VOUT-.t69 two_stage_opamp_dummy_magic_29_0.cap_res_X.t92 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X265 VOUT+.t79 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t83 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X266 VDDA.t23 two_stage_opamp_dummy_magic_29_0.Y.t37 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.t11 GNDA_2.t22 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X267 VOUT+.t80 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t82 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X268 GNDA_2.t281 a_11300_28630.t1 GNDA_2.t280 sky130_fd_pr__res_xhigh_po_0p35 l=6
X269 GNDA_2.t273 bgr_11_0.NFET_GATE_10uA.t12 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.t3 GNDA_2.t272 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X270 VOUT-.t70 two_stage_opamp_dummy_magic_29_0.cap_res_X.t91 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X271 two_stage_opamp_dummy_magic_29_0.Vb2.t2 GNDA_2.t138 GNDA_2.t140 GNDA_2.t139 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X272 two_stage_opamp_dummy_magic_29_0.VD3.t28 two_stage_opamp_dummy_magic_29_0.Vb2.t16 two_stage_opamp_dummy_magic_29_0.X.t13 two_stage_opamp_dummy_magic_29_0.VD3.t27 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X273 GNDA_2.t47 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t18 two_stage_opamp_dummy_magic_29_0.V_p_mir.t1 GNDA_2.t46 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X274 GNDA_2.t137 GNDA_2.t136 two_stage_opamp_dummy_magic_29_0.VD2.t2 GNDA_2.t24 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X275 GNDA_2.t39 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t19 two_stage_opamp_dummy_magic_29_0.V_source.t7 GNDA_2.t6 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X276 VOUT+.t81 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t81 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X277 bgr_11_0.1st_Vout_2.t16 bgr_11_0.cap_res2.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X278 bgr_11_0.V_TOP.t32 VDDA.t104 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X279 VOUT+.t82 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t80 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X280 VOUT-.t71 two_stage_opamp_dummy_magic_29_0.cap_res_X.t90 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X281 VOUT-.t72 two_stage_opamp_dummy_magic_29_0.cap_res_X.t89 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X282 VDDA.t181 two_stage_opamp_dummy_magic_29_0.Vb3.t12 two_stage_opamp_dummy_magic_29_0.VD3.t13 VDDA.t180 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X283 VOUT+.t83 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t79 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X284 VOUT+.t8 two_stage_opamp_dummy_magic_29_0.Y.t38 VDDA.t138 VDDA.t137 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X285 bgr_11_0.V_p_1.t2 bgr_11_0.Vin+.t6 bgr_11_0.1st_Vout_1.t3 GNDA_2.t176 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=1 ps=5.8 w=2.5 l=0.2
X286 VOUT+.t84 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t78 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X287 VOUT-.t73 two_stage_opamp_dummy_magic_29_0.cap_res_X.t88 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X288 VOUT-.t10 a_13940_76.t0 GNDA_2.t209 sky130_fd_pr__res_xhigh_po_0p35 l=2.63
X289 VDDA.t63 a_6540_22450.t14 bgr_11_0.1st_Vout_2.t2 VDDA.t62 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X290 two_stage_opamp_dummy_magic_29_0.err_amp_mir.t1 VDDA.t336 VDDA.t338 VDDA.t337 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=1 ps=5.8 w=2.5 l=0.15
X291 two_stage_opamp_dummy_magic_29_0.VD1.t15 two_stage_opamp_dummy_magic_29_0.Vb1.t20 two_stage_opamp_dummy_magic_29_0.X.t0 GNDA_2.t3 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X292 bgr_11_0.1st_Vout_1.t15 bgr_11_0.cap_res1.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X293 GNDA_2.t53 two_stage_opamp_dummy_magic_29_0.err_amp_mir.t2 two_stage_opamp_dummy_magic_29_0.err_amp_mir.t3 GNDA_2.t52 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X294 two_stage_opamp_dummy_magic_29_0.V_source.t22 two_stage_opamp_dummy_magic_29_0.err_amp_out.t4 GNDA_2.t224 GNDA_2.t223 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X295 VOUT+.t18 GNDA_2.t133 GNDA_2.t135 GNDA_2.t134 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=2.8 ps=14.8 w=7 l=0.6
X296 VOUT+.t85 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t77 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X297 VOUT+.t86 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t76 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X298 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.t0 a_3830_76.t0 GNDA_2.t51 sky130_fd_pr__res_xhigh_po_0p35 l=2.63
X299 VOUT+.t87 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t75 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X300 VOUT+.t88 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t74 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X301 bgr_11_0.1st_Vout_2.t17 bgr_11_0.cap_res2.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X302 GNDA_2.t132 GNDA_2.t129 GNDA_2.t131 GNDA_2.t130 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0 ps=0 w=1 l=0.15
X303 GNDA_2.t181 two_stage_opamp_dummy_magic_29_0.X.t34 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.t7 VDDA.t76 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X304 VOUT+.t89 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t73 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X305 two_stage_opamp_dummy_magic_29_0.VD3.t8 two_stage_opamp_dummy_magic_29_0.VD3.t6 two_stage_opamp_dummy_magic_29_0.X.t2 two_stage_opamp_dummy_magic_29_0.VD3.t7 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X306 VOUT-.t74 two_stage_opamp_dummy_magic_29_0.cap_res_X.t87 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X307 two_stage_opamp_dummy_magic_29_0.X.t10 two_stage_opamp_dummy_magic_29_0.Vb1.t21 two_stage_opamp_dummy_magic_29_0.VD1.t14 GNDA_2.t177 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X308 VDDA.t94 two_stage_opamp_dummy_magic_29_0.X.t35 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.t10 GNDA_2.t202 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X309 bgr_11_0.1st_Vout_1.t16 bgr_11_0.cap_res1.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X310 a_5700_30088.t1 a_5820_28824.t1 GNDA_2.t189 sky130_fd_pr__res_xhigh_po_0p35 l=4.28
X311 VDDA.t55 two_stage_opamp_dummy_magic_29_0.X.t36 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.t9 GNDA_2.t62 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X312 VOUT+.t90 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t72 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X313 bgr_11_0.1st_Vout_2.t18 bgr_11_0.cap_res2.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X314 VDDA.t243 bgr_11_0.PFET_GATE_10uA.t15 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.t2 VDDA.t242 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X315 VOUT+.t91 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t71 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X316 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.t6 VDDA.t333 VDDA.t335 VDDA.t334 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X317 VOUT-.t75 two_stage_opamp_dummy_magic_29_0.cap_res_X.t86 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X318 two_stage_opamp_dummy_magic_29_0.VD1.t5 GNDA_2.t127 GNDA_2.t128 GNDA_2.t24 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X319 VOUT-.t76 two_stage_opamp_dummy_magic_29_0.cap_res_X.t85 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X320 a_6540_22450.t8 a_6540_22450.t7 VDDA.t163 VDDA.t162 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X321 VOUT+.t92 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t70 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X322 two_stage_opamp_dummy_magic_29_0.V_err_gate.t5 two_stage_opamp_dummy_magic_29_0.V_tot.t4 two_stage_opamp_dummy_magic_29_0.V_err_mir_p.t1 VDDA.t372 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X323 two_stage_opamp_dummy_magic_29_0.Y.t9 two_stage_opamp_dummy_magic_29_0.Vb1.t22 two_stage_opamp_dummy_magic_29_0.VD2.t11 GNDA_2.t3 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X324 VOUT-.t77 two_stage_opamp_dummy_magic_29_0.cap_res_X.t84 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X325 bgr_11_0.1st_Vout_1.t17 bgr_11_0.cap_res1.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X326 VOUT-.t78 two_stage_opamp_dummy_magic_29_0.cap_res_X.t83 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X327 bgr_11_0.1st_Vout_2.t19 bgr_11_0.cap_res2.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X328 VOUT+.t93 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t69 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X329 GNDA_2.t73 GNDA_2.t74 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t3 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X330 VOUT+.t94 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t68 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X331 VOUT-.t14 two_stage_opamp_dummy_magic_29_0.X.t37 VDDA.t176 VDDA.t175 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X332 VOUT+.t95 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t67 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X333 VOUT-.t79 two_stage_opamp_dummy_magic_29_0.cap_res_X.t82 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X334 VOUT+.t96 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t66 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X335 GNDA_2.t240 two_stage_opamp_dummy_magic_29_0.Y.t39 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.t12 VDDA.t174 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X336 VOUT+.t97 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t65 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X337 VDDA.t404 GNDA_2.t124 GNDA_2.t126 GNDA_2.t125 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=1.2 ps=6.8 w=3 l=0.15
X338 bgr_11_0.1st_Vout_2.t20 bgr_11_0.cap_res2.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X339 VDDA.t24 two_stage_opamp_dummy_magic_29_0.Y.t40 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.t10 GNDA_2.t23 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X340 GNDA_2.t123 GNDA_2.t120 GNDA_2.t122 GNDA_2.t121 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=0 ps=0 w=2.5 l=0.15
X341 two_stage_opamp_dummy_magic_29_0.V_source.t35 VIN+.t2 two_stage_opamp_dummy_magic_29_0.VD2.t18 GNDA_2.t24 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X342 VOUT-.t80 two_stage_opamp_dummy_magic_29_0.cap_res_X.t81 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X343 GNDA_2.t40 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t20 two_stage_opamp_dummy_magic_29_0.V_source.t8 GNDA_2.t6 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X344 VOUT-.t81 two_stage_opamp_dummy_magic_29_0.cap_res_X.t80 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X345 bgr_11_0.START_UP.t2 bgr_11_0.V_TOP.t33 VDDA.t106 VDDA.t105 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X346 VDDA.t332 VDDA.t330 VDDA.t332 VDDA.t331 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0 ps=0 w=1 l=0.15
X347 VOUT+.t98 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t64 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X348 bgr_11_0.1st_Vout_1.t18 bgr_11_0.cap_res1.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X349 VDDA.t16 bgr_11_0.V_mir1.t15 bgr_11_0.1st_Vout_1.t1 VDDA.t15 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X350 VDDA.t241 bgr_11_0.PFET_GATE_10uA.t16 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t9 VDDA.t240 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X351 bgr_11_0.cap_res2.t0 bgr_11_0.PFET_GATE_10uA.t0 GNDA_2.t188 sky130_fd_pr__res_high_po_0p35 l=2.05
X352 VOUT+.t99 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t63 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X353 bgr_11_0.V_TOP.t34 VDDA.t409 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X354 two_stage_opamp_dummy_magic_29_0.Vb3.t7 two_stage_opamp_dummy_magic_29_0.Vb2.t17 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.t10 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.t9 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X355 VOUT+.t2 two_stage_opamp_dummy_magic_29_0.Y.t41 VDDA.t54 VDDA.t53 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X356 GNDA_2.t73 GNDA_2.t85 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t2 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X357 VOUT-.t82 two_stage_opamp_dummy_magic_29_0.cap_res_X.t79 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X358 VOUT-.t83 two_stage_opamp_dummy_magic_29_0.cap_res_X.t78 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X359 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.t13 bgr_11_0.PFET_GATE_10uA.t17 VDDA.t239 VDDA.t238 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X360 GNDA_2.t219 two_stage_opamp_dummy_magic_29_0.X.t38 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.t6 VDDA.t128 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X361 GNDA_2.t179 two_stage_opamp_dummy_magic_29_0.X.t39 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.t5 VDDA.t74 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X362 VOUT+.t100 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t62 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X363 VOUT+.t101 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t61 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X364 two_stage_opamp_dummy_magic_29_0.Vb1.t8 two_stage_opamp_dummy_magic_29_0.Vb1.t7 two_stage_opamp_dummy_magic_29_0.Vb1_2.t1 GNDA_2.t106 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X365 a_6350_30238.t1 a_6470_28630.t1 GNDA_2.t16 sky130_fd_pr__res_xhigh_po_0p35 l=6
X366 two_stage_opamp_dummy_magic_29_0.VD4.t29 two_stage_opamp_dummy_magic_29_0.Vb2.t18 two_stage_opamp_dummy_magic_29_0.Y.t16 two_stage_opamp_dummy_magic_29_0.VD4.t28 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X367 VDDA.t92 two_stage_opamp_dummy_magic_29_0.X.t40 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.t8 GNDA_2.t198 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X368 bgr_11_0.1st_Vout_2.t4 a_6540_22450.t15 VDDA.t187 VDDA.t186 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X369 VDDA.t71 bgr_11_0.1st_Vout_1.t19 bgr_11_0.V_TOP.t4 VDDA.t70 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X370 VOUT+.t102 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t60 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X371 VOUT-.t84 two_stage_opamp_dummy_magic_29_0.cap_res_X.t77 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X372 VOUT-.t85 two_stage_opamp_dummy_magic_29_0.cap_res_X.t76 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X373 VOUT+.t103 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t59 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X374 VOUT-.t86 two_stage_opamp_dummy_magic_29_0.cap_res_X.t75 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X375 VOUT+.t104 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t58 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X376 VDDA.t65 bgr_11_0.V_mir1.t16 bgr_11_0.1st_Vout_1.t2 VDDA.t64 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X377 two_stage_opamp_dummy_magic_29_0.Y.t8 two_stage_opamp_dummy_magic_29_0.Vb1.t23 two_stage_opamp_dummy_magic_29_0.VD2.t10 GNDA_2.t170 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X378 VDDA.t179 two_stage_opamp_dummy_magic_29_0.Vb3.t13 two_stage_opamp_dummy_magic_29_0.VD4.t7 VDDA.t178 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X379 VDDA.t26 two_stage_opamp_dummy_magic_29_0.V_err_gate.t7 two_stage_opamp_dummy_magic_29_0.V_err_mir_p.t3 VDDA.t25 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X380 two_stage_opamp_dummy_magic_29_0.Y.t11 two_stage_opamp_dummy_magic_29_0.Vb1.t24 two_stage_opamp_dummy_magic_29_0.VD2.t9 GNDA_2.t3 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X381 VOUT-.t87 two_stage_opamp_dummy_magic_29_0.cap_res_X.t74 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X382 bgr_11_0.V_TOP.t35 VDDA.t410 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X383 VOUT-.t15 two_stage_opamp_dummy_magic_29_0.X.t41 VDDA.t199 VDDA.t198 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X384 VOUT-.t3 two_stage_opamp_dummy_magic_29_0.X.t42 VDDA.t57 VDDA.t56 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X385 VOUT+.t105 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t57 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X386 GNDA_2.t76 GNDA_2.t119 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t1 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X387 a_12070_30088.t1 a_11950_28880.t1 GNDA_2.t230 sky130_fd_pr__res_xhigh_po_0p35 l=4
X388 two_stage_opamp_dummy_magic_29_0.VD3.t15 VDDA.t327 VDDA.t329 VDDA.t328 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X389 GNDA_2.t269 VDDA.t324 VDDA.t326 VDDA.t325 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X390 GNDA_2.t218 two_stage_opamp_dummy_magic_29_0.Y.t42 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.t11 VDDA.t125 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X391 two_stage_opamp_dummy_magic_29_0.X.t18 two_stage_opamp_dummy_magic_29_0.Vb2.t19 two_stage_opamp_dummy_magic_29_0.VD3.t26 two_stage_opamp_dummy_magic_29_0.VD3.t25 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X392 VDDA.t386 bgr_11_0.V_TOP.t36 bgr_11_0.Vin+.t0 VDDA.t385 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X393 VOUT-.t88 two_stage_opamp_dummy_magic_29_0.cap_res_X.t73 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X394 GNDA_2.t118 GNDA_2.t116 two_stage_opamp_dummy_magic_29_0.Vb3.t0 GNDA_2.t117 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X395 VOUT-.t89 two_stage_opamp_dummy_magic_29_0.cap_res_X.t72 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X396 VDDA.t109 two_stage_opamp_dummy_magic_29_0.Y.t43 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.t9 GNDA_2.t208 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X397 two_stage_opamp_dummy_magic_29_0.V_source.t34 VIN+.t3 two_stage_opamp_dummy_magic_29_0.VD2.t21 GNDA_2.t229 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X398 VOUT+.t106 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t56 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X399 VOUT+.t107 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t55 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X400 VOUT+.t108 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t54 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X401 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t1 GNDA_2.t114 GNDA_2.t115 GNDA_2.t24 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X402 VOUT-.t90 two_stage_opamp_dummy_magic_29_0.cap_res_X.t71 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X403 GNDA_2.t200 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t21 two_stage_opamp_dummy_magic_29_0.V_source.t17 GNDA_2.t6 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X404 bgr_11_0.V_TOP.t5 bgr_11_0.START_UP.t6 bgr_11_0.Vin-.t7 VDDA.t152 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X405 VOUT-.t91 two_stage_opamp_dummy_magic_29_0.cap_res_X.t70 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X406 VOUT-.t92 two_stage_opamp_dummy_magic_29_0.cap_res_X.t69 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X407 a_6540_22450.t6 a_6540_22450.t5 VDDA.t38 VDDA.t37 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X408 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.t8 VDDA.t321 VDDA.t323 VDDA.t322 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X409 VOUT+.t109 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t53 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X410 bgr_11_0.1st_Vout_1.t20 bgr_11_0.cap_res1.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X411 VDDA.t320 VDDA.t318 bgr_11_0.V_TOP.t10 VDDA.t319 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X412 VOUT+.t11 VDDA.t315 VDDA.t317 VDDA.t316 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=2.4 ps=12.8 w=6 l=0.15
X413 VOUT+.t110 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t52 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X414 VOUT+.t12 two_stage_opamp_dummy_magic_29_0.Y.t44 VDDA.t371 VDDA.t370 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X415 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref.t1 bgr_11_0.V_TOP.t37 VDDA.t388 VDDA.t387 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X416 VOUT+.t111 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t51 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X417 VOUT-.t93 two_stage_opamp_dummy_magic_29_0.cap_res_X.t68 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X418 GNDA_2.t113 GNDA_2.t111 VOUT-.t5 GNDA_2.t112 sky130_fd_pr__nfet_01v8 ad=2.8 pd=14.8 as=1.4 ps=7.4 w=7 l=0.6
X419 GNDA_2.t249 two_stage_opamp_dummy_magic_29_0.X.t43 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.t4 VDDA.t185 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X420 GNDA_2.t110 GNDA_2.t108 VDDA.t403 GNDA_2.t109 sky130_fd_pr__nfet_01v8 ad=1.2 pd=6.8 as=0.6 ps=3.4 w=3 l=0.15
X421 VOUT+.t112 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t50 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X422 VOUT-.t94 two_stage_opamp_dummy_magic_29_0.cap_res_X.t67 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X423 VDDA_2.t2 VDDA_2.t0 two_stage_opamp_dummy_magic_29_0.Vb1.t2 VDDA_2.t1 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X424 VDDA.t237 bgr_11_0.PFET_GATE_10uA.t18 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t8 VDDA.t236 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X425 VOUT-.t95 two_stage_opamp_dummy_magic_29_0.cap_res_X.t66 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X426 VOUT-.t96 two_stage_opamp_dummy_magic_29_0.cap_res_X.t65 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X427 GNDA_2.t107 GNDA_2.t105 two_stage_opamp_dummy_magic_29_0.Vb1.t0 GNDA_2.t106 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X428 VDDA.t61 two_stage_opamp_dummy_magic_29_0.Vb3.t14 two_stage_opamp_dummy_magic_29_0.VD4.t2 VDDA.t60 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X429 two_stage_opamp_dummy_magic_29_0.V_source.t26 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t22 GNDA_2.t243 GNDA_2.t6 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X430 bgr_11_0.PFET_GATE_10uA.t7 bgr_11_0.1st_Vout_2.t21 VDDA.t209 VDDA.t208 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X431 VDDA.t364 two_stage_opamp_dummy_magic_29_0.X.t44 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.t7 GNDA_2.t271 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X432 VOUT+.t113 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t49 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X433 two_stage_opamp_dummy_magic_29_0.V_source.t2 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t23 GNDA_2.t13 GNDA_2.t6 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X434 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t7 bgr_11_0.PFET_GATE_10uA.t19 VDDA.t235 VDDA.t234 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X435 bgr_11_0.1st_Vout_1.t21 bgr_11_0.cap_res1.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X436 VOUT-.t97 two_stage_opamp_dummy_magic_29_0.cap_res_X.t64 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X437 VOUT+.t114 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t48 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X438 VOUT+.t3 a_3830_76.t1 GNDA_2.t171 sky130_fd_pr__res_xhigh_po_0p35 l=2.63
X439 VOUT-.t98 two_stage_opamp_dummy_magic_29_0.cap_res_X.t63 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X440 two_stage_opamp_dummy_magic_29_0.Y.t12 two_stage_opamp_dummy_magic_29_0.Vb1.t25 two_stage_opamp_dummy_magic_29_0.VD2.t8 GNDA_2.t25 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X441 GNDA_2.t28 bgr_11_0.NFET_GATE_10uA.t13 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.t3 GNDA_2.t27 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X442 VDDA.t146 bgr_11_0.V_TOP.t38 bgr_11_0.START_UP.t1 VDDA.t145 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X443 bgr_11_0.Vin-.t2 bgr_11_0.V_TOP.t39 VDDA.t148 VDDA.t147 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X444 VOUT-.t99 two_stage_opamp_dummy_magic_29_0.cap_res_X.t62 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X445 bgr_11_0.1st_Vout_1.t22 bgr_11_0.cap_res1.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X446 VOUT-.t13 two_stage_opamp_dummy_magic_29_0.X.t45 VDDA.t168 VDDA.t167 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X447 VOUT-.t100 two_stage_opamp_dummy_magic_29_0.cap_res_X.t61 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X448 VOUT+.t115 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t47 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X449 VOUT-.t101 two_stage_opamp_dummy_magic_29_0.cap_res_X.t60 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X450 GNDA_2.t285 two_stage_opamp_dummy_magic_29_0.Y.t45 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.t10 VDDA.t398 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X451 VOUT-.t102 two_stage_opamp_dummy_magic_29_0.cap_res_X.t59 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X452 two_stage_opamp_dummy_magic_29_0.Y.t0 two_stage_opamp_dummy_magic_29_0.VD4.t32 two_stage_opamp_dummy_magic_29_0.VD4.t34 two_stage_opamp_dummy_magic_29_0.VD4.t33 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X453 VOUT-.t6 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.t7 GNDA_2.t19 GNDA_2.t18 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X454 GNDA_2.t268 VDDA.t412 bgr_11_0.V_TOP.t8 GNDA_2.t267 sky130_fd_pr__nfet_01v8 ad=1.01 pd=6.15 as=1 ps=5.8 w=2.5 l=5
X455 two_stage_opamp_dummy_magic_29_0.V_source.t33 VIN+.t4 two_stage_opamp_dummy_magic_29_0.VD2.t20 GNDA_2.t43 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X456 bgr_11_0.1st_Vout_1.t23 bgr_11_0.cap_res1.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X457 a_14420_3878.t0 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.t14 GNDA_2.t279 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X458 GNDA_2.t251 bgr_11_0.NFET_GATE_10uA.t14 two_stage_opamp_dummy_magic_29_0.V_err_gate.t1 GNDA_2.t250 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X459 GNDA_2.t197 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t24 two_stage_opamp_dummy_magic_29_0.V_source.t16 GNDA_2.t6 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X460 VOUT+.t116 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t46 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X461 bgr_11_0.V_TOP.t40 VDDA.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X462 VOUT+.t117 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t45 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X463 bgr_11_0.1st_Vout_2.t0 a_6540_22450.t16 VDDA.t14 VDDA.t13 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X464 two_stage_opamp_dummy_magic_29_0.VD4.t10 VDDA.t312 VDDA.t314 VDDA.t313 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X465 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.t3 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.t1 two_stage_opamp_dummy_magic_29_0.Vb3.t6 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.t2 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X466 VOUT+.t118 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t44 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X467 two_stage_opamp_dummy_magic_29_0.VD3.t11 two_stage_opamp_dummy_magic_29_0.Vb3.t15 VDDA.t96 VDDA.t95 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X468 VOUT-.t103 two_stage_opamp_dummy_magic_29_0.cap_res_X.t58 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X469 VOUT+.t119 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t43 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X470 bgr_11_0.V_p_1.t1 VDDA.t413 GNDA_2.t264 GNDA_2.t263 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=1.01 ps=6.15 w=2.5 l=5
X471 VOUT-.t104 two_stage_opamp_dummy_magic_29_0.cap_res_X.t57 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X472 VOUT-.t105 two_stage_opamp_dummy_magic_29_0.cap_res_X.t56 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X473 VOUT-.t106 two_stage_opamp_dummy_magic_29_0.cap_res_X.t55 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X474 VOUT+.t17 two_stage_opamp_dummy_magic_29_0.Y.t46 VDDA.t400 VDDA.t399 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X475 bgr_11_0.NFET_GATE_10uA.t3 bgr_11_0.PFET_GATE_10uA.t20 VDDA.t233 VDDA.t232 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X476 GNDA_2.t104 GNDA_2.t103 two_stage_opamp_dummy_magic_29_0.err_amp_out.t1 GNDA_2.t52 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=0.5 ps=2.9 w=2.5 l=0.15
X477 VOUT+.t120 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t42 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X478 VOUT-.t107 two_stage_opamp_dummy_magic_29_0.cap_res_X.t54 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X479 two_stage_opamp_dummy_magic_29_0.Vb3.t4 bgr_11_0.NFET_GATE_10uA.t15 GNDA_2.t45 GNDA_2.t44 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X480 VDDA.t311 VDDA.t309 GNDA_2.t266 VDDA.t310 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X481 bgr_11_0.1st_Vout_2.t22 bgr_11_0.cap_res2.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X482 bgr_11_0.V_mir1.t6 bgr_11_0.V_mir1.t5 VDDA.t2 VDDA.t1 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X483 two_stage_opamp_dummy_magic_29_0.Y.t18 two_stage_opamp_dummy_magic_29_0.Vb2.t20 two_stage_opamp_dummy_magic_29_0.VD4.t27 two_stage_opamp_dummy_magic_29_0.VD4.t26 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X484 bgr_11_0.1st_Vout_2.t6 bgr_11_0.V_CUR_REF_REG.t3 bgr_11_0.V_p_2.t1 GNDA_2.t270 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=0.5 ps=2.9 w=2.5 l=0.2
X485 GNDA_2.t42 two_stage_opamp_dummy_magic_29_0.X.t46 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.t3 VDDA.t43 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X486 VOUT+.t121 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t41 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X487 VOUT-.t108 two_stage_opamp_dummy_magic_29_0.cap_res_X.t53 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X488 VOUT+.t122 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t40 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X489 bgr_11_0.1st_Vout_1.t24 bgr_11_0.cap_res1.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X490 two_stage_opamp_dummy_magic_29_0.V_source.t20 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t25 GNDA_2.t207 GNDA_2.t6 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X491 VDDA.t402 GNDA_2.t100 GNDA_2.t102 GNDA_2.t101 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=1.2 ps=6.8 w=3 l=0.15
X492 VOUT+.t123 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t39 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X493 VOUT-.t109 two_stage_opamp_dummy_magic_29_0.cap_res_X.t52 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X494 two_stage_opamp_dummy_magic_29_0.VD4.t0 two_stage_opamp_dummy_magic_29_0.Vb3.t16 VDDA.t4 VDDA.t3 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X495 bgr_11_0.1st_Vout_2.t23 bgr_11_0.cap_res2.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X496 VOUT+.t124 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t38 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X497 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.t2 bgr_11_0.NFET_GATE_10uA.t16 GNDA_2.t12 GNDA_2.t11 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X498 VOUT-.t110 two_stage_opamp_dummy_magic_29_0.cap_res_X.t51 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X499 VOUT-.t111 two_stage_opamp_dummy_magic_29_0.cap_res_X.t50 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X500 two_stage_opamp_dummy_magic_29_0.Y.t6 two_stage_opamp_dummy_magic_29_0.Vb1.t26 two_stage_opamp_dummy_magic_29_0.VD2.t7 GNDA_2.t183 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X501 VOUT-.t112 two_stage_opamp_dummy_magic_29_0.cap_res_X.t49 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X502 GNDA_2.t73 GNDA_2.t98 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t0 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X503 GNDA_2.t255 bgr_11_0.NFET_GATE_10uA.t17 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.t1 GNDA_2.t254 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X504 VDDA.t308 VDDA.t306 two_stage_opamp_dummy_magic_29_0.err_amp_out.t2 VDDA.t307 sky130_fd_pr__pfet_01v8 ad=1 pd=5.8 as=0.5 ps=2.9 w=2.5 l=0.15
X505 VDDA.t305 VDDA.t303 VOUT+.t10 VDDA.t304 sky130_fd_pr__pfet_01v8 ad=2.4 pd=12.8 as=1.2 ps=6.4 w=6 l=0.15
X506 VOUT-.t16 two_stage_opamp_dummy_magic_29_0.X.t47 VDDA.t203 VDDA.t202 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X507 VOUT-.t113 two_stage_opamp_dummy_magic_29_0.cap_res_X.t48 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X508 two_stage_opamp_dummy_magic_29_0.Vb1_2.t0 two_stage_opamp_dummy_magic_29_0.Vb1.t5 two_stage_opamp_dummy_magic_29_0.Vb1.t6 GNDA_2.t106 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X509 VDDA.t157 two_stage_opamp_dummy_magic_29_0.Vb3.t17 two_stage_opamp_dummy_magic_29_0.VD3.t12 VDDA.t156 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X510 VOUT-.t114 two_stage_opamp_dummy_magic_29_0.cap_res_X.t47 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X511 bgr_11_0.1st_Vout_2.t24 bgr_11_0.cap_res2.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X512 two_stage_opamp_dummy_magic_29_0.V_source.t24 VIN-.t4 two_stage_opamp_dummy_magic_29_0.VD1.t20 GNDA_2.t235 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X513 two_stage_opamp_dummy_magic_29_0.VD4.t3 two_stage_opamp_dummy_magic_29_0.Vb3.t18 VDDA.t80 VDDA.t79 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X514 VOUT+.t125 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t37 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X515 VOUT-.t115 two_stage_opamp_dummy_magic_29_0.cap_res_X.t46 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X516 bgr_11_0.1st_Vout_1.t25 bgr_11_0.cap_res1.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X517 GNDA_2.t10 bgr_11_0.NFET_GATE_10uA.t18 two_stage_opamp_dummy_magic_29_0.Vb2.t0 GNDA_2.t9 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X518 VOUT+.t126 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t36 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X519 bgr_11_0.1st_Vout_2.t25 bgr_11_0.cap_res2.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X520 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.t2 bgr_11_0.NFET_GATE_10uA.t19 GNDA_2.t31 GNDA_2.t30 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X521 bgr_11_0.PFET_GATE_10uA.t6 bgr_11_0.1st_Vout_2.t26 VDDA.t207 VDDA.t206 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X522 VOUT+.t127 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t35 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X523 VDDA.t86 two_stage_opamp_dummy_magic_29_0.Vb3.t19 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.t0 VDDA.t85 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X524 two_stage_opamp_dummy_magic_29_0.V_source.t32 VIN+.t5 two_stage_opamp_dummy_magic_29_0.VD2.t1 GNDA_2.t50 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X525 VOUT-.t116 two_stage_opamp_dummy_magic_29_0.cap_res_X.t45 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X526 VOUT-.t117 two_stage_opamp_dummy_magic_29_0.cap_res_X.t44 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X527 two_stage_opamp_dummy_magic_29_0.V_source.t19 VIN-.t5 two_stage_opamp_dummy_magic_29_0.VD1.t9 GNDA_2.t61 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X528 VOUT-.t118 two_stage_opamp_dummy_magic_29_0.cap_res_X.t43 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X529 bgr_11_0.1st_Vout_1.t26 bgr_11_0.cap_res1.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X530 VOUT-.t119 two_stage_opamp_dummy_magic_29_0.cap_res_X.t42 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X531 two_stage_opamp_dummy_magic_29_0.Y.t15 two_stage_opamp_dummy_magic_29_0.Vb2.t21 two_stage_opamp_dummy_magic_29_0.VD4.t25 two_stage_opamp_dummy_magic_29_0.VD4.t24 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X532 VOUT+.t128 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t34 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X533 VOUT+.t129 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t33 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X534 bgr_11_0.1st_Vout_2.t27 bgr_11_0.cap_res2.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X535 GNDA_2.t73 GNDA_2.t99 bgr_11_0.Vin-.t4 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X536 VOUT+.t130 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t32 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X537 VOUT-.t120 two_stage_opamp_dummy_magic_29_0.cap_res_X.t41 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X538 bgr_11_0.1st_Vout_2.t5 a_6540_22450.t17 VDDA.t195 VDDA.t194 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X539 bgr_11_0.1st_Vout_1.t27 bgr_11_0.cap_res1.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X540 bgr_11_0.V_TOP.t0 bgr_11_0.1st_Vout_1.t28 VDDA.t6 VDDA.t5 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X541 two_stage_opamp_dummy_magic_29_0.VD4.t9 two_stage_opamp_dummy_magic_29_0.Vb3.t20 VDDA.t201 VDDA.t200 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X542 VOUT+.t131 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t31 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X543 VOUT+.t132 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t30 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X544 GNDA_2.t265 VDDA.t300 VDDA.t302 VDDA.t301 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X545 VOUT-.t121 two_stage_opamp_dummy_magic_29_0.cap_res_X.t40 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X546 bgr_11_0.1st_Vout_1.t4 bgr_11_0.V_mir1.t17 VDDA.t159 VDDA.t158 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X547 two_stage_opamp_dummy_magic_29_0.X.t9 two_stage_opamp_dummy_magic_29_0.Vb1.t27 two_stage_opamp_dummy_magic_29_0.VD1.t13 GNDA_2.t15 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X548 VOUT-.t122 two_stage_opamp_dummy_magic_29_0.cap_res_X.t39 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X549 VOUT-.t123 two_stage_opamp_dummy_magic_29_0.cap_res_X.t38 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X550 VOUT-.t124 two_stage_opamp_dummy_magic_29_0.cap_res_X.t37 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X551 VDDA.t299 VDDA.t297 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.t5 VDDA.t298 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X552 VOUT-.t125 two_stage_opamp_dummy_magic_29_0.cap_res_X.t36 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X553 two_stage_opamp_dummy_magic_29_0.V_source.t27 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t26 GNDA_2.t247 GNDA_2.t6 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X554 bgr_11_0.PFET_GATE_10uA.t1 VDDA.t414 GNDA_2.t262 GNDA_2.t261 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=1 ps=5.8 w=2.5 l=5
X555 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.t1 bgr_11_0.PFET_GATE_10uA.t21 VDDA.t231 VDDA.t230 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X556 VDDA.t205 two_stage_opamp_dummy_magic_29_0.Vb3.t21 two_stage_opamp_dummy_magic_29_0.VD3.t14 VDDA.t204 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X557 VOUT+.t1 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.t8 GNDA_2.t60 GNDA_2.t59 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X558 VOUT+.t133 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t29 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X559 VOUT+.t134 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t28 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X560 VOUT+.t135 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t27 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X561 two_stage_opamp_dummy_magic_29_0.Y.t4 GNDA_2.t95 GNDA_2.t97 GNDA_2.t96 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X562 VOUT+.t136 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t26 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X563 bgr_11_0.V_TOP.t41 VDDA.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X564 two_stage_opamp_dummy_magic_29_0.V_err_p.t2 two_stage_opamp_dummy_magic_29_0.V_err_gate.t8 VDDA.t28 VDDA.t27 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X565 VDDA.t296 VDDA.t294 bgr_11_0.PFET_GATE_10uA.t9 VDDA.t295 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.2
X566 VDDA.t150 bgr_11_0.V_TOP.t42 bgr_11_0.START_UP.t0 VDDA.t149 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X567 two_stage_opamp_dummy_magic_29_0.X.t5 two_stage_opamp_dummy_magic_29_0.Vb1.t28 two_stage_opamp_dummy_magic_29_0.VD1.t12 GNDA_2.t3 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X568 VOUT+.t137 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t25 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X569 VOUT-.t18 VDDA.t291 VDDA.t293 VDDA.t292 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=2.4 ps=12.8 w=6 l=0.15
X570 two_stage_opamp_dummy_magic_29_0.VD4.t23 two_stage_opamp_dummy_magic_29_0.Vb2.t22 two_stage_opamp_dummy_magic_29_0.Y.t13 two_stage_opamp_dummy_magic_29_0.VD4.t22 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X571 VOUT-.t126 two_stage_opamp_dummy_magic_29_0.cap_res_X.t35 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X572 two_stage_opamp_dummy_magic_29_0.VD3.t24 two_stage_opamp_dummy_magic_29_0.Vb2.t23 two_stage_opamp_dummy_magic_29_0.X.t19 two_stage_opamp_dummy_magic_29_0.VD3.t23 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X573 VOUT+.t138 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t24 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X574 VOUT+.t139 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t23 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X575 two_stage_opamp_dummy_magic_29_0.V_source.t14 VIN-.t6 two_stage_opamp_dummy_magic_29_0.VD1.t7 GNDA_2.t164 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X576 a_14540_3878.t0 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.t0 GNDA_2.t167 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X577 a_6540_22450.t4 a_6540_22450.t3 VDDA.t189 VDDA.t188 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X578 VOUT-.t127 two_stage_opamp_dummy_magic_29_0.cap_res_X.t34 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X579 bgr_11_0.V_TOP.t43 VDDA.t151 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X580 VOUT+.t140 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t22 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X581 GNDA_2.t206 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t27 two_stage_opamp_dummy_magic_29_0.V_source.t18 GNDA_2.t205 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X582 VDDA.t100 two_stage_opamp_dummy_magic_29_0.Vb3.t22 two_stage_opamp_dummy_magic_29_0.VD4.t4 VDDA.t99 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X583 GNDA_2.t94 GNDA_2.t92 VDDA.t401 GNDA_2.t93 sky130_fd_pr__nfet_01v8 ad=1.2 pd=6.8 as=0.6 ps=3.4 w=3 l=0.15
X584 a_11420_30238.t0 a_11300_28630.t0 GNDA_2.t34 sky130_fd_pr__res_xhigh_po_0p35 l=6
X585 VDDA.t394 two_stage_opamp_dummy_magic_29_0.Vb3.t23 two_stage_opamp_dummy_magic_29_0.VD3.t37 VDDA.t393 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X586 two_stage_opamp_dummy_magic_29_0.V_source.t31 VIN+.t6 two_stage_opamp_dummy_magic_29_0.VD2.t19 GNDA_2.t24 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X587 VOUT+.t141 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t21 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X588 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t0 VIN-.t7 two_stage_opamp_dummy_magic_29_0.V_p_mir.t2 GNDA_2.t24 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X589 two_stage_opamp_dummy_magic_29_0.V_source.t6 VIN-.t8 two_stage_opamp_dummy_magic_29_0.VD1.t2 GNDA_2.t24 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X590 VOUT-.t128 two_stage_opamp_dummy_magic_29_0.cap_res_X.t33 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X591 VDDA.t229 bgr_11_0.PFET_GATE_10uA.t22 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t6 VDDA.t228 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X592 GNDA_2.t217 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.t9 VOUT+.t7 GNDA_2.t216 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X593 VOUT-.t129 two_stage_opamp_dummy_magic_29_0.cap_res_X.t32 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X594 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t5 bgr_11_0.PFET_GATE_10uA.t23 VDDA.t227 VDDA.t226 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X595 VOUT+.t142 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t20 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X596 bgr_11_0.V_TOP.t44 VDDA.t171 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X597 VOUT-.t130 two_stage_opamp_dummy_magic_29_0.cap_res_X.t31 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X598 VOUT-.t131 two_stage_opamp_dummy_magic_29_0.cap_res_X.t30 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X599 bgr_11_0.1st_Vout_1.t5 bgr_11_0.V_mir1.t18 VDDA.t161 VDDA.t160 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X600 VOUT+.t143 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X601 VOUT+.t144 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X602 two_stage_opamp_dummy_magic_29_0.VD4.t21 two_stage_opamp_dummy_magic_29_0.Vb2.t24 two_stage_opamp_dummy_magic_29_0.Y.t20 two_stage_opamp_dummy_magic_29_0.VD4.t20 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X603 VOUT-.t4 GNDA_2.t89 GNDA_2.t91 GNDA_2.t90 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=2.8 ps=14.8 w=7 l=0.6
X604 bgr_11_0.V_mir1.t0 bgr_11_0.Vin-.t8 bgr_11_0.V_p_1.t0 GNDA_2.t201 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=0.5 ps=2.9 w=2.5 l=0.2
X605 VOUT-.t132 two_stage_opamp_dummy_magic_29_0.cap_res_X.t29 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X606 VDDA.t290 VDDA.t287 VDDA.t289 VDDA.t288 sky130_fd_pr__pfet_01v8 ad=0.72 pd=4.4 as=0 ps=0 w=1.8 l=0.2
X607 VOUT-.t133 two_stage_opamp_dummy_magic_29_0.cap_res_X.t28 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X608 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.t12 bgr_11_0.PFET_GATE_10uA.t24 VDDA.t225 VDDA.t224 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X609 VOUT+.t145 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X610 VDDA.t223 bgr_11_0.PFET_GATE_10uA.t25 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.t11 VDDA.t222 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X611 VOUT-.t134 two_stage_opamp_dummy_magic_29_0.cap_res_X.t27 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X612 VOUT-.t135 two_stage_opamp_dummy_magic_29_0.cap_res_X.t26 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X613 VDDA.t286 VDDA.t284 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.t15 VDDA.t285 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X614 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.t8 two_stage_opamp_dummy_magic_29_0.Y.t47 VDDA.t166 GNDA_2.t237 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X615 two_stage_opamp_dummy_magic_29_0.X.t23 two_stage_opamp_dummy_magic_29_0.VD3.t3 two_stage_opamp_dummy_magic_29_0.VD3.t5 two_stage_opamp_dummy_magic_29_0.VD3.t4 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X616 VOUT+.t146 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X617 VOUT+.t147 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X618 two_stage_opamp_dummy_magic_29_0.X.t3 two_stage_opamp_dummy_magic_29_0.Vb1.t29 two_stage_opamp_dummy_magic_29_0.VD1.t11 GNDA_2.t41 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X619 VOUT+.t148 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X620 VOUT-.t136 two_stage_opamp_dummy_magic_29_0.cap_res_X.t25 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X621 two_stage_opamp_dummy_magic_29_0.V_source.t0 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t28 GNDA_2.t7 GNDA_2.t6 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X622 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref.t0 bgr_11_0.V_TOP.t45 VDDA.t173 VDDA.t172 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X623 bgr_11_0.V_TOP.t46 VDDA.t107 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X624 GNDA_2.t175 a_5820_28824.t0 GNDA_2.t174 sky130_fd_pr__res_xhigh_po_0p35 l=4.28
X625 bgr_11_0.V_TOP.t1 bgr_11_0.1st_Vout_1.t29 VDDA.t34 VDDA.t33 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X626 two_stage_opamp_dummy_magic_29_0.VD4.t19 two_stage_opamp_dummy_magic_29_0.Vb2.t25 two_stage_opamp_dummy_magic_29_0.Y.t19 two_stage_opamp_dummy_magic_29_0.VD4.t18 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X627 a_3110_3878.t1 two_stage_opamp_dummy_magic_29_0.V_tot.t0 GNDA_2.t182 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X628 VOUT-.t137 two_stage_opamp_dummy_magic_29_0.cap_res_X.t24 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X629 two_stage_opamp_dummy_magic_29_0.VD3.t2 two_stage_opamp_dummy_magic_29_0.Vb3.t24 VDDA.t51 VDDA.t50 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X630 two_stage_opamp_dummy_magic_29_0.V_err_gate.t4 VDDA.t281 VDDA.t283 VDDA.t282 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=1 ps=5.8 w=2.5 l=0.15
X631 two_stage_opamp_dummy_magic_29_0.V_err_p.t1 two_stage_opamp_dummy_magic_29_0.V_tot.t5 two_stage_opamp_dummy_magic_29_0.err_amp_mir.t4 VDDA.t375 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X632 two_stage_opamp_dummy_magic_29_0.X.t22 two_stage_opamp_dummy_magic_29_0.Vb1.t30 two_stage_opamp_dummy_magic_29_0.VD1.t10 GNDA_2.t3 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X633 GNDA_2.t287 two_stage_opamp_dummy_magic_29_0.err_amp_out.t5 two_stage_opamp_dummy_magic_29_0.V_source.t40 GNDA_2.t286 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X634 VDDA.t183 two_stage_opamp_dummy_magic_29_0.Vb3.t25 two_stage_opamp_dummy_magic_29_0.VD4.t8 VDDA.t182 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X635 bgr_11_0.V_TOP.t2 bgr_11_0.1st_Vout_1.t30 VDDA.t67 VDDA.t66 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X636 bgr_11_0.1st_Vout_2.t28 bgr_11_0.cap_res2.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X637 two_stage_opamp_dummy_magic_29_0.Vb2.t10 two_stage_opamp_dummy_magic_29_0.Vb2_2.t0 two_stage_opamp_dummy_magic_29_0.Vb2_2.t2 two_stage_opamp_dummy_magic_29_0.Vb2_2.t1 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X638 VOUT-.t138 two_stage_opamp_dummy_magic_29_0.cap_res_X.t23 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X639 VDDA.t280 VDDA.t278 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref.t5 VDDA.t279 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.8 as=0.6 ps=3.4 w=3 l=0.5
X640 VDDA.t274 VDDA.t272 VDDA.t274 VDDA.t273 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0 ps=0 w=3.5 l=0.2
X641 VDDA.t277 VDDA.t275 GNDA_2.t260 VDDA.t276 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X642 two_stage_opamp_dummy_magic_29_0.Vb3.t3 bgr_11_0.NFET_GATE_10uA.t20 GNDA_2.t5 GNDA_2.t4 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X643 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.t6 two_stage_opamp_dummy_magic_29_0.X.t48 VDDA.t184 GNDA_2.t248 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X644 GNDA_2.t88 GNDA_2.t86 two_stage_opamp_dummy_magic_29_0.X.t7 GNDA_2.t87 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X645 VOUT-.t139 two_stage_opamp_dummy_magic_29_0.cap_res_X.t22 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X646 bgr_11_0.1st_Vout_1.t31 bgr_11_0.cap_res1.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X647 two_stage_opamp_dummy_magic_29_0.V_source.t23 two_stage_opamp_dummy_magic_29_0.Vb1.t31 two_stage_opamp_dummy_magic_29_0.Vb1_2.t4 GNDA_2.t256 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.6 ps=3.8 w=1.5 l=3
X648 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.t5 two_stage_opamp_dummy_magic_29_0.X.t49 VDDA.t177 GNDA_2.t244 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X649 VOUT+.t149 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X650 VOUT+.t150 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X651 two_stage_opamp_dummy_magic_29_0.VD4.t17 two_stage_opamp_dummy_magic_29_0.Vb2.t26 two_stage_opamp_dummy_magic_29_0.Y.t22 two_stage_opamp_dummy_magic_29_0.VD4.t16 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X652 two_stage_opamp_dummy_magic_29_0.V_source.t9 VIN-.t9 two_stage_opamp_dummy_magic_29_0.VD1.t3 GNDA_2.t24 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X653 VOUT+.t151 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X654 bgr_11_0.Vin-.t6 bgr_11_0.START_UP.t7 bgr_11_0.V_TOP.t7 VDDA.t164 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X655 VDDA.t271 VDDA.t269 two_stage_opamp_dummy_magic_29_0.Vb2_2.t6 VDDA.t270 sky130_fd_pr__pfet_01v8 ad=0.72 pd=4.4 as=0.36 ps=2.2 w=1.8 l=0.2
X656 VDDA.t268 VDDA.t266 two_stage_opamp_dummy_magic_29_0.V_err_gate.t3 VDDA.t267 sky130_fd_pr__pfet_01v8 ad=1 pd=5.8 as=0.5 ps=2.9 w=2.5 l=0.15
X657 VOUT+.t152 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X658 GNDA_2.t84 GNDA_2.t83 two_stage_opamp_dummy_magic_29_0.Y.t3 GNDA_2.t3 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X659 bgr_11_0.V_mir1.t4 bgr_11_0.V_mir1.t3 VDDA.t47 VDDA.t46 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X660 VOUT-.t140 two_stage_opamp_dummy_magic_29_0.cap_res_X.t21 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X661 bgr_11_0.V_p_2.t0 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref.t9 a_6540_22450.t0 GNDA_2.t165 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=1 ps=5.8 w=2.5 l=0.2
X662 two_stage_opamp_dummy_magic_29_0.X.t14 two_stage_opamp_dummy_magic_29_0.Vb2.t27 two_stage_opamp_dummy_magic_29_0.VD3.t22 two_stage_opamp_dummy_magic_29_0.VD3.t21 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X663 VDDA.t265 VDDA.t263 VOUT-.t17 VDDA.t264 sky130_fd_pr__pfet_01v8 ad=2.4 pd=12.8 as=1.2 ps=6.4 w=6 l=0.15
X664 VOUT+.t153 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X665 VDDA.t170 two_stage_opamp_dummy_magic_29_0.Vb3.t26 two_stage_opamp_dummy_magic_29_0.VD4.t6 VDDA.t169 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X666 bgr_11_0.V_TOP.t9 VDDA.t260 VDDA.t262 VDDA.t261 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.2
X667 two_stage_opamp_dummy_magic_29_0.VD1.t8 VIN-.t10 two_stage_opamp_dummy_magic_29_0.V_source.t15 GNDA_2.t177 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X668 VOUT-.t141 two_stage_opamp_dummy_magic_29_0.cap_res_X.t20 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X669 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.t9 two_stage_opamp_dummy_magic_29_0.Y.t48 GNDA_2.t20 VDDA.t21 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X670 bgr_11_0.V_TOP.t47 VDDA.t108 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X671 two_stage_opamp_dummy_magic_29_0.cap_res_X.t143 two_stage_opamp_dummy_magic_29_0.X.t8 GNDA_2.t184 sky130_fd_pr__res_high_po_1p41 l=1.41
X672 VDDA.t120 bgr_11_0.V_TOP.t48 bgr_11_0.Vin-.t1 VDDA.t119 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X673 VOUT+.t154 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X674 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.t7 two_stage_opamp_dummy_magic_29_0.Y.t49 VDDA.t22 GNDA_2.t21 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X675 two_stage_opamp_dummy_magic_29_0.Vb1.t11 bgr_11_0.PFET_GATE_10uA.t26 VDDA_2.t8 VDDA_2.t7 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X676 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t4 bgr_11_0.PFET_GATE_10uA.t27 VDDA.t221 VDDA.t220 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X677 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.t6 two_stage_opamp_dummy_magic_29_0.Y.t50 VDDA.t139 GNDA_2.t226 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X678 two_stage_opamp_dummy_magic_29_0.VD3.t10 two_stage_opamp_dummy_magic_29_0.Vb3.t27 VDDA.t90 VDDA.t89 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X679 two_stage_opamp_dummy_magic_29_0.V_p_mir.t0 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t29 GNDA_2.t234 GNDA_2.t233 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X680 two_stage_opamp_dummy_magic_29_0.VD2.t17 VIN+.t7 two_stage_opamp_dummy_magic_29_0.V_source.t30 GNDA_2.t24 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X681 two_stage_opamp_dummy_magic_29_0.V_source.t1 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t30 GNDA_2.t8 GNDA_2.t6 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X682 GNDA_2.t17 a_6470_28630.t0 GNDA_2.t16 sky130_fd_pr__res_xhigh_po_0p35 l=6
X683 VOUT-.t142 two_stage_opamp_dummy_magic_29_0.cap_res_X.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X684 GNDA_2.t82 GNDA_2.t80 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.t0 GNDA_2.t81 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X685 VDDA.t30 a_6540_22450.t18 bgr_11_0.1st_Vout_2.t1 VDDA.t29 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X686 bgr_11_0.1st_Vout_2.t29 bgr_11_0.cap_res2.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X687 VOUT-.t143 two_stage_opamp_dummy_magic_29_0.cap_res_X.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X688 VOUT+.t155 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X689 VOUT-.t144 two_stage_opamp_dummy_magic_29_0.cap_res_X.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X690 GNDA_2.t173 bgr_11_0.NFET_GATE_10uA.t21 two_stage_opamp_dummy_magic_29_0.Vb2.t4 GNDA_2.t172 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X691 VOUT-.t145 two_stage_opamp_dummy_magic_29_0.cap_res_X.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X692 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.t0 GNDA_2.t77 GNDA_2.t79 GNDA_2.t78 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X693 GNDA_2.t259 VDDA.t415 bgr_11_0.V_p_2.t2 GNDA_2.t258 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=1 ps=5.8 w=2.5 l=5
X694 bgr_11_0.V_mir1.t2 bgr_11_0.V_mir1.t1 VDDA.t193 VDDA.t192 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X695 VDDA.t141 two_stage_opamp_dummy_magic_29_0.Y.t51 VOUT+.t9 VDDA.t140 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X696 VOUT-.t146 two_stage_opamp_dummy_magic_29_0.cap_res_X.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X697 two_stage_opamp_dummy_magic_29_0.Y.t21 two_stage_opamp_dummy_magic_29_0.Vb2.t28 two_stage_opamp_dummy_magic_29_0.VD4.t15 two_stage_opamp_dummy_magic_29_0.VD4.t14 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X698 VOUT+.t156 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X699 two_stage_opamp_dummy_magic_29_0.X.t21 two_stage_opamp_dummy_magic_29_0.Vb2.t29 two_stage_opamp_dummy_magic_29_0.VD3.t20 two_stage_opamp_dummy_magic_29_0.VD3.t19 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X700 VOUT-.t147 two_stage_opamp_dummy_magic_29_0.cap_res_X.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X701 VOUT+.t157 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X702 VOUT-.t148 two_stage_opamp_dummy_magic_29_0.cap_res_X.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X703 two_stage_opamp_dummy_magic_29_0.err_amp_mir.t0 GNDA_2.t70 GNDA_2.t71 GNDA_2.t52 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=1 ps=5.8 w=2.5 l=0.15
X704 two_stage_opamp_dummy_magic_29_0.X.t6 GNDA_2.t68 GNDA_2.t69 GNDA_2.t3 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X705 bgr_11_0.PFET_GATE_10uA.t8 VDDA.t257 VDDA.t259 VDDA.t258 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.2
X706 a_14540_3878.t1 two_stage_opamp_dummy_magic_29_0.V_tot.t1 GNDA_2.t193 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X707 VOUT-.t149 two_stage_opamp_dummy_magic_29_0.cap_res_X.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X708 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.t2 two_stage_opamp_dummy_magic_29_0.X.t50 GNDA_2.t203 VDDA.t97 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X709 VOUT-.t150 two_stage_opamp_dummy_magic_29_0.cap_res_X.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X710 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.t1 two_stage_opamp_dummy_magic_29_0.X.t51 GNDA_2.t213 VDDA.t118 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X711 a_12070_30088.t0 bgr_11_0.V_CUR_REF_REG.t0 GNDA_2.t14 sky130_fd_pr__res_xhigh_po_0p35 l=4
X712 two_stage_opamp_dummy_magic_29_0.VD3.t0 two_stage_opamp_dummy_magic_29_0.Vb3.t28 VDDA.t12 VDDA.t11 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X713 VOUT+.t158 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X714 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.t4 two_stage_opamp_dummy_magic_29_0.X.t52 VDDA.t91 GNDA_2.t192 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X715 VOUT-.t151 two_stage_opamp_dummy_magic_29_0.cap_res_X.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X716 bgr_11_0.1st_Vout_2.t30 bgr_11_0.cap_res2.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X717 GNDA_2.t67 GNDA_2.t65 bgr_11_0.NFET_GATE_10uA.t0 GNDA_2.t66 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X718 bgr_11_0.Vin-.t0 bgr_11_0.V_TOP.t49 VDDA.t122 VDDA.t121 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X719 VOUT+.t159 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X720 VOUT-.t152 two_stage_opamp_dummy_magic_29_0.cap_res_X.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X721 two_stage_opamp_dummy_magic_29_0.V_err_mir_p.t2 two_stage_opamp_dummy_magic_29_0.V_err_gate.t9 VDDA.t374 VDDA.t373 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X722 VDDA.t115 a_6540_22450.t1 a_6540_22450.t2 VDDA.t114 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X723 two_stage_opamp_dummy_magic_29_0.VD2.t6 two_stage_opamp_dummy_magic_29_0.Vb1.t32 two_stage_opamp_dummy_magic_29_0.Y.t23 GNDA_2.t3 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X724 VOUT-.t153 two_stage_opamp_dummy_magic_29_0.cap_res_X.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X725 VOUT-.t154 two_stage_opamp_dummy_magic_29_0.cap_res_X.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X726 VOUT-.t155 two_stage_opamp_dummy_magic_29_0.cap_res_X.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X727 bgr_11_0.1st_Vout_2.t31 bgr_11_0.cap_res2.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X728 two_stage_opamp_dummy_magic_29_0.Vb2_2.t7 two_stage_opamp_dummy_magic_29_0.Vb2.t30 VDDA.t135 VDDA.t134 sky130_fd_pr__pfet_01v8 ad=0.36 pd=2.2 as=0.36 ps=2.2 w=1.8 l=0.2
X729 VDDA.t133 two_stage_opamp_dummy_magic_29_0.X.t53 VOUT-.t12 VDDA.t132 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X730 bgr_11_0.V_CUR_REF_REG.t2 VDDA.t254 VDDA.t256 VDDA.t255 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X731 VDDA.t42 two_stage_opamp_dummy_magic_29_0.X.t54 VOUT-.t0 VDDA.t41 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X732 VOUT-.t156 two_stage_opamp_dummy_magic_29_0.cap_res_X.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X733 two_stage_opamp_dummy_magic_29_0.Vb3.t2 bgr_11_0.NFET_GATE_10uA.t22 GNDA_2.t246 GNDA_2.t245 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X734 VDDA.t219 bgr_11_0.PFET_GATE_10uA.t28 bgr_11_0.V_CUR_REF_REG.t1 VDDA.t218 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X735 GNDA_2.t2 bgr_11_0.NFET_GATE_10uA.t23 two_stage_opamp_dummy_magic_29_0.Vb3.t1 GNDA_2.t1 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X736 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.t8 two_stage_opamp_dummy_magic_29_0.Y.t52 GNDA_2.t227 VDDA.t142 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X737 VOUT-.t157 two_stage_opamp_dummy_magic_29_0.cap_res_X.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X738 bgr_11_0.1st_Vout_1.t32 bgr_11_0.cap_res1.t0 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X739 two_stage_opamp_dummy_magic_29_0.VD3.t18 two_stage_opamp_dummy_magic_29_0.Vb2.t31 two_stage_opamp_dummy_magic_29_0.X.t12 two_stage_opamp_dummy_magic_29_0.VD3.t17 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X740 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.t7 two_stage_opamp_dummy_magic_29_0.Y.t53 GNDA_2.t204 VDDA.t98 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X741 VOUT+.t160 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X742 a_5700_30088.t0 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref.t4 GNDA_2.t166 sky130_fd_pr__res_xhigh_po_0p35 l=4.28
X743 VOUT+.t161 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X744 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.t5 two_stage_opamp_dummy_magic_29_0.Y.t54 VDDA.t31 GNDA_2.t26 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X745 bgr_11_0.1st_Vout_2.t32 bgr_11_0.cap_res2.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X746 two_stage_opamp_dummy_magic_29_0.VD2.t4 VIN+.t8 two_stage_opamp_dummy_magic_29_0.V_source.t29 GNDA_2.t170 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X747 two_stage_opamp_dummy_magic_29_0.Y.t14 two_stage_opamp_dummy_magic_29_0.Vb2.t32 two_stage_opamp_dummy_magic_29_0.VD4.t13 two_stage_opamp_dummy_magic_29_0.VD4.t12 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X748 two_stage_opamp_dummy_magic_29_0.VD2.t16 VIN+.t9 two_stage_opamp_dummy_magic_29_0.V_source.t28 GNDA_2.t24 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X749 two_stage_opamp_dummy_magic_29_0.V_p_mir.t3 VIN+.t10 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t3 GNDA_2.t24 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X750 VOUT-.t158 two_stage_opamp_dummy_magic_29_0.cap_res_X.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X751 VOUT-.t159 two_stage_opamp_dummy_magic_29_0.cap_res_X.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X752 VOUT-.t160 two_stage_opamp_dummy_magic_29_0.cap_res_X.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X753 two_stage_opamp_dummy_magic_29_0.V_source.t38 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t31 GNDA_2.t257 GNDA_2.t6 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X754 a_3230_3878.t1 two_stage_opamp_dummy_magic_29_0.V_tot.t2 GNDA_2.t214 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X755 VOUT-.t161 two_stage_opamp_dummy_magic_29_0.cap_res_X.t0 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
R0 bgr_11_0.1st_Vout_2.n9 bgr_11_0.1st_Vout_2.t15 362.341
R1 bgr_11_0.1st_Vout_2.n7 bgr_11_0.1st_Vout_2.t14 355.094
R2 bgr_11_0.1st_Vout_2.n4 bgr_11_0.1st_Vout_2.n10 302.183
R3 bgr_11_0.1st_Vout_2.n7 bgr_11_0.1st_Vout_2.n6 302.183
R4 bgr_11_0.1st_Vout_2.n12 bgr_11_0.1st_Vout_2.n5 297.683
R5 bgr_11_0.1st_Vout_2.n11 bgr_11_0.1st_Vout_2.t26 194.809
R6 bgr_11_0.1st_Vout_2.n11 bgr_11_0.1st_Vout_2.t9 194.809
R7 bgr_11_0.1st_Vout_2.n8 bgr_11_0.1st_Vout_2.t21 194.809
R8 bgr_11_0.1st_Vout_2.n8 bgr_11_0.1st_Vout_2.t7 194.809
R9 bgr_11_0.1st_Vout_2.n4 bgr_11_0.1st_Vout_2.n11 166.03
R10 bgr_11_0.1st_Vout_2.n3 bgr_11_0.1st_Vout_2.n8 166.03
R11 bgr_11_0.1st_Vout_2.t6 bgr_11_0.1st_Vout_2.n12 49.5021
R12 bgr_11_0.1st_Vout_2.n10 bgr_11_0.1st_Vout_2.t2 39.4005
R13 bgr_11_0.1st_Vout_2.n10 bgr_11_0.1st_Vout_2.t0 39.4005
R14 bgr_11_0.1st_Vout_2.n6 bgr_11_0.1st_Vout_2.t1 39.4005
R15 bgr_11_0.1st_Vout_2.n6 bgr_11_0.1st_Vout_2.t4 39.4005
R16 bgr_11_0.1st_Vout_2.n5 bgr_11_0.1st_Vout_2.t3 39.4005
R17 bgr_11_0.1st_Vout_2.n5 bgr_11_0.1st_Vout_2.t5 39.4005
R18 bgr_11_0.1st_Vout_2.n9 bgr_11_0.1st_Vout_2.n0 35.7185
R19 bgr_11_0.1st_Vout_2.n1 bgr_11_0.1st_Vout_2.t32 4.8295
R20 bgr_11_0.1st_Vout_2.n1 bgr_11_0.1st_Vout_2.t12 4.8295
R21 bgr_11_0.1st_Vout_2.n2 bgr_11_0.1st_Vout_2.t13 4.8295
R22 bgr_11_0.1st_Vout_2.n2 bgr_11_0.1st_Vout_2.t19 4.8295
R23 bgr_11_0.1st_Vout_2.n2 bgr_11_0.1st_Vout_2.t30 4.8295
R24 bgr_11_0.1st_Vout_2.n2 bgr_11_0.1st_Vout_2.t11 4.8295
R25 bgr_11_0.1st_Vout_2.n0 bgr_11_0.1st_Vout_2.t23 4.8295
R26 bgr_11_0.1st_Vout_2.n0 bgr_11_0.1st_Vout_2.t28 4.8295
R27 bgr_11_0.1st_Vout_2.n0 bgr_11_0.1st_Vout_2.t8 4.8295
R28 bgr_11_0.1st_Vout_2.n1 bgr_11_0.1st_Vout_2.t27 4.5005
R29 bgr_11_0.1st_Vout_2.n1 bgr_11_0.1st_Vout_2.t20 4.5005
R30 bgr_11_0.1st_Vout_2.n2 bgr_11_0.1st_Vout_2.t31 4.5005
R31 bgr_11_0.1st_Vout_2.n2 bgr_11_0.1st_Vout_2.t25 4.5005
R32 bgr_11_0.1st_Vout_2.n2 bgr_11_0.1st_Vout_2.t24 4.5005
R33 bgr_11_0.1st_Vout_2.n2 bgr_11_0.1st_Vout_2.t18 4.5005
R34 bgr_11_0.1st_Vout_2.n0 bgr_11_0.1st_Vout_2.t17 4.5005
R35 bgr_11_0.1st_Vout_2.n0 bgr_11_0.1st_Vout_2.t10 4.5005
R36 bgr_11_0.1st_Vout_2.n0 bgr_11_0.1st_Vout_2.t29 4.5005
R37 bgr_11_0.1st_Vout_2.n0 bgr_11_0.1st_Vout_2.t22 4.5005
R38 bgr_11_0.1st_Vout_2.n0 bgr_11_0.1st_Vout_2.t16 4.5005
R39 bgr_11_0.1st_Vout_2.n12 bgr_11_0.1st_Vout_2.n3 4.5005
R40 bgr_11_0.1st_Vout_2.n4 bgr_11_0.1st_Vout_2.n9 2.90725
R41 bgr_11_0.1st_Vout_2.n0 bgr_11_0.1st_Vout_2.n2 2.2095
R42 bgr_11_0.1st_Vout_2.n3 bgr_11_0.1st_Vout_2.n4 1.1255
R43 bgr_11_0.1st_Vout_2.n3 bgr_11_0.1st_Vout_2.n7 1.1255
R44 bgr_11_0.1st_Vout_2.n2 bgr_11_0.1st_Vout_2.n1 0.8935
R45 bgr_11_0.PFET_GATE_10uA.n14 bgr_11_0.PFET_GATE_10uA.t26 614.04
R46 bgr_11_0.PFET_GATE_10uA.n4 bgr_11_0.PFET_GATE_10uA.n0 510.991
R47 bgr_11_0.PFET_GATE_10uA bgr_11_0.PFET_GATE_10uA.n25 509.226
R48 bgr_11_0.PFET_GATE_10uA.n22 bgr_11_0.PFET_GATE_10uA.t22 369.534
R49 bgr_11_0.PFET_GATE_10uA.n19 bgr_11_0.PFET_GATE_10uA.t27 369.534
R50 bgr_11_0.PFET_GATE_10uA.n16 bgr_11_0.PFET_GATE_10uA.t11 369.534
R51 bgr_11_0.PFET_GATE_10uA.n15 bgr_11_0.PFET_GATE_10uA.t10 369.534
R52 bgr_11_0.PFET_GATE_10uA.n2 bgr_11_0.PFET_GATE_10uA.t25 369.534
R53 bgr_11_0.PFET_GATE_10uA.n1 bgr_11_0.PFET_GATE_10uA.t24 369.534
R54 bgr_11_0.PFET_GATE_10uA.n12 bgr_11_0.PFET_GATE_10uA.n11 301.933
R55 bgr_11_0.PFET_GATE_10uA.n10 bgr_11_0.PFET_GATE_10uA.n9 301.933
R56 bgr_11_0.PFET_GATE_10uA.n8 bgr_11_0.PFET_GATE_10uA.n7 301.933
R57 bgr_11_0.PFET_GATE_10uA.n6 bgr_11_0.PFET_GATE_10uA.n5 301.933
R58 bgr_11_0.PFET_GATE_10uA.n0 bgr_11_0.PFET_GATE_10uA.t20 249.034
R59 bgr_11_0.PFET_GATE_10uA.n0 bgr_11_0.PFET_GATE_10uA.t28 249.034
R60 bgr_11_0.PFET_GATE_10uA.n22 bgr_11_0.PFET_GATE_10uA.t12 192.8
R61 bgr_11_0.PFET_GATE_10uA.n23 bgr_11_0.PFET_GATE_10uA.t16 192.8
R62 bgr_11_0.PFET_GATE_10uA.n24 bgr_11_0.PFET_GATE_10uA.t23 192.8
R63 bgr_11_0.PFET_GATE_10uA.n21 bgr_11_0.PFET_GATE_10uA.t14 192.8
R64 bgr_11_0.PFET_GATE_10uA.n20 bgr_11_0.PFET_GATE_10uA.t19 192.8
R65 bgr_11_0.PFET_GATE_10uA.n19 bgr_11_0.PFET_GATE_10uA.t18 192.8
R66 bgr_11_0.PFET_GATE_10uA.n16 bgr_11_0.PFET_GATE_10uA.t21 192.8
R67 bgr_11_0.PFET_GATE_10uA.n15 bgr_11_0.PFET_GATE_10uA.t15 192.8
R68 bgr_11_0.PFET_GATE_10uA.n2 bgr_11_0.PFET_GATE_10uA.t17 192.8
R69 bgr_11_0.PFET_GATE_10uA.n1 bgr_11_0.PFET_GATE_10uA.t13 192.8
R70 bgr_11_0.PFET_GATE_10uA.n21 bgr_11_0.PFET_GATE_10uA.n20 176.733
R71 bgr_11_0.PFET_GATE_10uA.n20 bgr_11_0.PFET_GATE_10uA.n19 176.733
R72 bgr_11_0.PFET_GATE_10uA.n23 bgr_11_0.PFET_GATE_10uA.n22 176.733
R73 bgr_11_0.PFET_GATE_10uA.n24 bgr_11_0.PFET_GATE_10uA.n23 176.733
R74 bgr_11_0.PFET_GATE_10uA.n18 bgr_11_0.PFET_GATE_10uA.n17 166.343
R75 bgr_11_0.PFET_GATE_10uA.n4 bgr_11_0.PFET_GATE_10uA.n3 166.343
R76 bgr_11_0.PFET_GATE_10uA.n13 bgr_11_0.PFET_GATE_10uA.t0 119.118
R77 bgr_11_0.PFET_GATE_10uA.n6 bgr_11_0.PFET_GATE_10uA.t1 104.474
R78 bgr_11_0.PFET_GATE_10uA.n17 bgr_11_0.PFET_GATE_10uA.n16 56.2338
R79 bgr_11_0.PFET_GATE_10uA.n17 bgr_11_0.PFET_GATE_10uA.n15 56.2338
R80 bgr_11_0.PFET_GATE_10uA.n3 bgr_11_0.PFET_GATE_10uA.n2 56.2338
R81 bgr_11_0.PFET_GATE_10uA.n3 bgr_11_0.PFET_GATE_10uA.n1 56.2338
R82 bgr_11_0.PFET_GATE_10uA.n25 bgr_11_0.PFET_GATE_10uA.n21 56.2338
R83 bgr_11_0.PFET_GATE_10uA.n25 bgr_11_0.PFET_GATE_10uA.n24 56.2338
R84 bgr_11_0.PFET_GATE_10uA.n11 bgr_11_0.PFET_GATE_10uA.t4 39.4005
R85 bgr_11_0.PFET_GATE_10uA.n11 bgr_11_0.PFET_GATE_10uA.t8 39.4005
R86 bgr_11_0.PFET_GATE_10uA.n9 bgr_11_0.PFET_GATE_10uA.t3 39.4005
R87 bgr_11_0.PFET_GATE_10uA.n9 bgr_11_0.PFET_GATE_10uA.t6 39.4005
R88 bgr_11_0.PFET_GATE_10uA.n7 bgr_11_0.PFET_GATE_10uA.t5 39.4005
R89 bgr_11_0.PFET_GATE_10uA.n7 bgr_11_0.PFET_GATE_10uA.t7 39.4005
R90 bgr_11_0.PFET_GATE_10uA.n5 bgr_11_0.PFET_GATE_10uA.t9 39.4005
R91 bgr_11_0.PFET_GATE_10uA.n5 bgr_11_0.PFET_GATE_10uA.t2 39.4005
R92 bgr_11_0.PFET_GATE_10uA.n18 bgr_11_0.PFET_GATE_10uA.n14 10.3755
R93 bgr_11_0.PFET_GATE_10uA.n13 bgr_11_0.PFET_GATE_10uA.n12 6.15675
R94 bgr_11_0.PFET_GATE_10uA bgr_11_0.PFET_GATE_10uA.n4 2.28175
R95 bgr_11_0.PFET_GATE_10uA bgr_11_0.PFET_GATE_10uA.n18 2.28175
R96 bgr_11_0.PFET_GATE_10uA.n14 bgr_11_0.PFET_GATE_10uA.n13 1.54738
R97 bgr_11_0.PFET_GATE_10uA.n8 bgr_11_0.PFET_GATE_10uA.n6 1.1255
R98 bgr_11_0.PFET_GATE_10uA.n10 bgr_11_0.PFET_GATE_10uA.n8 1.1255
R99 bgr_11_0.PFET_GATE_10uA.n12 bgr_11_0.PFET_GATE_10uA.n10 1.1255
R100 VDDA.n762 VDDA.t303 1231.74
R101 VDDA.n765 VDDA.t315 1231.74
R102 VDDA.n627 VDDA.t263 1231.74
R103 VDDA.n630 VDDA.t291 1231.74
R104 VDDA.n644 VDDA.t306 858.933
R105 VDDA.n689 VDDA.t281 858.933
R106 VDDA.n684 VDDA.t266 858.933
R107 VDDA.n188 VDDA.t336 858.933
R108 VDDA.t296 VDDA.n315 708.125
R109 VDDA.n338 VDDA.t296 708.125
R110 VDDA.n335 VDDA.t259 708.125
R111 VDDA.t259 VDDA.n316 708.125
R112 VDDA.t344 VDDA.n295 708.125
R113 VDDA.n348 VDDA.t344 708.125
R114 VDDA.n345 VDDA.t262 708.125
R115 VDDA.t262 VDDA.n296 708.125
R116 VDDA.t350 VDDA.n425 676.966
R117 VDDA.n655 VDDA.t272 661.375
R118 VDDA.n658 VDDA.t321 661.375
R119 VDDA.n706 VDDA.t352 661.375
R120 VDDA.n703 VDDA.t312 661.375
R121 VDDA.n202 VDDA.t361 661.375
R122 VDDA.n205 VDDA.t327 661.375
R123 VDDA.n337 VDDA.t295 657.76
R124 VDDA.n347 VDDA.t343 657.76
R125 VDDA.t298 VDDA.n455 648.726
R126 VDDA.n456 VDDA.t334 648.726
R127 VDDA.t285 VDDA.n442 648.726
R128 VDDA.n443 VDDA.t359 648.726
R129 VDDA.n426 VDDA.t319 643.038
R130 VDDA.n452 VDDA.t346 642.992
R131 VDDA.t331 VDDA.n451 642.992
R132 VDDA.n439 VDDA.t255 642.992
R133 VDDA.t340 VDDA.n438 642.992
R134 VDDA.n234 VDDA.t275 589.076
R135 VDDA.n237 VDDA.t300 589.076
R136 VDDA.n742 VDDA.t309 589.076
R137 VDDA.n739 VDDA.t324 589.076
R138 VDDA.n377 VDDA.n375 587.407
R139 VDDA.n381 VDDA.n378 587.407
R140 VDDA.n407 VDDA.n406 587.407
R141 VDDA.n402 VDDA.n368 587.407
R142 VDDA.n406 VDDA.n405 585
R143 VDDA.n404 VDDA.n402 585
R144 VDDA.n388 VDDA.n377 585
R145 VDDA.n385 VDDA.n378 585
R146 VDDA.t258 VDDA.n336 540.818
R147 VDDA.t261 VDDA.n346 540.818
R148 VDDA.n671 VDDA.t269 456.526
R149 VDDA.n668 VDDA.t287 456.526
R150 VDDA.n445 VDDA.t330 441.2
R151 VDDA.n453 VDDA.t345 441.2
R152 VDDA.n436 VDDA.t339 441.2
R153 VDDA.n440 VDDA.t254 441.2
R154 VDDA.n454 VDDA.t297 418.368
R155 VDDA.n457 VDDA.t333 418.368
R156 VDDA.n441 VDDA.t284 418.368
R157 VDDA.n444 VDDA.t358 418.368
R158 VDDA.n427 VDDA.t318 413.084
R159 VDDA.n424 VDDA.t349 413.084
R160 VDDA.t295 VDDA.t212 407.144
R161 VDDA.t212 VDDA.t29 407.144
R162 VDDA.t29 VDDA.t186 407.144
R163 VDDA.t186 VDDA.t376 407.144
R164 VDDA.t376 VDDA.t162 407.144
R165 VDDA.t162 VDDA.t216 407.144
R166 VDDA.t216 VDDA.t208 407.144
R167 VDDA.t208 VDDA.t126 407.144
R168 VDDA.t126 VDDA.t194 407.144
R169 VDDA.t194 VDDA.t114 407.144
R170 VDDA.t114 VDDA.t37 407.144
R171 VDDA.t37 VDDA.t214 407.144
R172 VDDA.t214 VDDA.t206 407.144
R173 VDDA.t206 VDDA.t62 407.144
R174 VDDA.t62 VDDA.t13 407.144
R175 VDDA.t13 VDDA.t77 407.144
R176 VDDA.t77 VDDA.t188 407.144
R177 VDDA.t188 VDDA.t210 407.144
R178 VDDA.t210 VDDA.t258 407.144
R179 VDDA.t343 VDDA.t33 407.144
R180 VDDA.t33 VDDA.t196 407.144
R181 VDDA.t196 VDDA.t1 407.144
R182 VDDA.t1 VDDA.t190 407.144
R183 VDDA.t190 VDDA.t160 407.144
R184 VDDA.t160 VDDA.t70 407.144
R185 VDDA.t70 VDDA.t5 407.144
R186 VDDA.t5 VDDA.t39 407.144
R187 VDDA.t39 VDDA.t46 407.144
R188 VDDA.t46 VDDA.t15 407.144
R189 VDDA.t15 VDDA.t7 407.144
R190 VDDA.t7 VDDA.t68 407.144
R191 VDDA.t68 VDDA.t66 407.144
R192 VDDA.t66 VDDA.t365 407.144
R193 VDDA.t365 VDDA.t192 407.144
R194 VDDA.t192 VDDA.t64 407.144
R195 VDDA.t64 VDDA.t158 407.144
R196 VDDA.t158 VDDA.t154 407.144
R197 VDDA.t154 VDDA.t261 407.144
R198 VDDA.n670 VDDA.t270 397.784
R199 VDDA.t288 VDDA.n669 397.784
R200 VDDA.t252 VDDA.t298 373.214
R201 VDDA.t242 VDDA.t252 373.214
R202 VDDA.t230 VDDA.t242 373.214
R203 VDDA.t250 VDDA.t230 373.214
R204 VDDA.t334 VDDA.t250 373.214
R205 VDDA.t228 VDDA.t331 373.214
R206 VDDA.t248 VDDA.t228 373.214
R207 VDDA.t240 VDDA.t248 373.214
R208 VDDA.t226 VDDA.t240 373.214
R209 VDDA.t244 VDDA.t226 373.214
R210 VDDA.t234 VDDA.t244 373.214
R211 VDDA.t236 VDDA.t234 373.214
R212 VDDA.t220 VDDA.t236 373.214
R213 VDDA.t346 VDDA.t220 373.214
R214 VDDA.t224 VDDA.t285 373.214
R215 VDDA.t246 VDDA.t224 373.214
R216 VDDA.t238 VDDA.t246 373.214
R217 VDDA.t222 VDDA.t238 373.214
R218 VDDA.t359 VDDA.t222 373.214
R219 VDDA.t232 VDDA.t340 373.214
R220 VDDA.t218 VDDA.t232 373.214
R221 VDDA.t255 VDDA.t218 373.214
R222 VDDA.t319 VDDA.t152 373.214
R223 VDDA.t152 VDDA.t164 373.214
R224 VDDA.t164 VDDA.t350 373.214
R225 VDDA.n340 VDDA.t294 370.168
R226 VDDA.n333 VDDA.t257 370.168
R227 VDDA.n350 VDDA.t342 370.168
R228 VDDA.n343 VDDA.t260 370.168
R229 VDDA.n359 VDDA.t278 360.868
R230 VDDA.n413 VDDA.t355 360.868
R231 VDDA.n452 VDDA.t348 354.154
R232 VDDA.n451 VDDA.t332 354.154
R233 VDDA.n439 VDDA.t256 354.154
R234 VDDA.n438 VDDA.t341 354.154
R235 VDDA.n426 VDDA.t320 354.063
R236 VDDA.n425 VDDA.t351 347.224
R237 VDDA.t276 VDDA.n235 343.882
R238 VDDA.n236 VDDA.t301 343.882
R239 VDDA.n741 VDDA.t310 343.882
R240 VDDA.t325 VDDA.n740 343.882
R241 VDDA.n464 VDDA.n450 336.341
R242 VDDA.n465 VDDA.n449 336.341
R243 VDDA.n466 VDDA.n448 336.341
R244 VDDA.n467 VDDA.n447 336.341
R245 VDDA.n468 VDDA.n446 336.341
R246 VDDA.n477 VDDA.n437 336.341
R247 VDDA.n455 VDDA.t299 331.901
R248 VDDA.n456 VDDA.t335 331.901
R249 VDDA.n442 VDDA.t286 331.901
R250 VDDA.n443 VDDA.t360 331.901
R251 VDDA.n332 VDDA.n331 299.231
R252 VDDA.n330 VDDA.n329 299.231
R253 VDDA.n328 VDDA.n327 299.231
R254 VDDA.n326 VDDA.n325 299.231
R255 VDDA.n324 VDDA.n323 299.231
R256 VDDA.n322 VDDA.n321 299.231
R257 VDDA.n320 VDDA.n319 299.231
R258 VDDA.n318 VDDA.n317 299.231
R259 VDDA.n314 VDDA.n313 299.231
R260 VDDA.n312 VDDA.n311 299.231
R261 VDDA.n310 VDDA.n309 299.231
R262 VDDA.n308 VDDA.n307 299.231
R263 VDDA.n306 VDDA.n305 299.231
R264 VDDA.n304 VDDA.n303 299.231
R265 VDDA.n302 VDDA.n301 299.231
R266 VDDA.n300 VDDA.n299 299.231
R267 VDDA.n298 VDDA.n297 299.231
R268 VDDA.n294 VDDA.n293 299.231
R269 VDDA.n459 VDDA.n458 299.053
R270 VDDA.n461 VDDA.n460 299.053
R271 VDDA.n472 VDDA.n471 299.053
R272 VDDA.n474 VDDA.n473 299.053
R273 VDDA.n643 VDDA.t307 282.788
R274 VDDA.n688 VDDA.t282 282.788
R275 VDDA.t270 VDDA.t134 259.091
R276 VDDA.t134 VDDA.t288 259.091
R277 VDDA.t387 VDDA.t279 251.471
R278 VDDA.t145 VDDA.t387 251.471
R279 VDDA.t380 VDDA.t145 251.471
R280 VDDA.t119 VDDA.t380 251.471
R281 VDDA.t147 VDDA.t119 251.471
R282 VDDA.t407 VDDA.t147 251.471
R283 VDDA.t383 VDDA.t407 251.471
R284 VDDA.t367 VDDA.t383 251.471
R285 VDDA.t172 VDDA.t367 251.471
R286 VDDA.t385 VDDA.t172 251.471
R287 VDDA.t102 VDDA.t385 251.471
R288 VDDA.t405 VDDA.t102 251.471
R289 VDDA.t121 VDDA.t405 251.471
R290 VDDA.t149 VDDA.t121 251.471
R291 VDDA.t105 VDDA.t149 251.471
R292 VDDA.t396 VDDA.t105 251.471
R293 VDDA.t356 VDDA.t396 251.471
R294 VDDA.n409 VDDA.n408 238.367
R295 VDDA.n336 VDDA.n335 238.367
R296 VDDA.n336 VDDA.n316 238.367
R297 VDDA.n346 VDDA.n345 238.367
R298 VDDA.n346 VDDA.n296 238.367
R299 VDDA.t279 VDDA.n393 237.5
R300 VDDA.n410 VDDA.t356 237.5
R301 VDDA.n187 VDDA.n186 222.524
R302 VDDA.n647 VDDA.n646 222.524
R303 VDDA.n687 VDDA.t337 221.121
R304 VDDA.t267 VDDA.n687 221.121
R305 VDDA.t76 VDDA.t276 217.708
R306 VDDA.t118 VDDA.t76 217.708
R307 VDDA.t74 VDDA.t118 217.708
R308 VDDA.t97 VDDA.t74 217.708
R309 VDDA.t128 VDDA.t97 217.708
R310 VDDA.t75 VDDA.t128 217.708
R311 VDDA.t185 VDDA.t75 217.708
R312 VDDA.t113 VDDA.t185 217.708
R313 VDDA.t43 VDDA.t113 217.708
R314 VDDA.t32 VDDA.t43 217.708
R315 VDDA.t301 VDDA.t32 217.708
R316 VDDA.t310 VDDA.t112 217.708
R317 VDDA.t112 VDDA.t98 217.708
R318 VDDA.t98 VDDA.t125 217.708
R319 VDDA.t125 VDDA.t165 217.708
R320 VDDA.t165 VDDA.t398 217.708
R321 VDDA.t398 VDDA.t52 217.708
R322 VDDA.t52 VDDA.t0 217.708
R323 VDDA.t0 VDDA.t21 217.708
R324 VDDA.t21 VDDA.t174 217.708
R325 VDDA.t174 VDDA.t142 217.708
R326 VDDA.t142 VDDA.t325 217.708
R327 VDDA.t273 VDDA.n656 213.131
R328 VDDA.n657 VDDA.t322 213.131
R329 VDDA.n705 VDDA.t353 213.131
R330 VDDA.t313 VDDA.n704 213.131
R331 VDDA.t362 VDDA.n203 213.131
R332 VDDA.n204 VDDA.t328 213.131
R333 VDDA.n398 VDDA.n396 185
R334 VDDA.n405 VDDA.n395 185
R335 VDDA.n410 VDDA.n395 185
R336 VDDA.n404 VDDA.n403 185
R337 VDDA.n401 VDDA.n370 185
R338 VDDA.n412 VDDA.n411 185
R339 VDDA.n411 VDDA.n410 185
R340 VDDA.n392 VDDA.n391 185
R341 VDDA.n393 VDDA.n392 185
R342 VDDA.n389 VDDA.n374 185
R343 VDDA.n388 VDDA.n387 185
R344 VDDA.n386 VDDA.n385 185
R345 VDDA.n380 VDDA.n379 185
R346 VDDA.n382 VDDA.n373 185
R347 VDDA.n393 VDDA.n373 185
R348 VDDA.t307 VDDA.t378 180.173
R349 VDDA.t378 VDDA.t27 180.173
R350 VDDA.t27 VDDA.t58 180.173
R351 VDDA.t58 VDDA.t375 180.173
R352 VDDA.t375 VDDA.t337 180.173
R353 VDDA.t372 VDDA.t267 180.173
R354 VDDA.t373 VDDA.t372 180.173
R355 VDDA.t25 VDDA.t373 180.173
R356 VDDA.t72 VDDA.t25 180.173
R357 VDDA.t282 VDDA.t72 180.173
R358 VDDA.n670 VDDA.t271 168.139
R359 VDDA.n669 VDDA.t290 168.139
R360 VDDA.n667 VDDA.n666 150.643
R361 VDDA.n396 VDDA.n395 150
R362 VDDA.n403 VDDA.n395 150
R363 VDDA.n411 VDDA.n370 150
R364 VDDA.n392 VDDA.n374 150
R365 VDDA.n387 VDDA.n386 150
R366 VDDA.n379 VDDA.n373 150
R367 VDDA.t85 VDDA.t273 146.155
R368 VDDA.t322 VDDA.t85 146.155
R369 VDDA.t353 VDDA.t116 146.155
R370 VDDA.t116 VDDA.t169 146.155
R371 VDDA.t169 VDDA.t200 146.155
R372 VDDA.t200 VDDA.t60 146.155
R373 VDDA.t60 VDDA.t3 146.155
R374 VDDA.t3 VDDA.t178 146.155
R375 VDDA.t178 VDDA.t9 146.155
R376 VDDA.t9 VDDA.t182 146.155
R377 VDDA.t182 VDDA.t79 146.155
R378 VDDA.t79 VDDA.t99 146.155
R379 VDDA.t99 VDDA.t313 146.155
R380 VDDA.t11 VDDA.t362 146.155
R381 VDDA.t393 VDDA.t11 146.155
R382 VDDA.t95 VDDA.t393 146.155
R383 VDDA.t180 VDDA.t95 146.155
R384 VDDA.t83 VDDA.t180 146.155
R385 VDDA.t35 VDDA.t83 146.155
R386 VDDA.t89 VDDA.t35 146.155
R387 VDDA.t204 VDDA.t89 146.155
R388 VDDA.t50 VDDA.t204 146.155
R389 VDDA.t156 VDDA.t50 146.155
R390 VDDA.t328 VDDA.t156 146.155
R391 VDDA.n414 VDDA.n367 141.712
R392 VDDA.n415 VDDA.n366 141.712
R393 VDDA.n416 VDDA.n365 141.712
R394 VDDA.n417 VDDA.n364 141.712
R395 VDDA.n418 VDDA.n363 141.712
R396 VDDA.n419 VDDA.n362 141.712
R397 VDDA.n420 VDDA.n361 141.712
R398 VDDA.n421 VDDA.n360 141.712
R399 VDDA.n235 VDDA.t277 136.701
R400 VDDA.n236 VDDA.t302 136.701
R401 VDDA.n741 VDDA.t311 136.701
R402 VDDA.n740 VDDA.t326 136.701
R403 VDDA.t280 VDDA.n377 123.126
R404 VDDA.n378 VDDA.t280 123.126
R405 VDDA.n406 VDDA.t357 123.126
R406 VDDA.n402 VDDA.t357 123.126
R407 VDDA.t304 VDDA.n763 122.829
R408 VDDA.n764 VDDA.t316 122.829
R409 VDDA.t264 VDDA.n628 122.829
R410 VDDA.n629 VDDA.t292 122.829
R411 VDDA.n643 VDDA.t308 113.26
R412 VDDA.n688 VDDA.t283 113.26
R413 VDDA.n686 VDDA.t268 113.26
R414 VDDA.n686 VDDA.t338 113.26
R415 VDDA.n689 VDDA.n688 82.7434
R416 VDDA.n644 VDDA.n643 82.7434
R417 VDDA.t391 VDDA.t304 81.6411
R418 VDDA.t110 VDDA.t391 81.6411
R419 VDDA.t370 VDDA.t110 81.6411
R420 VDDA.t389 VDDA.t370 81.6411
R421 VDDA.t399 VDDA.t389 81.6411
R422 VDDA.t123 VDDA.t399 81.6411
R423 VDDA.t137 VDDA.t123 81.6411
R424 VDDA.t140 VDDA.t137 81.6411
R425 VDDA.t53 VDDA.t140 81.6411
R426 VDDA.t19 VDDA.t53 81.6411
R427 VDDA.t316 VDDA.t19 81.6411
R428 VDDA.t175 VDDA.t264 81.6411
R429 VDDA.t41 VDDA.t175 81.6411
R430 VDDA.t56 VDDA.t41 81.6411
R431 VDDA.t132 VDDA.t56 81.6411
R432 VDDA.t198 VDDA.t132 81.6411
R433 VDDA.t44 VDDA.t198 81.6411
R434 VDDA.t167 VDDA.t44 81.6411
R435 VDDA.t48 VDDA.t167 81.6411
R436 VDDA.t202 VDDA.t48 81.6411
R437 VDDA.t129 VDDA.t202 81.6411
R438 VDDA.t292 VDDA.t129 81.6411
R439 VDDA.n656 VDDA.t274 76.2576
R440 VDDA.n657 VDDA.t323 76.2576
R441 VDDA.n705 VDDA.t354 76.2576
R442 VDDA.n704 VDDA.t314 76.2576
R443 VDDA.n203 VDDA.t363 76.2576
R444 VDDA.n204 VDDA.t329 76.2576
R445 VDDA.n702 VDDA.n701 71.388
R446 VDDA.n700 VDDA.n699 71.388
R447 VDDA.n698 VDDA.n697 71.388
R448 VDDA.n696 VDDA.n695 71.388
R449 VDDA.n694 VDDA.n693 71.388
R450 VDDA.n193 VDDA.n192 71.388
R451 VDDA.n195 VDDA.n194 71.388
R452 VDDA.n197 VDDA.n196 71.388
R453 VDDA.n199 VDDA.n198 71.388
R454 VDDA.n201 VDDA.n200 71.388
R455 VDDA.n654 VDDA.n653 68.4557
R456 VDDA.n410 VDDA.n409 65.8183
R457 VDDA.n410 VDDA.n394 65.8183
R458 VDDA.n393 VDDA.n371 65.8183
R459 VDDA.n393 VDDA.n372 65.8183
R460 VDDA.n687 VDDA.n686 61.6672
R461 VDDA.n685 VDDA.n684 60.8005
R462 VDDA.n685 VDDA.n188 60.8005
R463 VDDA.n284 VDDA.t412 58.8005
R464 VDDA.n283 VDDA.t414 58.8005
R465 VDDA.n403 VDDA.n394 53.3664
R466 VDDA.n409 VDDA.n396 53.3664
R467 VDDA.n394 VDDA.n370 53.3664
R468 VDDA.n374 VDDA.n371 53.3664
R469 VDDA.n386 VDDA.n372 53.3664
R470 VDDA.n387 VDDA.n371 53.3664
R471 VDDA.n379 VDDA.n372 53.3664
R472 VDDA.n283 VDDA.t415 49.1638
R473 VDDA.n285 VDDA.t413 48.5162
R474 VDDA.n763 VDDA.t305 40.9789
R475 VDDA.n764 VDDA.t317 40.9789
R476 VDDA.n628 VDDA.t265 40.9789
R477 VDDA.n629 VDDA.t293 40.9789
R478 VDDA.n450 VDDA.t221 39.4005
R479 VDDA.n450 VDDA.t347 39.4005
R480 VDDA.n449 VDDA.t235 39.4005
R481 VDDA.n449 VDDA.t237 39.4005
R482 VDDA.n448 VDDA.t227 39.4005
R483 VDDA.n448 VDDA.t245 39.4005
R484 VDDA.n447 VDDA.t249 39.4005
R485 VDDA.n447 VDDA.t241 39.4005
R486 VDDA.t332 VDDA.n446 39.4005
R487 VDDA.n446 VDDA.t229 39.4005
R488 VDDA.n437 VDDA.t233 39.4005
R489 VDDA.n437 VDDA.t219 39.4005
R490 VDDA.n458 VDDA.t231 39.4005
R491 VDDA.n458 VDDA.t251 39.4005
R492 VDDA.n460 VDDA.t253 39.4005
R493 VDDA.n460 VDDA.t243 39.4005
R494 VDDA.n471 VDDA.t239 39.4005
R495 VDDA.n471 VDDA.t223 39.4005
R496 VDDA.n473 VDDA.t225 39.4005
R497 VDDA.n473 VDDA.t247 39.4005
R498 VDDA.n331 VDDA.t189 39.4005
R499 VDDA.n331 VDDA.t211 39.4005
R500 VDDA.n329 VDDA.t14 39.4005
R501 VDDA.n329 VDDA.t78 39.4005
R502 VDDA.n327 VDDA.t207 39.4005
R503 VDDA.n327 VDDA.t63 39.4005
R504 VDDA.n325 VDDA.t38 39.4005
R505 VDDA.n325 VDDA.t215 39.4005
R506 VDDA.n323 VDDA.t195 39.4005
R507 VDDA.n323 VDDA.t115 39.4005
R508 VDDA.n321 VDDA.t209 39.4005
R509 VDDA.n321 VDDA.t127 39.4005
R510 VDDA.n319 VDDA.t163 39.4005
R511 VDDA.n319 VDDA.t217 39.4005
R512 VDDA.n317 VDDA.t187 39.4005
R513 VDDA.n317 VDDA.t377 39.4005
R514 VDDA.n313 VDDA.t213 39.4005
R515 VDDA.n313 VDDA.t30 39.4005
R516 VDDA.n311 VDDA.t159 39.4005
R517 VDDA.n311 VDDA.t155 39.4005
R518 VDDA.n309 VDDA.t193 39.4005
R519 VDDA.n309 VDDA.t65 39.4005
R520 VDDA.n307 VDDA.t67 39.4005
R521 VDDA.n307 VDDA.t366 39.4005
R522 VDDA.n305 VDDA.t8 39.4005
R523 VDDA.n305 VDDA.t69 39.4005
R524 VDDA.n303 VDDA.t47 39.4005
R525 VDDA.n303 VDDA.t16 39.4005
R526 VDDA.n301 VDDA.t6 39.4005
R527 VDDA.n301 VDDA.t40 39.4005
R528 VDDA.n299 VDDA.t161 39.4005
R529 VDDA.n299 VDDA.t71 39.4005
R530 VDDA.n297 VDDA.t2 39.4005
R531 VDDA.n297 VDDA.t191 39.4005
R532 VDDA.n293 VDDA.t34 39.4005
R533 VDDA.n293 VDDA.t197 39.4005
R534 VDDA.n181 VDDA.n180 38.2695
R535 VDDA.n754 VDDA.n753 38.2695
R536 VDDA.n756 VDDA.n755 38.2695
R537 VDDA.n758 VDDA.n757 38.2695
R538 VDDA.n760 VDDA.n759 38.2695
R539 VDDA.n246 VDDA.n245 38.2695
R540 VDDA.n619 VDDA.n618 38.2695
R541 VDDA.n621 VDDA.n620 38.2695
R542 VDDA.n623 VDDA.n622 38.2695
R543 VDDA.n625 VDDA.n624 38.2695
R544 VDDA.n220 VDDA.n218 26.8887
R545 VDDA.n724 VDDA.n722 26.8887
R546 VDDA.n228 VDDA.n227 26.7741
R547 VDDA.n226 VDDA.n225 26.7741
R548 VDDA.n224 VDDA.n223 26.7741
R549 VDDA.n222 VDDA.n221 26.7741
R550 VDDA.n220 VDDA.n219 26.7741
R551 VDDA.n724 VDDA.n723 26.7741
R552 VDDA.n726 VDDA.n725 26.7741
R553 VDDA.n728 VDDA.n727 26.7741
R554 VDDA.n730 VDDA.n729 26.7741
R555 VDDA.n732 VDDA.n731 26.7741
R556 VDDA.n453 VDDA.n452 24.9931
R557 VDDA.n451 VDDA.n445 24.9931
R558 VDDA.n440 VDDA.n439 24.9931
R559 VDDA.n438 VDDA.n436 24.9931
R560 VDDA.n48 VDDA.t369 24.1029
R561 VDDA.n427 VDDA.n426 22.9536
R562 VDDA.n413 VDDA.n412 22.8576
R563 VDDA.n382 VDDA.n359 22.8576
R564 VDDA.n666 VDDA.t135 21.8894
R565 VDDA.n666 VDDA.t289 21.8894
R566 VDDA.n425 VDDA.n424 20.4312
R567 VDDA.n186 VDDA.t374 15.7605
R568 VDDA.n186 VDDA.t26 15.7605
R569 VDDA.n646 VDDA.t28 15.7605
R570 VDDA.n646 VDDA.t59 15.7605
R571 VDDA.n686 VDDA.n685 13.9641
R572 VDDA.n367 VDDA.t106 13.1338
R573 VDDA.n367 VDDA.t397 13.1338
R574 VDDA.n366 VDDA.t122 13.1338
R575 VDDA.n366 VDDA.t150 13.1338
R576 VDDA.n365 VDDA.t103 13.1338
R577 VDDA.n365 VDDA.t406 13.1338
R578 VDDA.n364 VDDA.t173 13.1338
R579 VDDA.n364 VDDA.t386 13.1338
R580 VDDA.n363 VDDA.t384 13.1338
R581 VDDA.n363 VDDA.t368 13.1338
R582 VDDA.n362 VDDA.t148 13.1338
R583 VDDA.n362 VDDA.t408 13.1338
R584 VDDA.n361 VDDA.t381 13.1338
R585 VDDA.n361 VDDA.t120 13.1338
R586 VDDA.n360 VDDA.t388 13.1338
R587 VDDA.n360 VDDA.t146 13.1338
R588 VDDA.n424 VDDA.n423 11.37
R589 VDDA.n428 VDDA.n427 11.37
R590 VDDA.t274 VDDA.n654 11.2576
R591 VDDA.n654 VDDA.t86 11.2576
R592 VDDA.n701 VDDA.t80 11.2576
R593 VDDA.n701 VDDA.t100 11.2576
R594 VDDA.n699 VDDA.t10 11.2576
R595 VDDA.n699 VDDA.t183 11.2576
R596 VDDA.n697 VDDA.t4 11.2576
R597 VDDA.n697 VDDA.t179 11.2576
R598 VDDA.n695 VDDA.t201 11.2576
R599 VDDA.n695 VDDA.t61 11.2576
R600 VDDA.n693 VDDA.t117 11.2576
R601 VDDA.n693 VDDA.t170 11.2576
R602 VDDA.n192 VDDA.t51 11.2576
R603 VDDA.n192 VDDA.t157 11.2576
R604 VDDA.n194 VDDA.t90 11.2576
R605 VDDA.n194 VDDA.t205 11.2576
R606 VDDA.n196 VDDA.t84 11.2576
R607 VDDA.n196 VDDA.t36 11.2576
R608 VDDA.n198 VDDA.t96 11.2576
R609 VDDA.n198 VDDA.t181 11.2576
R610 VDDA.n200 VDDA.t12 11.2576
R611 VDDA.n200 VDDA.t394 11.2576
R612 VDDA.n414 VDDA.n413 11.0575
R613 VDDA.n469 VDDA.n445 10.87
R614 VDDA.n478 VDDA.n436 10.87
R615 VDDA.n476 VDDA.n440 10.87
R616 VDDA.n463 VDDA.n453 10.87
R617 VDDA.n422 VDDA.n359 10.87
R618 VDDA.n645 VDDA.n644 10.8696
R619 VDDA.n690 VDDA.n689 10.869
R620 VDDA.n391 VDDA.n390 9.50883
R621 VDDA.n383 VDDA.n382 9.50883
R622 VDDA.n408 VDDA.n397 9.50883
R623 VDDA.n412 VDDA.n369 9.50883
R624 VDDA.n339 VDDA.n315 9.50883
R625 VDDA.n349 VDDA.n295 9.50883
R626 VDDA.n401 VDDA.n369 9.3005
R627 VDDA.n404 VDDA.n400 9.3005
R628 VDDA.n405 VDDA.n399 9.3005
R629 VDDA.n398 VDDA.n397 9.3005
R630 VDDA.n383 VDDA.n380 9.3005
R631 VDDA.n385 VDDA.n384 9.3005
R632 VDDA.n388 VDDA.n376 9.3005
R633 VDDA.n390 VDDA.n389 9.3005
R634 VDDA.n339 VDDA.n338 9.3005
R635 VDDA.n349 VDDA.n348 9.3005
R636 VDDA.n684 VDDA.n683 9.3005
R637 VDDA.n683 VDDA.n188 9.3005
R638 VDDA.n405 VDDA.n398 9.14336
R639 VDDA.n405 VDDA.n404 9.14336
R640 VDDA.n404 VDDA.n401 9.14336
R641 VDDA.n389 VDDA.n388 9.14336
R642 VDDA.n388 VDDA.n385 9.14336
R643 VDDA.n385 VDDA.n380 9.14336
R644 VDDA.n227 VDDA.t131 8.0005
R645 VDDA.n227 VDDA.t402 8.0005
R646 VDDA.n225 VDDA.t73 8.0005
R647 VDDA.n225 VDDA.t364 8.0005
R648 VDDA.n223 VDDA.t91 8.0005
R649 VDDA.n223 VDDA.t92 8.0005
R650 VDDA.n221 VDDA.t184 8.0005
R651 VDDA.n221 VDDA.t94 8.0005
R652 VDDA.n219 VDDA.t177 8.0005
R653 VDDA.n219 VDDA.t55 8.0005
R654 VDDA.n218 VDDA.t401 8.0005
R655 VDDA.n218 VDDA.t93 8.0005
R656 VDDA.n722 VDDA.t22 8.0005
R657 VDDA.n722 VDDA.t404 8.0005
R658 VDDA.n723 VDDA.t166 8.0005
R659 VDDA.n723 VDDA.t23 8.0005
R660 VDDA.n725 VDDA.t153 8.0005
R661 VDDA.n725 VDDA.t136 8.0005
R662 VDDA.n727 VDDA.t31 8.0005
R663 VDDA.n727 VDDA.t109 8.0005
R664 VDDA.n729 VDDA.t139 8.0005
R665 VDDA.n729 VDDA.t24 8.0005
R666 VDDA.n731 VDDA.t403 8.0005
R667 VDDA.n731 VDDA.t411 8.0005
R668 VDDA.n180 VDDA.t54 6.56717
R669 VDDA.n180 VDDA.t20 6.56717
R670 VDDA.n753 VDDA.t138 6.56717
R671 VDDA.n753 VDDA.t141 6.56717
R672 VDDA.n755 VDDA.t400 6.56717
R673 VDDA.n755 VDDA.t124 6.56717
R674 VDDA.n757 VDDA.t371 6.56717
R675 VDDA.n757 VDDA.t390 6.56717
R676 VDDA.n759 VDDA.t392 6.56717
R677 VDDA.n759 VDDA.t111 6.56717
R678 VDDA.n245 VDDA.t203 6.56717
R679 VDDA.n245 VDDA.t130 6.56717
R680 VDDA.n618 VDDA.t168 6.56717
R681 VDDA.n618 VDDA.t49 6.56717
R682 VDDA.n620 VDDA.t199 6.56717
R683 VDDA.n620 VDDA.t45 6.56717
R684 VDDA.n622 VDDA.t57 6.56717
R685 VDDA.n622 VDDA.t133 6.56717
R686 VDDA.n624 VDDA.t176 6.56717
R687 VDDA.n624 VDDA.t42 6.56717
R688 VDDA.n408 VDDA.n407 5.33286
R689 VDDA.n412 VDDA.n368 5.33286
R690 VDDA.n391 VDDA.n375 5.33286
R691 VDDA.n382 VDDA.n381 5.33286
R692 VDDA.n457 VDDA.n456 4.98383
R693 VDDA.n455 VDDA.n454 4.98383
R694 VDDA.n444 VDDA.n443 4.98383
R695 VDDA.n442 VDDA.n441 4.98383
R696 VDDA.n703 VDDA.n702 4.8755
R697 VDDA.n202 VDDA.n201 4.8755
R698 VDDA.n772 VDDA.n771 4.58383
R699 VDDA.n615 VDDA.n611 4.58383
R700 VDDA.n48 VDDA.n47 4.5005
R701 VDDA.n49 VDDA.n41 4.5005
R702 VDDA.n53 VDDA.n50 4.5005
R703 VDDA.n54 VDDA.n40 4.5005
R704 VDDA.n58 VDDA.n57 4.5005
R705 VDDA.n59 VDDA.n39 4.5005
R706 VDDA.n63 VDDA.n60 4.5005
R707 VDDA.n64 VDDA.n38 4.5005
R708 VDDA.n68 VDDA.n67 4.5005
R709 VDDA.n69 VDDA.n37 4.5005
R710 VDDA.n73 VDDA.n70 4.5005
R711 VDDA.n74 VDDA.n36 4.5005
R712 VDDA.n78 VDDA.n77 4.5005
R713 VDDA.n79 VDDA.n35 4.5005
R714 VDDA.n83 VDDA.n80 4.5005
R715 VDDA.n84 VDDA.n34 4.5005
R716 VDDA.n88 VDDA.n87 4.5005
R717 VDDA.n89 VDDA.n33 4.5005
R718 VDDA.n93 VDDA.n90 4.5005
R719 VDDA.n94 VDDA.n32 4.5005
R720 VDDA.n98 VDDA.n97 4.5005
R721 VDDA.n289 VDDA.n288 4.5005
R722 VDDA.n355 VDDA.n354 4.5005
R723 VDDA.n432 VDDA.n431 4.5005
R724 VDDA.n482 VDDA.n481 4.5005
R725 VDDA.n485 VDDA.n274 4.5005
R726 VDDA.n488 VDDA.n486 4.5005
R727 VDDA.n489 VDDA.n273 4.5005
R728 VDDA.n493 VDDA.n492 4.5005
R729 VDDA.n494 VDDA.n272 4.5005
R730 VDDA.n498 VDDA.n495 4.5005
R731 VDDA.n499 VDDA.n271 4.5005
R732 VDDA.n503 VDDA.n502 4.5005
R733 VDDA.n504 VDDA.n270 4.5005
R734 VDDA.n508 VDDA.n505 4.5005
R735 VDDA.n509 VDDA.n269 4.5005
R736 VDDA.n513 VDDA.n512 4.5005
R737 VDDA.n514 VDDA.n268 4.5005
R738 VDDA.n518 VDDA.n515 4.5005
R739 VDDA.n519 VDDA.n267 4.5005
R740 VDDA.n523 VDDA.n522 4.5005
R741 VDDA.n524 VDDA.n266 4.5005
R742 VDDA.n528 VDDA.n525 4.5005
R743 VDDA.n529 VDDA.n265 4.5005
R744 VDDA.n533 VDDA.n532 4.5005
R745 VDDA.n676 VDDA.n650 4.5005
R746 VDDA.n661 VDDA.n652 4.5005
R747 VDDA.n137 VDDA.n136 4.5005
R748 VDDA.n138 VDDA.n131 4.5005
R749 VDDA.n142 VDDA.n141 4.5005
R750 VDDA.n143 VDDA.n128 4.5005
R751 VDDA.n145 VDDA.n144 4.5005
R752 VDDA.n146 VDDA.n127 4.5005
R753 VDDA.n150 VDDA.n149 4.5005
R754 VDDA.n151 VDDA.n124 4.5005
R755 VDDA.n153 VDDA.n152 4.5005
R756 VDDA.n154 VDDA.n123 4.5005
R757 VDDA.n158 VDDA.n157 4.5005
R758 VDDA.n159 VDDA.n120 4.5005
R759 VDDA.n161 VDDA.n160 4.5005
R760 VDDA.n162 VDDA.n119 4.5005
R761 VDDA.n166 VDDA.n165 4.5005
R762 VDDA.n167 VDDA.n116 4.5005
R763 VDDA.n169 VDDA.n168 4.5005
R764 VDDA.n170 VDDA.n115 4.5005
R765 VDDA.n174 VDDA.n173 4.5005
R766 VDDA.n175 VDDA.n114 4.5005
R767 VDDA.n773 VDDA.n772 4.5005
R768 VDDA.n767 VDDA.n177 4.5005
R769 VDDA.n769 VDDA.n768 4.5005
R770 VDDA.n768 VDDA.n767 4.5005
R771 VDDA.n707 VDDA.n706 4.5005
R772 VDDA.n713 VDDA.n183 4.5005
R773 VDDA.n716 VDDA.n715 4.5005
R774 VDDA.n719 VDDA.n718 4.5005
R775 VDDA.n711 VDDA.n691 4.5005
R776 VDDA.n712 VDDA.n185 4.5005
R777 VDDA.n712 VDDA.n711 4.5005
R778 VDDA.n680 VDDA.n648 4.5005
R779 VDDA.n683 VDDA.n682 4.5005
R780 VDDA.n206 VDDA.n205 4.5005
R781 VDDA.n207 VDDA.n191 4.5005
R782 VDDA.n214 VDDA.n213 4.5005
R783 VDDA.n217 VDDA.n216 4.5005
R784 VDDA.n632 VDDA.n209 4.5005
R785 VDDA.n634 VDDA.n633 4.5005
R786 VDDA.n633 VDDA.n632 4.5005
R787 VDDA.n612 VDDA.n248 4.5005
R788 VDDA.n604 VDDA.n549 4.5005
R789 VDDA.n603 VDDA.n550 4.5005
R790 VDDA.n600 VDDA.n551 4.5005
R791 VDDA.n599 VDDA.n552 4.5005
R792 VDDA.n596 VDDA.n553 4.5005
R793 VDDA.n595 VDDA.n554 4.5005
R794 VDDA.n592 VDDA.n555 4.5005
R795 VDDA.n591 VDDA.n556 4.5005
R796 VDDA.n588 VDDA.n557 4.5005
R797 VDDA.n587 VDDA.n558 4.5005
R798 VDDA.n584 VDDA.n559 4.5005
R799 VDDA.n583 VDDA.n560 4.5005
R800 VDDA.n580 VDDA.n561 4.5005
R801 VDDA.n579 VDDA.n562 4.5005
R802 VDDA.n576 VDDA.n563 4.5005
R803 VDDA.n575 VDDA.n564 4.5005
R804 VDDA.n572 VDDA.n565 4.5005
R805 VDDA.n571 VDDA.n566 4.5005
R806 VDDA.n568 VDDA.n567 4.5005
R807 VDDA.n250 VDDA.n249 4.5005
R808 VDDA.n611 VDDA.n610 4.5005
R809 VDDA.n338 VDDA.n337 4.48641
R810 VDDA.n337 VDDA.n315 4.48641
R811 VDDA.n348 VDDA.n347 4.48641
R812 VDDA.n347 VDDA.n295 4.48641
R813 VDDA.n407 VDDA.n398 3.75335
R814 VDDA.n401 VDDA.n368 3.75335
R815 VDDA.n389 VDDA.n375 3.75335
R816 VDDA.n381 VDDA.n380 3.75335
R817 VDDA.n135 VDDA.n112 3.50398
R818 VDDA.n607 VDDA.n547 3.50398
R819 VDDA.n100 VDDA.n99 3.48334
R820 VDDA.n535 VDDA.n534 3.48334
R821 VDDA.n47 VDDA.n29 3.43627
R822 VDDA.n334 VDDA.n333 3.41464
R823 VDDA.n344 VDDA.n343 3.41464
R824 VDDA.n31 VDDA.n30 3.4105
R825 VDDA.n97 VDDA.n96 3.4105
R826 VDDA.n95 VDDA.n94 3.4105
R827 VDDA.n93 VDDA.n92 3.4105
R828 VDDA.n91 VDDA.n33 3.4105
R829 VDDA.n87 VDDA.n86 3.4105
R830 VDDA.n85 VDDA.n84 3.4105
R831 VDDA.n83 VDDA.n82 3.4105
R832 VDDA.n81 VDDA.n35 3.4105
R833 VDDA.n77 VDDA.n76 3.4105
R834 VDDA.n75 VDDA.n74 3.4105
R835 VDDA.n73 VDDA.n72 3.4105
R836 VDDA.n71 VDDA.n37 3.4105
R837 VDDA.n67 VDDA.n66 3.4105
R838 VDDA.n65 VDDA.n64 3.4105
R839 VDDA.n63 VDDA.n62 3.4105
R840 VDDA.n61 VDDA.n39 3.4105
R841 VDDA.n57 VDDA.n56 3.4105
R842 VDDA.n55 VDDA.n54 3.4105
R843 VDDA.n53 VDDA.n52 3.4105
R844 VDDA.n51 VDDA.n41 3.4105
R845 VDDA.n264 VDDA.n263 3.4105
R846 VDDA.n532 VDDA.n531 3.4105
R847 VDDA.n530 VDDA.n529 3.4105
R848 VDDA.n528 VDDA.n527 3.4105
R849 VDDA.n526 VDDA.n266 3.4105
R850 VDDA.n522 VDDA.n521 3.4105
R851 VDDA.n520 VDDA.n519 3.4105
R852 VDDA.n518 VDDA.n517 3.4105
R853 VDDA.n516 VDDA.n268 3.4105
R854 VDDA.n512 VDDA.n511 3.4105
R855 VDDA.n510 VDDA.n509 3.4105
R856 VDDA.n508 VDDA.n507 3.4105
R857 VDDA.n506 VDDA.n270 3.4105
R858 VDDA.n502 VDDA.n501 3.4105
R859 VDDA.n500 VDDA.n499 3.4105
R860 VDDA.n498 VDDA.n497 3.4105
R861 VDDA.n496 VDDA.n272 3.4105
R862 VDDA.n492 VDDA.n491 3.4105
R863 VDDA.n490 VDDA.n489 3.4105
R864 VDDA.n488 VDDA.n487 3.4105
R865 VDDA.n114 VDDA.n113 3.4105
R866 VDDA.n173 VDDA.n172 3.4105
R867 VDDA.n171 VDDA.n170 3.4105
R868 VDDA.n169 VDDA.n118 3.4105
R869 VDDA.n117 VDDA.n116 3.4105
R870 VDDA.n165 VDDA.n164 3.4105
R871 VDDA.n163 VDDA.n162 3.4105
R872 VDDA.n161 VDDA.n122 3.4105
R873 VDDA.n121 VDDA.n120 3.4105
R874 VDDA.n157 VDDA.n156 3.4105
R875 VDDA.n155 VDDA.n154 3.4105
R876 VDDA.n153 VDDA.n126 3.4105
R877 VDDA.n125 VDDA.n124 3.4105
R878 VDDA.n149 VDDA.n148 3.4105
R879 VDDA.n147 VDDA.n146 3.4105
R880 VDDA.n145 VDDA.n130 3.4105
R881 VDDA.n129 VDDA.n128 3.4105
R882 VDDA.n141 VDDA.n140 3.4105
R883 VDDA.n139 VDDA.n138 3.4105
R884 VDDA.n137 VDDA.n134 3.4105
R885 VDDA.n133 VDDA.n132 3.4105
R886 VDDA.n774 VDDA.n773 3.4105
R887 VDDA.n251 VDDA.n250 3.4105
R888 VDDA.n569 VDDA.n568 3.4105
R889 VDDA.n571 VDDA.n570 3.4105
R890 VDDA.n573 VDDA.n572 3.4105
R891 VDDA.n575 VDDA.n574 3.4105
R892 VDDA.n577 VDDA.n576 3.4105
R893 VDDA.n579 VDDA.n578 3.4105
R894 VDDA.n581 VDDA.n580 3.4105
R895 VDDA.n583 VDDA.n582 3.4105
R896 VDDA.n585 VDDA.n584 3.4105
R897 VDDA.n587 VDDA.n586 3.4105
R898 VDDA.n589 VDDA.n588 3.4105
R899 VDDA.n591 VDDA.n590 3.4105
R900 VDDA.n593 VDDA.n592 3.4105
R901 VDDA.n595 VDDA.n594 3.4105
R902 VDDA.n597 VDDA.n596 3.4105
R903 VDDA.n599 VDDA.n598 3.4105
R904 VDDA.n601 VDDA.n600 3.4105
R905 VDDA.n603 VDDA.n602 3.4105
R906 VDDA.n605 VDDA.n604 3.4105
R907 VDDA.n606 VDDA.n548 3.4105
R908 VDDA.n610 VDDA.n609 3.4105
R909 VDDA.n609 VDDA.n608 3.4105
R910 VDDA.n536 VDDA.n535 3.4105
R911 VDDA.n775 VDDA.n774 3.4105
R912 VDDA.n101 VDDA.n100 3.4105
R913 VDDA.n890 VDDA.n17 3.4105
R914 VDDA.n890 VDDA.n16 3.4105
R915 VDDA.n890 VDDA.n18 3.4105
R916 VDDA.n890 VDDA.n889 3.4105
R917 VDDA.n889 VDDA.n794 3.4105
R918 VDDA.n791 VDDA.n16 3.4105
R919 VDDA.n859 VDDA.n791 3.4105
R920 VDDA.n856 VDDA.n791 3.4105
R921 VDDA.n861 VDDA.n791 3.4105
R922 VDDA.n855 VDDA.n791 3.4105
R923 VDDA.n863 VDDA.n791 3.4105
R924 VDDA.n854 VDDA.n791 3.4105
R925 VDDA.n865 VDDA.n791 3.4105
R926 VDDA.n853 VDDA.n791 3.4105
R927 VDDA.n867 VDDA.n791 3.4105
R928 VDDA.n852 VDDA.n791 3.4105
R929 VDDA.n869 VDDA.n791 3.4105
R930 VDDA.n851 VDDA.n791 3.4105
R931 VDDA.n871 VDDA.n791 3.4105
R932 VDDA.n850 VDDA.n791 3.4105
R933 VDDA.n873 VDDA.n791 3.4105
R934 VDDA.n849 VDDA.n791 3.4105
R935 VDDA.n875 VDDA.n791 3.4105
R936 VDDA.n848 VDDA.n791 3.4105
R937 VDDA.n877 VDDA.n791 3.4105
R938 VDDA.n847 VDDA.n791 3.4105
R939 VDDA.n879 VDDA.n791 3.4105
R940 VDDA.n846 VDDA.n791 3.4105
R941 VDDA.n881 VDDA.n791 3.4105
R942 VDDA.n845 VDDA.n791 3.4105
R943 VDDA.n883 VDDA.n791 3.4105
R944 VDDA.n844 VDDA.n791 3.4105
R945 VDDA.n885 VDDA.n791 3.4105
R946 VDDA.n843 VDDA.n791 3.4105
R947 VDDA.n887 VDDA.n791 3.4105
R948 VDDA.n842 VDDA.n791 3.4105
R949 VDDA.n791 VDDA.n18 3.4105
R950 VDDA.n889 VDDA.n791 3.4105
R951 VDDA.n797 VDDA.n16 3.4105
R952 VDDA.n859 VDDA.n797 3.4105
R953 VDDA.n856 VDDA.n797 3.4105
R954 VDDA.n861 VDDA.n797 3.4105
R955 VDDA.n855 VDDA.n797 3.4105
R956 VDDA.n863 VDDA.n797 3.4105
R957 VDDA.n854 VDDA.n797 3.4105
R958 VDDA.n865 VDDA.n797 3.4105
R959 VDDA.n853 VDDA.n797 3.4105
R960 VDDA.n867 VDDA.n797 3.4105
R961 VDDA.n852 VDDA.n797 3.4105
R962 VDDA.n869 VDDA.n797 3.4105
R963 VDDA.n851 VDDA.n797 3.4105
R964 VDDA.n871 VDDA.n797 3.4105
R965 VDDA.n850 VDDA.n797 3.4105
R966 VDDA.n873 VDDA.n797 3.4105
R967 VDDA.n849 VDDA.n797 3.4105
R968 VDDA.n875 VDDA.n797 3.4105
R969 VDDA.n848 VDDA.n797 3.4105
R970 VDDA.n877 VDDA.n797 3.4105
R971 VDDA.n847 VDDA.n797 3.4105
R972 VDDA.n879 VDDA.n797 3.4105
R973 VDDA.n846 VDDA.n797 3.4105
R974 VDDA.n881 VDDA.n797 3.4105
R975 VDDA.n845 VDDA.n797 3.4105
R976 VDDA.n883 VDDA.n797 3.4105
R977 VDDA.n844 VDDA.n797 3.4105
R978 VDDA.n885 VDDA.n797 3.4105
R979 VDDA.n843 VDDA.n797 3.4105
R980 VDDA.n887 VDDA.n797 3.4105
R981 VDDA.n842 VDDA.n797 3.4105
R982 VDDA.n797 VDDA.n18 3.4105
R983 VDDA.n889 VDDA.n797 3.4105
R984 VDDA.n790 VDDA.n16 3.4105
R985 VDDA.n859 VDDA.n790 3.4105
R986 VDDA.n856 VDDA.n790 3.4105
R987 VDDA.n861 VDDA.n790 3.4105
R988 VDDA.n855 VDDA.n790 3.4105
R989 VDDA.n863 VDDA.n790 3.4105
R990 VDDA.n854 VDDA.n790 3.4105
R991 VDDA.n865 VDDA.n790 3.4105
R992 VDDA.n853 VDDA.n790 3.4105
R993 VDDA.n867 VDDA.n790 3.4105
R994 VDDA.n852 VDDA.n790 3.4105
R995 VDDA.n869 VDDA.n790 3.4105
R996 VDDA.n851 VDDA.n790 3.4105
R997 VDDA.n871 VDDA.n790 3.4105
R998 VDDA.n850 VDDA.n790 3.4105
R999 VDDA.n873 VDDA.n790 3.4105
R1000 VDDA.n849 VDDA.n790 3.4105
R1001 VDDA.n875 VDDA.n790 3.4105
R1002 VDDA.n848 VDDA.n790 3.4105
R1003 VDDA.n877 VDDA.n790 3.4105
R1004 VDDA.n847 VDDA.n790 3.4105
R1005 VDDA.n879 VDDA.n790 3.4105
R1006 VDDA.n846 VDDA.n790 3.4105
R1007 VDDA.n881 VDDA.n790 3.4105
R1008 VDDA.n845 VDDA.n790 3.4105
R1009 VDDA.n883 VDDA.n790 3.4105
R1010 VDDA.n844 VDDA.n790 3.4105
R1011 VDDA.n885 VDDA.n790 3.4105
R1012 VDDA.n843 VDDA.n790 3.4105
R1013 VDDA.n887 VDDA.n790 3.4105
R1014 VDDA.n842 VDDA.n790 3.4105
R1015 VDDA.n790 VDDA.n18 3.4105
R1016 VDDA.n889 VDDA.n790 3.4105
R1017 VDDA.n800 VDDA.n16 3.4105
R1018 VDDA.n859 VDDA.n800 3.4105
R1019 VDDA.n856 VDDA.n800 3.4105
R1020 VDDA.n861 VDDA.n800 3.4105
R1021 VDDA.n855 VDDA.n800 3.4105
R1022 VDDA.n863 VDDA.n800 3.4105
R1023 VDDA.n854 VDDA.n800 3.4105
R1024 VDDA.n865 VDDA.n800 3.4105
R1025 VDDA.n853 VDDA.n800 3.4105
R1026 VDDA.n867 VDDA.n800 3.4105
R1027 VDDA.n852 VDDA.n800 3.4105
R1028 VDDA.n869 VDDA.n800 3.4105
R1029 VDDA.n851 VDDA.n800 3.4105
R1030 VDDA.n871 VDDA.n800 3.4105
R1031 VDDA.n850 VDDA.n800 3.4105
R1032 VDDA.n873 VDDA.n800 3.4105
R1033 VDDA.n849 VDDA.n800 3.4105
R1034 VDDA.n875 VDDA.n800 3.4105
R1035 VDDA.n848 VDDA.n800 3.4105
R1036 VDDA.n877 VDDA.n800 3.4105
R1037 VDDA.n847 VDDA.n800 3.4105
R1038 VDDA.n879 VDDA.n800 3.4105
R1039 VDDA.n846 VDDA.n800 3.4105
R1040 VDDA.n881 VDDA.n800 3.4105
R1041 VDDA.n845 VDDA.n800 3.4105
R1042 VDDA.n883 VDDA.n800 3.4105
R1043 VDDA.n844 VDDA.n800 3.4105
R1044 VDDA.n885 VDDA.n800 3.4105
R1045 VDDA.n843 VDDA.n800 3.4105
R1046 VDDA.n887 VDDA.n800 3.4105
R1047 VDDA.n842 VDDA.n800 3.4105
R1048 VDDA.n800 VDDA.n18 3.4105
R1049 VDDA.n889 VDDA.n800 3.4105
R1050 VDDA.n789 VDDA.n16 3.4105
R1051 VDDA.n859 VDDA.n789 3.4105
R1052 VDDA.n856 VDDA.n789 3.4105
R1053 VDDA.n861 VDDA.n789 3.4105
R1054 VDDA.n855 VDDA.n789 3.4105
R1055 VDDA.n863 VDDA.n789 3.4105
R1056 VDDA.n854 VDDA.n789 3.4105
R1057 VDDA.n865 VDDA.n789 3.4105
R1058 VDDA.n853 VDDA.n789 3.4105
R1059 VDDA.n867 VDDA.n789 3.4105
R1060 VDDA.n852 VDDA.n789 3.4105
R1061 VDDA.n869 VDDA.n789 3.4105
R1062 VDDA.n851 VDDA.n789 3.4105
R1063 VDDA.n871 VDDA.n789 3.4105
R1064 VDDA.n850 VDDA.n789 3.4105
R1065 VDDA.n873 VDDA.n789 3.4105
R1066 VDDA.n849 VDDA.n789 3.4105
R1067 VDDA.n875 VDDA.n789 3.4105
R1068 VDDA.n848 VDDA.n789 3.4105
R1069 VDDA.n877 VDDA.n789 3.4105
R1070 VDDA.n847 VDDA.n789 3.4105
R1071 VDDA.n879 VDDA.n789 3.4105
R1072 VDDA.n846 VDDA.n789 3.4105
R1073 VDDA.n881 VDDA.n789 3.4105
R1074 VDDA.n845 VDDA.n789 3.4105
R1075 VDDA.n883 VDDA.n789 3.4105
R1076 VDDA.n844 VDDA.n789 3.4105
R1077 VDDA.n885 VDDA.n789 3.4105
R1078 VDDA.n843 VDDA.n789 3.4105
R1079 VDDA.n887 VDDA.n789 3.4105
R1080 VDDA.n842 VDDA.n789 3.4105
R1081 VDDA.n789 VDDA.n18 3.4105
R1082 VDDA.n889 VDDA.n789 3.4105
R1083 VDDA.n803 VDDA.n16 3.4105
R1084 VDDA.n859 VDDA.n803 3.4105
R1085 VDDA.n856 VDDA.n803 3.4105
R1086 VDDA.n861 VDDA.n803 3.4105
R1087 VDDA.n855 VDDA.n803 3.4105
R1088 VDDA.n863 VDDA.n803 3.4105
R1089 VDDA.n854 VDDA.n803 3.4105
R1090 VDDA.n865 VDDA.n803 3.4105
R1091 VDDA.n853 VDDA.n803 3.4105
R1092 VDDA.n867 VDDA.n803 3.4105
R1093 VDDA.n852 VDDA.n803 3.4105
R1094 VDDA.n869 VDDA.n803 3.4105
R1095 VDDA.n851 VDDA.n803 3.4105
R1096 VDDA.n871 VDDA.n803 3.4105
R1097 VDDA.n850 VDDA.n803 3.4105
R1098 VDDA.n873 VDDA.n803 3.4105
R1099 VDDA.n849 VDDA.n803 3.4105
R1100 VDDA.n875 VDDA.n803 3.4105
R1101 VDDA.n848 VDDA.n803 3.4105
R1102 VDDA.n877 VDDA.n803 3.4105
R1103 VDDA.n847 VDDA.n803 3.4105
R1104 VDDA.n879 VDDA.n803 3.4105
R1105 VDDA.n846 VDDA.n803 3.4105
R1106 VDDA.n881 VDDA.n803 3.4105
R1107 VDDA.n845 VDDA.n803 3.4105
R1108 VDDA.n883 VDDA.n803 3.4105
R1109 VDDA.n844 VDDA.n803 3.4105
R1110 VDDA.n885 VDDA.n803 3.4105
R1111 VDDA.n843 VDDA.n803 3.4105
R1112 VDDA.n887 VDDA.n803 3.4105
R1113 VDDA.n842 VDDA.n803 3.4105
R1114 VDDA.n803 VDDA.n18 3.4105
R1115 VDDA.n889 VDDA.n803 3.4105
R1116 VDDA.n788 VDDA.n16 3.4105
R1117 VDDA.n859 VDDA.n788 3.4105
R1118 VDDA.n856 VDDA.n788 3.4105
R1119 VDDA.n861 VDDA.n788 3.4105
R1120 VDDA.n855 VDDA.n788 3.4105
R1121 VDDA.n863 VDDA.n788 3.4105
R1122 VDDA.n854 VDDA.n788 3.4105
R1123 VDDA.n865 VDDA.n788 3.4105
R1124 VDDA.n853 VDDA.n788 3.4105
R1125 VDDA.n867 VDDA.n788 3.4105
R1126 VDDA.n852 VDDA.n788 3.4105
R1127 VDDA.n869 VDDA.n788 3.4105
R1128 VDDA.n851 VDDA.n788 3.4105
R1129 VDDA.n871 VDDA.n788 3.4105
R1130 VDDA.n850 VDDA.n788 3.4105
R1131 VDDA.n873 VDDA.n788 3.4105
R1132 VDDA.n849 VDDA.n788 3.4105
R1133 VDDA.n875 VDDA.n788 3.4105
R1134 VDDA.n848 VDDA.n788 3.4105
R1135 VDDA.n877 VDDA.n788 3.4105
R1136 VDDA.n847 VDDA.n788 3.4105
R1137 VDDA.n879 VDDA.n788 3.4105
R1138 VDDA.n846 VDDA.n788 3.4105
R1139 VDDA.n881 VDDA.n788 3.4105
R1140 VDDA.n845 VDDA.n788 3.4105
R1141 VDDA.n883 VDDA.n788 3.4105
R1142 VDDA.n844 VDDA.n788 3.4105
R1143 VDDA.n885 VDDA.n788 3.4105
R1144 VDDA.n843 VDDA.n788 3.4105
R1145 VDDA.n887 VDDA.n788 3.4105
R1146 VDDA.n842 VDDA.n788 3.4105
R1147 VDDA.n788 VDDA.n18 3.4105
R1148 VDDA.n889 VDDA.n788 3.4105
R1149 VDDA.n806 VDDA.n16 3.4105
R1150 VDDA.n859 VDDA.n806 3.4105
R1151 VDDA.n856 VDDA.n806 3.4105
R1152 VDDA.n861 VDDA.n806 3.4105
R1153 VDDA.n855 VDDA.n806 3.4105
R1154 VDDA.n863 VDDA.n806 3.4105
R1155 VDDA.n854 VDDA.n806 3.4105
R1156 VDDA.n865 VDDA.n806 3.4105
R1157 VDDA.n853 VDDA.n806 3.4105
R1158 VDDA.n867 VDDA.n806 3.4105
R1159 VDDA.n852 VDDA.n806 3.4105
R1160 VDDA.n869 VDDA.n806 3.4105
R1161 VDDA.n851 VDDA.n806 3.4105
R1162 VDDA.n871 VDDA.n806 3.4105
R1163 VDDA.n850 VDDA.n806 3.4105
R1164 VDDA.n873 VDDA.n806 3.4105
R1165 VDDA.n849 VDDA.n806 3.4105
R1166 VDDA.n875 VDDA.n806 3.4105
R1167 VDDA.n848 VDDA.n806 3.4105
R1168 VDDA.n877 VDDA.n806 3.4105
R1169 VDDA.n847 VDDA.n806 3.4105
R1170 VDDA.n879 VDDA.n806 3.4105
R1171 VDDA.n846 VDDA.n806 3.4105
R1172 VDDA.n881 VDDA.n806 3.4105
R1173 VDDA.n845 VDDA.n806 3.4105
R1174 VDDA.n883 VDDA.n806 3.4105
R1175 VDDA.n844 VDDA.n806 3.4105
R1176 VDDA.n885 VDDA.n806 3.4105
R1177 VDDA.n843 VDDA.n806 3.4105
R1178 VDDA.n887 VDDA.n806 3.4105
R1179 VDDA.n842 VDDA.n806 3.4105
R1180 VDDA.n806 VDDA.n18 3.4105
R1181 VDDA.n889 VDDA.n806 3.4105
R1182 VDDA.n787 VDDA.n16 3.4105
R1183 VDDA.n859 VDDA.n787 3.4105
R1184 VDDA.n856 VDDA.n787 3.4105
R1185 VDDA.n861 VDDA.n787 3.4105
R1186 VDDA.n855 VDDA.n787 3.4105
R1187 VDDA.n863 VDDA.n787 3.4105
R1188 VDDA.n854 VDDA.n787 3.4105
R1189 VDDA.n865 VDDA.n787 3.4105
R1190 VDDA.n853 VDDA.n787 3.4105
R1191 VDDA.n867 VDDA.n787 3.4105
R1192 VDDA.n852 VDDA.n787 3.4105
R1193 VDDA.n869 VDDA.n787 3.4105
R1194 VDDA.n851 VDDA.n787 3.4105
R1195 VDDA.n871 VDDA.n787 3.4105
R1196 VDDA.n850 VDDA.n787 3.4105
R1197 VDDA.n873 VDDA.n787 3.4105
R1198 VDDA.n849 VDDA.n787 3.4105
R1199 VDDA.n875 VDDA.n787 3.4105
R1200 VDDA.n848 VDDA.n787 3.4105
R1201 VDDA.n877 VDDA.n787 3.4105
R1202 VDDA.n847 VDDA.n787 3.4105
R1203 VDDA.n879 VDDA.n787 3.4105
R1204 VDDA.n846 VDDA.n787 3.4105
R1205 VDDA.n881 VDDA.n787 3.4105
R1206 VDDA.n845 VDDA.n787 3.4105
R1207 VDDA.n883 VDDA.n787 3.4105
R1208 VDDA.n844 VDDA.n787 3.4105
R1209 VDDA.n885 VDDA.n787 3.4105
R1210 VDDA.n843 VDDA.n787 3.4105
R1211 VDDA.n887 VDDA.n787 3.4105
R1212 VDDA.n842 VDDA.n787 3.4105
R1213 VDDA.n787 VDDA.n18 3.4105
R1214 VDDA.n889 VDDA.n787 3.4105
R1215 VDDA.n809 VDDA.n16 3.4105
R1216 VDDA.n859 VDDA.n809 3.4105
R1217 VDDA.n856 VDDA.n809 3.4105
R1218 VDDA.n861 VDDA.n809 3.4105
R1219 VDDA.n855 VDDA.n809 3.4105
R1220 VDDA.n863 VDDA.n809 3.4105
R1221 VDDA.n854 VDDA.n809 3.4105
R1222 VDDA.n865 VDDA.n809 3.4105
R1223 VDDA.n853 VDDA.n809 3.4105
R1224 VDDA.n867 VDDA.n809 3.4105
R1225 VDDA.n852 VDDA.n809 3.4105
R1226 VDDA.n869 VDDA.n809 3.4105
R1227 VDDA.n851 VDDA.n809 3.4105
R1228 VDDA.n871 VDDA.n809 3.4105
R1229 VDDA.n850 VDDA.n809 3.4105
R1230 VDDA.n873 VDDA.n809 3.4105
R1231 VDDA.n849 VDDA.n809 3.4105
R1232 VDDA.n875 VDDA.n809 3.4105
R1233 VDDA.n848 VDDA.n809 3.4105
R1234 VDDA.n877 VDDA.n809 3.4105
R1235 VDDA.n847 VDDA.n809 3.4105
R1236 VDDA.n879 VDDA.n809 3.4105
R1237 VDDA.n846 VDDA.n809 3.4105
R1238 VDDA.n881 VDDA.n809 3.4105
R1239 VDDA.n845 VDDA.n809 3.4105
R1240 VDDA.n883 VDDA.n809 3.4105
R1241 VDDA.n844 VDDA.n809 3.4105
R1242 VDDA.n885 VDDA.n809 3.4105
R1243 VDDA.n843 VDDA.n809 3.4105
R1244 VDDA.n887 VDDA.n809 3.4105
R1245 VDDA.n842 VDDA.n809 3.4105
R1246 VDDA.n809 VDDA.n18 3.4105
R1247 VDDA.n889 VDDA.n809 3.4105
R1248 VDDA.n786 VDDA.n16 3.4105
R1249 VDDA.n859 VDDA.n786 3.4105
R1250 VDDA.n856 VDDA.n786 3.4105
R1251 VDDA.n861 VDDA.n786 3.4105
R1252 VDDA.n855 VDDA.n786 3.4105
R1253 VDDA.n863 VDDA.n786 3.4105
R1254 VDDA.n854 VDDA.n786 3.4105
R1255 VDDA.n865 VDDA.n786 3.4105
R1256 VDDA.n853 VDDA.n786 3.4105
R1257 VDDA.n867 VDDA.n786 3.4105
R1258 VDDA.n852 VDDA.n786 3.4105
R1259 VDDA.n869 VDDA.n786 3.4105
R1260 VDDA.n851 VDDA.n786 3.4105
R1261 VDDA.n871 VDDA.n786 3.4105
R1262 VDDA.n850 VDDA.n786 3.4105
R1263 VDDA.n873 VDDA.n786 3.4105
R1264 VDDA.n849 VDDA.n786 3.4105
R1265 VDDA.n875 VDDA.n786 3.4105
R1266 VDDA.n848 VDDA.n786 3.4105
R1267 VDDA.n877 VDDA.n786 3.4105
R1268 VDDA.n847 VDDA.n786 3.4105
R1269 VDDA.n879 VDDA.n786 3.4105
R1270 VDDA.n846 VDDA.n786 3.4105
R1271 VDDA.n881 VDDA.n786 3.4105
R1272 VDDA.n845 VDDA.n786 3.4105
R1273 VDDA.n883 VDDA.n786 3.4105
R1274 VDDA.n844 VDDA.n786 3.4105
R1275 VDDA.n885 VDDA.n786 3.4105
R1276 VDDA.n843 VDDA.n786 3.4105
R1277 VDDA.n887 VDDA.n786 3.4105
R1278 VDDA.n842 VDDA.n786 3.4105
R1279 VDDA.n786 VDDA.n18 3.4105
R1280 VDDA.n889 VDDA.n786 3.4105
R1281 VDDA.n812 VDDA.n16 3.4105
R1282 VDDA.n859 VDDA.n812 3.4105
R1283 VDDA.n856 VDDA.n812 3.4105
R1284 VDDA.n861 VDDA.n812 3.4105
R1285 VDDA.n855 VDDA.n812 3.4105
R1286 VDDA.n863 VDDA.n812 3.4105
R1287 VDDA.n854 VDDA.n812 3.4105
R1288 VDDA.n865 VDDA.n812 3.4105
R1289 VDDA.n853 VDDA.n812 3.4105
R1290 VDDA.n867 VDDA.n812 3.4105
R1291 VDDA.n852 VDDA.n812 3.4105
R1292 VDDA.n869 VDDA.n812 3.4105
R1293 VDDA.n851 VDDA.n812 3.4105
R1294 VDDA.n871 VDDA.n812 3.4105
R1295 VDDA.n850 VDDA.n812 3.4105
R1296 VDDA.n873 VDDA.n812 3.4105
R1297 VDDA.n849 VDDA.n812 3.4105
R1298 VDDA.n875 VDDA.n812 3.4105
R1299 VDDA.n848 VDDA.n812 3.4105
R1300 VDDA.n877 VDDA.n812 3.4105
R1301 VDDA.n847 VDDA.n812 3.4105
R1302 VDDA.n879 VDDA.n812 3.4105
R1303 VDDA.n846 VDDA.n812 3.4105
R1304 VDDA.n881 VDDA.n812 3.4105
R1305 VDDA.n845 VDDA.n812 3.4105
R1306 VDDA.n883 VDDA.n812 3.4105
R1307 VDDA.n844 VDDA.n812 3.4105
R1308 VDDA.n885 VDDA.n812 3.4105
R1309 VDDA.n843 VDDA.n812 3.4105
R1310 VDDA.n887 VDDA.n812 3.4105
R1311 VDDA.n842 VDDA.n812 3.4105
R1312 VDDA.n812 VDDA.n18 3.4105
R1313 VDDA.n889 VDDA.n812 3.4105
R1314 VDDA.n785 VDDA.n16 3.4105
R1315 VDDA.n859 VDDA.n785 3.4105
R1316 VDDA.n856 VDDA.n785 3.4105
R1317 VDDA.n861 VDDA.n785 3.4105
R1318 VDDA.n855 VDDA.n785 3.4105
R1319 VDDA.n863 VDDA.n785 3.4105
R1320 VDDA.n854 VDDA.n785 3.4105
R1321 VDDA.n865 VDDA.n785 3.4105
R1322 VDDA.n853 VDDA.n785 3.4105
R1323 VDDA.n867 VDDA.n785 3.4105
R1324 VDDA.n852 VDDA.n785 3.4105
R1325 VDDA.n869 VDDA.n785 3.4105
R1326 VDDA.n851 VDDA.n785 3.4105
R1327 VDDA.n871 VDDA.n785 3.4105
R1328 VDDA.n850 VDDA.n785 3.4105
R1329 VDDA.n873 VDDA.n785 3.4105
R1330 VDDA.n849 VDDA.n785 3.4105
R1331 VDDA.n875 VDDA.n785 3.4105
R1332 VDDA.n848 VDDA.n785 3.4105
R1333 VDDA.n877 VDDA.n785 3.4105
R1334 VDDA.n847 VDDA.n785 3.4105
R1335 VDDA.n879 VDDA.n785 3.4105
R1336 VDDA.n846 VDDA.n785 3.4105
R1337 VDDA.n881 VDDA.n785 3.4105
R1338 VDDA.n845 VDDA.n785 3.4105
R1339 VDDA.n883 VDDA.n785 3.4105
R1340 VDDA.n844 VDDA.n785 3.4105
R1341 VDDA.n885 VDDA.n785 3.4105
R1342 VDDA.n843 VDDA.n785 3.4105
R1343 VDDA.n887 VDDA.n785 3.4105
R1344 VDDA.n842 VDDA.n785 3.4105
R1345 VDDA.n785 VDDA.n18 3.4105
R1346 VDDA.n889 VDDA.n785 3.4105
R1347 VDDA.n815 VDDA.n16 3.4105
R1348 VDDA.n859 VDDA.n815 3.4105
R1349 VDDA.n856 VDDA.n815 3.4105
R1350 VDDA.n861 VDDA.n815 3.4105
R1351 VDDA.n855 VDDA.n815 3.4105
R1352 VDDA.n863 VDDA.n815 3.4105
R1353 VDDA.n854 VDDA.n815 3.4105
R1354 VDDA.n865 VDDA.n815 3.4105
R1355 VDDA.n853 VDDA.n815 3.4105
R1356 VDDA.n867 VDDA.n815 3.4105
R1357 VDDA.n852 VDDA.n815 3.4105
R1358 VDDA.n869 VDDA.n815 3.4105
R1359 VDDA.n851 VDDA.n815 3.4105
R1360 VDDA.n871 VDDA.n815 3.4105
R1361 VDDA.n850 VDDA.n815 3.4105
R1362 VDDA.n873 VDDA.n815 3.4105
R1363 VDDA.n849 VDDA.n815 3.4105
R1364 VDDA.n875 VDDA.n815 3.4105
R1365 VDDA.n848 VDDA.n815 3.4105
R1366 VDDA.n877 VDDA.n815 3.4105
R1367 VDDA.n847 VDDA.n815 3.4105
R1368 VDDA.n879 VDDA.n815 3.4105
R1369 VDDA.n846 VDDA.n815 3.4105
R1370 VDDA.n881 VDDA.n815 3.4105
R1371 VDDA.n845 VDDA.n815 3.4105
R1372 VDDA.n883 VDDA.n815 3.4105
R1373 VDDA.n844 VDDA.n815 3.4105
R1374 VDDA.n885 VDDA.n815 3.4105
R1375 VDDA.n843 VDDA.n815 3.4105
R1376 VDDA.n887 VDDA.n815 3.4105
R1377 VDDA.n842 VDDA.n815 3.4105
R1378 VDDA.n815 VDDA.n18 3.4105
R1379 VDDA.n889 VDDA.n815 3.4105
R1380 VDDA.n784 VDDA.n16 3.4105
R1381 VDDA.n859 VDDA.n784 3.4105
R1382 VDDA.n856 VDDA.n784 3.4105
R1383 VDDA.n861 VDDA.n784 3.4105
R1384 VDDA.n855 VDDA.n784 3.4105
R1385 VDDA.n863 VDDA.n784 3.4105
R1386 VDDA.n854 VDDA.n784 3.4105
R1387 VDDA.n865 VDDA.n784 3.4105
R1388 VDDA.n853 VDDA.n784 3.4105
R1389 VDDA.n867 VDDA.n784 3.4105
R1390 VDDA.n852 VDDA.n784 3.4105
R1391 VDDA.n869 VDDA.n784 3.4105
R1392 VDDA.n851 VDDA.n784 3.4105
R1393 VDDA.n871 VDDA.n784 3.4105
R1394 VDDA.n850 VDDA.n784 3.4105
R1395 VDDA.n873 VDDA.n784 3.4105
R1396 VDDA.n849 VDDA.n784 3.4105
R1397 VDDA.n875 VDDA.n784 3.4105
R1398 VDDA.n848 VDDA.n784 3.4105
R1399 VDDA.n877 VDDA.n784 3.4105
R1400 VDDA.n847 VDDA.n784 3.4105
R1401 VDDA.n879 VDDA.n784 3.4105
R1402 VDDA.n846 VDDA.n784 3.4105
R1403 VDDA.n881 VDDA.n784 3.4105
R1404 VDDA.n845 VDDA.n784 3.4105
R1405 VDDA.n883 VDDA.n784 3.4105
R1406 VDDA.n844 VDDA.n784 3.4105
R1407 VDDA.n885 VDDA.n784 3.4105
R1408 VDDA.n843 VDDA.n784 3.4105
R1409 VDDA.n887 VDDA.n784 3.4105
R1410 VDDA.n842 VDDA.n784 3.4105
R1411 VDDA.n784 VDDA.n18 3.4105
R1412 VDDA.n889 VDDA.n784 3.4105
R1413 VDDA.n818 VDDA.n16 3.4105
R1414 VDDA.n859 VDDA.n818 3.4105
R1415 VDDA.n856 VDDA.n818 3.4105
R1416 VDDA.n861 VDDA.n818 3.4105
R1417 VDDA.n855 VDDA.n818 3.4105
R1418 VDDA.n863 VDDA.n818 3.4105
R1419 VDDA.n854 VDDA.n818 3.4105
R1420 VDDA.n865 VDDA.n818 3.4105
R1421 VDDA.n853 VDDA.n818 3.4105
R1422 VDDA.n867 VDDA.n818 3.4105
R1423 VDDA.n852 VDDA.n818 3.4105
R1424 VDDA.n869 VDDA.n818 3.4105
R1425 VDDA.n851 VDDA.n818 3.4105
R1426 VDDA.n871 VDDA.n818 3.4105
R1427 VDDA.n850 VDDA.n818 3.4105
R1428 VDDA.n873 VDDA.n818 3.4105
R1429 VDDA.n849 VDDA.n818 3.4105
R1430 VDDA.n875 VDDA.n818 3.4105
R1431 VDDA.n848 VDDA.n818 3.4105
R1432 VDDA.n877 VDDA.n818 3.4105
R1433 VDDA.n847 VDDA.n818 3.4105
R1434 VDDA.n879 VDDA.n818 3.4105
R1435 VDDA.n846 VDDA.n818 3.4105
R1436 VDDA.n881 VDDA.n818 3.4105
R1437 VDDA.n845 VDDA.n818 3.4105
R1438 VDDA.n883 VDDA.n818 3.4105
R1439 VDDA.n844 VDDA.n818 3.4105
R1440 VDDA.n885 VDDA.n818 3.4105
R1441 VDDA.n843 VDDA.n818 3.4105
R1442 VDDA.n887 VDDA.n818 3.4105
R1443 VDDA.n842 VDDA.n818 3.4105
R1444 VDDA.n818 VDDA.n18 3.4105
R1445 VDDA.n889 VDDA.n818 3.4105
R1446 VDDA.n783 VDDA.n16 3.4105
R1447 VDDA.n859 VDDA.n783 3.4105
R1448 VDDA.n856 VDDA.n783 3.4105
R1449 VDDA.n861 VDDA.n783 3.4105
R1450 VDDA.n855 VDDA.n783 3.4105
R1451 VDDA.n863 VDDA.n783 3.4105
R1452 VDDA.n854 VDDA.n783 3.4105
R1453 VDDA.n865 VDDA.n783 3.4105
R1454 VDDA.n853 VDDA.n783 3.4105
R1455 VDDA.n867 VDDA.n783 3.4105
R1456 VDDA.n852 VDDA.n783 3.4105
R1457 VDDA.n869 VDDA.n783 3.4105
R1458 VDDA.n851 VDDA.n783 3.4105
R1459 VDDA.n871 VDDA.n783 3.4105
R1460 VDDA.n850 VDDA.n783 3.4105
R1461 VDDA.n873 VDDA.n783 3.4105
R1462 VDDA.n849 VDDA.n783 3.4105
R1463 VDDA.n875 VDDA.n783 3.4105
R1464 VDDA.n848 VDDA.n783 3.4105
R1465 VDDA.n877 VDDA.n783 3.4105
R1466 VDDA.n847 VDDA.n783 3.4105
R1467 VDDA.n879 VDDA.n783 3.4105
R1468 VDDA.n846 VDDA.n783 3.4105
R1469 VDDA.n881 VDDA.n783 3.4105
R1470 VDDA.n845 VDDA.n783 3.4105
R1471 VDDA.n883 VDDA.n783 3.4105
R1472 VDDA.n844 VDDA.n783 3.4105
R1473 VDDA.n885 VDDA.n783 3.4105
R1474 VDDA.n843 VDDA.n783 3.4105
R1475 VDDA.n887 VDDA.n783 3.4105
R1476 VDDA.n842 VDDA.n783 3.4105
R1477 VDDA.n783 VDDA.n18 3.4105
R1478 VDDA.n889 VDDA.n783 3.4105
R1479 VDDA.n821 VDDA.n16 3.4105
R1480 VDDA.n859 VDDA.n821 3.4105
R1481 VDDA.n856 VDDA.n821 3.4105
R1482 VDDA.n861 VDDA.n821 3.4105
R1483 VDDA.n855 VDDA.n821 3.4105
R1484 VDDA.n863 VDDA.n821 3.4105
R1485 VDDA.n854 VDDA.n821 3.4105
R1486 VDDA.n865 VDDA.n821 3.4105
R1487 VDDA.n853 VDDA.n821 3.4105
R1488 VDDA.n867 VDDA.n821 3.4105
R1489 VDDA.n852 VDDA.n821 3.4105
R1490 VDDA.n869 VDDA.n821 3.4105
R1491 VDDA.n851 VDDA.n821 3.4105
R1492 VDDA.n871 VDDA.n821 3.4105
R1493 VDDA.n850 VDDA.n821 3.4105
R1494 VDDA.n873 VDDA.n821 3.4105
R1495 VDDA.n849 VDDA.n821 3.4105
R1496 VDDA.n875 VDDA.n821 3.4105
R1497 VDDA.n848 VDDA.n821 3.4105
R1498 VDDA.n877 VDDA.n821 3.4105
R1499 VDDA.n847 VDDA.n821 3.4105
R1500 VDDA.n879 VDDA.n821 3.4105
R1501 VDDA.n846 VDDA.n821 3.4105
R1502 VDDA.n881 VDDA.n821 3.4105
R1503 VDDA.n845 VDDA.n821 3.4105
R1504 VDDA.n883 VDDA.n821 3.4105
R1505 VDDA.n844 VDDA.n821 3.4105
R1506 VDDA.n885 VDDA.n821 3.4105
R1507 VDDA.n843 VDDA.n821 3.4105
R1508 VDDA.n887 VDDA.n821 3.4105
R1509 VDDA.n842 VDDA.n821 3.4105
R1510 VDDA.n821 VDDA.n18 3.4105
R1511 VDDA.n889 VDDA.n821 3.4105
R1512 VDDA.n782 VDDA.n16 3.4105
R1513 VDDA.n859 VDDA.n782 3.4105
R1514 VDDA.n856 VDDA.n782 3.4105
R1515 VDDA.n861 VDDA.n782 3.4105
R1516 VDDA.n855 VDDA.n782 3.4105
R1517 VDDA.n863 VDDA.n782 3.4105
R1518 VDDA.n854 VDDA.n782 3.4105
R1519 VDDA.n865 VDDA.n782 3.4105
R1520 VDDA.n853 VDDA.n782 3.4105
R1521 VDDA.n867 VDDA.n782 3.4105
R1522 VDDA.n852 VDDA.n782 3.4105
R1523 VDDA.n869 VDDA.n782 3.4105
R1524 VDDA.n851 VDDA.n782 3.4105
R1525 VDDA.n871 VDDA.n782 3.4105
R1526 VDDA.n850 VDDA.n782 3.4105
R1527 VDDA.n873 VDDA.n782 3.4105
R1528 VDDA.n849 VDDA.n782 3.4105
R1529 VDDA.n875 VDDA.n782 3.4105
R1530 VDDA.n848 VDDA.n782 3.4105
R1531 VDDA.n877 VDDA.n782 3.4105
R1532 VDDA.n847 VDDA.n782 3.4105
R1533 VDDA.n879 VDDA.n782 3.4105
R1534 VDDA.n846 VDDA.n782 3.4105
R1535 VDDA.n881 VDDA.n782 3.4105
R1536 VDDA.n845 VDDA.n782 3.4105
R1537 VDDA.n883 VDDA.n782 3.4105
R1538 VDDA.n844 VDDA.n782 3.4105
R1539 VDDA.n885 VDDA.n782 3.4105
R1540 VDDA.n843 VDDA.n782 3.4105
R1541 VDDA.n887 VDDA.n782 3.4105
R1542 VDDA.n842 VDDA.n782 3.4105
R1543 VDDA.n782 VDDA.n18 3.4105
R1544 VDDA.n889 VDDA.n782 3.4105
R1545 VDDA.n824 VDDA.n16 3.4105
R1546 VDDA.n859 VDDA.n824 3.4105
R1547 VDDA.n856 VDDA.n824 3.4105
R1548 VDDA.n861 VDDA.n824 3.4105
R1549 VDDA.n855 VDDA.n824 3.4105
R1550 VDDA.n863 VDDA.n824 3.4105
R1551 VDDA.n854 VDDA.n824 3.4105
R1552 VDDA.n865 VDDA.n824 3.4105
R1553 VDDA.n853 VDDA.n824 3.4105
R1554 VDDA.n867 VDDA.n824 3.4105
R1555 VDDA.n852 VDDA.n824 3.4105
R1556 VDDA.n869 VDDA.n824 3.4105
R1557 VDDA.n851 VDDA.n824 3.4105
R1558 VDDA.n871 VDDA.n824 3.4105
R1559 VDDA.n850 VDDA.n824 3.4105
R1560 VDDA.n873 VDDA.n824 3.4105
R1561 VDDA.n849 VDDA.n824 3.4105
R1562 VDDA.n875 VDDA.n824 3.4105
R1563 VDDA.n848 VDDA.n824 3.4105
R1564 VDDA.n877 VDDA.n824 3.4105
R1565 VDDA.n847 VDDA.n824 3.4105
R1566 VDDA.n879 VDDA.n824 3.4105
R1567 VDDA.n846 VDDA.n824 3.4105
R1568 VDDA.n881 VDDA.n824 3.4105
R1569 VDDA.n845 VDDA.n824 3.4105
R1570 VDDA.n883 VDDA.n824 3.4105
R1571 VDDA.n844 VDDA.n824 3.4105
R1572 VDDA.n885 VDDA.n824 3.4105
R1573 VDDA.n843 VDDA.n824 3.4105
R1574 VDDA.n887 VDDA.n824 3.4105
R1575 VDDA.n842 VDDA.n824 3.4105
R1576 VDDA.n824 VDDA.n18 3.4105
R1577 VDDA.n889 VDDA.n824 3.4105
R1578 VDDA.n781 VDDA.n16 3.4105
R1579 VDDA.n859 VDDA.n781 3.4105
R1580 VDDA.n856 VDDA.n781 3.4105
R1581 VDDA.n861 VDDA.n781 3.4105
R1582 VDDA.n855 VDDA.n781 3.4105
R1583 VDDA.n863 VDDA.n781 3.4105
R1584 VDDA.n854 VDDA.n781 3.4105
R1585 VDDA.n865 VDDA.n781 3.4105
R1586 VDDA.n853 VDDA.n781 3.4105
R1587 VDDA.n867 VDDA.n781 3.4105
R1588 VDDA.n852 VDDA.n781 3.4105
R1589 VDDA.n869 VDDA.n781 3.4105
R1590 VDDA.n851 VDDA.n781 3.4105
R1591 VDDA.n871 VDDA.n781 3.4105
R1592 VDDA.n850 VDDA.n781 3.4105
R1593 VDDA.n873 VDDA.n781 3.4105
R1594 VDDA.n849 VDDA.n781 3.4105
R1595 VDDA.n875 VDDA.n781 3.4105
R1596 VDDA.n848 VDDA.n781 3.4105
R1597 VDDA.n877 VDDA.n781 3.4105
R1598 VDDA.n847 VDDA.n781 3.4105
R1599 VDDA.n879 VDDA.n781 3.4105
R1600 VDDA.n846 VDDA.n781 3.4105
R1601 VDDA.n881 VDDA.n781 3.4105
R1602 VDDA.n845 VDDA.n781 3.4105
R1603 VDDA.n883 VDDA.n781 3.4105
R1604 VDDA.n844 VDDA.n781 3.4105
R1605 VDDA.n885 VDDA.n781 3.4105
R1606 VDDA.n843 VDDA.n781 3.4105
R1607 VDDA.n887 VDDA.n781 3.4105
R1608 VDDA.n842 VDDA.n781 3.4105
R1609 VDDA.n781 VDDA.n18 3.4105
R1610 VDDA.n889 VDDA.n781 3.4105
R1611 VDDA.n827 VDDA.n16 3.4105
R1612 VDDA.n859 VDDA.n827 3.4105
R1613 VDDA.n856 VDDA.n827 3.4105
R1614 VDDA.n861 VDDA.n827 3.4105
R1615 VDDA.n855 VDDA.n827 3.4105
R1616 VDDA.n863 VDDA.n827 3.4105
R1617 VDDA.n854 VDDA.n827 3.4105
R1618 VDDA.n865 VDDA.n827 3.4105
R1619 VDDA.n853 VDDA.n827 3.4105
R1620 VDDA.n867 VDDA.n827 3.4105
R1621 VDDA.n852 VDDA.n827 3.4105
R1622 VDDA.n869 VDDA.n827 3.4105
R1623 VDDA.n851 VDDA.n827 3.4105
R1624 VDDA.n871 VDDA.n827 3.4105
R1625 VDDA.n850 VDDA.n827 3.4105
R1626 VDDA.n873 VDDA.n827 3.4105
R1627 VDDA.n849 VDDA.n827 3.4105
R1628 VDDA.n875 VDDA.n827 3.4105
R1629 VDDA.n848 VDDA.n827 3.4105
R1630 VDDA.n877 VDDA.n827 3.4105
R1631 VDDA.n847 VDDA.n827 3.4105
R1632 VDDA.n879 VDDA.n827 3.4105
R1633 VDDA.n846 VDDA.n827 3.4105
R1634 VDDA.n881 VDDA.n827 3.4105
R1635 VDDA.n845 VDDA.n827 3.4105
R1636 VDDA.n883 VDDA.n827 3.4105
R1637 VDDA.n844 VDDA.n827 3.4105
R1638 VDDA.n885 VDDA.n827 3.4105
R1639 VDDA.n843 VDDA.n827 3.4105
R1640 VDDA.n887 VDDA.n827 3.4105
R1641 VDDA.n842 VDDA.n827 3.4105
R1642 VDDA.n827 VDDA.n18 3.4105
R1643 VDDA.n889 VDDA.n827 3.4105
R1644 VDDA.n780 VDDA.n16 3.4105
R1645 VDDA.n859 VDDA.n780 3.4105
R1646 VDDA.n856 VDDA.n780 3.4105
R1647 VDDA.n861 VDDA.n780 3.4105
R1648 VDDA.n855 VDDA.n780 3.4105
R1649 VDDA.n863 VDDA.n780 3.4105
R1650 VDDA.n854 VDDA.n780 3.4105
R1651 VDDA.n865 VDDA.n780 3.4105
R1652 VDDA.n853 VDDA.n780 3.4105
R1653 VDDA.n867 VDDA.n780 3.4105
R1654 VDDA.n852 VDDA.n780 3.4105
R1655 VDDA.n869 VDDA.n780 3.4105
R1656 VDDA.n851 VDDA.n780 3.4105
R1657 VDDA.n871 VDDA.n780 3.4105
R1658 VDDA.n850 VDDA.n780 3.4105
R1659 VDDA.n873 VDDA.n780 3.4105
R1660 VDDA.n849 VDDA.n780 3.4105
R1661 VDDA.n875 VDDA.n780 3.4105
R1662 VDDA.n848 VDDA.n780 3.4105
R1663 VDDA.n877 VDDA.n780 3.4105
R1664 VDDA.n847 VDDA.n780 3.4105
R1665 VDDA.n879 VDDA.n780 3.4105
R1666 VDDA.n846 VDDA.n780 3.4105
R1667 VDDA.n881 VDDA.n780 3.4105
R1668 VDDA.n845 VDDA.n780 3.4105
R1669 VDDA.n883 VDDA.n780 3.4105
R1670 VDDA.n844 VDDA.n780 3.4105
R1671 VDDA.n885 VDDA.n780 3.4105
R1672 VDDA.n843 VDDA.n780 3.4105
R1673 VDDA.n887 VDDA.n780 3.4105
R1674 VDDA.n842 VDDA.n780 3.4105
R1675 VDDA.n780 VDDA.n18 3.4105
R1676 VDDA.n889 VDDA.n780 3.4105
R1677 VDDA.n830 VDDA.n16 3.4105
R1678 VDDA.n859 VDDA.n830 3.4105
R1679 VDDA.n856 VDDA.n830 3.4105
R1680 VDDA.n861 VDDA.n830 3.4105
R1681 VDDA.n855 VDDA.n830 3.4105
R1682 VDDA.n863 VDDA.n830 3.4105
R1683 VDDA.n854 VDDA.n830 3.4105
R1684 VDDA.n865 VDDA.n830 3.4105
R1685 VDDA.n853 VDDA.n830 3.4105
R1686 VDDA.n867 VDDA.n830 3.4105
R1687 VDDA.n852 VDDA.n830 3.4105
R1688 VDDA.n869 VDDA.n830 3.4105
R1689 VDDA.n851 VDDA.n830 3.4105
R1690 VDDA.n871 VDDA.n830 3.4105
R1691 VDDA.n850 VDDA.n830 3.4105
R1692 VDDA.n873 VDDA.n830 3.4105
R1693 VDDA.n849 VDDA.n830 3.4105
R1694 VDDA.n875 VDDA.n830 3.4105
R1695 VDDA.n848 VDDA.n830 3.4105
R1696 VDDA.n877 VDDA.n830 3.4105
R1697 VDDA.n847 VDDA.n830 3.4105
R1698 VDDA.n879 VDDA.n830 3.4105
R1699 VDDA.n846 VDDA.n830 3.4105
R1700 VDDA.n881 VDDA.n830 3.4105
R1701 VDDA.n845 VDDA.n830 3.4105
R1702 VDDA.n883 VDDA.n830 3.4105
R1703 VDDA.n844 VDDA.n830 3.4105
R1704 VDDA.n885 VDDA.n830 3.4105
R1705 VDDA.n843 VDDA.n830 3.4105
R1706 VDDA.n887 VDDA.n830 3.4105
R1707 VDDA.n842 VDDA.n830 3.4105
R1708 VDDA.n830 VDDA.n18 3.4105
R1709 VDDA.n889 VDDA.n830 3.4105
R1710 VDDA.n779 VDDA.n16 3.4105
R1711 VDDA.n859 VDDA.n779 3.4105
R1712 VDDA.n856 VDDA.n779 3.4105
R1713 VDDA.n861 VDDA.n779 3.4105
R1714 VDDA.n855 VDDA.n779 3.4105
R1715 VDDA.n863 VDDA.n779 3.4105
R1716 VDDA.n854 VDDA.n779 3.4105
R1717 VDDA.n865 VDDA.n779 3.4105
R1718 VDDA.n853 VDDA.n779 3.4105
R1719 VDDA.n867 VDDA.n779 3.4105
R1720 VDDA.n852 VDDA.n779 3.4105
R1721 VDDA.n869 VDDA.n779 3.4105
R1722 VDDA.n851 VDDA.n779 3.4105
R1723 VDDA.n871 VDDA.n779 3.4105
R1724 VDDA.n850 VDDA.n779 3.4105
R1725 VDDA.n873 VDDA.n779 3.4105
R1726 VDDA.n849 VDDA.n779 3.4105
R1727 VDDA.n875 VDDA.n779 3.4105
R1728 VDDA.n848 VDDA.n779 3.4105
R1729 VDDA.n877 VDDA.n779 3.4105
R1730 VDDA.n847 VDDA.n779 3.4105
R1731 VDDA.n879 VDDA.n779 3.4105
R1732 VDDA.n846 VDDA.n779 3.4105
R1733 VDDA.n881 VDDA.n779 3.4105
R1734 VDDA.n845 VDDA.n779 3.4105
R1735 VDDA.n883 VDDA.n779 3.4105
R1736 VDDA.n844 VDDA.n779 3.4105
R1737 VDDA.n885 VDDA.n779 3.4105
R1738 VDDA.n843 VDDA.n779 3.4105
R1739 VDDA.n887 VDDA.n779 3.4105
R1740 VDDA.n842 VDDA.n779 3.4105
R1741 VDDA.n779 VDDA.n18 3.4105
R1742 VDDA.n889 VDDA.n779 3.4105
R1743 VDDA.n833 VDDA.n16 3.4105
R1744 VDDA.n859 VDDA.n833 3.4105
R1745 VDDA.n856 VDDA.n833 3.4105
R1746 VDDA.n861 VDDA.n833 3.4105
R1747 VDDA.n855 VDDA.n833 3.4105
R1748 VDDA.n863 VDDA.n833 3.4105
R1749 VDDA.n854 VDDA.n833 3.4105
R1750 VDDA.n865 VDDA.n833 3.4105
R1751 VDDA.n853 VDDA.n833 3.4105
R1752 VDDA.n867 VDDA.n833 3.4105
R1753 VDDA.n852 VDDA.n833 3.4105
R1754 VDDA.n869 VDDA.n833 3.4105
R1755 VDDA.n851 VDDA.n833 3.4105
R1756 VDDA.n871 VDDA.n833 3.4105
R1757 VDDA.n850 VDDA.n833 3.4105
R1758 VDDA.n873 VDDA.n833 3.4105
R1759 VDDA.n849 VDDA.n833 3.4105
R1760 VDDA.n875 VDDA.n833 3.4105
R1761 VDDA.n848 VDDA.n833 3.4105
R1762 VDDA.n877 VDDA.n833 3.4105
R1763 VDDA.n847 VDDA.n833 3.4105
R1764 VDDA.n879 VDDA.n833 3.4105
R1765 VDDA.n846 VDDA.n833 3.4105
R1766 VDDA.n881 VDDA.n833 3.4105
R1767 VDDA.n845 VDDA.n833 3.4105
R1768 VDDA.n883 VDDA.n833 3.4105
R1769 VDDA.n844 VDDA.n833 3.4105
R1770 VDDA.n885 VDDA.n833 3.4105
R1771 VDDA.n843 VDDA.n833 3.4105
R1772 VDDA.n887 VDDA.n833 3.4105
R1773 VDDA.n842 VDDA.n833 3.4105
R1774 VDDA.n833 VDDA.n18 3.4105
R1775 VDDA.n889 VDDA.n833 3.4105
R1776 VDDA.n778 VDDA.n16 3.4105
R1777 VDDA.n859 VDDA.n778 3.4105
R1778 VDDA.n856 VDDA.n778 3.4105
R1779 VDDA.n861 VDDA.n778 3.4105
R1780 VDDA.n855 VDDA.n778 3.4105
R1781 VDDA.n863 VDDA.n778 3.4105
R1782 VDDA.n854 VDDA.n778 3.4105
R1783 VDDA.n865 VDDA.n778 3.4105
R1784 VDDA.n853 VDDA.n778 3.4105
R1785 VDDA.n867 VDDA.n778 3.4105
R1786 VDDA.n852 VDDA.n778 3.4105
R1787 VDDA.n869 VDDA.n778 3.4105
R1788 VDDA.n851 VDDA.n778 3.4105
R1789 VDDA.n871 VDDA.n778 3.4105
R1790 VDDA.n850 VDDA.n778 3.4105
R1791 VDDA.n873 VDDA.n778 3.4105
R1792 VDDA.n849 VDDA.n778 3.4105
R1793 VDDA.n875 VDDA.n778 3.4105
R1794 VDDA.n848 VDDA.n778 3.4105
R1795 VDDA.n877 VDDA.n778 3.4105
R1796 VDDA.n847 VDDA.n778 3.4105
R1797 VDDA.n879 VDDA.n778 3.4105
R1798 VDDA.n846 VDDA.n778 3.4105
R1799 VDDA.n881 VDDA.n778 3.4105
R1800 VDDA.n845 VDDA.n778 3.4105
R1801 VDDA.n883 VDDA.n778 3.4105
R1802 VDDA.n844 VDDA.n778 3.4105
R1803 VDDA.n885 VDDA.n778 3.4105
R1804 VDDA.n843 VDDA.n778 3.4105
R1805 VDDA.n887 VDDA.n778 3.4105
R1806 VDDA.n842 VDDA.n778 3.4105
R1807 VDDA.n778 VDDA.n18 3.4105
R1808 VDDA.n889 VDDA.n778 3.4105
R1809 VDDA.n836 VDDA.n16 3.4105
R1810 VDDA.n859 VDDA.n836 3.4105
R1811 VDDA.n856 VDDA.n836 3.4105
R1812 VDDA.n861 VDDA.n836 3.4105
R1813 VDDA.n855 VDDA.n836 3.4105
R1814 VDDA.n863 VDDA.n836 3.4105
R1815 VDDA.n854 VDDA.n836 3.4105
R1816 VDDA.n865 VDDA.n836 3.4105
R1817 VDDA.n853 VDDA.n836 3.4105
R1818 VDDA.n867 VDDA.n836 3.4105
R1819 VDDA.n852 VDDA.n836 3.4105
R1820 VDDA.n869 VDDA.n836 3.4105
R1821 VDDA.n851 VDDA.n836 3.4105
R1822 VDDA.n871 VDDA.n836 3.4105
R1823 VDDA.n850 VDDA.n836 3.4105
R1824 VDDA.n873 VDDA.n836 3.4105
R1825 VDDA.n849 VDDA.n836 3.4105
R1826 VDDA.n875 VDDA.n836 3.4105
R1827 VDDA.n848 VDDA.n836 3.4105
R1828 VDDA.n877 VDDA.n836 3.4105
R1829 VDDA.n847 VDDA.n836 3.4105
R1830 VDDA.n879 VDDA.n836 3.4105
R1831 VDDA.n846 VDDA.n836 3.4105
R1832 VDDA.n881 VDDA.n836 3.4105
R1833 VDDA.n845 VDDA.n836 3.4105
R1834 VDDA.n883 VDDA.n836 3.4105
R1835 VDDA.n844 VDDA.n836 3.4105
R1836 VDDA.n885 VDDA.n836 3.4105
R1837 VDDA.n843 VDDA.n836 3.4105
R1838 VDDA.n887 VDDA.n836 3.4105
R1839 VDDA.n842 VDDA.n836 3.4105
R1840 VDDA.n836 VDDA.n18 3.4105
R1841 VDDA.n889 VDDA.n836 3.4105
R1842 VDDA.n777 VDDA.n16 3.4105
R1843 VDDA.n859 VDDA.n777 3.4105
R1844 VDDA.n856 VDDA.n777 3.4105
R1845 VDDA.n861 VDDA.n777 3.4105
R1846 VDDA.n855 VDDA.n777 3.4105
R1847 VDDA.n863 VDDA.n777 3.4105
R1848 VDDA.n854 VDDA.n777 3.4105
R1849 VDDA.n865 VDDA.n777 3.4105
R1850 VDDA.n853 VDDA.n777 3.4105
R1851 VDDA.n867 VDDA.n777 3.4105
R1852 VDDA.n852 VDDA.n777 3.4105
R1853 VDDA.n869 VDDA.n777 3.4105
R1854 VDDA.n851 VDDA.n777 3.4105
R1855 VDDA.n871 VDDA.n777 3.4105
R1856 VDDA.n850 VDDA.n777 3.4105
R1857 VDDA.n873 VDDA.n777 3.4105
R1858 VDDA.n849 VDDA.n777 3.4105
R1859 VDDA.n875 VDDA.n777 3.4105
R1860 VDDA.n848 VDDA.n777 3.4105
R1861 VDDA.n877 VDDA.n777 3.4105
R1862 VDDA.n847 VDDA.n777 3.4105
R1863 VDDA.n879 VDDA.n777 3.4105
R1864 VDDA.n846 VDDA.n777 3.4105
R1865 VDDA.n881 VDDA.n777 3.4105
R1866 VDDA.n845 VDDA.n777 3.4105
R1867 VDDA.n883 VDDA.n777 3.4105
R1868 VDDA.n844 VDDA.n777 3.4105
R1869 VDDA.n885 VDDA.n777 3.4105
R1870 VDDA.n843 VDDA.n777 3.4105
R1871 VDDA.n887 VDDA.n777 3.4105
R1872 VDDA.n842 VDDA.n777 3.4105
R1873 VDDA.n777 VDDA.n18 3.4105
R1874 VDDA.n889 VDDA.n777 3.4105
R1875 VDDA.n839 VDDA.n16 3.4105
R1876 VDDA.n859 VDDA.n839 3.4105
R1877 VDDA.n856 VDDA.n839 3.4105
R1878 VDDA.n861 VDDA.n839 3.4105
R1879 VDDA.n855 VDDA.n839 3.4105
R1880 VDDA.n863 VDDA.n839 3.4105
R1881 VDDA.n854 VDDA.n839 3.4105
R1882 VDDA.n865 VDDA.n839 3.4105
R1883 VDDA.n853 VDDA.n839 3.4105
R1884 VDDA.n867 VDDA.n839 3.4105
R1885 VDDA.n852 VDDA.n839 3.4105
R1886 VDDA.n869 VDDA.n839 3.4105
R1887 VDDA.n851 VDDA.n839 3.4105
R1888 VDDA.n871 VDDA.n839 3.4105
R1889 VDDA.n850 VDDA.n839 3.4105
R1890 VDDA.n873 VDDA.n839 3.4105
R1891 VDDA.n849 VDDA.n839 3.4105
R1892 VDDA.n875 VDDA.n839 3.4105
R1893 VDDA.n848 VDDA.n839 3.4105
R1894 VDDA.n877 VDDA.n839 3.4105
R1895 VDDA.n847 VDDA.n839 3.4105
R1896 VDDA.n879 VDDA.n839 3.4105
R1897 VDDA.n846 VDDA.n839 3.4105
R1898 VDDA.n881 VDDA.n839 3.4105
R1899 VDDA.n845 VDDA.n839 3.4105
R1900 VDDA.n883 VDDA.n839 3.4105
R1901 VDDA.n844 VDDA.n839 3.4105
R1902 VDDA.n885 VDDA.n839 3.4105
R1903 VDDA.n843 VDDA.n839 3.4105
R1904 VDDA.n887 VDDA.n839 3.4105
R1905 VDDA.n842 VDDA.n839 3.4105
R1906 VDDA.n839 VDDA.n18 3.4105
R1907 VDDA.n889 VDDA.n839 3.4105
R1908 VDDA.n776 VDDA.n16 3.4105
R1909 VDDA.n859 VDDA.n776 3.4105
R1910 VDDA.n856 VDDA.n776 3.4105
R1911 VDDA.n861 VDDA.n776 3.4105
R1912 VDDA.n855 VDDA.n776 3.4105
R1913 VDDA.n863 VDDA.n776 3.4105
R1914 VDDA.n854 VDDA.n776 3.4105
R1915 VDDA.n865 VDDA.n776 3.4105
R1916 VDDA.n853 VDDA.n776 3.4105
R1917 VDDA.n867 VDDA.n776 3.4105
R1918 VDDA.n852 VDDA.n776 3.4105
R1919 VDDA.n869 VDDA.n776 3.4105
R1920 VDDA.n851 VDDA.n776 3.4105
R1921 VDDA.n871 VDDA.n776 3.4105
R1922 VDDA.n850 VDDA.n776 3.4105
R1923 VDDA.n873 VDDA.n776 3.4105
R1924 VDDA.n849 VDDA.n776 3.4105
R1925 VDDA.n875 VDDA.n776 3.4105
R1926 VDDA.n848 VDDA.n776 3.4105
R1927 VDDA.n877 VDDA.n776 3.4105
R1928 VDDA.n847 VDDA.n776 3.4105
R1929 VDDA.n879 VDDA.n776 3.4105
R1930 VDDA.n846 VDDA.n776 3.4105
R1931 VDDA.n881 VDDA.n776 3.4105
R1932 VDDA.n845 VDDA.n776 3.4105
R1933 VDDA.n883 VDDA.n776 3.4105
R1934 VDDA.n844 VDDA.n776 3.4105
R1935 VDDA.n885 VDDA.n776 3.4105
R1936 VDDA.n843 VDDA.n776 3.4105
R1937 VDDA.n887 VDDA.n776 3.4105
R1938 VDDA.n842 VDDA.n776 3.4105
R1939 VDDA.n776 VDDA.n18 3.4105
R1940 VDDA.n889 VDDA.n776 3.4105
R1941 VDDA.n888 VDDA.n859 3.4105
R1942 VDDA.n888 VDDA.n856 3.4105
R1943 VDDA.n888 VDDA.n861 3.4105
R1944 VDDA.n888 VDDA.n855 3.4105
R1945 VDDA.n888 VDDA.n863 3.4105
R1946 VDDA.n888 VDDA.n854 3.4105
R1947 VDDA.n888 VDDA.n865 3.4105
R1948 VDDA.n888 VDDA.n853 3.4105
R1949 VDDA.n888 VDDA.n867 3.4105
R1950 VDDA.n888 VDDA.n852 3.4105
R1951 VDDA.n888 VDDA.n869 3.4105
R1952 VDDA.n888 VDDA.n851 3.4105
R1953 VDDA.n888 VDDA.n871 3.4105
R1954 VDDA.n888 VDDA.n850 3.4105
R1955 VDDA.n888 VDDA.n873 3.4105
R1956 VDDA.n888 VDDA.n849 3.4105
R1957 VDDA.n888 VDDA.n875 3.4105
R1958 VDDA.n888 VDDA.n848 3.4105
R1959 VDDA.n888 VDDA.n877 3.4105
R1960 VDDA.n888 VDDA.n847 3.4105
R1961 VDDA.n888 VDDA.n879 3.4105
R1962 VDDA.n888 VDDA.n846 3.4105
R1963 VDDA.n888 VDDA.n881 3.4105
R1964 VDDA.n888 VDDA.n845 3.4105
R1965 VDDA.n888 VDDA.n883 3.4105
R1966 VDDA.n888 VDDA.n844 3.4105
R1967 VDDA.n888 VDDA.n885 3.4105
R1968 VDDA.n888 VDDA.n843 3.4105
R1969 VDDA.n888 VDDA.n887 3.4105
R1970 VDDA.n888 VDDA.n842 3.4105
R1971 VDDA.n888 VDDA.n18 3.4105
R1972 VDDA.n889 VDDA.n888 3.4105
R1973 VDDA.n335 VDDA.n334 3.11118
R1974 VDDA.n345 VDDA.n344 3.11118
R1975 VDDA.n334 VDDA.n316 3.04304
R1976 VDDA.n344 VDDA.n296 3.04304
R1977 VDDA.n238 VDDA.n234 2.96402
R1978 VDDA.n743 VDDA.n739 2.96402
R1979 VDDA.n669 VDDA.n668 2.8255
R1980 VDDA.n671 VDDA.n670 2.8255
R1981 VDDA.n237 VDDA.n236 2.423
R1982 VDDA.n235 VDDA.n234 2.423
R1983 VDDA.n740 VDDA.n739 2.423
R1984 VDDA.n742 VDDA.n741 2.423
R1985 VDDA.n709 VDDA.n707 2.3971
R1986 VDDA.n640 VDDA.n206 2.39632
R1987 VDDA.n136 VDDA.n135 2.30736
R1988 VDDA.n549 VDDA.n547 2.30736
R1989 VDDA.n99 VDDA.n98 2.30612
R1990 VDDA.n534 VDDA.n533 2.30612
R1991 VDDA.n238 VDDA.n237 2.27652
R1992 VDDA.n743 VDDA.n742 2.27652
R1993 VDDA.n290 VDDA.n282 2.26187
R1994 VDDA.n356 VDDA.n280 2.26187
R1995 VDDA.n433 VDDA.n278 2.26187
R1996 VDDA.n483 VDDA.n276 2.26187
R1997 VDDA.n660 VDDA.n651 2.26187
R1998 VDDA.n662 VDDA.n660 2.26187
R1999 VDDA.n749 VDDA.n748 2.26187
R2000 VDDA.n736 VDDA.n714 2.26187
R2001 VDDA.n720 VDDA.n717 2.26187
R2002 VDDA.n721 VDDA.n720 2.26187
R2003 VDDA.n639 VDDA.n638 2.26187
R2004 VDDA.n231 VDDA.n230 2.26187
R2005 VDDA.n614 VDDA.n613 2.26187
R2006 VDDA.n613 VDDA.n247 2.26187
R2007 VDDA.n287 VDDA.n282 2.26187
R2008 VDDA.n232 VDDA.n231 2.26187
R2009 VDDA.n243 VDDA.n242 2.26187
R2010 VDDA.n678 VDDA.n677 2.26187
R2011 VDDA.n291 VDDA.n281 2.24063
R2012 VDDA.n357 VDDA.n279 2.24063
R2013 VDDA.n434 VDDA.n277 2.24063
R2014 VDDA.n484 VDDA.n275 2.24063
R2015 VDDA.n679 VDDA.n678 2.24063
R2016 VDDA.n673 VDDA.n649 2.24063
R2017 VDDA.n675 VDDA.n674 2.24063
R2018 VDDA.n665 VDDA.n664 2.24063
R2019 VDDA.n770 VDDA.n769 2.24063
R2020 VDDA.n179 VDDA.n178 2.24063
R2021 VDDA.n747 VDDA.n182 2.24063
R2022 VDDA.n738 VDDA.n737 2.24063
R2023 VDDA.n708 VDDA.n185 2.24063
R2024 VDDA.n692 VDDA.n184 2.24063
R2025 VDDA.n682 VDDA.n681 2.24063
R2026 VDDA.n648 VDDA.n189 2.24063
R2027 VDDA.n637 VDDA.n190 2.24063
R2028 VDDA.n240 VDDA.n239 2.24063
R2029 VDDA.n242 VDDA.n241 2.24063
R2030 VDDA.n230 VDDA.n229 2.24063
R2031 VDDA.n635 VDDA.n634 2.24063
R2032 VDDA.n211 VDDA.n210 2.24063
R2033 VDDA.n287 VDDA.n286 2.24063
R2034 VDDA.n292 VDDA.n280 2.24063
R2035 VDDA.n353 VDDA.n352 2.24063
R2036 VDDA.n358 VDDA.n278 2.24063
R2037 VDDA.n430 VDDA.n429 2.24063
R2038 VDDA.n435 VDDA.n276 2.24063
R2039 VDDA.n480 VDDA.n479 2.24063
R2040 VDDA.n663 VDDA.n662 2.24063
R2041 VDDA.n771 VDDA.n176 2.24063
R2042 VDDA.n750 VDDA.n749 2.24063
R2043 VDDA.n752 VDDA.n751 2.24063
R2044 VDDA.n746 VDDA.n714 2.24063
R2045 VDDA.n745 VDDA.n744 2.24063
R2046 VDDA.n735 VDDA.n717 2.24063
R2047 VDDA.n734 VDDA.n733 2.24063
R2048 VDDA.n710 VDDA.n709 2.24063
R2049 VDDA.n640 VDDA.n639 2.24063
R2050 VDDA.n642 VDDA.n641 2.24063
R2051 VDDA.n244 VDDA.n212 2.24063
R2052 VDDA.n233 VDDA.n215 2.24063
R2053 VDDA.n636 VDDA.n208 2.24063
R2054 VDDA.n615 VDDA.n614 2.24063
R2055 VDDA.n617 VDDA.n616 2.24063
R2056 VDDA.n765 VDDA.n764 1.97758
R2057 VDDA.n763 VDDA.n762 1.97758
R2058 VDDA.n630 VDDA.n629 1.97758
R2059 VDDA.n628 VDDA.n627 1.97758
R2060 VDDA.n333 VDDA.n332 1.90331
R2061 VDDA.n658 VDDA.n657 1.888
R2062 VDDA.n656 VDDA.n655 1.888
R2063 VDDA.n704 VDDA.n703 1.888
R2064 VDDA.n706 VDDA.n705 1.888
R2065 VDDA.n205 VDDA.n204 1.888
R2066 VDDA.n203 VDDA.n202 1.888
R2067 VDDA.n766 VDDA.n765 1.88069
R2068 VDDA.n762 VDDA.n761 1.88069
R2069 VDDA.n631 VDDA.n630 1.88069
R2070 VDDA.n627 VDDA.n626 1.88069
R2071 VDDA.n341 VDDA.n340 1.77831
R2072 VDDA.n343 VDDA.n342 1.77831
R2073 VDDA.n351 VDDA.n350 1.77831
R2074 VDDA.n274 VDDA.n262 1.73971
R2075 VDDA.n536 VDDA.n262 1.70624
R2076 VDDA.n792 VDDA.n0 1.70567
R2077 VDDA.n793 VDDA.n17 1.70567
R2078 VDDA.n795 VDDA.n792 1.70567
R2079 VDDA.n796 VDDA.n17 1.70567
R2080 VDDA.n798 VDDA.n792 1.70567
R2081 VDDA.n799 VDDA.n17 1.70567
R2082 VDDA.n801 VDDA.n792 1.70567
R2083 VDDA.n802 VDDA.n17 1.70567
R2084 VDDA.n804 VDDA.n792 1.70567
R2085 VDDA.n805 VDDA.n17 1.70567
R2086 VDDA.n807 VDDA.n792 1.70567
R2087 VDDA.n808 VDDA.n17 1.70567
R2088 VDDA.n810 VDDA.n792 1.70567
R2089 VDDA.n811 VDDA.n17 1.70567
R2090 VDDA.n813 VDDA.n792 1.70567
R2091 VDDA.n814 VDDA.n17 1.70567
R2092 VDDA.n816 VDDA.n792 1.70567
R2093 VDDA.n817 VDDA.n17 1.70567
R2094 VDDA.n819 VDDA.n792 1.70567
R2095 VDDA.n820 VDDA.n17 1.70567
R2096 VDDA.n822 VDDA.n792 1.70567
R2097 VDDA.n823 VDDA.n17 1.70567
R2098 VDDA.n825 VDDA.n792 1.70567
R2099 VDDA.n826 VDDA.n17 1.70567
R2100 VDDA.n828 VDDA.n792 1.70567
R2101 VDDA.n829 VDDA.n17 1.70567
R2102 VDDA.n831 VDDA.n792 1.70567
R2103 VDDA.n832 VDDA.n17 1.70567
R2104 VDDA.n834 VDDA.n792 1.70567
R2105 VDDA.n835 VDDA.n17 1.70567
R2106 VDDA.n837 VDDA.n792 1.70567
R2107 VDDA.n838 VDDA.n17 1.70567
R2108 VDDA.n840 VDDA.n792 1.70567
R2109 VDDA.n890 VDDA.n15 1.70566
R2110 VDDA.n890 VDDA.n14 1.70566
R2111 VDDA.n890 VDDA.n13 1.70566
R2112 VDDA.n890 VDDA.n12 1.70566
R2113 VDDA.n890 VDDA.n11 1.70566
R2114 VDDA.n890 VDDA.n10 1.70566
R2115 VDDA.n890 VDDA.n9 1.70566
R2116 VDDA.n890 VDDA.n8 1.70566
R2117 VDDA.n890 VDDA.n7 1.70566
R2118 VDDA.n890 VDDA.n6 1.70566
R2119 VDDA.n890 VDDA.n5 1.70566
R2120 VDDA.n890 VDDA.n4 1.70566
R2121 VDDA.n890 VDDA.n3 1.70566
R2122 VDDA.n890 VDDA.n2 1.70566
R2123 VDDA.n890 VDDA.n1 1.70566
R2124 VDDA.n858 VDDA.n794 1.70566
R2125 VDDA.n860 VDDA.n794 1.70566
R2126 VDDA.n862 VDDA.n794 1.70566
R2127 VDDA.n864 VDDA.n794 1.70566
R2128 VDDA.n866 VDDA.n794 1.70566
R2129 VDDA.n868 VDDA.n794 1.70566
R2130 VDDA.n870 VDDA.n794 1.70566
R2131 VDDA.n872 VDDA.n794 1.70566
R2132 VDDA.n874 VDDA.n794 1.70566
R2133 VDDA.n876 VDDA.n794 1.70566
R2134 VDDA.n878 VDDA.n794 1.70566
R2135 VDDA.n880 VDDA.n794 1.70566
R2136 VDDA.n882 VDDA.n794 1.70566
R2137 VDDA.n884 VDDA.n794 1.70566
R2138 VDDA.n886 VDDA.n794 1.70566
R2139 VDDA.n841 VDDA.n794 1.70566
R2140 VDDA.n888 VDDA.n857 1.70566
R2141 VDDA.n608 VDDA.n538 1.69337
R2142 VDDA.n608 VDDA.n539 1.69337
R2143 VDDA.n608 VDDA.n541 1.69337
R2144 VDDA.n608 VDDA.n542 1.69337
R2145 VDDA.n608 VDDA.n544 1.69337
R2146 VDDA.n608 VDDA.n545 1.69337
R2147 VDDA.n608 VDDA.n607 1.69337
R2148 VDDA.n536 VDDA.n253 1.69337
R2149 VDDA.n536 VDDA.n254 1.69337
R2150 VDDA.n536 VDDA.n256 1.69337
R2151 VDDA.n536 VDDA.n257 1.69337
R2152 VDDA.n536 VDDA.n259 1.69337
R2153 VDDA.n536 VDDA.n260 1.69337
R2154 VDDA.n775 VDDA.n103 1.69337
R2155 VDDA.n775 VDDA.n104 1.69337
R2156 VDDA.n775 VDDA.n106 1.69337
R2157 VDDA.n775 VDDA.n107 1.69337
R2158 VDDA.n775 VDDA.n109 1.69337
R2159 VDDA.n775 VDDA.n110 1.69337
R2160 VDDA.n775 VDDA.n112 1.69337
R2161 VDDA.n101 VDDA.n20 1.69337
R2162 VDDA.n101 VDDA.n21 1.69337
R2163 VDDA.n101 VDDA.n23 1.69337
R2164 VDDA.n101 VDDA.n24 1.69337
R2165 VDDA.n101 VDDA.n26 1.69337
R2166 VDDA.n101 VDDA.n27 1.69337
R2167 VDDA.n101 VDDA.n29 1.69337
R2168 VDDA.n608 VDDA.n537 1.6924
R2169 VDDA.n608 VDDA.n540 1.6924
R2170 VDDA.n608 VDDA.n543 1.6924
R2171 VDDA.n608 VDDA.n546 1.6924
R2172 VDDA.n536 VDDA.n252 1.6924
R2173 VDDA.n536 VDDA.n255 1.6924
R2174 VDDA.n536 VDDA.n258 1.6924
R2175 VDDA.n536 VDDA.n261 1.6924
R2176 VDDA.n775 VDDA.n102 1.6924
R2177 VDDA.n775 VDDA.n105 1.6924
R2178 VDDA.n775 VDDA.n108 1.6924
R2179 VDDA.n775 VDDA.n111 1.6924
R2180 VDDA.n101 VDDA.n19 1.6924
R2181 VDDA.n101 VDDA.n22 1.6924
R2182 VDDA.n101 VDDA.n25 1.6924
R2183 VDDA.n101 VDDA.n28 1.6924
R2184 VDDA.n459 VDDA.n457 1.68456
R2185 VDDA.n655 VDDA.n653 1.63212
R2186 VDDA.n668 VDDA.n667 1.63212
R2187 VDDA.n475 VDDA.n441 1.56997
R2188 VDDA.n470 VDDA.n444 1.56997
R2189 VDDA.n462 VDDA.n454 1.56997
R2190 VDDA.n659 VDDA.n658 1.56962
R2191 VDDA.n672 VDDA.n671 1.56962
R2192 VDDA.n286 VDDA.n285 1.26222
R2193 VDDA.n889 VDDA.n775 1.17314
R2194 VDDA.n747 VDDA.n746 1.14633
R2195 VDDA.n633 VDDA.n244 1.14633
R2196 VDDA.n737 VDDA.n735 1.06821
R2197 VDDA.n241 VDDA.n233 1.06821
R2198 VDDA.n292 VDDA.n291 0.943208
R2199 VDDA.n645 VDDA.n642 0.932792
R2200 VDDA.n711 VDDA.n690 0.932792
R2201 VDDA.n767 VDDA.n766 0.885917
R2202 VDDA.n626 VDDA.n617 0.885917
R2203 VDDA.n429 VDDA.n428 0.880708
R2204 VDDA.n352 VDDA.n351 0.865083
R2205 VDDA.n479 VDDA.n478 0.807792
R2206 VDDA.n284 VDDA.n283 0.75233
R2207 VDDA.n358 VDDA.n357 0.672375
R2208 VDDA.n285 VDDA.n284 0.648711
R2209 VDDA.n750 VDDA.n712 0.495292
R2210 VDDA.n637 VDDA.n636 0.495292
R2211 VDDA.n485 VDDA.n484 0.448417
R2212 VDDA.n680 VDDA.n679 0.417167
R2213 VDDA.n707 VDDA.n694 0.3755
R2214 VDDA.n696 VDDA.n694 0.3755
R2215 VDDA.n698 VDDA.n696 0.3755
R2216 VDDA.n700 VDDA.n698 0.3755
R2217 VDDA.n702 VDDA.n700 0.3755
R2218 VDDA.n201 VDDA.n199 0.3755
R2219 VDDA.n199 VDDA.n197 0.3755
R2220 VDDA.n197 VDDA.n195 0.3755
R2221 VDDA.n195 VDDA.n193 0.3755
R2222 VDDA.n206 VDDA.n193 0.3755
R2223 VDDA.n342 VDDA.n341 0.333833
R2224 VDDA.n423 VDDA.n422 0.328625
R2225 VDDA.n229 VDDA.n228 0.323417
R2226 VDDA.n733 VDDA.n732 0.323417
R2227 VDDA.n476 VDDA.n475 0.292167
R2228 VDDA.n470 VDDA.n469 0.292167
R2229 VDDA.n463 VDDA.n462 0.292167
R2230 VDDA.n435 VDDA.n434 0.292167
R2231 VDDA.n239 VDDA.n238 0.266125
R2232 VDDA.n744 VDDA.n743 0.266125
R2233 VDDA.n761 VDDA.n752 0.266125
R2234 VDDA.n632 VDDA.n631 0.266125
R2235 VDDA.n340 VDDA.n339 0.2505
R2236 VDDA.n350 VDDA.n349 0.2505
R2237 VDDA.n428 VDDA.n423 0.229667
R2238 VDDA.n663 VDDA.n659 0.214042
R2239 VDDA.n673 VDDA.n672 0.214042
R2240 VDDA.n390 VDDA.n376 0.208833
R2241 VDDA.n384 VDDA.n376 0.208833
R2242 VDDA.n384 VDDA.n383 0.208833
R2243 VDDA.n399 VDDA.n397 0.208833
R2244 VDDA.n400 VDDA.n399 0.208833
R2245 VDDA.n400 VDDA.n369 0.208833
R2246 VDDA.n422 VDDA.n421 0.188
R2247 VDDA.n421 VDDA.n420 0.188
R2248 VDDA.n420 VDDA.n419 0.188
R2249 VDDA.n419 VDDA.n418 0.188
R2250 VDDA.n418 VDDA.n417 0.188
R2251 VDDA.n417 VDDA.n416 0.188
R2252 VDDA.n416 VDDA.n415 0.188
R2253 VDDA.n415 VDDA.n414 0.188
R2254 VDDA.n647 VDDA.n645 0.172375
R2255 VDDA.n682 VDDA.n647 0.172375
R2256 VDDA.n648 VDDA.n187 0.172375
R2257 VDDA.n690 VDDA.n187 0.172375
R2258 VDDA.t382 VDDA.t395 0.1603
R2259 VDDA.t87 VDDA.t108 0.1603
R2260 VDDA.t143 VDDA.t379 0.1603
R2261 VDDA.t17 VDDA.t409 0.1603
R2262 VDDA.t104 VDDA.t101 0.1603
R2263 VDDA.n43 VDDA.t82 0.159278
R2264 VDDA.n44 VDDA.t144 0.159278
R2265 VDDA.n45 VDDA.t88 0.159278
R2266 VDDA.n46 VDDA.t151 0.159278
R2267 VDDA.n53 VDDA.n41 0.146333
R2268 VDDA.n54 VDDA.n53 0.146333
R2269 VDDA.n57 VDDA.n54 0.146333
R2270 VDDA.n67 VDDA.n64 0.146333
R2271 VDDA.n67 VDDA.n37 0.146333
R2272 VDDA.n73 VDDA.n37 0.146333
R2273 VDDA.n83 VDDA.n35 0.146333
R2274 VDDA.n84 VDDA.n83 0.146333
R2275 VDDA.n87 VDDA.n84 0.146333
R2276 VDDA.n97 VDDA.n94 0.146333
R2277 VDDA.n97 VDDA.n31 0.146333
R2278 VDDA.n488 VDDA.n274 0.146333
R2279 VDDA.n489 VDDA.n488 0.146333
R2280 VDDA.n492 VDDA.n489 0.146333
R2281 VDDA.n502 VDDA.n499 0.146333
R2282 VDDA.n502 VDDA.n270 0.146333
R2283 VDDA.n508 VDDA.n270 0.146333
R2284 VDDA.n518 VDDA.n268 0.146333
R2285 VDDA.n519 VDDA.n518 0.146333
R2286 VDDA.n522 VDDA.n519 0.146333
R2287 VDDA.n532 VDDA.n529 0.146333
R2288 VDDA.n532 VDDA.n264 0.146333
R2289 VDDA.n137 VDDA.n132 0.146333
R2290 VDDA.n138 VDDA.n137 0.146333
R2291 VDDA.n141 VDDA.n138 0.146333
R2292 VDDA.n149 VDDA.n146 0.146333
R2293 VDDA.n149 VDDA.n124 0.146333
R2294 VDDA.n153 VDDA.n124 0.146333
R2295 VDDA.n161 VDDA.n120 0.146333
R2296 VDDA.n162 VDDA.n161 0.146333
R2297 VDDA.n165 VDDA.n162 0.146333
R2298 VDDA.n173 VDDA.n170 0.146333
R2299 VDDA.n173 VDDA.n114 0.146333
R2300 VDDA.n773 VDDA.n114 0.146333
R2301 VDDA.n604 VDDA.n548 0.146333
R2302 VDDA.n604 VDDA.n603 0.146333
R2303 VDDA.n603 VDDA.n600 0.146333
R2304 VDDA.n595 VDDA.n592 0.146333
R2305 VDDA.n592 VDDA.n591 0.146333
R2306 VDDA.n591 VDDA.n588 0.146333
R2307 VDDA.n583 VDDA.n580 0.146333
R2308 VDDA.n580 VDDA.n579 0.146333
R2309 VDDA.n579 VDDA.n576 0.146333
R2310 VDDA.n571 VDDA.n568 0.146333
R2311 VDDA.n568 VDDA.n250 0.146333
R2312 VDDA.n610 VDDA.n250 0.146333
R2313 VDDA.n46 VDDA.t18 0.1368
R2314 VDDA.n46 VDDA.t382 0.1368
R2315 VDDA.n45 VDDA.t410 0.1368
R2316 VDDA.n45 VDDA.t87 0.1368
R2317 VDDA.n44 VDDA.t171 0.1368
R2318 VDDA.n44 VDDA.t143 0.1368
R2319 VDDA.n43 VDDA.t81 0.1368
R2320 VDDA.n43 VDDA.t17 0.1368
R2321 VDDA.n42 VDDA.t107 0.1368
R2322 VDDA.n42 VDDA.t104 0.1368
R2323 VDDA.n536 VDDA.n101 0.136024
R2324 VDDA.n47 VDDA.n41 0.135917
R2325 VDDA.n57 VDDA.n39 0.135917
R2326 VDDA.n64 VDDA.n63 0.135917
R2327 VDDA.n74 VDDA.n73 0.135917
R2328 VDDA.n77 VDDA.n35 0.135917
R2329 VDDA.n87 VDDA.n33 0.135917
R2330 VDDA.n94 VDDA.n93 0.135917
R2331 VDDA.n492 VDDA.n272 0.135917
R2332 VDDA.n499 VDDA.n498 0.135917
R2333 VDDA.n509 VDDA.n508 0.135917
R2334 VDDA.n512 VDDA.n268 0.135917
R2335 VDDA.n522 VDDA.n266 0.135917
R2336 VDDA.n529 VDDA.n528 0.135917
R2337 VDDA.n141 VDDA.n128 0.135917
R2338 VDDA.n146 VDDA.n145 0.135917
R2339 VDDA.n154 VDDA.n153 0.135917
R2340 VDDA.n157 VDDA.n120 0.135917
R2341 VDDA.n165 VDDA.n116 0.135917
R2342 VDDA.n170 VDDA.n169 0.135917
R2343 VDDA.n600 VDDA.n599 0.135917
R2344 VDDA.n596 VDDA.n595 0.135917
R2345 VDDA.n588 VDDA.n587 0.135917
R2346 VDDA.n584 VDDA.n583 0.135917
R2347 VDDA.n576 VDDA.n575 0.135917
R2348 VDDA.n572 VDDA.n571 0.135917
R2349 VDDA.n63 VDDA.n39 0.1255
R2350 VDDA.n77 VDDA.n74 0.1255
R2351 VDDA.n93 VDDA.n33 0.1255
R2352 VDDA.n478 VDDA.n477 0.1255
R2353 VDDA.n477 VDDA.n476 0.1255
R2354 VDDA.n351 VDDA.n294 0.1255
R2355 VDDA.n298 VDDA.n294 0.1255
R2356 VDDA.n300 VDDA.n298 0.1255
R2357 VDDA.n302 VDDA.n300 0.1255
R2358 VDDA.n304 VDDA.n302 0.1255
R2359 VDDA.n306 VDDA.n304 0.1255
R2360 VDDA.n308 VDDA.n306 0.1255
R2361 VDDA.n310 VDDA.n308 0.1255
R2362 VDDA.n312 VDDA.n310 0.1255
R2363 VDDA.n342 VDDA.n312 0.1255
R2364 VDDA.n341 VDDA.n314 0.1255
R2365 VDDA.n318 VDDA.n314 0.1255
R2366 VDDA.n320 VDDA.n318 0.1255
R2367 VDDA.n322 VDDA.n320 0.1255
R2368 VDDA.n324 VDDA.n322 0.1255
R2369 VDDA.n326 VDDA.n324 0.1255
R2370 VDDA.n328 VDDA.n326 0.1255
R2371 VDDA.n330 VDDA.n328 0.1255
R2372 VDDA.n332 VDDA.n330 0.1255
R2373 VDDA.n498 VDDA.n272 0.1255
R2374 VDDA.n512 VDDA.n509 0.1255
R2375 VDDA.n528 VDDA.n266 0.1255
R2376 VDDA.n659 VDDA.n653 0.1255
R2377 VDDA.n672 VDDA.n667 0.1255
R2378 VDDA.n145 VDDA.n128 0.1255
R2379 VDDA.n157 VDDA.n154 0.1255
R2380 VDDA.n169 VDDA.n116 0.1255
R2381 VDDA.n599 VDDA.n596 0.1255
R2382 VDDA.n587 VDDA.n584 0.1255
R2383 VDDA.n575 VDDA.n572 0.1255
R2384 VDDA.n475 VDDA.n474 0.115083
R2385 VDDA.n474 VDDA.n472 0.115083
R2386 VDDA.n472 VDDA.n470 0.115083
R2387 VDDA.n468 VDDA.n467 0.115083
R2388 VDDA.n467 VDDA.n466 0.115083
R2389 VDDA.n466 VDDA.n465 0.115083
R2390 VDDA.n465 VDDA.n464 0.115083
R2391 VDDA.n462 VDDA.n461 0.115083
R2392 VDDA.n461 VDDA.n459 0.115083
R2393 VDDA.n222 VDDA.n220 0.115083
R2394 VDDA.n224 VDDA.n222 0.115083
R2395 VDDA.n226 VDDA.n224 0.115083
R2396 VDDA.n228 VDDA.n226 0.115083
R2397 VDDA.n732 VDDA.n730 0.115083
R2398 VDDA.n730 VDDA.n728 0.115083
R2399 VDDA.n728 VDDA.n726 0.115083
R2400 VDDA.n726 VDDA.n724 0.115083
R2401 VDDA.n761 VDDA.n760 0.115083
R2402 VDDA.n760 VDDA.n758 0.115083
R2403 VDDA.n758 VDDA.n756 0.115083
R2404 VDDA.n756 VDDA.n754 0.115083
R2405 VDDA.n754 VDDA.n181 0.115083
R2406 VDDA.n766 VDDA.n181 0.115083
R2407 VDDA.n626 VDDA.n625 0.115083
R2408 VDDA.n625 VDDA.n623 0.115083
R2409 VDDA.n623 VDDA.n621 0.115083
R2410 VDDA.n621 VDDA.n619 0.115083
R2411 VDDA.n619 VDDA.n246 0.115083
R2412 VDDA.n631 VDDA.n246 0.115083
R2413 VDDA.n675 VDDA.n665 0.09425
R2414 VDDA.n682 VDDA.n648 0.0838333
R2415 VDDA.n50 VDDA.n49 0.0734167
R2416 VDDA.n50 VDDA.n40 0.0734167
R2417 VDDA.n58 VDDA.n40 0.0734167
R2418 VDDA.n68 VDDA.n38 0.0734167
R2419 VDDA.n69 VDDA.n68 0.0734167
R2420 VDDA.n70 VDDA.n69 0.0734167
R2421 VDDA.n80 VDDA.n79 0.0734167
R2422 VDDA.n80 VDDA.n34 0.0734167
R2423 VDDA.n88 VDDA.n34 0.0734167
R2424 VDDA.n98 VDDA.n32 0.0734167
R2425 VDDA.n486 VDDA.n485 0.0734167
R2426 VDDA.n486 VDDA.n273 0.0734167
R2427 VDDA.n493 VDDA.n273 0.0734167
R2428 VDDA.n503 VDDA.n271 0.0734167
R2429 VDDA.n504 VDDA.n503 0.0734167
R2430 VDDA.n505 VDDA.n504 0.0734167
R2431 VDDA.n515 VDDA.n514 0.0734167
R2432 VDDA.n515 VDDA.n267 0.0734167
R2433 VDDA.n523 VDDA.n267 0.0734167
R2434 VDDA.n533 VDDA.n265 0.0734167
R2435 VDDA.n136 VDDA.n131 0.0734167
R2436 VDDA.n142 VDDA.n131 0.0734167
R2437 VDDA.n150 VDDA.n127 0.0734167
R2438 VDDA.n151 VDDA.n150 0.0734167
R2439 VDDA.n152 VDDA.n151 0.0734167
R2440 VDDA.n160 VDDA.n159 0.0734167
R2441 VDDA.n160 VDDA.n119 0.0734167
R2442 VDDA.n166 VDDA.n119 0.0734167
R2443 VDDA.n174 VDDA.n115 0.0734167
R2444 VDDA.n175 VDDA.n174 0.0734167
R2445 VDDA.n772 VDDA.n175 0.0734167
R2446 VDDA.n550 VDDA.n549 0.0734167
R2447 VDDA.n551 VDDA.n550 0.0734167
R2448 VDDA.n555 VDDA.n554 0.0734167
R2449 VDDA.n556 VDDA.n555 0.0734167
R2450 VDDA.n557 VDDA.n556 0.0734167
R2451 VDDA.n561 VDDA.n560 0.0734167
R2452 VDDA.n562 VDDA.n561 0.0734167
R2453 VDDA.n563 VDDA.n562 0.0734167
R2454 VDDA.n567 VDDA.n566 0.0734167
R2455 VDDA.n567 VDDA.n249 0.0734167
R2456 VDDA.n611 VDDA.n249 0.0734167
R2457 VDDA.n99 VDDA.n31 0.0721864
R2458 VDDA.n534 VDDA.n264 0.0721864
R2459 VDDA.n487 VDDA.n262 0.0683791
R2460 VDDA.n49 VDDA.n48 0.0682083
R2461 VDDA.n59 VDDA.n58 0.0682083
R2462 VDDA.n60 VDDA.n38 0.0682083
R2463 VDDA.n70 VDDA.n36 0.0682083
R2464 VDDA.n79 VDDA.n78 0.0682083
R2465 VDDA.n89 VDDA.n88 0.0682083
R2466 VDDA.n90 VDDA.n32 0.0682083
R2467 VDDA.n469 VDDA.n468 0.0682083
R2468 VDDA.n464 VDDA.n463 0.0682083
R2469 VDDA.n494 VDDA.n493 0.0682083
R2470 VDDA.n495 VDDA.n271 0.0682083
R2471 VDDA.n505 VDDA.n269 0.0682083
R2472 VDDA.n514 VDDA.n513 0.0682083
R2473 VDDA.n524 VDDA.n523 0.0682083
R2474 VDDA.n525 VDDA.n265 0.0682083
R2475 VDDA.n143 VDDA.n142 0.0682083
R2476 VDDA.n144 VDDA.n127 0.0682083
R2477 VDDA.n152 VDDA.n123 0.0682083
R2478 VDDA.n159 VDDA.n158 0.0682083
R2479 VDDA.n167 VDDA.n166 0.0682083
R2480 VDDA.n168 VDDA.n115 0.0682083
R2481 VDDA.n552 VDDA.n551 0.0682083
R2482 VDDA.n554 VDDA.n553 0.0682083
R2483 VDDA.n558 VDDA.n557 0.0682083
R2484 VDDA.n560 VDDA.n559 0.0682083
R2485 VDDA.n564 VDDA.n563 0.0682083
R2486 VDDA.n566 VDDA.n565 0.0682083
R2487 VDDA.n135 VDDA.n132 0.0672139
R2488 VDDA.n548 VDDA.n547 0.0672139
R2489 VDDA.n60 VDDA.n59 0.063
R2490 VDDA.n78 VDDA.n36 0.063
R2491 VDDA.n90 VDDA.n89 0.063
R2492 VDDA.n495 VDDA.n494 0.063
R2493 VDDA.n513 VDDA.n269 0.063
R2494 VDDA.n525 VDDA.n524 0.063
R2495 VDDA.n144 VDDA.n143 0.063
R2496 VDDA.n158 VDDA.n123 0.063
R2497 VDDA.n168 VDDA.n167 0.063
R2498 VDDA.n553 VDDA.n552 0.063
R2499 VDDA.n559 VDDA.n558 0.063
R2500 VDDA.n565 VDDA.n564 0.063
R2501 VDDA.n52 VDDA.n51 0.0553333
R2502 VDDA.n56 VDDA.n55 0.0553333
R2503 VDDA.n66 VDDA.n65 0.0553333
R2504 VDDA.n72 VDDA.n71 0.0553333
R2505 VDDA.n82 VDDA.n81 0.0553333
R2506 VDDA.n86 VDDA.n85 0.0553333
R2507 VDDA.n96 VDDA.n95 0.0553333
R2508 VDDA.n100 VDDA.n30 0.0553333
R2509 VDDA.n491 VDDA.n490 0.0553333
R2510 VDDA.n501 VDDA.n500 0.0553333
R2511 VDDA.n507 VDDA.n506 0.0553333
R2512 VDDA.n517 VDDA.n516 0.0553333
R2513 VDDA.n521 VDDA.n520 0.0553333
R2514 VDDA.n531 VDDA.n530 0.0553333
R2515 VDDA.n535 VDDA.n263 0.0553333
R2516 VDDA.n134 VDDA.n133 0.0553333
R2517 VDDA.n140 VDDA.n139 0.0553333
R2518 VDDA.n148 VDDA.n147 0.0553333
R2519 VDDA.n126 VDDA.n125 0.0553333
R2520 VDDA.n122 VDDA.n121 0.0553333
R2521 VDDA.n164 VDDA.n163 0.0553333
R2522 VDDA.n172 VDDA.n171 0.0553333
R2523 VDDA.n774 VDDA.n113 0.0553333
R2524 VDDA.n606 VDDA.n605 0.0553333
R2525 VDDA.n602 VDDA.n601 0.0553333
R2526 VDDA.n594 VDDA.n593 0.0553333
R2527 VDDA.n590 VDDA.n589 0.0553333
R2528 VDDA.n582 VDDA.n581 0.0553333
R2529 VDDA.n578 VDDA.n577 0.0553333
R2530 VDDA.n570 VDDA.n569 0.0553333
R2531 VDDA.n609 VDDA.n251 0.0553333
R2532 VDDA.n62 VDDA.n61 0.0475
R2533 VDDA.n76 VDDA.n75 0.0475
R2534 VDDA.n92 VDDA.n91 0.0475
R2535 VDDA.n497 VDDA.n496 0.0475
R2536 VDDA.n511 VDDA.n510 0.0475
R2537 VDDA.n527 VDDA.n526 0.0475
R2538 VDDA.n130 VDDA.n129 0.0475
R2539 VDDA.n156 VDDA.n155 0.0475
R2540 VDDA.n118 VDDA.n117 0.0475
R2541 VDDA.n598 VDDA.n597 0.0475
R2542 VDDA.n586 VDDA.n585 0.0475
R2543 VDDA.n574 VDDA.n573 0.0475
R2544 VDDA.n681 VDDA.n189 0.0429747
R2545 VDDA.n769 VDDA.n178 0.0421667
R2546 VDDA.n692 VDDA.n185 0.0421667
R2547 VDDA.n634 VDDA.n210 0.0421667
R2548 VDDA.n775 VDDA.n101 0.0286392
R2549 VDDA.n608 VDDA.n536 0.0284871
R2550 VDDA.n55 VDDA.n28 0.028198
R2551 VDDA.n71 VDDA.n25 0.028198
R2552 VDDA.n85 VDDA.n22 0.028198
R2553 VDDA.n30 VDDA.n19 0.028198
R2554 VDDA.n490 VDDA.n261 0.028198
R2555 VDDA.n506 VDDA.n258 0.028198
R2556 VDDA.n520 VDDA.n255 0.028198
R2557 VDDA.n263 VDDA.n252 0.028198
R2558 VDDA.n139 VDDA.n111 0.028198
R2559 VDDA.n125 VDDA.n108 0.028198
R2560 VDDA.n163 VDDA.n105 0.028198
R2561 VDDA.n113 VDDA.n102 0.028198
R2562 VDDA.n602 VDDA.n546 0.028198
R2563 VDDA.n590 VDDA.n543 0.028198
R2564 VDDA.n578 VDDA.n540 0.028198
R2565 VDDA.n537 VDDA.n251 0.028198
R2566 VDDA.n569 VDDA.n537 0.028198
R2567 VDDA.n581 VDDA.n540 0.028198
R2568 VDDA.n593 VDDA.n543 0.028198
R2569 VDDA.n605 VDDA.n546 0.028198
R2570 VDDA.n531 VDDA.n252 0.028198
R2571 VDDA.n517 VDDA.n255 0.028198
R2572 VDDA.n501 VDDA.n258 0.028198
R2573 VDDA.n487 VDDA.n261 0.028198
R2574 VDDA.n172 VDDA.n102 0.028198
R2575 VDDA.n122 VDDA.n105 0.028198
R2576 VDDA.n148 VDDA.n108 0.028198
R2577 VDDA.n134 VDDA.n111 0.028198
R2578 VDDA.n96 VDDA.n19 0.028198
R2579 VDDA.n82 VDDA.n22 0.028198
R2580 VDDA.n66 VDDA.n25 0.028198
R2581 VDDA.n52 VDDA.n28 0.028198
R2582 VDDA.n51 VDDA.n29 0.0262697
R2583 VDDA.n61 VDDA.n27 0.0262697
R2584 VDDA.n65 VDDA.n26 0.0262697
R2585 VDDA.n75 VDDA.n24 0.0262697
R2586 VDDA.n81 VDDA.n23 0.0262697
R2587 VDDA.n91 VDDA.n21 0.0262697
R2588 VDDA.n95 VDDA.n20 0.0262697
R2589 VDDA.n496 VDDA.n260 0.0262697
R2590 VDDA.n500 VDDA.n259 0.0262697
R2591 VDDA.n510 VDDA.n257 0.0262697
R2592 VDDA.n516 VDDA.n256 0.0262697
R2593 VDDA.n526 VDDA.n254 0.0262697
R2594 VDDA.n530 VDDA.n253 0.0262697
R2595 VDDA.n133 VDDA.n112 0.0262697
R2596 VDDA.n129 VDDA.n110 0.0262697
R2597 VDDA.n147 VDDA.n109 0.0262697
R2598 VDDA.n155 VDDA.n107 0.0262697
R2599 VDDA.n121 VDDA.n106 0.0262697
R2600 VDDA.n117 VDDA.n104 0.0262697
R2601 VDDA.n171 VDDA.n103 0.0262697
R2602 VDDA.n607 VDDA.n606 0.0262697
R2603 VDDA.n598 VDDA.n545 0.0262697
R2604 VDDA.n594 VDDA.n544 0.0262697
R2605 VDDA.n586 VDDA.n542 0.0262697
R2606 VDDA.n582 VDDA.n541 0.0262697
R2607 VDDA.n574 VDDA.n539 0.0262697
R2608 VDDA.n570 VDDA.n538 0.0262697
R2609 VDDA.n573 VDDA.n538 0.0262697
R2610 VDDA.n577 VDDA.n539 0.0262697
R2611 VDDA.n585 VDDA.n541 0.0262697
R2612 VDDA.n589 VDDA.n542 0.0262697
R2613 VDDA.n597 VDDA.n544 0.0262697
R2614 VDDA.n601 VDDA.n545 0.0262697
R2615 VDDA.n527 VDDA.n253 0.0262697
R2616 VDDA.n521 VDDA.n254 0.0262697
R2617 VDDA.n511 VDDA.n256 0.0262697
R2618 VDDA.n507 VDDA.n257 0.0262697
R2619 VDDA.n497 VDDA.n259 0.0262697
R2620 VDDA.n491 VDDA.n260 0.0262697
R2621 VDDA.n118 VDDA.n103 0.0262697
R2622 VDDA.n164 VDDA.n104 0.0262697
R2623 VDDA.n156 VDDA.n106 0.0262697
R2624 VDDA.n126 VDDA.n107 0.0262697
R2625 VDDA.n130 VDDA.n109 0.0262697
R2626 VDDA.n140 VDDA.n110 0.0262697
R2627 VDDA.n92 VDDA.n20 0.0262697
R2628 VDDA.n86 VDDA.n21 0.0262697
R2629 VDDA.n76 VDDA.n23 0.0262697
R2630 VDDA.n72 VDDA.n24 0.0262697
R2631 VDDA.n62 VDDA.n26 0.0262697
R2632 VDDA.n56 VDDA.n27 0.0262697
R2633 VDDA.n479 VDDA.n275 0.0217373
R2634 VDDA.n429 VDDA.n277 0.0217373
R2635 VDDA.n352 VDDA.n279 0.0217373
R2636 VDDA.n286 VDDA.n281 0.0217373
R2637 VDDA.n290 VDDA.n289 0.0217373
R2638 VDDA.n356 VDDA.n355 0.0217373
R2639 VDDA.n433 VDDA.n432 0.0217373
R2640 VDDA.n483 VDDA.n482 0.0217373
R2641 VDDA.n288 VDDA.n281 0.0217373
R2642 VDDA.n291 VDDA.n290 0.0217373
R2643 VDDA.n354 VDDA.n279 0.0217373
R2644 VDDA.n357 VDDA.n356 0.0217373
R2645 VDDA.n431 VDDA.n277 0.0217373
R2646 VDDA.n434 VDDA.n433 0.0217373
R2647 VDDA.n481 VDDA.n275 0.0217373
R2648 VDDA.n484 VDDA.n483 0.0217373
R2649 VDDA.n664 VDDA.n663 0.0217373
R2650 VDDA.n660 VDDA.n652 0.0217373
R2651 VDDA.n674 VDDA.n650 0.0217373
R2652 VDDA.n665 VDDA.n651 0.0217373
R2653 VDDA.n679 VDDA.n649 0.0217373
R2654 VDDA.n683 VDDA.n189 0.0217373
R2655 VDDA.n678 VDDA.n650 0.0217373
R2656 VDDA.n676 VDDA.n649 0.0217373
R2657 VDDA.n674 VDDA.n673 0.0217373
R2658 VDDA.n664 VDDA.n652 0.0217373
R2659 VDDA.n661 VDDA.n651 0.0217373
R2660 VDDA.n733 VDDA.n721 0.0217373
R2661 VDDA.n744 VDDA.n738 0.0217373
R2662 VDDA.n771 VDDA.n770 0.0217373
R2663 VDDA.n768 VDDA.n179 0.0217373
R2664 VDDA.n752 VDDA.n182 0.0217373
R2665 VDDA.n770 VDDA.n177 0.0217373
R2666 VDDA.n179 VDDA.n177 0.0217373
R2667 VDDA.n709 VDDA.n708 0.0217373
R2668 VDDA.n712 VDDA.n184 0.0217373
R2669 VDDA.n748 VDDA.n183 0.0217373
R2670 VDDA.n736 VDDA.n715 0.0217373
R2671 VDDA.n720 VDDA.n718 0.0217373
R2672 VDDA.n713 VDDA.n182 0.0217373
R2673 VDDA.n748 VDDA.n747 0.0217373
R2674 VDDA.n738 VDDA.n716 0.0217373
R2675 VDDA.n737 VDDA.n736 0.0217373
R2676 VDDA.n721 VDDA.n719 0.0217373
R2677 VDDA.n642 VDDA.n190 0.0217373
R2678 VDDA.n708 VDDA.n691 0.0217373
R2679 VDDA.n691 VDDA.n184 0.0217373
R2680 VDDA.n681 VDDA.n680 0.0217373
R2681 VDDA.n638 VDDA.n191 0.0217373
R2682 VDDA.n636 VDDA.n635 0.0217373
R2683 VDDA.n633 VDDA.n211 0.0217373
R2684 VDDA.n240 VDDA.n213 0.0217373
R2685 VDDA.n230 VDDA.n216 0.0217373
R2686 VDDA.n207 VDDA.n190 0.0217373
R2687 VDDA.n638 VDDA.n637 0.0217373
R2688 VDDA.n242 VDDA.n214 0.0217373
R2689 VDDA.n241 VDDA.n240 0.0217373
R2690 VDDA.n231 VDDA.n217 0.0217373
R2691 VDDA.n617 VDDA.n247 0.0217373
R2692 VDDA.n635 VDDA.n209 0.0217373
R2693 VDDA.n211 VDDA.n209 0.0217373
R2694 VDDA.n613 VDDA.n248 0.0217373
R2695 VDDA.n612 VDDA.n247 0.0217373
R2696 VDDA.n481 VDDA.n276 0.0217373
R2697 VDDA.n431 VDDA.n278 0.0217373
R2698 VDDA.n354 VDDA.n280 0.0217373
R2699 VDDA.n288 VDDA.n282 0.0217373
R2700 VDDA.n289 VDDA.n287 0.0217373
R2701 VDDA.n355 VDDA.n353 0.0217373
R2702 VDDA.n432 VDDA.n430 0.0217373
R2703 VDDA.n482 VDDA.n480 0.0217373
R2704 VDDA.n353 VDDA.n292 0.0217373
R2705 VDDA.n430 VDDA.n358 0.0217373
R2706 VDDA.n480 VDDA.n435 0.0217373
R2707 VDDA.n217 VDDA.n215 0.0217373
R2708 VDDA.n214 VDDA.n212 0.0217373
R2709 VDDA.n677 VDDA.n675 0.0217373
R2710 VDDA.n677 VDDA.n676 0.0217373
R2711 VDDA.n662 VDDA.n661 0.0217373
R2712 VDDA.n719 VDDA.n717 0.0217373
R2713 VDDA.n716 VDDA.n714 0.0217373
R2714 VDDA.n749 VDDA.n713 0.0217373
R2715 VDDA.n767 VDDA.n176 0.0217373
R2716 VDDA.n178 VDDA.n176 0.0217373
R2717 VDDA.n751 VDDA.n183 0.0217373
R2718 VDDA.n745 VDDA.n715 0.0217373
R2719 VDDA.n734 VDDA.n718 0.0217373
R2720 VDDA.n751 VDDA.n750 0.0217373
R2721 VDDA.n746 VDDA.n745 0.0217373
R2722 VDDA.n735 VDDA.n734 0.0217373
R2723 VDDA.n639 VDDA.n207 0.0217373
R2724 VDDA.n711 VDDA.n710 0.0217373
R2725 VDDA.n710 VDDA.n692 0.0217373
R2726 VDDA.n641 VDDA.n191 0.0217373
R2727 VDDA.n243 VDDA.n213 0.0217373
R2728 VDDA.n232 VDDA.n216 0.0217373
R2729 VDDA.n641 VDDA.n640 0.0217373
R2730 VDDA.n244 VDDA.n243 0.0217373
R2731 VDDA.n239 VDDA.n212 0.0217373
R2732 VDDA.n233 VDDA.n232 0.0217373
R2733 VDDA.n229 VDDA.n215 0.0217373
R2734 VDDA.n614 VDDA.n612 0.0217373
R2735 VDDA.n632 VDDA.n208 0.0217373
R2736 VDDA.n210 VDDA.n208 0.0217373
R2737 VDDA.n616 VDDA.n248 0.0217373
R2738 VDDA.n616 VDDA.n615 0.0217373
R2739 VDDA VDDA.n890 0.0164359
R2740 VDDA.n889 VDDA.n792 0.00186893
R2741 VDDA.n792 VDDA.n18 0.00186893
R2742 VDDA.n842 VDDA.n841 0.00168433
R2743 VDDA.n842 VDDA.n1 0.00168433
R2744 VDDA.n886 VDDA.n843 0.00168433
R2745 VDDA.n843 VDDA.n2 0.00168433
R2746 VDDA.n884 VDDA.n844 0.00168433
R2747 VDDA.n844 VDDA.n3 0.00168433
R2748 VDDA.n882 VDDA.n845 0.00168433
R2749 VDDA.n845 VDDA.n4 0.00168433
R2750 VDDA.n880 VDDA.n846 0.00168433
R2751 VDDA.n846 VDDA.n5 0.00168433
R2752 VDDA.n878 VDDA.n847 0.00168433
R2753 VDDA.n847 VDDA.n6 0.00168433
R2754 VDDA.n876 VDDA.n848 0.00168433
R2755 VDDA.n848 VDDA.n7 0.00168433
R2756 VDDA.n874 VDDA.n849 0.00168433
R2757 VDDA.n849 VDDA.n8 0.00168433
R2758 VDDA.n872 VDDA.n850 0.00168433
R2759 VDDA.n850 VDDA.n9 0.00168433
R2760 VDDA.n870 VDDA.n851 0.00168433
R2761 VDDA.n851 VDDA.n10 0.00168433
R2762 VDDA.n868 VDDA.n852 0.00168433
R2763 VDDA.n852 VDDA.n11 0.00168433
R2764 VDDA.n866 VDDA.n853 0.00168433
R2765 VDDA.n853 VDDA.n12 0.00168433
R2766 VDDA.n864 VDDA.n854 0.00168433
R2767 VDDA.n854 VDDA.n13 0.00168433
R2768 VDDA.n862 VDDA.n855 0.00168433
R2769 VDDA.n855 VDDA.n14 0.00168433
R2770 VDDA.n860 VDDA.n856 0.00168433
R2771 VDDA.n856 VDDA.n15 0.00168433
R2772 VDDA.n858 VDDA.n16 0.00168433
R2773 VDDA.n857 VDDA.n17 0.00168433
R2774 VDDA.n859 VDDA.n15 0.00168433
R2775 VDDA.n861 VDDA.n14 0.00168433
R2776 VDDA.n863 VDDA.n13 0.00168433
R2777 VDDA.n865 VDDA.n12 0.00168433
R2778 VDDA.n867 VDDA.n11 0.00168433
R2779 VDDA.n869 VDDA.n10 0.00168433
R2780 VDDA.n871 VDDA.n9 0.00168433
R2781 VDDA.n873 VDDA.n8 0.00168433
R2782 VDDA.n875 VDDA.n7 0.00168433
R2783 VDDA.n877 VDDA.n6 0.00168433
R2784 VDDA.n879 VDDA.n5 0.00168433
R2785 VDDA.n881 VDDA.n4 0.00168433
R2786 VDDA.n883 VDDA.n3 0.00168433
R2787 VDDA.n885 VDDA.n2 0.00168433
R2788 VDDA.n887 VDDA.n1 0.00168433
R2789 VDDA.n859 VDDA.n858 0.00168433
R2790 VDDA.n861 VDDA.n860 0.00168433
R2791 VDDA.n863 VDDA.n862 0.00168433
R2792 VDDA.n865 VDDA.n864 0.00168433
R2793 VDDA.n867 VDDA.n866 0.00168433
R2794 VDDA.n869 VDDA.n868 0.00168433
R2795 VDDA.n871 VDDA.n870 0.00168433
R2796 VDDA.n873 VDDA.n872 0.00168433
R2797 VDDA.n875 VDDA.n874 0.00168433
R2798 VDDA.n877 VDDA.n876 0.00168433
R2799 VDDA.n879 VDDA.n878 0.00168433
R2800 VDDA.n881 VDDA.n880 0.00168433
R2801 VDDA.n883 VDDA.n882 0.00168433
R2802 VDDA.n885 VDDA.n884 0.00168433
R2803 VDDA.n887 VDDA.n886 0.00168433
R2804 VDDA.n841 VDDA.n18 0.00168433
R2805 VDDA.n857 VDDA.n16 0.00168433
R2806 VDDA.n794 VDDA.n0 0.00166081
R2807 VDDA.n793 VDDA.n791 0.00166081
R2808 VDDA.n797 VDDA.n795 0.00166081
R2809 VDDA.n796 VDDA.n790 0.00166081
R2810 VDDA.n800 VDDA.n798 0.00166081
R2811 VDDA.n799 VDDA.n789 0.00166081
R2812 VDDA.n803 VDDA.n801 0.00166081
R2813 VDDA.n802 VDDA.n788 0.00166081
R2814 VDDA.n806 VDDA.n804 0.00166081
R2815 VDDA.n805 VDDA.n787 0.00166081
R2816 VDDA.n809 VDDA.n807 0.00166081
R2817 VDDA.n808 VDDA.n786 0.00166081
R2818 VDDA.n812 VDDA.n810 0.00166081
R2819 VDDA.n811 VDDA.n785 0.00166081
R2820 VDDA.n815 VDDA.n813 0.00166081
R2821 VDDA.n814 VDDA.n784 0.00166081
R2822 VDDA.n818 VDDA.n816 0.00166081
R2823 VDDA.n817 VDDA.n783 0.00166081
R2824 VDDA.n821 VDDA.n819 0.00166081
R2825 VDDA.n820 VDDA.n782 0.00166081
R2826 VDDA.n824 VDDA.n822 0.00166081
R2827 VDDA.n823 VDDA.n781 0.00166081
R2828 VDDA.n827 VDDA.n825 0.00166081
R2829 VDDA.n826 VDDA.n780 0.00166081
R2830 VDDA.n830 VDDA.n828 0.00166081
R2831 VDDA.n829 VDDA.n779 0.00166081
R2832 VDDA.n833 VDDA.n831 0.00166081
R2833 VDDA.n832 VDDA.n778 0.00166081
R2834 VDDA.n836 VDDA.n834 0.00166081
R2835 VDDA.n835 VDDA.n777 0.00166081
R2836 VDDA.n839 VDDA.n837 0.00166081
R2837 VDDA.n838 VDDA.n776 0.00166081
R2838 VDDA.n888 VDDA.n840 0.00166081
R2839 VDDA.n890 VDDA.n0 0.00166081
R2840 VDDA.n794 VDDA.n793 0.00166081
R2841 VDDA.n795 VDDA.n791 0.00166081
R2842 VDDA.n797 VDDA.n796 0.00166081
R2843 VDDA.n798 VDDA.n790 0.00166081
R2844 VDDA.n800 VDDA.n799 0.00166081
R2845 VDDA.n801 VDDA.n789 0.00166081
R2846 VDDA.n803 VDDA.n802 0.00166081
R2847 VDDA.n804 VDDA.n788 0.00166081
R2848 VDDA.n806 VDDA.n805 0.00166081
R2849 VDDA.n807 VDDA.n787 0.00166081
R2850 VDDA.n809 VDDA.n808 0.00166081
R2851 VDDA.n810 VDDA.n786 0.00166081
R2852 VDDA.n812 VDDA.n811 0.00166081
R2853 VDDA.n813 VDDA.n785 0.00166081
R2854 VDDA.n815 VDDA.n814 0.00166081
R2855 VDDA.n816 VDDA.n784 0.00166081
R2856 VDDA.n818 VDDA.n817 0.00166081
R2857 VDDA.n819 VDDA.n783 0.00166081
R2858 VDDA.n821 VDDA.n820 0.00166081
R2859 VDDA.n822 VDDA.n782 0.00166081
R2860 VDDA.n824 VDDA.n823 0.00166081
R2861 VDDA.n825 VDDA.n781 0.00166081
R2862 VDDA.n827 VDDA.n826 0.00166081
R2863 VDDA.n828 VDDA.n780 0.00166081
R2864 VDDA.n830 VDDA.n829 0.00166081
R2865 VDDA.n831 VDDA.n779 0.00166081
R2866 VDDA.n833 VDDA.n832 0.00166081
R2867 VDDA.n834 VDDA.n778 0.00166081
R2868 VDDA.n836 VDDA.n835 0.00166081
R2869 VDDA.n837 VDDA.n777 0.00166081
R2870 VDDA.n839 VDDA.n838 0.00166081
R2871 VDDA.n840 VDDA.n776 0.00166081
R2872 VDDA.t82 VDDA.n42 0.00152174
R2873 VDDA.t144 VDDA.n43 0.00152174
R2874 VDDA.t88 VDDA.n44 0.00152174
R2875 VDDA.t151 VDDA.n45 0.00152174
R2876 VDDA.t369 VDDA.n46 0.00152174
R2877 VOUT+.n197 VOUT+.t3 110.386
R2878 VOUT+.n47 VOUT+.n46 34.9935
R2879 VOUT+.n45 VOUT+.n44 34.9935
R2880 VOUT+.n59 VOUT+.n58 34.9935
R2881 VOUT+.n55 VOUT+.n54 34.9935
R2882 VOUT+.n52 VOUT+.n51 34.9935
R2883 VOUT+.n49 VOUT+.n48 34.9935
R2884 VOUT+.n2 VOUT+.n1 9.73997
R2885 VOUT+.n6 VOUT+.n5 9.73997
R2886 VOUT+.n9 VOUT+.n8 9.73997
R2887 VOUT+.n7 VOUT+.n6 6.64633
R2888 VOUT+.n7 VOUT+.n2 6.64633
R2889 VOUT+.n46 VOUT+.t0 6.56717
R2890 VOUT+.n46 VOUT+.t11 6.56717
R2891 VOUT+.n44 VOUT+.t10 6.56717
R2892 VOUT+.n44 VOUT+.t16 6.56717
R2893 VOUT+.n58 VOUT+.t5 6.56717
R2894 VOUT+.n58 VOUT+.t12 6.56717
R2895 VOUT+.n54 VOUT+.t15 6.56717
R2896 VOUT+.n54 VOUT+.t17 6.56717
R2897 VOUT+.n51 VOUT+.t6 6.56717
R2898 VOUT+.n51 VOUT+.t8 6.56717
R2899 VOUT+.n48 VOUT+.t9 6.56717
R2900 VOUT+.n48 VOUT+.t2 6.56717
R2901 VOUT+.n57 VOUT+.n45 6.3755
R2902 VOUT+.n50 VOUT+.n47 6.3755
R2903 VOUT+.n9 VOUT+.n7 6.02133
R2904 VOUT+.n59 VOUT+.n57 5.813
R2905 VOUT+.n56 VOUT+.n55 5.813
R2906 VOUT+.n53 VOUT+.n52 5.813
R2907 VOUT+.n50 VOUT+.n49 5.813
R2908 VOUT+.n60 VOUT+.n36 5.063
R2909 VOUT+.n63 VOUT+.n43 5.063
R2910 VOUT+.n134 VOUT+.t140 4.8295
R2911 VOUT+.n135 VOUT+.t50 4.8295
R2912 VOUT+.n136 VOUT+.t88 4.8295
R2913 VOUT+.n149 VOUT+.t33 4.8295
R2914 VOUT+.n151 VOUT+.t83 4.8295
R2915 VOUT+.n152 VOUT+.t71 4.8295
R2916 VOUT+.n154 VOUT+.t107 4.8295
R2917 VOUT+.n155 VOUT+.t79 4.8295
R2918 VOUT+.n157 VOUT+.t63 4.8295
R2919 VOUT+.n158 VOUT+.t38 4.8295
R2920 VOUT+.n160 VOUT+.t104 4.8295
R2921 VOUT+.n161 VOUT+.t74 4.8295
R2922 VOUT+.n163 VOUT+.t59 4.8295
R2923 VOUT+.n164 VOUT+.t27 4.8295
R2924 VOUT+.n166 VOUT+.t156 4.8295
R2925 VOUT+.n167 VOUT+.t134 4.8295
R2926 VOUT+.n169 VOUT+.t55 4.8295
R2927 VOUT+.n170 VOUT+.t21 4.8295
R2928 VOUT+.n172 VOUT+.t153 4.8295
R2929 VOUT+.n173 VOUT+.t129 4.8295
R2930 VOUT+.n175 VOUT+.t115 4.8295
R2931 VOUT+.n176 VOUT+.t95 4.8295
R2932 VOUT+.n97 VOUT+.t58 4.8295
R2933 VOUT+.n111 VOUT+.t155 4.8295
R2934 VOUT+.n113 VOUT+.t142 4.8295
R2935 VOUT+.n114 VOUT+.t117 4.8295
R2936 VOUT+.n116 VOUT+.t30 4.8295
R2937 VOUT+.n117 VOUT+.t149 4.8295
R2938 VOUT+.n119 VOUT+.t98 4.8295
R2939 VOUT+.n120 VOUT+.t102 4.8295
R2940 VOUT+.n122 VOUT+.t62 4.8295
R2941 VOUT+.n123 VOUT+.t36 4.8295
R2942 VOUT+.n125 VOUT+.t19 4.8295
R2943 VOUT+.n126 VOUT+.t147 4.8295
R2944 VOUT+.n128 VOUT+.t67 4.8295
R2945 VOUT+.n129 VOUT+.t44 4.8295
R2946 VOUT+.n131 VOUT+.t112 4.8295
R2947 VOUT+.n132 VOUT+.t86 4.8295
R2948 VOUT+.n178 VOUT+.t51 4.8295
R2949 VOUT+.n141 VOUT+.t53 4.8154
R2950 VOUT+.n140 VOUT+.t92 4.8154
R2951 VOUT+.n138 VOUT+.t108 4.8154
R2952 VOUT+.n137 VOUT+.t144 4.8154
R2953 VOUT+.n143 VOUT+.t25 4.806
R2954 VOUT+.n142 VOUT+.t152 4.806
R2955 VOUT+.n139 VOUT+.t125 4.806
R2956 VOUT+.n110 VOUT+.t60 4.806
R2957 VOUT+.n109 VOUT+.t65 4.806
R2958 VOUT+.n108 VOUT+.t109 4.806
R2959 VOUT+.n107 VOUT+.t84 4.806
R2960 VOUT+.n106 VOUT+.t122 4.806
R2961 VOUT+.n105 VOUT+.t157 4.806
R2962 VOUT+.n104 VOUT+.t138 4.806
R2963 VOUT+.n103 VOUT+.t29 4.806
R2964 VOUT+.n102 VOUT+.t70 4.806
R2965 VOUT+.n101 VOUT+.t114 4.806
R2966 VOUT+.n100 VOUT+.t93 4.806
R2967 VOUT+.n99 VOUT+.t126 4.806
R2968 VOUT+.n134 VOUT+.t121 4.5005
R2969 VOUT+.n135 VOUT+.t103 4.5005
R2970 VOUT+.n136 VOUT+.t137 4.5005
R2971 VOUT+.n137 VOUT+.t111 4.5005
R2972 VOUT+.n138 VOUT+.t68 4.5005
R2973 VOUT+.n139 VOUT+.t97 4.5005
R2974 VOUT+.n140 VOUT+.t54 4.5005
R2975 VOUT+.n141 VOUT+.t154 4.5005
R2976 VOUT+.n142 VOUT+.t119 4.5005
R2977 VOUT+.n143 VOUT+.t141 4.5005
R2978 VOUT+.n144 VOUT+.t105 4.5005
R2979 VOUT+.n145 VOUT+.t61 4.5005
R2980 VOUT+.n146 VOUT+.t89 4.5005
R2981 VOUT+.n147 VOUT+.t46 4.5005
R2982 VOUT+.n148 VOUT+.t41 4.5005
R2983 VOUT+.n150 VOUT+.t76 4.5005
R2984 VOUT+.n149 VOUT+.t145 4.5005
R2985 VOUT+.n151 VOUT+.t77 4.5005
R2986 VOUT+.n153 VOUT+.t113 4.5005
R2987 VOUT+.n152 VOUT+.t32 4.5005
R2988 VOUT+.n154 VOUT+.t78 4.5005
R2989 VOUT+.n156 VOUT+.t80 4.5005
R2990 VOUT+.n155 VOUT+.t23 4.5005
R2991 VOUT+.n157 VOUT+.t35 4.5005
R2992 VOUT+.n159 VOUT+.t37 4.5005
R2993 VOUT+.n158 VOUT+.t132 4.5005
R2994 VOUT+.n160 VOUT+.t73 4.5005
R2995 VOUT+.n162 VOUT+.t75 4.5005
R2996 VOUT+.n161 VOUT+.t160 4.5005
R2997 VOUT+.n163 VOUT+.t26 4.5005
R2998 VOUT+.n165 VOUT+.t28 4.5005
R2999 VOUT+.n164 VOUT+.t127 4.5005
R3000 VOUT+.n166 VOUT+.t133 4.5005
R3001 VOUT+.n168 VOUT+.t135 4.5005
R3002 VOUT+.n167 VOUT+.t91 4.5005
R3003 VOUT+.n169 VOUT+.t20 4.5005
R3004 VOUT+.n171 VOUT+.t22 4.5005
R3005 VOUT+.n170 VOUT+.t123 4.5005
R3006 VOUT+.n172 VOUT+.t128 4.5005
R3007 VOUT+.n174 VOUT+.t130 4.5005
R3008 VOUT+.n173 VOUT+.t82 4.5005
R3009 VOUT+.n175 VOUT+.t94 4.5005
R3010 VOUT+.n177 VOUT+.t96 4.5005
R3011 VOUT+.n176 VOUT+.t40 4.5005
R3012 VOUT+.n98 VOUT+.t99 4.5005
R3013 VOUT+.n97 VOUT+.t159 4.5005
R3014 VOUT+.n99 VOUT+.t90 4.5005
R3015 VOUT+.n100 VOUT+.t48 4.5005
R3016 VOUT+.n101 VOUT+.t69 4.5005
R3017 VOUT+.n102 VOUT+.t24 4.5005
R3018 VOUT+.n103 VOUT+.t136 4.5005
R3019 VOUT+.n104 VOUT+.t100 4.5005
R3020 VOUT+.n105 VOUT+.t120 4.5005
R3021 VOUT+.n106 VOUT+.t81 4.5005
R3022 VOUT+.n107 VOUT+.t42 4.5005
R3023 VOUT+.n108 VOUT+.t64 4.5005
R3024 VOUT+.n109 VOUT+.t161 4.5005
R3025 VOUT+.n110 VOUT+.t158 4.5005
R3026 VOUT+.n112 VOUT+.t56 4.5005
R3027 VOUT+.n111 VOUT+.t124 4.5005
R3028 VOUT+.n113 VOUT+.t116 4.5005
R3029 VOUT+.n115 VOUT+.t118 4.5005
R3030 VOUT+.n114 VOUT+.t66 4.5005
R3031 VOUT+.n116 VOUT+.t150 4.5005
R3032 VOUT+.n118 VOUT+.t151 4.5005
R3033 VOUT+.n117 VOUT+.t106 4.5005
R3034 VOUT+.n119 VOUT+.t57 4.5005
R3035 VOUT+.n121 VOUT+.t110 4.5005
R3036 VOUT+.n120 VOUT+.t47 4.5005
R3037 VOUT+.n122 VOUT+.t34 4.5005
R3038 VOUT+.n124 VOUT+.t39 4.5005
R3039 VOUT+.n123 VOUT+.t131 4.5005
R3040 VOUT+.n125 VOUT+.t146 4.5005
R3041 VOUT+.n127 VOUT+.t148 4.5005
R3042 VOUT+.n126 VOUT+.t101 4.5005
R3043 VOUT+.n128 VOUT+.t43 4.5005
R3044 VOUT+.n130 VOUT+.t45 4.5005
R3045 VOUT+.n129 VOUT+.t139 4.5005
R3046 VOUT+.n131 VOUT+.t85 4.5005
R3047 VOUT+.n133 VOUT+.t87 4.5005
R3048 VOUT+.n132 VOUT+.t31 4.5005
R3049 VOUT+.n180 VOUT+.t49 4.5005
R3050 VOUT+.n179 VOUT+.t52 4.5005
R3051 VOUT+.n178 VOUT+.t143 4.5005
R3052 VOUT+.n181 VOUT+.t72 4.5005
R3053 VOUT+.n60 VOUT+.n37 4.5005
R3054 VOUT+.n61 VOUT+.n40 4.5005
R3055 VOUT+.n62 VOUT+.n41 4.5005
R3056 VOUT+.n64 VOUT+.n63 4.5005
R3057 VOUT+.n87 VOUT+.n86 4.5005
R3058 VOUT+.n83 VOUT+.n80 4.5005
R3059 VOUT+.n87 VOUT+.n80 4.5005
R3060 VOUT+.n88 VOUT+.n32 4.5005
R3061 VOUT+.n88 VOUT+.n34 4.5005
R3062 VOUT+.n88 VOUT+.n87 4.5005
R3063 VOUT+.n186 VOUT+.n91 4.5005
R3064 VOUT+.n187 VOUT+.n186 4.5005
R3065 VOUT+.n187 VOUT+.n28 4.5005
R3066 VOUT+.n188 VOUT+.n27 4.5005
R3067 VOUT+.n188 VOUT+.n187 4.5005
R3068 VOUT+.n192 VOUT+.n191 4.5005
R3069 VOUT+.n191 VOUT+.n19 4.5005
R3070 VOUT+.n22 VOUT+.n19 4.5005
R3071 VOUT+.n194 VOUT+.n19 4.5005
R3072 VOUT+.n196 VOUT+.n19 4.5005
R3073 VOUT+.n195 VOUT+.n22 4.5005
R3074 VOUT+.n195 VOUT+.n194 4.5005
R3075 VOUT+.n196 VOUT+.n195 4.5005
R3076 VOUT+.n1 VOUT+.t7 3.42907
R3077 VOUT+.n1 VOUT+.t18 3.42907
R3078 VOUT+.n5 VOUT+.t14 3.42907
R3079 VOUT+.n5 VOUT+.t1 3.42907
R3080 VOUT+.n8 VOUT+.t13 3.42907
R3081 VOUT+.n8 VOUT+.t4 3.42907
R3082 VOUT+.n85 VOUT+.n33 2.26725
R3083 VOUT+.n81 VOUT+.n31 2.24601
R3084 VOUT+.n190 VOUT+.n189 2.24601
R3085 VOUT+.n24 VOUT+.n21 2.24601
R3086 VOUT+.n185 VOUT+.n184 2.24477
R3087 VOUT+.n30 VOUT+.n25 2.24477
R3088 VOUT+.n88 VOUT+.n33 2.24063
R3089 VOUT+.n188 VOUT+.n26 2.24063
R3090 VOUT+.n195 VOUT+.n23 2.24063
R3091 VOUT+.n80 VOUT+.n79 2.24063
R3092 VOUT+.n186 VOUT+.n89 2.24063
R3093 VOUT+.n90 VOUT+.n28 2.24063
R3094 VOUT+.n193 VOUT+.n192 2.24063
R3095 VOUT+.n192 VOUT+.n20 2.24063
R3096 VOUT+.n86 VOUT+.n84 2.23934
R3097 VOUT+.n86 VOUT+.n82 2.23934
R3098 VOUT+.n6 VOUT+.n4 1.83719
R3099 VOUT+.n10 VOUT+.n9 1.72967
R3100 VOUT+.n17 VOUT+.n2 1.72967
R3101 VOUT+.n78 VOUT+.n77 1.5005
R3102 VOUT+.n76 VOUT+.n35 1.5005
R3103 VOUT+.n75 VOUT+.n74 1.5005
R3104 VOUT+.n73 VOUT+.n38 1.5005
R3105 VOUT+.n72 VOUT+.n71 1.5005
R3106 VOUT+.n70 VOUT+.n39 1.5005
R3107 VOUT+.n69 VOUT+.n68 1.5005
R3108 VOUT+.n67 VOUT+.n42 1.5005
R3109 VOUT+.n18 VOUT+.n17 1.5005
R3110 VOUT+.n16 VOUT+.n0 1.5005
R3111 VOUT+.n15 VOUT+.n14 1.5005
R3112 VOUT+.n13 VOUT+.n3 1.5005
R3113 VOUT+.n12 VOUT+.n11 1.5005
R3114 VOUT+.n64 VOUT+.n59 1.313
R3115 VOUT+.n55 VOUT+.n41 1.313
R3116 VOUT+.n52 VOUT+.n40 1.313
R3117 VOUT+.n49 VOUT+.n37 1.313
R3118 VOUT+.n45 VOUT+.n43 1.313
R3119 VOUT+.n47 VOUT+.n36 1.313
R3120 VOUT+.n187 VOUT+.n29 1.1455
R3121 VOUT+.n95 VOUT+.n94 1.13717
R3122 VOUT+.n96 VOUT+.n92 1.13717
R3123 VOUT+.n183 VOUT+.n182 1.13717
R3124 VOUT+.n93 VOUT+.n30 1.13717
R3125 VOUT+.n94 VOUT+.n27 1.13717
R3126 VOUT+.n92 VOUT+.n91 1.13717
R3127 VOUT+.n184 VOUT+.n183 1.13717
R3128 VOUT+.n87 VOUT+.n78 0.859875
R3129 VOUT+.n66 VOUT+.n43 0.715216
R3130 VOUT+.n65 VOUT+.n64 0.65675
R3131 VOUT+.n69 VOUT+.n41 0.65675
R3132 VOUT+.n71 VOUT+.n40 0.65675
R3133 VOUT+.n75 VOUT+.n37 0.65675
R3134 VOUT+.n77 VOUT+.n36 0.65675
R3135 VOUT+.n95 VOUT+.n29 0.585
R3136 VOUT+.n67 VOUT+.n66 0.564601
R3137 VOUT+.n61 VOUT+.n60 0.563
R3138 VOUT+.n62 VOUT+.n61 0.563
R3139 VOUT+.n63 VOUT+.n62 0.563
R3140 VOUT+.n57 VOUT+.n56 0.563
R3141 VOUT+.n56 VOUT+.n53 0.563
R3142 VOUT+.n53 VOUT+.n50 0.563
R3143 VOUT+.n197 VOUT+.n196 0.557792
R3144 VOUT+.n192 VOUT+.n188 0.5455
R3145 VOUT+.n138 VOUT+.n137 0.3295
R3146 VOUT+.n139 VOUT+.n138 0.3295
R3147 VOUT+.n140 VOUT+.n139 0.3295
R3148 VOUT+.n141 VOUT+.n140 0.3295
R3149 VOUT+.n142 VOUT+.n141 0.3295
R3150 VOUT+.n143 VOUT+.n142 0.3295
R3151 VOUT+.n144 VOUT+.n143 0.3295
R3152 VOUT+.n145 VOUT+.n144 0.3295
R3153 VOUT+.n146 VOUT+.n145 0.3295
R3154 VOUT+.n147 VOUT+.n146 0.3295
R3155 VOUT+.n148 VOUT+.n147 0.3295
R3156 VOUT+.n150 VOUT+.n148 0.3295
R3157 VOUT+.n150 VOUT+.n149 0.3295
R3158 VOUT+.n153 VOUT+.n151 0.3295
R3159 VOUT+.n153 VOUT+.n152 0.3295
R3160 VOUT+.n156 VOUT+.n154 0.3295
R3161 VOUT+.n156 VOUT+.n155 0.3295
R3162 VOUT+.n159 VOUT+.n157 0.3295
R3163 VOUT+.n159 VOUT+.n158 0.3295
R3164 VOUT+.n162 VOUT+.n160 0.3295
R3165 VOUT+.n162 VOUT+.n161 0.3295
R3166 VOUT+.n165 VOUT+.n163 0.3295
R3167 VOUT+.n165 VOUT+.n164 0.3295
R3168 VOUT+.n168 VOUT+.n166 0.3295
R3169 VOUT+.n168 VOUT+.n167 0.3295
R3170 VOUT+.n171 VOUT+.n169 0.3295
R3171 VOUT+.n171 VOUT+.n170 0.3295
R3172 VOUT+.n174 VOUT+.n172 0.3295
R3173 VOUT+.n174 VOUT+.n173 0.3295
R3174 VOUT+.n177 VOUT+.n175 0.3295
R3175 VOUT+.n177 VOUT+.n176 0.3295
R3176 VOUT+.n98 VOUT+.n97 0.3295
R3177 VOUT+.n100 VOUT+.n99 0.3295
R3178 VOUT+.n101 VOUT+.n100 0.3295
R3179 VOUT+.n102 VOUT+.n101 0.3295
R3180 VOUT+.n103 VOUT+.n102 0.3295
R3181 VOUT+.n104 VOUT+.n103 0.3295
R3182 VOUT+.n105 VOUT+.n104 0.3295
R3183 VOUT+.n106 VOUT+.n105 0.3295
R3184 VOUT+.n107 VOUT+.n106 0.3295
R3185 VOUT+.n108 VOUT+.n107 0.3295
R3186 VOUT+.n109 VOUT+.n108 0.3295
R3187 VOUT+.n110 VOUT+.n109 0.3295
R3188 VOUT+.n112 VOUT+.n110 0.3295
R3189 VOUT+.n112 VOUT+.n111 0.3295
R3190 VOUT+.n115 VOUT+.n113 0.3295
R3191 VOUT+.n115 VOUT+.n114 0.3295
R3192 VOUT+.n118 VOUT+.n116 0.3295
R3193 VOUT+.n118 VOUT+.n117 0.3295
R3194 VOUT+.n121 VOUT+.n119 0.3295
R3195 VOUT+.n121 VOUT+.n120 0.3295
R3196 VOUT+.n124 VOUT+.n122 0.3295
R3197 VOUT+.n124 VOUT+.n123 0.3295
R3198 VOUT+.n127 VOUT+.n125 0.3295
R3199 VOUT+.n127 VOUT+.n126 0.3295
R3200 VOUT+.n130 VOUT+.n128 0.3295
R3201 VOUT+.n130 VOUT+.n129 0.3295
R3202 VOUT+.n133 VOUT+.n131 0.3295
R3203 VOUT+.n133 VOUT+.n132 0.3295
R3204 VOUT+.n180 VOUT+.n179 0.3295
R3205 VOUT+.n179 VOUT+.n178 0.3295
R3206 VOUT+.n12 VOUT+.n4 0.314966
R3207 VOUT+.n181 VOUT+.n180 0.313833
R3208 VOUT+.n146 VOUT+.n134 0.306
R3209 VOUT+.n145 VOUT+.n135 0.306
R3210 VOUT+.n144 VOUT+.n136 0.306
R3211 VOUT+.n153 VOUT+.n150 0.2825
R3212 VOUT+.n156 VOUT+.n153 0.2825
R3213 VOUT+.n159 VOUT+.n156 0.2825
R3214 VOUT+.n162 VOUT+.n159 0.2825
R3215 VOUT+.n165 VOUT+.n162 0.2825
R3216 VOUT+.n168 VOUT+.n165 0.2825
R3217 VOUT+.n171 VOUT+.n168 0.2825
R3218 VOUT+.n174 VOUT+.n171 0.2825
R3219 VOUT+.n177 VOUT+.n174 0.2825
R3220 VOUT+.n112 VOUT+.n98 0.2825
R3221 VOUT+.n115 VOUT+.n112 0.2825
R3222 VOUT+.n118 VOUT+.n115 0.2825
R3223 VOUT+.n121 VOUT+.n118 0.2825
R3224 VOUT+.n124 VOUT+.n121 0.2825
R3225 VOUT+.n127 VOUT+.n124 0.2825
R3226 VOUT+.n130 VOUT+.n127 0.2825
R3227 VOUT+.n133 VOUT+.n130 0.2825
R3228 VOUT+.n179 VOUT+.n133 0.2825
R3229 VOUT+.n179 VOUT+.n177 0.2825
R3230 VOUT+.n186 VOUT+.n88 0.2455
R3231 VOUT+ VOUT+.n197 0.198417
R3232 VOUT+ VOUT+.n18 0.182792
R3233 VOUT+.n182 VOUT+.n181 0.138367
R3234 VOUT+.n10 VOUT+.n4 0.0891864
R3235 VOUT+.n65 VOUT+.n42 0.0577917
R3236 VOUT+.n69 VOUT+.n42 0.0577917
R3237 VOUT+.n70 VOUT+.n69 0.0577917
R3238 VOUT+.n71 VOUT+.n70 0.0577917
R3239 VOUT+.n71 VOUT+.n38 0.0577917
R3240 VOUT+.n75 VOUT+.n38 0.0577917
R3241 VOUT+.n76 VOUT+.n75 0.0577917
R3242 VOUT+.n77 VOUT+.n76 0.0577917
R3243 VOUT+.n68 VOUT+.n67 0.0577917
R3244 VOUT+.n68 VOUT+.n39 0.0577917
R3245 VOUT+.n72 VOUT+.n39 0.0577917
R3246 VOUT+.n73 VOUT+.n72 0.0577917
R3247 VOUT+.n74 VOUT+.n73 0.0577917
R3248 VOUT+.n74 VOUT+.n35 0.0577917
R3249 VOUT+.n78 VOUT+.n35 0.0577917
R3250 VOUT+.n66 VOUT+.n65 0.054517
R3251 VOUT+.n194 VOUT+.n24 0.047375
R3252 VOUT+.n189 VOUT+.n22 0.047375
R3253 VOUT+.n187 VOUT+.n30 0.0421667
R3254 VOUT+.n87 VOUT+.n81 0.0421667
R3255 VOUT+.n11 VOUT+.n10 0.0421667
R3256 VOUT+.n11 VOUT+.n3 0.0421667
R3257 VOUT+.n15 VOUT+.n3 0.0421667
R3258 VOUT+.n16 VOUT+.n15 0.0421667
R3259 VOUT+.n17 VOUT+.n16 0.0421667
R3260 VOUT+.n13 VOUT+.n12 0.0421667
R3261 VOUT+.n14 VOUT+.n13 0.0421667
R3262 VOUT+.n14 VOUT+.n0 0.0421667
R3263 VOUT+.n18 VOUT+.n0 0.0421667
R3264 VOUT+.n82 VOUT+.n81 0.0243161
R3265 VOUT+.n84 VOUT+.n32 0.0243161
R3266 VOUT+.n84 VOUT+.n83 0.0243161
R3267 VOUT+.n82 VOUT+.n34 0.0243161
R3268 VOUT+.n184 VOUT+.n26 0.0217373
R3269 VOUT+.n83 VOUT+.n33 0.0217373
R3270 VOUT+.n91 VOUT+.n26 0.0217373
R3271 VOUT+.n191 VOUT+.n23 0.0217373
R3272 VOUT+.n189 VOUT+.n23 0.0217373
R3273 VOUT+.n89 VOUT+.n30 0.0217373
R3274 VOUT+.n91 VOUT+.n90 0.0217373
R3275 VOUT+.n79 VOUT+.n32 0.0217373
R3276 VOUT+.n79 VOUT+.n34 0.0217373
R3277 VOUT+.n89 VOUT+.n27 0.0217373
R3278 VOUT+.n90 VOUT+.n27 0.0217373
R3279 VOUT+.n196 VOUT+.n20 0.0217373
R3280 VOUT+.n194 VOUT+.n193 0.0217373
R3281 VOUT+.n193 VOUT+.n22 0.0217373
R3282 VOUT+.n24 VOUT+.n20 0.0217373
R3283 VOUT+.n96 VOUT+.n95 0.0161667
R3284 VOUT+.n182 VOUT+.n96 0.0161667
R3285 VOUT+.n94 VOUT+.n93 0.0161667
R3286 VOUT+.n94 VOUT+.n92 0.0161667
R3287 VOUT+.n183 VOUT+.n92 0.0161667
R3288 VOUT+.n185 VOUT+.n28 0.0134654
R3289 VOUT+.n188 VOUT+.n25 0.0134654
R3290 VOUT+.n186 VOUT+.n185 0.0134654
R3291 VOUT+.n28 VOUT+.n25 0.0134654
R3292 VOUT+.n85 VOUT+.n80 0.0109778
R3293 VOUT+.n88 VOUT+.n31 0.0109778
R3294 VOUT+.n190 VOUT+.n19 0.0109778
R3295 VOUT+.n195 VOUT+.n21 0.0109778
R3296 VOUT+.n86 VOUT+.n85 0.0109778
R3297 VOUT+.n80 VOUT+.n31 0.0109778
R3298 VOUT+.n192 VOUT+.n190 0.0109778
R3299 VOUT+.n21 VOUT+.n19 0.0109778
R3300 VOUT+.n93 VOUT+.n29 0.00872683
R3301 two_stage_opamp_dummy_magic_29_0.cap_res_Y two_stage_opamp_dummy_magic_29_0.cap_res_Y.t0 49.895
R3302 two_stage_opamp_dummy_magic_29_0.cap_res_Y two_stage_opamp_dummy_magic_29_0.cap_res_Y.t74 0.9405
R3303 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t17 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t129 0.1603
R3304 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t130 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t91 0.1603
R3305 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t85 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t79 0.1603
R3306 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t139 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t83 0.1603
R3307 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t84 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t55 0.1603
R3308 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t30 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t124 0.1603
R3309 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t127 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t99 0.1603
R3310 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t2 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t88 0.1603
R3311 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t89 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t58 0.1603
R3312 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t35 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t135 0.1603
R3313 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t136 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t103 0.1603
R3314 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t71 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t28 0.1603
R3315 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t29 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t6 0.1603
R3316 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t39 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t141 0.1603
R3317 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t142 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t107 0.1603
R3318 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t80 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t33 0.1603
R3319 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t34 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t9 0.1603
R3320 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t122 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t67 0.1603
R3321 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t68 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t47 0.1603
R3322 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t19 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t111 0.1603
R3323 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t113 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t90 0.1603
R3324 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t131 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t76 0.1603
R3325 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t77 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t50 0.1603
R3326 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t23 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t118 0.1603
R3327 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t119 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t95 0.1603
R3328 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t61 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t15 0.1603
R3329 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t16 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t143 0.1603
R3330 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t31 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t126 0.1603
R3331 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t128 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t100 0.1603
R3332 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t115 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t60 0.1603
R3333 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t105 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t64 0.1603
R3334 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t56 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t13 0.1603
R3335 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t12 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t132 0.1603
R3336 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t96 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t45 0.1603
R3337 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t46 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t20 0.1603
R3338 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t38 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t7 0.1603
R3339 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t72 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t36 0.1603
R3340 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t114 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t69 0.1603
R3341 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t93 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t48 0.1603
R3342 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t138 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t92 0.1603
R3343 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t26 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t133 0.1603
R3344 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t62 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t24 0.1603
R3345 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t42 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t5 0.1603
R3346 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t81 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t40 0.1603
R3347 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t120 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t78 0.1603
R3348 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t98 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t53 0.1603
R3349 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t1 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t97 0.1603
R3350 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t4 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t102 0.1603
R3351 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t3 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t104 0.1603
R3352 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t116 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t121 0.1603
R3353 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t41 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t22 0.1603
R3354 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t73 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t41 0.1603
R3355 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t59 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t112 0.1603
R3356 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t101 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t59 0.1603
R3357 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t51 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t18 0.1603
R3358 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t94 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t54 0.1603
R3359 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t65 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t37 0.1603
R3360 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t108 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t70 0.1603
R3361 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t8 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t109 0.1603
R3362 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t43 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t10 0.1603
R3363 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t21 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t137 0.1603
R3364 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t25 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t57 0.1603
R3365 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t74 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t25 0.1603
R3366 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t106 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n17 0.159278
R3367 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t44 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n18 0.159278
R3368 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t11 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n19 0.159278
R3369 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t52 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n20 0.159278
R3370 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t123 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n21 0.159278
R3371 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t14 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n22 0.159278
R3372 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t117 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n23 0.159278
R3373 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t75 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n24 0.159278
R3374 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t110 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n25 0.159278
R3375 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t66 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n26 0.159278
R3376 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t32 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n27 0.159278
R3377 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t140 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n28 0.159278
R3378 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t27 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n29 0.159278
R3379 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t134 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n30 0.159278
R3380 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t87 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n31 0.159278
R3381 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t125 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n32 0.159278
R3382 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t82 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n33 0.159278
R3383 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t49 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n34 0.159278
R3384 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t86 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n35 0.159278
R3385 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n36 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t17 0.1368
R3386 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n35 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t130 0.1368
R3387 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n35 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t85 0.1368
R3388 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n34 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t139 0.1368
R3389 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n34 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t84 0.1368
R3390 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n33 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t30 0.1368
R3391 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n33 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t127 0.1368
R3392 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n32 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t2 0.1368
R3393 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n32 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t89 0.1368
R3394 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n31 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t35 0.1368
R3395 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n31 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t136 0.1368
R3396 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n30 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t71 0.1368
R3397 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n30 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t29 0.1368
R3398 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n29 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t39 0.1368
R3399 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n29 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t142 0.1368
R3400 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n28 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t80 0.1368
R3401 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n28 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t34 0.1368
R3402 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n27 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t122 0.1368
R3403 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n27 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t68 0.1368
R3404 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n26 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t19 0.1368
R3405 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n26 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t113 0.1368
R3406 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n25 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t131 0.1368
R3407 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n25 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t77 0.1368
R3408 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n24 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t23 0.1368
R3409 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n24 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t119 0.1368
R3410 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n23 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t61 0.1368
R3411 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n23 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t16 0.1368
R3412 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n22 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t31 0.1368
R3413 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n22 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t128 0.1368
R3414 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n21 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t115 0.1368
R3415 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n21 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t105 0.1368
R3416 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n20 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t56 0.1368
R3417 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n20 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t12 0.1368
R3418 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n19 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t96 0.1368
R3419 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n19 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t46 0.1368
R3420 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n18 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t38 0.1368
R3421 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n17 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t3 0.1368
R3422 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t121 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n36 0.1368
R3423 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n37 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t116 0.1368
R3424 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n6 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t72 0.114322
R3425 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n0 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t51 0.114322
R3426 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n7 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n6 0.1133
R3427 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n8 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n7 0.1133
R3428 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n9 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n8 0.1133
R3429 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n10 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n9 0.1133
R3430 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n11 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n10 0.1133
R3431 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n12 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n11 0.1133
R3432 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n13 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n12 0.1133
R3433 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n14 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n13 0.1133
R3434 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n15 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n14 0.1133
R3435 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n16 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n15 0.1133
R3436 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n18 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n16 0.1133
R3437 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n38 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n37 0.1133
R3438 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n1 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n0 0.1133
R3439 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n2 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n1 0.1133
R3440 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n3 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n2 0.1133
R3441 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n4 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n3 0.1133
R3442 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n5 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n4 0.1133
R3443 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n39 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n5 0.1133
R3444 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n39 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n38 0.1133
R3445 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n6 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t114 0.00152174
R3446 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n7 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t93 0.00152174
R3447 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n8 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t138 0.00152174
R3448 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n9 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t26 0.00152174
R3449 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n10 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t62 0.00152174
R3450 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n11 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t42 0.00152174
R3451 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n12 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t81 0.00152174
R3452 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n13 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t120 0.00152174
R3453 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n14 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t98 0.00152174
R3454 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n15 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t1 0.00152174
R3455 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n16 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t4 0.00152174
R3456 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n17 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t63 0.00152174
R3457 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n18 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t106 0.00152174
R3458 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n19 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t44 0.00152174
R3459 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n20 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t11 0.00152174
R3460 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n21 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t52 0.00152174
R3461 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n22 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t123 0.00152174
R3462 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n23 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t14 0.00152174
R3463 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n24 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t117 0.00152174
R3464 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n25 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t75 0.00152174
R3465 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n26 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t110 0.00152174
R3466 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n27 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t66 0.00152174
R3467 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n28 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t32 0.00152174
R3468 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n29 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t140 0.00152174
R3469 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n30 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t27 0.00152174
R3470 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n31 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t134 0.00152174
R3471 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n32 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t87 0.00152174
R3472 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n33 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t125 0.00152174
R3473 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n34 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t82 0.00152174
R3474 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n35 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t49 0.00152174
R3475 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n36 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t86 0.00152174
R3476 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n37 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t73 0.00152174
R3477 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n38 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t101 0.00152174
R3478 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n0 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t94 0.00152174
R3479 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n1 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t65 0.00152174
R3480 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n2 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t108 0.00152174
R3481 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n3 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t8 0.00152174
R3482 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n4 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t43 0.00152174
R3483 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n5 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t21 0.00152174
R3484 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t57 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n39 0.00152174
R3485 GNDA_2.n5256 GNDA_2.n130 554309
R3486 GNDA_2.n5256 GNDA_2.n131 438167
R3487 GNDA_2.n4319 GNDA_2.n1083 396244
R3488 GNDA_2.n4318 GNDA_2.n333 247185
R3489 GNDA_2.n5257 GNDA_2.n129 235669
R3490 GNDA_2.n4462 GNDA_2.n4461 215632
R3491 GNDA_2.n4319 GNDA_2.n1082 204995
R3492 GNDA_2.n4319 GNDA_2.n300 191583
R3493 GNDA_2.n4463 GNDA_2.n131 182270
R3494 GNDA_2.n4462 GNDA_2.n300 151067
R3495 GNDA_2.n5256 GNDA_2.n5255 132026
R3496 GNDA_2.n4318 GNDA_2.n4317 132026
R3497 GNDA_2.n1787 GNDA_2.n1083 105027
R3498 GNDA_2.n1790 GNDA_2.n1083 71214.8
R3499 GNDA_2.n5257 GNDA_2.n130 70780.9
R3500 GNDA_2.n4319 GNDA_2.t196 55812.1
R3501 GNDA_2.n4466 GNDA_2.n4462 52153.2
R3502 GNDA_2.t188 GNDA_2.n5256 28014.9
R3503 GNDA_2.t284 GNDA_2.n4318 28013.4
R3504 GNDA_2.n4321 GNDA_2.n333 23717.9
R3505 GNDA_2.n1081 GNDA_2.n300 21706.7
R3506 GNDA_2.n4466 GNDA_2.n4465 18170.4
R3507 GNDA_2.n3129 GNDA_2.n128 17109.1
R3508 GNDA_2.n4325 GNDA_2.n1081 16116.7
R3509 GNDA_2.n4320 GNDA_2.n1081 13566.7
R3510 GNDA_2.n1788 GNDA_2.n1082 13527.3
R3511 GNDA_2.n1789 GNDA_2.n1788 13460.8
R3512 GNDA_2.n4323 GNDA_2.n4321 13200
R3513 GNDA_2.n4326 GNDA_2.n1081 13111.6
R3514 GNDA_2.n1082 GNDA_2.n129 12640.3
R3515 GNDA_2.n4465 GNDA_2.n4464 11163
R3516 GNDA_2.n4347 GNDA_2.n301 11032
R3517 GNDA_2.n4347 GNDA_2.n334 11032
R3518 GNDA_2.n4361 GNDA_2.n334 10933.5
R3519 GNDA_2.n4361 GNDA_2.n301 10933.5
R3520 GNDA_2.n4460 GNDA_2.n303 10884.2
R3521 GNDA_2.n4404 GNDA_2.n303 10884.2
R3522 GNDA_2.n4404 GNDA_2.n302 10441
R3523 GNDA_2.n4460 GNDA_2.n302 10441
R3524 GNDA_2.n4321 GNDA_2.n4320 10046.7
R3525 GNDA_2.n4335 GNDA_2.n383 9850
R3526 GNDA_2.n4335 GNDA_2.n382 9751.5
R3527 GNDA_2.n1791 GNDA_2.n1790 9511.11
R3528 GNDA_2.n1791 GNDA_2.n129 9423.88
R3529 GNDA_2.n4344 GNDA_2.n383 9406.75
R3530 GNDA_2.n4344 GNDA_2.n382 9308.25
R3531 GNDA_2.n4407 GNDA_2.n4406 7292.48
R3532 GNDA_2.n3394 GNDA_2.n3393 7286.54
R3533 GNDA_2.n4463 GNDA_2.n130 6794.03
R3534 GNDA_2.n4464 GNDA_2.n4463 6475.77
R3535 GNDA_2.n4328 GNDA_2.n1078 5910
R3536 GNDA_2.n4465 GNDA_2.n131 5681.89
R3537 GNDA_2.n4332 GNDA_2.n1078 5466.75
R3538 GNDA_2.n4328 GNDA_2.n1077 5319
R3539 GNDA_2.n4332 GNDA_2.n1077 4875.75
R3540 GNDA_2.n1787 GNDA_2.n1084 4738.46
R3541 GNDA_2.n4319 GNDA_2.n1084 4538.62
R3542 GNDA_2.n4320 GNDA_2.n4319 4538.62
R3543 GNDA_2.n4363 GNDA_2.n4362 4375.56
R3544 GNDA_2.n1790 GNDA_2.n1789 4106.67
R3545 GNDA_2.t73 GNDA_2.n1791 4106.67
R3546 GNDA_2.n4368 GNDA_2.n347 3841.5
R3547 GNDA_2.n4370 GNDA_2.n347 3841.5
R3548 GNDA_2.n4368 GNDA_2.n348 3743
R3549 GNDA_2.n4370 GNDA_2.n348 3743
R3550 GNDA_2.n1677 GNDA_2.n1676 1684.55
R3551 GNDA_2.n4346 GNDA_2.n4345 1417.78
R3552 GNDA_2.n4334 GNDA_2.t6 1417.78
R3553 GNDA_2.t52 GNDA_2.n347 1319.17
R3554 GNDA_2.n3084 GNDA_2.n3077 1214.72
R3555 GNDA_2.n3112 GNDA_2.n3084 1214.72
R3556 GNDA_2.n3112 GNDA_2.n3111 1214.72
R3557 GNDA_2.n3111 GNDA_2.n3110 1214.72
R3558 GNDA_2.n3110 GNDA_2.n3087 1214.72
R3559 GNDA_2.n3104 GNDA_2.n3103 1214.72
R3560 GNDA_2.n3103 GNDA_2.n3102 1214.72
R3561 GNDA_2.n3102 GNDA_2.n3095 1214.72
R3562 GNDA_2.n3095 GNDA_2.n114 1214.72
R3563 GNDA_2.n5357 GNDA_2.n114 1214.72
R3564 GNDA_2.n3216 GNDA_2.n3215 1214.72
R3565 GNDA_2.n3215 GNDA_2.n3214 1214.72
R3566 GNDA_2.n3214 GNDA_2.n3183 1214.72
R3567 GNDA_2.n3208 GNDA_2.n3183 1214.72
R3568 GNDA_2.n3208 GNDA_2.n3207 1214.72
R3569 GNDA_2.n3204 GNDA_2.n3191 1214.72
R3570 GNDA_2.n3196 GNDA_2.n3191 1214.72
R3571 GNDA_2.n3197 GNDA_2.n3196 1214.72
R3572 GNDA_2.n3197 GNDA_2.n87 1214.72
R3573 GNDA_2.n5457 GNDA_2.n87 1214.72
R3574 GNDA_2.n4345 GNDA_2.t6 1148.89
R3575 GNDA_2.n4365 GNDA_2.n4364 1100
R3576 GNDA_2.n4369 GNDA_2.n4365 1075.56
R3577 GNDA_2.n4346 GNDA_2.t24 1075.56
R3578 GNDA_2.n4334 GNDA_2.n4333 1075.56
R3579 GNDA_2.n4464 GNDA_2.n4462 1068.57
R3580 GNDA_2.n4406 GNDA_2.n333 1038.4
R3581 GNDA_2.n1789 GNDA_2.n1787 1031.25
R3582 GNDA_2.n4362 GNDA_2.t24 1026.67
R3583 GNDA_2.t3 GNDA_2.n4363 1002.22
R3584 GNDA_2.t256 GNDA_2.n1080 855.557
R3585 GNDA_2.n1788 GNDA_2.n1084 854.477
R3586 GNDA_2.n3087 GNDA_2.t73 823.313
R3587 GNDA_2.n3207 GNDA_2.t73 823.313
R3588 GNDA_2.n4364 GNDA_2.t3 782.222
R3589 GNDA_2.n4333 GNDA_2.t106 782.222
R3590 GNDA_2.n5253 GNDA_2.t124 749.742
R3591 GNDA_2.n4467 GNDA_2.t108 749.742
R3592 GNDA_2.n4315 GNDA_2.t92 749.742
R3593 GNDA_2.n4409 GNDA_2.t100 747.734
R3594 GNDA_2.n2367 GNDA_2.t73 741.376
R3595 GNDA_2.n3381 GNDA_2.n3380 686.717
R3596 GNDA_2.n2839 GNDA_2.n2838 686.717
R3597 GNDA_2.n2831 GNDA_2.n2657 686.717
R3598 GNDA_2.n3372 GNDA_2.n1688 686.717
R3599 GNDA_2.n4360 GNDA_2.n4359 678.4
R3600 GNDA_2.n4360 GNDA_2.n349 678.4
R3601 GNDA_2.n4402 GNDA_2.n338 675.201
R3602 GNDA_2.n338 GNDA_2.n305 675.201
R3603 GNDA_2.n2206 GNDA_2.t16 671.187
R3604 GNDA_2.n2817 GNDA_2.n2816 669.307
R3605 GNDA_2.n2698 GNDA_2.n2697 669.307
R3606 GNDA_2.n569 GNDA_2.t120 659.367
R3607 GNDA_2.n568 GNDA_2.t149 659.367
R3608 GNDA_2.n343 GNDA_2.t103 659.367
R3609 GNDA_2.n4373 GNDA_2.t70 659.367
R3610 GNDA_2.n3066 GNDA_2.n2970 654.447
R3611 GNDA_2.n335 GNDA_2.n304 646.4
R3612 GNDA_2.n336 GNDA_2.n335 646.4
R3613 GNDA_2.n4343 GNDA_2.n4342 611.201
R3614 GNDA_2.n4343 GNDA_2.n384 604.801
R3615 GNDA_2.n2924 GNDA_2.n2923 585.001
R3616 GNDA_2.n2617 GNDA_2.n2616 585.001
R3617 GNDA_2.n1803 GNDA_2.n1802 585.001
R3618 GNDA_2.n2701 GNDA_2.n2700 585.001
R3619 GNDA_2.n2814 GNDA_2.n2813 585.001
R3620 GNDA_2.n1799 GNDA_2.n1798 585.001
R3621 GNDA_2.n3404 GNDA_2.n3403 585.001
R3622 GNDA_2.n1832 GNDA_2.n1831 585.001
R3623 GNDA_2.n3392 GNDA_2.n3391 585
R3624 GNDA_2.n3393 GNDA_2.n3392 585
R3625 GNDA_2.n3389 GNDA_2.n1678 585
R3626 GNDA_2.n1678 GNDA_2.n1677 585
R3627 GNDA_2.n1675 GNDA_2.n1674 585
R3628 GNDA_2.n2349 GNDA_2.n1673 585
R3629 GNDA_2.n2350 GNDA_2.n2349 585
R3630 GNDA_2.n2347 GNDA_2.n2346 585
R3631 GNDA_2.n2351 GNDA_2.n2347 585
R3632 GNDA_2.n2354 GNDA_2.n2353 585
R3633 GNDA_2.n2353 GNDA_2.n2352 585
R3634 GNDA_2.n2355 GNDA_2.n2345 585
R3635 GNDA_2.n2348 GNDA_2.n2345 585
R3636 GNDA_2.n2357 GNDA_2.n2356 585
R3637 GNDA_2.n2357 GNDA_2.n1691 585
R3638 GNDA_2.n2358 GNDA_2.n2344 585
R3639 GNDA_2.n2358 GNDA_2.n1690 585
R3640 GNDA_2.n2361 GNDA_2.n2360 585
R3641 GNDA_2.n2360 GNDA_2.n2359 585
R3642 GNDA_2.n2362 GNDA_2.n2342 585
R3643 GNDA_2.n2342 GNDA_2.n2341 585
R3644 GNDA_2.n2364 GNDA_2.n2363 585
R3645 GNDA_2.n2365 GNDA_2.n2364 585
R3646 GNDA_2.n2343 GNDA_2.n2340 585
R3647 GNDA_2.n2366 GNDA_2.n2340 585
R3648 GNDA_2.n2368 GNDA_2.n2338 585
R3649 GNDA_2.n2368 GNDA_2.n2367 585
R3650 GNDA_2.n3395 GNDA_2.n3394 585
R3651 GNDA_2.n2230 GNDA_2.n2229 585
R3652 GNDA_2.n2224 GNDA_2.n2167 585
R3653 GNDA_2.n2228 GNDA_2.n2167 585
R3654 GNDA_2.n2226 GNDA_2.n2225 585
R3655 GNDA_2.n2227 GNDA_2.n2226 585
R3656 GNDA_2.n2223 GNDA_2.n2169 585
R3657 GNDA_2.n2169 GNDA_2.n2168 585
R3658 GNDA_2.n2222 GNDA_2.n2221 585
R3659 GNDA_2.n2221 GNDA_2.n2220 585
R3660 GNDA_2.n2218 GNDA_2.n2170 585
R3661 GNDA_2.n2219 GNDA_2.n2218 585
R3662 GNDA_2.n2217 GNDA_2.n2172 585
R3663 GNDA_2.n2217 GNDA_2.n2216 585
R3664 GNDA_2.n2211 GNDA_2.n2171 585
R3665 GNDA_2.n2215 GNDA_2.n2171 585
R3666 GNDA_2.n2213 GNDA_2.n2212 585
R3667 GNDA_2.n2214 GNDA_2.n2213 585
R3668 GNDA_2.n2210 GNDA_2.n2174 585
R3669 GNDA_2.n2174 GNDA_2.n2173 585
R3670 GNDA_2.n2209 GNDA_2.n2208 585
R3671 GNDA_2.n2208 GNDA_2.n2207 585
R3672 GNDA_2.n2205 GNDA_2.n2175 585
R3673 GNDA_2.n2206 GNDA_2.n2205 585
R3674 GNDA_2.n2232 GNDA_2.n2166 585
R3675 GNDA_2.n5281 GNDA_2.n5280 585
R3676 GNDA_2.n5283 GNDA_2.n117 585
R3677 GNDA_2.n5275 GNDA_2.n118 585
R3678 GNDA_2.n5279 GNDA_2.n118 585
R3679 GNDA_2.n5277 GNDA_2.n5276 585
R3680 GNDA_2.n5278 GNDA_2.n5277 585
R3681 GNDA_2.n5274 GNDA_2.n120 585
R3682 GNDA_2.n120 GNDA_2.n119 585
R3683 GNDA_2.n5273 GNDA_2.n5272 585
R3684 GNDA_2.n5272 GNDA_2.n5271 585
R3685 GNDA_2.n5269 GNDA_2.n121 585
R3686 GNDA_2.n5270 GNDA_2.n5269 585
R3687 GNDA_2.n5268 GNDA_2.n123 585
R3688 GNDA_2.n5268 GNDA_2.n5267 585
R3689 GNDA_2.n5262 GNDA_2.n122 585
R3690 GNDA_2.n5266 GNDA_2.n122 585
R3691 GNDA_2.n5264 GNDA_2.n5263 585
R3692 GNDA_2.n5265 GNDA_2.n5264 585
R3693 GNDA_2.n5261 GNDA_2.n125 585
R3694 GNDA_2.n125 GNDA_2.n124 585
R3695 GNDA_2.n5260 GNDA_2.n5259 585
R3696 GNDA_2.n5259 GNDA_2.n5258 585
R3697 GNDA_2.n127 GNDA_2.n126 585
R3698 GNDA_2.n128 GNDA_2.n127 585
R3699 GNDA_2.n5358 GNDA_2.n113 585
R3700 GNDA_2.n5358 GNDA_2.n5357 585
R3701 GNDA_2.n3098 GNDA_2.n112 585
R3702 GNDA_2.n114 GNDA_2.n112 585
R3703 GNDA_2.n3099 GNDA_2.n3097 585
R3704 GNDA_2.n3097 GNDA_2.n3095 585
R3705 GNDA_2.n3100 GNDA_2.n3094 585
R3706 GNDA_2.n3102 GNDA_2.n3094 585
R3707 GNDA_2.n3093 GNDA_2.n3091 585
R3708 GNDA_2.n3103 GNDA_2.n3093 585
R3709 GNDA_2.n3106 GNDA_2.n3090 585
R3710 GNDA_2.n3104 GNDA_2.n3090 585
R3711 GNDA_2.n3107 GNDA_2.n3089 585
R3712 GNDA_2.n3089 GNDA_2.n3087 585
R3713 GNDA_2.n3108 GNDA_2.n3086 585
R3714 GNDA_2.n3110 GNDA_2.n3086 585
R3715 GNDA_2.n3085 GNDA_2.n3082 585
R3716 GNDA_2.n3111 GNDA_2.n3085 585
R3717 GNDA_2.n3114 GNDA_2.n3081 585
R3718 GNDA_2.n3112 GNDA_2.n3081 585
R3719 GNDA_2.n3115 GNDA_2.n3080 585
R3720 GNDA_2.n3084 GNDA_2.n3080 585
R3721 GNDA_2.n3116 GNDA_2.n3076 585
R3722 GNDA_2.n3077 GNDA_2.n3076 585
R3723 GNDA_2.n3117 GNDA_2.n3116 585
R3724 GNDA_2.n3117 GNDA_2.n3077 585
R3725 GNDA_2.n3115 GNDA_2.n3079 585
R3726 GNDA_2.n3084 GNDA_2.n3079 585
R3727 GNDA_2.n3114 GNDA_2.n3113 585
R3728 GNDA_2.n3113 GNDA_2.n3112 585
R3729 GNDA_2.n3083 GNDA_2.n3082 585
R3730 GNDA_2.n3111 GNDA_2.n3083 585
R3731 GNDA_2.n3109 GNDA_2.n3108 585
R3732 GNDA_2.n3110 GNDA_2.n3109 585
R3733 GNDA_2.n3107 GNDA_2.n3088 585
R3734 GNDA_2.n3088 GNDA_2.n3087 585
R3735 GNDA_2.n3106 GNDA_2.n3105 585
R3736 GNDA_2.n3105 GNDA_2.n3104 585
R3737 GNDA_2.n3092 GNDA_2.n3091 585
R3738 GNDA_2.n3103 GNDA_2.n3092 585
R3739 GNDA_2.n3101 GNDA_2.n3100 585
R3740 GNDA_2.n3102 GNDA_2.n3101 585
R3741 GNDA_2.n3099 GNDA_2.n3096 585
R3742 GNDA_2.n3096 GNDA_2.n3095 585
R3743 GNDA_2.n3098 GNDA_2.n115 585
R3744 GNDA_2.n115 GNDA_2.n114 585
R3745 GNDA_2.n5356 GNDA_2.n113 585
R3746 GNDA_2.n5357 GNDA_2.n5356 585
R3747 GNDA_2.n2461 GNDA_2.n2025 585
R3748 GNDA_2.n2463 GNDA_2.n2018 585
R3749 GNDA_2.n2464 GNDA_2.n2017 585
R3750 GNDA_2.n2467 GNDA_2.n2016 585
R3751 GNDA_2.n2468 GNDA_2.n2015 585
R3752 GNDA_2.n2471 GNDA_2.n2014 585
R3753 GNDA_2.n2472 GNDA_2.n2013 585
R3754 GNDA_2.n2475 GNDA_2.n2012 585
R3755 GNDA_2.n2476 GNDA_2.n2011 585
R3756 GNDA_2.n2477 GNDA_2.n2010 585
R3757 GNDA_2.n2009 GNDA_2.n2000 585
R3758 GNDA_2.n2483 GNDA_2.n2482 585
R3759 GNDA_2.n2482 GNDA_2.n2481 585
R3760 GNDA_2.n2002 GNDA_2.n2000 585
R3761 GNDA_2.n2478 GNDA_2.n2477 585
R3762 GNDA_2.n2479 GNDA_2.n2478 585
R3763 GNDA_2.n2476 GNDA_2.n2008 585
R3764 GNDA_2.n2475 GNDA_2.n2474 585
R3765 GNDA_2.n2473 GNDA_2.n2472 585
R3766 GNDA_2.n2471 GNDA_2.n2470 585
R3767 GNDA_2.n2469 GNDA_2.n2468 585
R3768 GNDA_2.n2467 GNDA_2.n2466 585
R3769 GNDA_2.n2465 GNDA_2.n2464 585
R3770 GNDA_2.n2463 GNDA_2.n2462 585
R3771 GNDA_2.n2461 GNDA_2.n2007 585
R3772 GNDA_2.n2479 GNDA_2.n2007 585
R3773 GNDA_2.n3337 GNDA_2.n1785 585
R3774 GNDA_2.n2405 GNDA_2.n1786 585
R3775 GNDA_2.n2406 GNDA_2.n2404 585
R3776 GNDA_2.n2401 GNDA_2.n2400 585
R3777 GNDA_2.n2412 GNDA_2.n2399 585
R3778 GNDA_2.n2413 GNDA_2.n2398 585
R3779 GNDA_2.n2414 GNDA_2.n2397 585
R3780 GNDA_2.n2395 GNDA_2.n2394 585
R3781 GNDA_2.n2419 GNDA_2.n2393 585
R3782 GNDA_2.n2420 GNDA_2.n2392 585
R3783 GNDA_2.n2391 GNDA_2.n2330 585
R3784 GNDA_2.n2453 GNDA_2.n2425 585
R3785 GNDA_2.n2425 GNDA_2.n2424 585
R3786 GNDA_2.n2422 GNDA_2.n2330 585
R3787 GNDA_2.n2421 GNDA_2.n2420 585
R3788 GNDA_2.n2419 GNDA_2.n2418 585
R3789 GNDA_2.n2417 GNDA_2.n2395 585
R3790 GNDA_2.n2415 GNDA_2.n2414 585
R3791 GNDA_2.n2413 GNDA_2.n2396 585
R3792 GNDA_2.n2412 GNDA_2.n2411 585
R3793 GNDA_2.n2409 GNDA_2.n2401 585
R3794 GNDA_2.n2407 GNDA_2.n2406 585
R3795 GNDA_2.n2405 GNDA_2.n2403 585
R3796 GNDA_2.n1785 GNDA_2.n1728 585
R3797 GNDA_2.n3330 GNDA_2.n1809 585
R3798 GNDA_2.n3328 GNDA_2.n3327 585
R3799 GNDA_2.n1811 GNDA_2.n1810 585
R3800 GNDA_2.n3321 GNDA_2.n3320 585
R3801 GNDA_2.n3318 GNDA_2.n1813 585
R3802 GNDA_2.n3316 GNDA_2.n3315 585
R3803 GNDA_2.n1815 GNDA_2.n1814 585
R3804 GNDA_2.n3309 GNDA_2.n3308 585
R3805 GNDA_2.n3306 GNDA_2.n1817 585
R3806 GNDA_2.n3304 GNDA_2.n3303 585
R3807 GNDA_2.n1819 GNDA_2.n1818 585
R3808 GNDA_2.n3297 GNDA_2.n3296 585
R3809 GNDA_2.n3298 GNDA_2.n3297 585
R3810 GNDA_2.n3300 GNDA_2.n1819 585
R3811 GNDA_2.n3303 GNDA_2.n3302 585
R3812 GNDA_2.n1817 GNDA_2.n1816 585
R3813 GNDA_2.n3310 GNDA_2.n3309 585
R3814 GNDA_2.n3312 GNDA_2.n1815 585
R3815 GNDA_2.n3315 GNDA_2.n3314 585
R3816 GNDA_2.n1813 GNDA_2.n1812 585
R3817 GNDA_2.n3322 GNDA_2.n3321 585
R3818 GNDA_2.n3324 GNDA_2.n1811 585
R3819 GNDA_2.n3327 GNDA_2.n3326 585
R3820 GNDA_2.n1809 GNDA_2.n1804 585
R3821 GNDA_2.n2533 GNDA_2.n1916 585
R3822 GNDA_2.n1925 GNDA_2.n1917 585
R3823 GNDA_2.n2529 GNDA_2.n2528 585
R3824 GNDA_2.n1924 GNDA_2.n1923 585
R3825 GNDA_2.n1929 GNDA_2.n1928 585
R3826 GNDA_2.n2521 GNDA_2.n2520 585
R3827 GNDA_2.n2519 GNDA_2.n2518 585
R3828 GNDA_2.n2517 GNDA_2.n1933 585
R3829 GNDA_2.n1932 GNDA_2.n1931 585
R3830 GNDA_2.n2511 GNDA_2.n2510 585
R3831 GNDA_2.n2509 GNDA_2.n2508 585
R3832 GNDA_2.n2507 GNDA_2.n1936 585
R3833 GNDA_2.n2507 GNDA_2.n2506 585
R3834 GNDA_2.n2508 GNDA_2.n1934 585
R3835 GNDA_2.n2512 GNDA_2.n2511 585
R3836 GNDA_2.n2514 GNDA_2.n1931 585
R3837 GNDA_2.n2517 GNDA_2.n2516 585
R3838 GNDA_2.n2518 GNDA_2.n1930 585
R3839 GNDA_2.n2522 GNDA_2.n2521 585
R3840 GNDA_2.n2524 GNDA_2.n1929 585
R3841 GNDA_2.n2525 GNDA_2.n1924 585
R3842 GNDA_2.n2528 GNDA_2.n2527 585
R3843 GNDA_2.n1926 GNDA_2.n1925 585
R3844 GNDA_2.n2102 GNDA_2.n1916 585
R3845 GNDA_2.n5458 GNDA_2.n86 585
R3846 GNDA_2.n5458 GNDA_2.n5457 585
R3847 GNDA_2.n3195 GNDA_2.n85 585
R3848 GNDA_2.n87 GNDA_2.n85 585
R3849 GNDA_2.n3199 GNDA_2.n3194 585
R3850 GNDA_2.n3197 GNDA_2.n3194 585
R3851 GNDA_2.n3200 GNDA_2.n3193 585
R3852 GNDA_2.n3196 GNDA_2.n3193 585
R3853 GNDA_2.n3201 GNDA_2.n3189 585
R3854 GNDA_2.n3191 GNDA_2.n3189 585
R3855 GNDA_2.n3205 GNDA_2.n3190 585
R3856 GNDA_2.n3205 GNDA_2.n3204 585
R3857 GNDA_2.n3206 GNDA_2.n3187 585
R3858 GNDA_2.n3207 GNDA_2.n3206 585
R3859 GNDA_2.n3210 GNDA_2.n3186 585
R3860 GNDA_2.n3208 GNDA_2.n3186 585
R3861 GNDA_2.n3211 GNDA_2.n3185 585
R3862 GNDA_2.n3185 GNDA_2.n3183 585
R3863 GNDA_2.n3212 GNDA_2.n3182 585
R3864 GNDA_2.n3214 GNDA_2.n3182 585
R3865 GNDA_2.n3181 GNDA_2.n2963 585
R3866 GNDA_2.n3215 GNDA_2.n3181 585
R3867 GNDA_2.n3218 GNDA_2.n2961 585
R3868 GNDA_2.n3216 GNDA_2.n2961 585
R3869 GNDA_2.n3218 GNDA_2.n3217 585
R3870 GNDA_2.n3217 GNDA_2.n3216 585
R3871 GNDA_2.n3180 GNDA_2.n2963 585
R3872 GNDA_2.n3215 GNDA_2.n3180 585
R3873 GNDA_2.n3213 GNDA_2.n3212 585
R3874 GNDA_2.n3214 GNDA_2.n3213 585
R3875 GNDA_2.n3211 GNDA_2.n3184 585
R3876 GNDA_2.n3184 GNDA_2.n3183 585
R3877 GNDA_2.n3210 GNDA_2.n3209 585
R3878 GNDA_2.n3209 GNDA_2.n3208 585
R3879 GNDA_2.n3188 GNDA_2.n3187 585
R3880 GNDA_2.n3207 GNDA_2.n3188 585
R3881 GNDA_2.n3203 GNDA_2.n3190 585
R3882 GNDA_2.n3204 GNDA_2.n3203 585
R3883 GNDA_2.n3202 GNDA_2.n3201 585
R3884 GNDA_2.n3202 GNDA_2.n3191 585
R3885 GNDA_2.n3200 GNDA_2.n3192 585
R3886 GNDA_2.n3196 GNDA_2.n3192 585
R3887 GNDA_2.n3199 GNDA_2.n3198 585
R3888 GNDA_2.n3198 GNDA_2.n3197 585
R3889 GNDA_2.n3195 GNDA_2.n88 585
R3890 GNDA_2.n88 GNDA_2.n87 585
R3891 GNDA_2.n5456 GNDA_2.n86 585
R3892 GNDA_2.n5457 GNDA_2.n5456 585
R3893 GNDA_2.n3221 GNDA_2.n3220 585
R3894 GNDA_2.n3222 GNDA_2.n3221 585
R3895 GNDA_2.n2959 GNDA_2.n2958 585
R3896 GNDA_2.n3223 GNDA_2.n2959 585
R3897 GNDA_2.n3226 GNDA_2.n3225 585
R3898 GNDA_2.n3225 GNDA_2.n3224 585
R3899 GNDA_2.n3227 GNDA_2.n2957 585
R3900 GNDA_2.n2957 GNDA_2.n2956 585
R3901 GNDA_2.n3229 GNDA_2.n3228 585
R3902 GNDA_2.n3230 GNDA_2.n3229 585
R3903 GNDA_2.n2955 GNDA_2.n2954 585
R3904 GNDA_2.n3231 GNDA_2.n2955 585
R3905 GNDA_2.n3234 GNDA_2.n3233 585
R3906 GNDA_2.n3233 GNDA_2.n3232 585
R3907 GNDA_2.n3235 GNDA_2.n2953 585
R3908 GNDA_2.n2953 GNDA_2.n2952 585
R3909 GNDA_2.n3237 GNDA_2.n3236 585
R3910 GNDA_2.n3238 GNDA_2.n3237 585
R3911 GNDA_2.n2950 GNDA_2.n2949 585
R3912 GNDA_2.n3239 GNDA_2.n2950 585
R3913 GNDA_2.n3242 GNDA_2.n3241 585
R3914 GNDA_2.n3241 GNDA_2.n3240 585
R3915 GNDA_2.n3243 GNDA_2.n2948 585
R3916 GNDA_2.n2951 GNDA_2.n2948 585
R3917 GNDA_2.n3156 GNDA_2.n3155 585
R3918 GNDA_2.n3155 GNDA_2.n3154 585
R3919 GNDA_2.n3157 GNDA_2.n3073 585
R3920 GNDA_2.n3073 GNDA_2.n3072 585
R3921 GNDA_2.n3159 GNDA_2.n3158 585
R3922 GNDA_2.n3160 GNDA_2.n3159 585
R3923 GNDA_2.n3074 GNDA_2.n3071 585
R3924 GNDA_2.n3161 GNDA_2.n3071 585
R3925 GNDA_2.n3163 GNDA_2.n3070 585
R3926 GNDA_2.n3163 GNDA_2.n3162 585
R3927 GNDA_2.n3165 GNDA_2.n3164 585
R3928 GNDA_2.n3164 GNDA_2.n2971 585
R3929 GNDA_2.n2969 GNDA_2.n2968 585
R3930 GNDA_2.n3169 GNDA_2.n2969 585
R3931 GNDA_2.n3172 GNDA_2.n3171 585
R3932 GNDA_2.n3171 GNDA_2.n3170 585
R3933 GNDA_2.n3173 GNDA_2.n2966 585
R3934 GNDA_2.n2966 GNDA_2.n2965 585
R3935 GNDA_2.n3175 GNDA_2.n3174 585
R3936 GNDA_2.n3176 GNDA_2.n3175 585
R3937 GNDA_2.n2967 GNDA_2.n2964 585
R3938 GNDA_2.n3177 GNDA_2.n2964 585
R3939 GNDA_2.n3179 GNDA_2.n2962 585
R3940 GNDA_2.n3179 GNDA_2.n3178 585
R3941 GNDA_2.n3128 GNDA_2.n3127 585
R3942 GNDA_2.n3129 GNDA_2.n3128 585
R3943 GNDA_2.n3132 GNDA_2.n3131 585
R3944 GNDA_2.n3131 GNDA_2.n3130 585
R3945 GNDA_2.n3133 GNDA_2.n3126 585
R3946 GNDA_2.n3126 GNDA_2.n3125 585
R3947 GNDA_2.n3135 GNDA_2.n3134 585
R3948 GNDA_2.n3136 GNDA_2.n3135 585
R3949 GNDA_2.n3124 GNDA_2.n3123 585
R3950 GNDA_2.n3137 GNDA_2.n3124 585
R3951 GNDA_2.n3140 GNDA_2.n3139 585
R3952 GNDA_2.n3139 GNDA_2.n3138 585
R3953 GNDA_2.n3141 GNDA_2.n3122 585
R3954 GNDA_2.n3122 GNDA_2.n3121 585
R3955 GNDA_2.n3143 GNDA_2.n3142 585
R3956 GNDA_2.n3144 GNDA_2.n3143 585
R3957 GNDA_2.n3120 GNDA_2.n3119 585
R3958 GNDA_2.n3145 GNDA_2.n3120 585
R3959 GNDA_2.n3148 GNDA_2.n3147 585
R3960 GNDA_2.n3147 GNDA_2.n3146 585
R3961 GNDA_2.n3149 GNDA_2.n3118 585
R3962 GNDA_2.n3118 GNDA_2.n3078 585
R3963 GNDA_2.n3151 GNDA_2.n3150 585
R3964 GNDA_2.n3152 GNDA_2.n3151 585
R3965 GNDA_2.n2973 GNDA_2.n2972 585
R3966 GNDA_2.n3168 GNDA_2.n3167 585
R3967 GNDA_2.t73 GNDA_2.n3168 585
R3968 GNDA_2.n1987 GNDA_2.n1986 585
R3969 GNDA_2.n1985 GNDA_2.n1943 585
R3970 GNDA_2.n1984 GNDA_2.n1983 585
R3971 GNDA_2.n1982 GNDA_2.n1981 585
R3972 GNDA_2.n1980 GNDA_2.n1979 585
R3973 GNDA_2.n1978 GNDA_2.n1977 585
R3974 GNDA_2.n1976 GNDA_2.n1975 585
R3975 GNDA_2.n1974 GNDA_2.n1973 585
R3976 GNDA_2.n1972 GNDA_2.n1971 585
R3977 GNDA_2.n1970 GNDA_2.n1969 585
R3978 GNDA_2.n1968 GNDA_2.n1967 585
R3979 GNDA_2.n1966 GNDA_2.n1965 585
R3980 GNDA_2.n2485 GNDA_2.n2484 585
R3981 GNDA_2.n2486 GNDA_2.n1996 585
R3982 GNDA_2.n2488 GNDA_2.n2487 585
R3983 GNDA_2.n2490 GNDA_2.n1994 585
R3984 GNDA_2.n2492 GNDA_2.n2491 585
R3985 GNDA_2.n2493 GNDA_2.n1993 585
R3986 GNDA_2.n2495 GNDA_2.n2494 585
R3987 GNDA_2.n2497 GNDA_2.n1991 585
R3988 GNDA_2.n2499 GNDA_2.n2498 585
R3989 GNDA_2.n2500 GNDA_2.n1990 585
R3990 GNDA_2.n2502 GNDA_2.n2501 585
R3991 GNDA_2.n2504 GNDA_2.n1937 585
R3992 GNDA_2.n2204 GNDA_2.n2203 585
R3993 GNDA_2.n2202 GNDA_2.n2201 585
R3994 GNDA_2.n2200 GNDA_2.n2177 585
R3995 GNDA_2.n2198 GNDA_2.n2197 585
R3996 GNDA_2.n2196 GNDA_2.n2178 585
R3997 GNDA_2.n2195 GNDA_2.n2194 585
R3998 GNDA_2.n2192 GNDA_2.n2179 585
R3999 GNDA_2.n2190 GNDA_2.n2189 585
R4000 GNDA_2.n2188 GNDA_2.n2180 585
R4001 GNDA_2.n2187 GNDA_2.n2186 585
R4002 GNDA_2.n2184 GNDA_2.n2182 585
R4003 GNDA_2.n2181 GNDA_2.n2001 585
R4004 GNDA_2.n5459 GNDA_2.n84 585
R4005 GNDA_2.n5459 GNDA_2.n83 585
R4006 GNDA_2.n5549 GNDA_2.n5548 585
R4007 GNDA_2.n5546 GNDA_2.n54 585
R4008 GNDA_2.n59 GNDA_2.n58 585
R4009 GNDA_2.n5541 GNDA_2.n5540 585
R4010 GNDA_2.n5539 GNDA_2.n5538 585
R4011 GNDA_2.n5465 GNDA_2.n63 585
R4012 GNDA_2.n5467 GNDA_2.n5466 585
R4013 GNDA_2.n5472 GNDA_2.n5471 585
R4014 GNDA_2.n5470 GNDA_2.n5463 585
R4015 GNDA_2.n5478 GNDA_2.n5477 585
R4016 GNDA_2.n5480 GNDA_2.n5479 585
R4017 GNDA_2.n5461 GNDA_2.n5460 585
R4018 GNDA_2.n5359 GNDA_2.n111 585
R4019 GNDA_2.n5359 GNDA_2.n83 585
R4020 GNDA_2.n5455 GNDA_2.n84 585
R4021 GNDA_2.n5455 GNDA_2.n83 585
R4022 GNDA_2.n5454 GNDA_2.n5453 585
R4023 GNDA_2.n5451 GNDA_2.n5450 585
R4024 GNDA_2.n5449 GNDA_2.n5448 585
R4025 GNDA_2.n5365 GNDA_2.n91 585
R4026 GNDA_2.n5367 GNDA_2.n5366 585
R4027 GNDA_2.n5371 GNDA_2.n5370 585
R4028 GNDA_2.n5373 GNDA_2.n5372 585
R4029 GNDA_2.n5380 GNDA_2.n5379 585
R4030 GNDA_2.n5378 GNDA_2.n5363 585
R4031 GNDA_2.n5386 GNDA_2.n5385 585
R4032 GNDA_2.n5388 GNDA_2.n5387 585
R4033 GNDA_2.n5361 GNDA_2.n5360 585
R4034 GNDA_2.n5355 GNDA_2.n111 585
R4035 GNDA_2.n5355 GNDA_2.n83 585
R4036 GNDA_2.n5354 GNDA_2.n5353 585
R4037 GNDA_2.n24 GNDA_2.n22 585
R4038 GNDA_2.n5554 GNDA_2.n5553 585
R4039 GNDA_2.n32 GNDA_2.n25 585
R4040 GNDA_2.n40 GNDA_2.n39 585
R4041 GNDA_2.n35 GNDA_2.n31 585
R4042 GNDA_2.n30 GNDA_2.n0 585
R4043 GNDA_2.n5288 GNDA_2.n1 585
R4044 GNDA_2.n5290 GNDA_2.n5289 585
R4045 GNDA_2.n5294 GNDA_2.n5293 585
R4046 GNDA_2.n5296 GNDA_2.n5295 585
R4047 GNDA_2.n5285 GNDA_2.n5284 585
R4048 GNDA_2.n3294 GNDA_2.n3293 585
R4049 GNDA_2.n3292 GNDA_2.n3291 585
R4050 GNDA_2.n3290 GNDA_2.n1823 585
R4051 GNDA_2.n3288 GNDA_2.n3287 585
R4052 GNDA_2.n3286 GNDA_2.n1824 585
R4053 GNDA_2.n3285 GNDA_2.n3284 585
R4054 GNDA_2.n3282 GNDA_2.n1825 585
R4055 GNDA_2.n3280 GNDA_2.n3279 585
R4056 GNDA_2.n3278 GNDA_2.n1826 585
R4057 GNDA_2.n3277 GNDA_2.n3276 585
R4058 GNDA_2.n3274 GNDA_2.n1827 585
R4059 GNDA_2.n3272 GNDA_2.n3271 585
R4060 GNDA_2.n2455 GNDA_2.n2454 585
R4061 GNDA_2.n2451 GNDA_2.n2426 585
R4062 GNDA_2.n2450 GNDA_2.n2449 585
R4063 GNDA_2.n2448 GNDA_2.n2447 585
R4064 GNDA_2.n2446 GNDA_2.n2428 585
R4065 GNDA_2.n2444 GNDA_2.n2443 585
R4066 GNDA_2.n2442 GNDA_2.n2429 585
R4067 GNDA_2.n2441 GNDA_2.n2440 585
R4068 GNDA_2.n2438 GNDA_2.n2430 585
R4069 GNDA_2.n2436 GNDA_2.n2435 585
R4070 GNDA_2.n2434 GNDA_2.n2432 585
R4071 GNDA_2.n2433 GNDA_2.n1820 585
R4072 GNDA_2.n2370 GNDA_2.n2369 585
R4073 GNDA_2.n2371 GNDA_2.n2337 585
R4074 GNDA_2.n2373 GNDA_2.n2372 585
R4075 GNDA_2.n2375 GNDA_2.n2335 585
R4076 GNDA_2.n2377 GNDA_2.n2376 585
R4077 GNDA_2.n2378 GNDA_2.n2334 585
R4078 GNDA_2.n2380 GNDA_2.n2379 585
R4079 GNDA_2.n2382 GNDA_2.n2332 585
R4080 GNDA_2.n2384 GNDA_2.n2383 585
R4081 GNDA_2.n2385 GNDA_2.n2331 585
R4082 GNDA_2.n2387 GNDA_2.n2386 585
R4083 GNDA_2.n2389 GNDA_2.n2329 585
R4084 GNDA_2.n2534 GNDA_2.n1915 585
R4085 GNDA_2.n2534 GNDA_2.n1914 585
R4086 GNDA_2.n2603 GNDA_2.n1845 585
R4087 GNDA_2.n2601 GNDA_2.n2600 585
R4088 GNDA_2.n1868 GNDA_2.n1849 585
R4089 GNDA_2.n2596 GNDA_2.n2595 585
R4090 GNDA_2.n1870 GNDA_2.n1867 585
R4091 GNDA_2.n1896 GNDA_2.n1895 585
R4092 GNDA_2.n1898 GNDA_2.n1897 585
R4093 GNDA_2.n1901 GNDA_2.n1900 585
R4094 GNDA_2.n1899 GNDA_2.n1889 585
R4095 GNDA_2.n1910 GNDA_2.n1909 585
R4096 GNDA_2.n1912 GNDA_2.n1911 585
R4097 GNDA_2.n2536 GNDA_2.n2535 585
R4098 GNDA_2.n2459 GNDA_2.n2328 585
R4099 GNDA_2.n2328 GNDA_2.n1914 585
R4100 GNDA_2.n2103 GNDA_2.n1915 585
R4101 GNDA_2.n2103 GNDA_2.n1914 585
R4102 GNDA_2.n2105 GNDA_2.n2104 585
R4103 GNDA_2.n2129 GNDA_2.n2107 585
R4104 GNDA_2.n2131 GNDA_2.n2130 585
R4105 GNDA_2.n2127 GNDA_2.n2126 585
R4106 GNDA_2.n2125 GNDA_2.n2124 585
R4107 GNDA_2.n2120 GNDA_2.n2119 585
R4108 GNDA_2.n2118 GNDA_2.n2117 585
R4109 GNDA_2.n2113 GNDA_2.n2112 585
R4110 GNDA_2.n2111 GNDA_2.n2028 585
R4111 GNDA_2.n2139 GNDA_2.n2138 585
R4112 GNDA_2.n2141 GNDA_2.n2140 585
R4113 GNDA_2.n2327 GNDA_2.n2143 585
R4114 GNDA_2.n2459 GNDA_2.n2458 585
R4115 GNDA_2.n2458 GNDA_2.n1914 585
R4116 GNDA_2.n2457 GNDA_2.n2326 585
R4117 GNDA_2.n2324 GNDA_2.n2323 585
R4118 GNDA_2.n2322 GNDA_2.n2321 585
R4119 GNDA_2.n2238 GNDA_2.n2146 585
R4120 GNDA_2.n2240 GNDA_2.n2239 585
R4121 GNDA_2.n2244 GNDA_2.n2243 585
R4122 GNDA_2.n2246 GNDA_2.n2245 585
R4123 GNDA_2.n2253 GNDA_2.n2252 585
R4124 GNDA_2.n2251 GNDA_2.n2236 585
R4125 GNDA_2.n2259 GNDA_2.n2258 585
R4126 GNDA_2.n2261 GNDA_2.n2260 585
R4127 GNDA_2.n2234 GNDA_2.n2233 585
R4128 GNDA_2.n2696 GNDA_2.n2688 585
R4129 GNDA_2.n2690 GNDA_2.n2687 585
R4130 GNDA_2.n2699 GNDA_2.n2687 585
R4131 GNDA_2.n2672 GNDA_2.n2671 585
R4132 GNDA_2.n2820 GNDA_2.n2819 585
R4133 GNDA_2.n2819 GNDA_2.n2818 585
R4134 GNDA_2.n2829 GNDA_2.n2659 585
R4135 GNDA_2.n2836 GNDA_2.n2658 585
R4136 GNDA_2.n2840 GNDA_2.n2658 585
R4137 GNDA_2.n2834 GNDA_2.n2833 585
R4138 GNDA_2.n3375 GNDA_2.n1686 585
R4139 GNDA_2.n3378 GNDA_2.n3377 585
R4140 GNDA_2.n3379 GNDA_2.n3378 585
R4141 GNDA_2.n3370 GNDA_2.n3369 585
R4142 GNDA_2.n3332 GNDA_2.n3331 585
R4143 GNDA_2.n3331 GNDA_2.n1808 585
R4144 GNDA_2.n2928 GNDA_2.n2927 585
R4145 GNDA_2.n2927 GNDA_2.n2926 585
R4146 GNDA_2.n2619 GNDA_2.n2615 585
R4147 GNDA_2.n2925 GNDA_2.n2615 585
R4148 GNDA_2.n2921 GNDA_2.n2920 585
R4149 GNDA_2.n2922 GNDA_2.n2921 585
R4150 GNDA_2.n2621 GNDA_2.n2618 585
R4151 GNDA_2.n2653 GNDA_2.n2618 585
R4152 GNDA_2.n2652 GNDA_2.n2651 585
R4153 GNDA_2.n2654 GNDA_2.n2652 585
R4154 GNDA_2.n2656 GNDA_2.n2647 585
R4155 GNDA_2.n2656 GNDA_2.n2655 585
R4156 GNDA_2.n2843 GNDA_2.n2842 585
R4157 GNDA_2.n2842 GNDA_2.n2841 585
R4158 GNDA_2.n2848 GNDA_2.n2646 585
R4159 GNDA_2.n2646 GNDA_2.n2645 585
R4160 GNDA_2.n2854 GNDA_2.n2853 585
R4161 GNDA_2.n2855 GNDA_2.n2854 585
R4162 GNDA_2.n2644 GNDA_2.n2643 585
R4163 GNDA_2.n2856 GNDA_2.n2644 585
R4164 GNDA_2.n2860 GNDA_2.n2859 585
R4165 GNDA_2.n2859 GNDA_2.n2858 585
R4166 GNDA_2.n2641 GNDA_2.n1807 585
R4167 GNDA_2.n2857 GNDA_2.n1807 585
R4168 GNDA_2.n3339 GNDA_2.n3338 585
R4169 GNDA_2.n3338 GNDA_2.n1784 585
R4170 GNDA_2.n3333 GNDA_2.n3332 585
R4171 GNDA_2.n3334 GNDA_2.n3333 585
R4172 GNDA_2.n2767 GNDA_2.n1805 585
R4173 GNDA_2.n2686 GNDA_2.n1805 585
R4174 GNDA_2.n2768 GNDA_2.n2703 585
R4175 GNDA_2.n2703 GNDA_2.n2702 585
R4176 GNDA_2.n2778 GNDA_2.n2777 585
R4177 GNDA_2.n2779 GNDA_2.n2778 585
R4178 GNDA_2.n2705 GNDA_2.n2685 585
R4179 GNDA_2.n2780 GNDA_2.n2685 585
R4180 GNDA_2.n2784 GNDA_2.n2783 585
R4181 GNDA_2.n2783 GNDA_2.n2782 585
R4182 GNDA_2.n2785 GNDA_2.n2680 585
R4183 GNDA_2.n2781 GNDA_2.n2680 585
R4184 GNDA_2.n2794 GNDA_2.n2793 585
R4185 GNDA_2.n2795 GNDA_2.n2794 585
R4186 GNDA_2.n2681 GNDA_2.n2679 585
R4187 GNDA_2.n2796 GNDA_2.n2679 585
R4188 GNDA_2.n2800 GNDA_2.n2799 585
R4189 GNDA_2.n2799 GNDA_2.n2798 585
R4190 GNDA_2.n2801 GNDA_2.n2673 585
R4191 GNDA_2.n2797 GNDA_2.n2673 585
R4192 GNDA_2.n2811 GNDA_2.n2810 585
R4193 GNDA_2.n2812 GNDA_2.n2811 585
R4194 GNDA_2.n2808 GNDA_2.n1783 585
R4195 GNDA_2.n2815 GNDA_2.n1783 585
R4196 GNDA_2.n3340 GNDA_2.n3339 585
R4197 GNDA_2.n3341 GNDA_2.n3340 585
R4198 GNDA_2.n1781 GNDA_2.n1727 585
R4199 GNDA_2.n3342 GNDA_2.n1727 585
R4200 GNDA_2.n3344 GNDA_2.n1725 585
R4201 GNDA_2.n3344 GNDA_2.n3343 585
R4202 GNDA_2.n3359 GNDA_2.n3358 585
R4203 GNDA_2.n3358 GNDA_2.n3357 585
R4204 GNDA_2.n3346 GNDA_2.n3345 585
R4205 GNDA_2.n3356 GNDA_2.n3345 585
R4206 GNDA_2.n3354 GNDA_2.n3353 585
R4207 GNDA_2.n3355 GNDA_2.n3354 585
R4208 GNDA_2.n3349 GNDA_2.n1692 585
R4209 GNDA_2.n1692 GNDA_2.n1687 585
R4210 GNDA_2.n3367 GNDA_2.n3366 585
R4211 GNDA_2.n3368 GNDA_2.n3367 585
R4212 GNDA_2.n1694 GNDA_2.n1693 585
R4213 GNDA_2.n1702 GNDA_2.n1693 585
R4214 GNDA_2.n1705 GNDA_2.n1704 585
R4215 GNDA_2.n1704 GNDA_2.n1703 585
R4216 GNDA_2.n1706 GNDA_2.n1669 585
R4217 GNDA_2.n1669 GNDA_2.n1667 585
R4218 GNDA_2.n3401 GNDA_2.n3400 585
R4219 GNDA_2.n3402 GNDA_2.n3401 585
R4220 GNDA_2.n3398 GNDA_2.n1670 585
R4221 GNDA_2.n1670 GNDA_2.n1668 585
R4222 GNDA_2.n3270 GNDA_2.n1828 585
R4223 GNDA_2.n3269 GNDA_2.n3268 585
R4224 GNDA_2.n1830 GNDA_2.n1829 585
R4225 GNDA_2.n2944 GNDA_2.n2943 585
R4226 GNDA_2.n2942 GNDA_2.n2612 585
R4227 GNDA_2.n2941 GNDA_2.n2940 585
R4228 GNDA_2.n2939 GNDA_2.n2938 585
R4229 GNDA_2.n2937 GNDA_2.n2936 585
R4230 GNDA_2.n2935 GNDA_2.n2934 585
R4231 GNDA_2.n2933 GNDA_2.n2932 585
R4232 GNDA_2.n2931 GNDA_2.n2930 585
R4233 GNDA_2.n3266 GNDA_2.n2607 585
R4234 GNDA_2.n1964 GNDA_2.n1963 585
R4235 GNDA_2.n1962 GNDA_2.n1961 585
R4236 GNDA_2.n1960 GNDA_2.n1959 585
R4237 GNDA_2.n1958 GNDA_2.n1957 585
R4238 GNDA_2.n1956 GNDA_2.n1955 585
R4239 GNDA_2.n1954 GNDA_2.n1953 585
R4240 GNDA_2.n1952 GNDA_2.n1951 585
R4241 GNDA_2.n1950 GNDA_2.n1949 585
R4242 GNDA_2.n1948 GNDA_2.n1947 585
R4243 GNDA_2.n1946 GNDA_2.n1945 585
R4244 GNDA_2.n1944 GNDA_2.n1846 585
R4245 GNDA_2.n3266 GNDA_2.n2606 585
R4246 GNDA_2.n3264 GNDA_2.n3263 585
R4247 GNDA_2.n3262 GNDA_2.n2947 585
R4248 GNDA_2.n3261 GNDA_2.n2946 585
R4249 GNDA_2.n3266 GNDA_2.n2946 585
R4250 GNDA_2.n3260 GNDA_2.n3259 585
R4251 GNDA_2.n3258 GNDA_2.n3257 585
R4252 GNDA_2.n3256 GNDA_2.n3255 585
R4253 GNDA_2.n3254 GNDA_2.n3253 585
R4254 GNDA_2.n3252 GNDA_2.n3251 585
R4255 GNDA_2.n3250 GNDA_2.n3249 585
R4256 GNDA_2.n3248 GNDA_2.n3247 585
R4257 GNDA_2.n3246 GNDA_2.n3245 585
R4258 GNDA_2.n3244 GNDA_2.n56 585
R4259 GNDA_2.n56 GNDA_2.n55 585
R4260 GNDA_2.n381 GNDA_2.n375 582.4
R4261 GNDA_2.n4355 GNDA_2.n4354 582.4
R4262 GNDA_2.n4327 GNDA_2.t256 562.222
R4263 GNDA_2.t16 GNDA_2.n117 557.13
R4264 GNDA_2.n351 GNDA_2.t155 548.082
R4265 GNDA_2.n372 GNDA_2.t141 546.375
R4266 GNDA_2.n4399 GNDA_2.t86 546.375
R4267 GNDA_2.n307 GNDA_2.t95 546.375
R4268 GNDA_2.n4472 GNDA_2.t157 524.808
R4269 GNDA_2.n4621 GNDA_2.t133 524.808
R4270 GNDA_2.n4209 GNDA_2.t89 524.808
R4271 GNDA_2.n4312 GNDA_2.t111 524.808
R4272 GNDA_2.n5357 GNDA_2.t73 512.884
R4273 GNDA_2.n5457 GNDA_2.t73 512.884
R4274 GNDA_2.n4431 GNDA_2.t83 509.2
R4275 GNDA_2.n4429 GNDA_2.t68 509.2
R4276 GNDA_2.n562 GNDA_2.t105 509.034
R4277 GNDA_2.n1075 GNDA_2.t143 509.034
R4278 GNDA_2.n4349 GNDA_2.t114 492.675
R4279 GNDA_2.n4352 GNDA_2.t136 492.675
R4280 GNDA_2.n376 GNDA_2.t127 492.675
R4281 GNDA_2.n379 GNDA_2.t153 492.675
R4282 GNDA_2.n2166 GNDA_2.t73 486.94
R4283 GNDA_2.n4337 GNDA_2.n4336 483.2
R4284 GNDA_2.n4336 GNDA_2.n387 476.8
R4285 GNDA_2.n1662 GNDA_2.t145 425.134
R4286 GNDA_2.n1652 GNDA_2.t129 425.134
R4287 GNDA_2.n1080 GNDA_2.t106 415.557
R4288 GNDA_2.n3405 GNDA_2.t138 409.067
R4289 GNDA_2.n1663 GNDA_2.t80 409.067
R4290 GNDA_2.n1658 GNDA_2.t116 409.067
R4291 GNDA_2.n1657 GNDA_2.t77 409.067
R4292 GNDA_2.n1653 GNDA_2.t161 409.067
R4293 GNDA_2.n1649 GNDA_2.t65 409.067
R4294 GNDA_2.n5258 GNDA_2.n128 394.817
R4295 GNDA_2.n5265 GNDA_2.n124 394.817
R4296 GNDA_2.n5266 GNDA_2.n5265 394.817
R4297 GNDA_2.n5267 GNDA_2.n5266 394.817
R4298 GNDA_2.n5271 GNDA_2.n5270 394.817
R4299 GNDA_2.n5271 GNDA_2.n119 394.817
R4300 GNDA_2.n5278 GNDA_2.n119 394.817
R4301 GNDA_2.n5279 GNDA_2.n5278 394.817
R4302 GNDA_2.n5280 GNDA_2.n5279 394.817
R4303 GNDA_2.n5280 GNDA_2.n117 394.817
R4304 GNDA_2.n2207 GNDA_2.n2206 394.817
R4305 GNDA_2.n2207 GNDA_2.n2173 394.817
R4306 GNDA_2.n2214 GNDA_2.n2173 394.817
R4307 GNDA_2.n2215 GNDA_2.n2214 394.817
R4308 GNDA_2.n2216 GNDA_2.n2215 394.817
R4309 GNDA_2.n2220 GNDA_2.n2219 394.817
R4310 GNDA_2.n2220 GNDA_2.n2168 394.817
R4311 GNDA_2.n2227 GNDA_2.n2168 394.817
R4312 GNDA_2.n2228 GNDA_2.n2227 394.817
R4313 GNDA_2.n2229 GNDA_2.n2228 394.817
R4314 GNDA_2.n2229 GNDA_2.n2166 394.817
R4315 GNDA_2.n2367 GNDA_2.n2366 394.817
R4316 GNDA_2.n2366 GNDA_2.n2365 394.817
R4317 GNDA_2.n2365 GNDA_2.n2341 394.817
R4318 GNDA_2.n2359 GNDA_2.n2341 394.817
R4319 GNDA_2.n2359 GNDA_2.n1690 394.817
R4320 GNDA_2.n2348 GNDA_2.n1691 394.817
R4321 GNDA_2.n2352 GNDA_2.n2348 394.817
R4322 GNDA_2.n2352 GNDA_2.n2351 394.817
R4323 GNDA_2.n2351 GNDA_2.n2350 394.817
R4324 GNDA_2.n2350 GNDA_2.n1675 394.817
R4325 GNDA_2.n3394 GNDA_2.n1675 394.817
R4326 GNDA_2.n3104 GNDA_2.t73 391.411
R4327 GNDA_2.n3204 GNDA_2.t73 391.411
R4328 GNDA_2.n4330 GNDA_2.n4329 384
R4329 GNDA_2.n5258 GNDA_2.n5257 377.269
R4330 GNDA_2.n4331 GNDA_2.n4330 355.2
R4331 GNDA_2.n4329 GNDA_2.n1079 345.601
R4332 GNDA_2.n1797 GNDA_2.t73 172.876
R4333 GNDA_2.n3335 GNDA_2.t73 172.876
R4334 GNDA_2.n1801 GNDA_2.t73 172.615
R4335 GNDA_2.t73 GNDA_2.n1689 172.615
R4336 GNDA_2.n4331 GNDA_2.n1079 316.8
R4337 GNDA_2.t106 GNDA_2.n1076 293.651
R4338 GNDA_2.t106 GNDA_2.n388 293.651
R4339 GNDA_2.n384 GNDA_2.n382 292.5
R4340 GNDA_2.n4322 GNDA_2.n382 292.5
R4341 GNDA_2.n369 GNDA_2.n334 292.5
R4342 GNDA_2.n4405 GNDA_2.n334 292.5
R4343 GNDA_2.n4404 GNDA_2.n4403 292.5
R4344 GNDA_2.n4405 GNDA_2.n4404 292.5
R4345 GNDA_2.n4342 GNDA_2.n383 292.5
R4346 GNDA_2.n4324 GNDA_2.n383 292.5
R4347 GNDA_2.n350 GNDA_2.n301 292.5
R4348 GNDA_2.n4461 GNDA_2.n301 292.5
R4349 GNDA_2.n4460 GNDA_2.n4459 292.5
R4350 GNDA_2.n4461 GNDA_2.n4460 292.5
R4351 GNDA_2.n4330 GNDA_2.n1078 292.5
R4352 GNDA_2.n1080 GNDA_2.n1078 292.5
R4353 GNDA_2.n4329 GNDA_2.n4328 292.5
R4354 GNDA_2.n4328 GNDA_2.n4327 292.5
R4355 GNDA_2.n1079 GNDA_2.n1077 292.5
R4356 GNDA_2.n1080 GNDA_2.n1077 292.5
R4357 GNDA_2.n4332 GNDA_2.n4331 292.5
R4358 GNDA_2.n4333 GNDA_2.n4332 292.5
R4359 GNDA_2.n4336 GNDA_2.n4335 292.5
R4360 GNDA_2.n4335 GNDA_2.n4334 292.5
R4361 GNDA_2.n4344 GNDA_2.n4343 292.5
R4362 GNDA_2.n4345 GNDA_2.n4344 292.5
R4363 GNDA_2.n4348 GNDA_2.n4347 292.5
R4364 GNDA_2.n4347 GNDA_2.n4346 292.5
R4365 GNDA_2.n4361 GNDA_2.n4360 292.5
R4366 GNDA_2.n4362 GNDA_2.n4361 292.5
R4367 GNDA_2.n338 GNDA_2.n303 292.5
R4368 GNDA_2.n4363 GNDA_2.n303 292.5
R4369 GNDA_2.n335 GNDA_2.n302 292.5
R4370 GNDA_2.n4364 GNDA_2.n302 292.5
R4371 GNDA_2.n4371 GNDA_2.n4370 292.5
R4372 GNDA_2.n4370 GNDA_2.n4369 292.5
R4373 GNDA_2.n348 GNDA_2.n345 292.5
R4374 GNDA_2.n4365 GNDA_2.n348 292.5
R4375 GNDA_2.n4368 GNDA_2.n4367 292.5
R4376 GNDA_2.n4369 GNDA_2.n4368 292.5
R4377 GNDA_2.n347 GNDA_2.n346 292.5
R4378 GNDA_2.n5267 GNDA_2.t73 267.598
R4379 GNDA_2.n2216 GNDA_2.t73 267.598
R4380 GNDA_2.t73 GNDA_2.n1690 267.598
R4381 GNDA_2.n3266 GNDA_2.n1838 264.301
R4382 GNDA_2.n3397 GNDA_2.n3396 264.301
R4383 GNDA_2.n2231 GNDA_2.n2165 264.301
R4384 GNDA_2.n5282 GNDA_2.n116 264.301
R4385 GNDA_2.n2929 GNDA_2.n2613 264.301
R4386 GNDA_2.n2605 GNDA_2.n2604 264.301
R4387 GNDA_2.n3391 GNDA_2.t49 260
R4388 GNDA_2.n3389 GNDA_2.t49 260
R4389 GNDA_2.n3221 GNDA_2.n2961 259.416
R4390 GNDA_2.n1987 GNDA_2.n1936 259.416
R4391 GNDA_2.n3296 GNDA_2.n3294 259.416
R4392 GNDA_2.n2454 GNDA_2.n2453 259.416
R4393 GNDA_2.n2484 GNDA_2.n2483 259.416
R4394 GNDA_2.n3155 GNDA_2.n3076 259.416
R4395 GNDA_2.n2205 GNDA_2.n2204 259.416
R4396 GNDA_2.n2369 GNDA_2.n2368 259.416
R4397 GNDA_2.n3128 GNDA_2.n127 259.416
R4398 GNDA_2.n5517 GNDA_2.n80 258.334
R4399 GNDA_2.n2573 GNDA_2.n2571 258.334
R4400 GNDA_2.n2899 GNDA_2.n2898 258.334
R4401 GNDA_2.n2752 GNDA_2.n2710 258.334
R4402 GNDA_2.n2084 GNDA_2.n2083 258.334
R4403 GNDA_2.n5427 GNDA_2.n5426 258.334
R4404 GNDA_2.n2300 GNDA_2.n2299 258.334
R4405 GNDA_2.n1763 GNDA_2.n1762 258.334
R4406 GNDA_2.n5335 GNDA_2.n5334 258.334
R4407 GNDA_2.t73 GNDA_2.n2970 257.779
R4408 GNDA_2.n2024 GNDA_2.n2023 254.34
R4409 GNDA_2.n2023 GNDA_2.n2022 254.34
R4410 GNDA_2.n2023 GNDA_2.n2021 254.34
R4411 GNDA_2.n2023 GNDA_2.n2020 254.34
R4412 GNDA_2.n2023 GNDA_2.n2019 254.34
R4413 GNDA_2.n2023 GNDA_2.n1999 254.34
R4414 GNDA_2.n2480 GNDA_2.n2479 254.34
R4415 GNDA_2.n2479 GNDA_2.n2003 254.34
R4416 GNDA_2.n2479 GNDA_2.n2004 254.34
R4417 GNDA_2.n2479 GNDA_2.n2005 254.34
R4418 GNDA_2.n2479 GNDA_2.n2006 254.34
R4419 GNDA_2.n3336 GNDA_2.n3335 254.34
R4420 GNDA_2.n3335 GNDA_2.n1796 254.34
R4421 GNDA_2.n3335 GNDA_2.n1795 254.34
R4422 GNDA_2.n3335 GNDA_2.n1794 254.34
R4423 GNDA_2.n3335 GNDA_2.n1793 254.34
R4424 GNDA_2.n3335 GNDA_2.n1792 254.34
R4425 GNDA_2.n2423 GNDA_2.n1689 254.34
R4426 GNDA_2.n2390 GNDA_2.n1689 254.34
R4427 GNDA_2.n2416 GNDA_2.n1689 254.34
R4428 GNDA_2.n2410 GNDA_2.n1689 254.34
R4429 GNDA_2.n2408 GNDA_2.n1689 254.34
R4430 GNDA_2.n2402 GNDA_2.n1689 254.34
R4431 GNDA_2.n3329 GNDA_2.n1797 254.34
R4432 GNDA_2.n3319 GNDA_2.n1797 254.34
R4433 GNDA_2.n3317 GNDA_2.n1797 254.34
R4434 GNDA_2.n3307 GNDA_2.n1797 254.34
R4435 GNDA_2.n3305 GNDA_2.n1797 254.34
R4436 GNDA_2.n3295 GNDA_2.n1797 254.34
R4437 GNDA_2.n3299 GNDA_2.n1801 254.34
R4438 GNDA_2.n3301 GNDA_2.n1801 254.34
R4439 GNDA_2.n3311 GNDA_2.n1801 254.34
R4440 GNDA_2.n3313 GNDA_2.n1801 254.34
R4441 GNDA_2.n3323 GNDA_2.n1801 254.34
R4442 GNDA_2.n3325 GNDA_2.n1801 254.34
R4443 GNDA_2.n2532 GNDA_2.n2531 254.34
R4444 GNDA_2.n2531 GNDA_2.n2530 254.34
R4445 GNDA_2.n2531 GNDA_2.n1922 254.34
R4446 GNDA_2.n2531 GNDA_2.n1921 254.34
R4447 GNDA_2.n2531 GNDA_2.n1920 254.34
R4448 GNDA_2.n2531 GNDA_2.n1919 254.34
R4449 GNDA_2.n2505 GNDA_2.n1927 254.34
R4450 GNDA_2.n2513 GNDA_2.n1927 254.34
R4451 GNDA_2.n2515 GNDA_2.n1927 254.34
R4452 GNDA_2.n2523 GNDA_2.n1927 254.34
R4453 GNDA_2.n2526 GNDA_2.n1927 254.34
R4454 GNDA_2.n2101 GNDA_2.n1927 254.34
R4455 GNDA_2.n1989 GNDA_2.n1988 254.34
R4456 GNDA_2.n1989 GNDA_2.n1942 254.34
R4457 GNDA_2.n1989 GNDA_2.n1941 254.34
R4458 GNDA_2.n1989 GNDA_2.n1940 254.34
R4459 GNDA_2.n1989 GNDA_2.n1939 254.34
R4460 GNDA_2.n1989 GNDA_2.n1938 254.34
R4461 GNDA_2.n1998 GNDA_2.n1989 254.34
R4462 GNDA_2.n2489 GNDA_2.n1989 254.34
R4463 GNDA_2.n1995 GNDA_2.n1989 254.34
R4464 GNDA_2.n2496 GNDA_2.n1989 254.34
R4465 GNDA_2.n1992 GNDA_2.n1989 254.34
R4466 GNDA_2.n2503 GNDA_2.n1989 254.34
R4467 GNDA_2.n2176 GNDA_2.n1989 254.34
R4468 GNDA_2.n2199 GNDA_2.n1989 254.34
R4469 GNDA_2.n2193 GNDA_2.n1989 254.34
R4470 GNDA_2.n2191 GNDA_2.n1989 254.34
R4471 GNDA_2.n2185 GNDA_2.n1989 254.34
R4472 GNDA_2.n2183 GNDA_2.n1989 254.34
R4473 GNDA_2.n5551 GNDA_2.n5550 254.34
R4474 GNDA_2.n5551 GNDA_2.n53 254.34
R4475 GNDA_2.n5551 GNDA_2.n52 254.34
R4476 GNDA_2.n5551 GNDA_2.n51 254.34
R4477 GNDA_2.n5551 GNDA_2.n50 254.34
R4478 GNDA_2.n5551 GNDA_2.n49 254.34
R4479 GNDA_2.n5551 GNDA_2.n48 254.34
R4480 GNDA_2.n5551 GNDA_2.n47 254.34
R4481 GNDA_2.n5551 GNDA_2.n46 254.34
R4482 GNDA_2.n5551 GNDA_2.n45 254.34
R4483 GNDA_2.n5551 GNDA_2.n44 254.34
R4484 GNDA_2.n5551 GNDA_2.n43 254.34
R4485 GNDA_2.n5551 GNDA_2.n42 254.34
R4486 GNDA_2.n5552 GNDA_2.n5551 254.34
R4487 GNDA_2.n5551 GNDA_2.n41 254.34
R4488 GNDA_2.n5551 GNDA_2.n29 254.34
R4489 GNDA_2.n5551 GNDA_2.n28 254.34
R4490 GNDA_2.n5551 GNDA_2.n27 254.34
R4491 GNDA_2.n1822 GNDA_2.n1800 254.34
R4492 GNDA_2.n3289 GNDA_2.n1800 254.34
R4493 GNDA_2.n3283 GNDA_2.n1800 254.34
R4494 GNDA_2.n3281 GNDA_2.n1800 254.34
R4495 GNDA_2.n3275 GNDA_2.n1800 254.34
R4496 GNDA_2.n3273 GNDA_2.n1800 254.34
R4497 GNDA_2.n2452 GNDA_2.n1800 254.34
R4498 GNDA_2.n2427 GNDA_2.n1800 254.34
R4499 GNDA_2.n2445 GNDA_2.n1800 254.34
R4500 GNDA_2.n2439 GNDA_2.n1800 254.34
R4501 GNDA_2.n2437 GNDA_2.n1800 254.34
R4502 GNDA_2.n2431 GNDA_2.n1800 254.34
R4503 GNDA_2.n2339 GNDA_2.n1800 254.34
R4504 GNDA_2.n2374 GNDA_2.n1800 254.34
R4505 GNDA_2.n2336 GNDA_2.n1800 254.34
R4506 GNDA_2.n2381 GNDA_2.n1800 254.34
R4507 GNDA_2.n2333 GNDA_2.n1800 254.34
R4508 GNDA_2.n2388 GNDA_2.n1800 254.34
R4509 GNDA_2.n2599 GNDA_2.n2598 254.34
R4510 GNDA_2.n2598 GNDA_2.n2597 254.34
R4511 GNDA_2.n2598 GNDA_2.n1866 254.34
R4512 GNDA_2.n2598 GNDA_2.n1865 254.34
R4513 GNDA_2.n2598 GNDA_2.n1864 254.34
R4514 GNDA_2.n2598 GNDA_2.n1863 254.34
R4515 GNDA_2.n2598 GNDA_2.n1862 254.34
R4516 GNDA_2.n2598 GNDA_2.n1861 254.34
R4517 GNDA_2.n2598 GNDA_2.n1860 254.34
R4518 GNDA_2.n2598 GNDA_2.n1859 254.34
R4519 GNDA_2.n2598 GNDA_2.n1858 254.34
R4520 GNDA_2.n2598 GNDA_2.n1857 254.34
R4521 GNDA_2.n2598 GNDA_2.n1856 254.34
R4522 GNDA_2.n2598 GNDA_2.n1855 254.34
R4523 GNDA_2.n2598 GNDA_2.n1854 254.34
R4524 GNDA_2.n2598 GNDA_2.n1853 254.34
R4525 GNDA_2.n2598 GNDA_2.n1852 254.34
R4526 GNDA_2.n2598 GNDA_2.n1851 254.34
R4527 GNDA_2.n3267 GNDA_2.n3266 254.34
R4528 GNDA_2.n3266 GNDA_2.n2945 254.34
R4529 GNDA_2.n3266 GNDA_2.n2611 254.34
R4530 GNDA_2.n3266 GNDA_2.n2610 254.34
R4531 GNDA_2.n3266 GNDA_2.n2609 254.34
R4532 GNDA_2.n3266 GNDA_2.n2608 254.34
R4533 GNDA_2.n3266 GNDA_2.n1839 254.34
R4534 GNDA_2.n3266 GNDA_2.n1840 254.34
R4535 GNDA_2.n3266 GNDA_2.n1841 254.34
R4536 GNDA_2.n3266 GNDA_2.n1842 254.34
R4537 GNDA_2.n3266 GNDA_2.n1843 254.34
R4538 GNDA_2.n3266 GNDA_2.n1844 254.34
R4539 GNDA_2.n3266 GNDA_2.n3265 254.34
R4540 GNDA_2.n3266 GNDA_2.n1834 254.34
R4541 GNDA_2.n3266 GNDA_2.n1835 254.34
R4542 GNDA_2.n3266 GNDA_2.n1836 254.34
R4543 GNDA_2.n3266 GNDA_2.n1837 254.34
R4544 GNDA_2.n2699 GNDA_2.n2698 250.349
R4545 GNDA_2.n2818 GNDA_2.n2817 250.349
R4546 GNDA_2.n3264 GNDA_2.n2948 249.663
R4547 GNDA_2.n1965 GNDA_2.n1964 249.663
R4548 GNDA_2.n3272 GNDA_2.n1828 249.663
R4549 GNDA_2.n3298 GNDA_2.n1820 249.663
R4550 GNDA_2.n2506 GNDA_2.n2504 249.663
R4551 GNDA_2.n3217 GNDA_2.n3179 249.663
R4552 GNDA_2.n2481 GNDA_2.n2001 249.663
R4553 GNDA_2.n2424 GNDA_2.n2389 249.663
R4554 GNDA_2.n3151 GNDA_2.n3117 249.663
R4555 GNDA_2.n4371 GNDA_2.n346 249.601
R4556 GNDA_2.n4367 GNDA_2.n346 249.601
R4557 GNDA_2.n3378 GNDA_2.n1686 246.25
R4558 GNDA_2.n3378 GNDA_2.n3369 246.25
R4559 GNDA_2.n2659 GNDA_2.n2658 246.25
R4560 GNDA_2.n2833 GNDA_2.n2658 246.25
R4561 GNDA_2.n3392 GNDA_2.n1678 246.25
R4562 GNDA_2.n2840 GNDA_2.n2839 241.643
R4563 GNDA_2.n2840 GNDA_2.n2657 241.643
R4564 GNDA_2.n3380 GNDA_2.n3379 241.643
R4565 GNDA_2.n3379 GNDA_2.n1688 241.643
R4566 GNDA_2.t29 GNDA_2.t130 227.873
R4567 GNDA_2.n3393 GNDA_2.t48 219.343
R4568 GNDA_2.n1677 GNDA_2.t48 219.343
R4569 GNDA_2.n4327 GNDA_2.n4326 207.779
R4570 GNDA_2.n2819 GNDA_2.n2672 197
R4571 GNDA_2.n2688 GNDA_2.n2687 197
R4572 GNDA_2.n5460 GNDA_2.n5459 197
R4573 GNDA_2.n2535 GNDA_2.n2534 197
R4574 GNDA_2.n3331 GNDA_2.n1807 197
R4575 GNDA_2.n3338 GNDA_2.n1783 197
R4576 GNDA_2.n2328 GNDA_2.n2327 197
R4577 GNDA_2.n5360 GNDA_2.n5359 197
R4578 GNDA_2.n2233 GNDA_2.n2232 197
R4579 GNDA_2.n3395 GNDA_2.n1670 197
R4580 GNDA_2.n5284 GNDA_2.n5283 197
R4581 GNDA_2.n5549 GNDA_2.n55 187.249
R4582 GNDA_2.n2606 GNDA_2.n1845 187.249
R4583 GNDA_2.n2927 GNDA_2.n2607 187.249
R4584 GNDA_2.n3333 GNDA_2.n1805 187.249
R4585 GNDA_2.n2104 GNDA_2.n2103 187.249
R4586 GNDA_2.n5455 GNDA_2.n5454 187.249
R4587 GNDA_2.n2458 GNDA_2.n2457 187.249
R4588 GNDA_2.n3340 GNDA_2.n1727 187.249
R4589 GNDA_2.n5355 GNDA_2.n5354 187.249
R4590 GNDA_2.n5519 GNDA_2.n80 185
R4591 GNDA_2.n5533 GNDA_2.n5532 185
R4592 GNDA_2.n5531 GNDA_2.n81 185
R4593 GNDA_2.n5530 GNDA_2.n5529 185
R4594 GNDA_2.n5528 GNDA_2.n5527 185
R4595 GNDA_2.n5526 GNDA_2.n5525 185
R4596 GNDA_2.n5524 GNDA_2.n5523 185
R4597 GNDA_2.n5522 GNDA_2.n5521 185
R4598 GNDA_2.n5520 GNDA_2.n57 185
R4599 GNDA_2.n5502 GNDA_2.n5501 185
R4600 GNDA_2.n5504 GNDA_2.n5503 185
R4601 GNDA_2.n5506 GNDA_2.n5505 185
R4602 GNDA_2.n5508 GNDA_2.n5507 185
R4603 GNDA_2.n5510 GNDA_2.n5509 185
R4604 GNDA_2.n5512 GNDA_2.n5511 185
R4605 GNDA_2.n5514 GNDA_2.n5513 185
R4606 GNDA_2.n5516 GNDA_2.n5515 185
R4607 GNDA_2.n5518 GNDA_2.n5517 185
R4608 GNDA_2.n5484 GNDA_2.n5483 185
R4609 GNDA_2.n5486 GNDA_2.n5485 185
R4610 GNDA_2.n5488 GNDA_2.n5487 185
R4611 GNDA_2.n5490 GNDA_2.n5489 185
R4612 GNDA_2.n5492 GNDA_2.n5491 185
R4613 GNDA_2.n5494 GNDA_2.n5493 185
R4614 GNDA_2.n5496 GNDA_2.n5495 185
R4615 GNDA_2.n5498 GNDA_2.n5497 185
R4616 GNDA_2.n5500 GNDA_2.n5499 185
R4617 GNDA_2.n5482 GNDA_2.n5481 185
R4618 GNDA_2.n5476 GNDA_2.n5475 185
R4619 GNDA_2.n5474 GNDA_2.n5473 185
R4620 GNDA_2.n5469 GNDA_2.n5468 185
R4621 GNDA_2.n5464 GNDA_2.n65 185
R4622 GNDA_2.n5537 GNDA_2.n5536 185
R4623 GNDA_2.n64 GNDA_2.n62 185
R4624 GNDA_2.n5543 GNDA_2.n5542 185
R4625 GNDA_2.n5545 GNDA_2.n5544 185
R4626 GNDA_2.n2574 GNDA_2.n2573 185
R4627 GNDA_2.n2575 GNDA_2.n1875 185
R4628 GNDA_2.n2577 GNDA_2.n2576 185
R4629 GNDA_2.n2579 GNDA_2.n1874 185
R4630 GNDA_2.n2582 GNDA_2.n2581 185
R4631 GNDA_2.n2583 GNDA_2.n1873 185
R4632 GNDA_2.n2585 GNDA_2.n2584 185
R4633 GNDA_2.n2587 GNDA_2.n1872 185
R4634 GNDA_2.n2588 GNDA_2.n1847 185
R4635 GNDA_2.n2555 GNDA_2.n1880 185
R4636 GNDA_2.n2558 GNDA_2.n2557 185
R4637 GNDA_2.n2559 GNDA_2.n1879 185
R4638 GNDA_2.n2561 GNDA_2.n2560 185
R4639 GNDA_2.n2563 GNDA_2.n1878 185
R4640 GNDA_2.n2566 GNDA_2.n2565 185
R4641 GNDA_2.n2567 GNDA_2.n1877 185
R4642 GNDA_2.n2569 GNDA_2.n2568 185
R4643 GNDA_2.n2571 GNDA_2.n1876 185
R4644 GNDA_2.n2539 GNDA_2.n2538 185
R4645 GNDA_2.n2541 GNDA_2.n1885 185
R4646 GNDA_2.n2543 GNDA_2.n2542 185
R4647 GNDA_2.n2544 GNDA_2.n1884 185
R4648 GNDA_2.n2546 GNDA_2.n2545 185
R4649 GNDA_2.n2548 GNDA_2.n1882 185
R4650 GNDA_2.n2550 GNDA_2.n2549 185
R4651 GNDA_2.n2551 GNDA_2.n1881 185
R4652 GNDA_2.n2553 GNDA_2.n2552 185
R4653 GNDA_2.n1888 GNDA_2.n1887 185
R4654 GNDA_2.n1908 GNDA_2.n1907 185
R4655 GNDA_2.n1905 GNDA_2.n1890 185
R4656 GNDA_2.n1903 GNDA_2.n1902 185
R4657 GNDA_2.n1894 GNDA_2.n1892 185
R4658 GNDA_2.n1893 GNDA_2.n1871 185
R4659 GNDA_2.n2594 GNDA_2.n2593 185
R4660 GNDA_2.n2591 GNDA_2.n1869 185
R4661 GNDA_2.n2590 GNDA_2.n1848 185
R4662 GNDA_2.n2900 GNDA_2.n2899 185
R4663 GNDA_2.n2902 GNDA_2.n2901 185
R4664 GNDA_2.n2904 GNDA_2.n2903 185
R4665 GNDA_2.n2906 GNDA_2.n2905 185
R4666 GNDA_2.n2908 GNDA_2.n2907 185
R4667 GNDA_2.n2910 GNDA_2.n2909 185
R4668 GNDA_2.n2912 GNDA_2.n2911 185
R4669 GNDA_2.n2913 GNDA_2.n2640 185
R4670 GNDA_2.n2915 GNDA_2.n2914 185
R4671 GNDA_2.n2882 GNDA_2.n2881 185
R4672 GNDA_2.n2884 GNDA_2.n2883 185
R4673 GNDA_2.n2886 GNDA_2.n2885 185
R4674 GNDA_2.n2888 GNDA_2.n2887 185
R4675 GNDA_2.n2890 GNDA_2.n2889 185
R4676 GNDA_2.n2892 GNDA_2.n2891 185
R4677 GNDA_2.n2894 GNDA_2.n2893 185
R4678 GNDA_2.n2896 GNDA_2.n2895 185
R4679 GNDA_2.n2898 GNDA_2.n2897 185
R4680 GNDA_2.n2864 GNDA_2.n2863 185
R4681 GNDA_2.n2866 GNDA_2.n2865 185
R4682 GNDA_2.n2868 GNDA_2.n2867 185
R4683 GNDA_2.n2870 GNDA_2.n2869 185
R4684 GNDA_2.n2872 GNDA_2.n2871 185
R4685 GNDA_2.n2874 GNDA_2.n2873 185
R4686 GNDA_2.n2876 GNDA_2.n2875 185
R4687 GNDA_2.n2878 GNDA_2.n2877 185
R4688 GNDA_2.n2880 GNDA_2.n2879 185
R4689 GNDA_2.n2862 GNDA_2.n2861 185
R4690 GNDA_2.n2852 GNDA_2.n2851 185
R4691 GNDA_2.n2850 GNDA_2.n2849 185
R4692 GNDA_2.n2847 GNDA_2.n2846 185
R4693 GNDA_2.n2845 GNDA_2.n2844 185
R4694 GNDA_2.n2650 GNDA_2.n2649 185
R4695 GNDA_2.n2648 GNDA_2.n2623 185
R4696 GNDA_2.n2919 GNDA_2.n2918 185
R4697 GNDA_2.n2622 GNDA_2.n2620 185
R4698 GNDA_2.n2752 GNDA_2.n2751 185
R4699 GNDA_2.n2754 GNDA_2.n2709 185
R4700 GNDA_2.n2757 GNDA_2.n2756 185
R4701 GNDA_2.n2758 GNDA_2.n2708 185
R4702 GNDA_2.n2760 GNDA_2.n2759 185
R4703 GNDA_2.n2762 GNDA_2.n2707 185
R4704 GNDA_2.n2765 GNDA_2.n2764 185
R4705 GNDA_2.n2766 GNDA_2.n2706 185
R4706 GNDA_2.n2771 GNDA_2.n2770 185
R4707 GNDA_2.n2734 GNDA_2.n2714 185
R4708 GNDA_2.n2736 GNDA_2.n2735 185
R4709 GNDA_2.n2738 GNDA_2.n2713 185
R4710 GNDA_2.n2741 GNDA_2.n2740 185
R4711 GNDA_2.n2742 GNDA_2.n2712 185
R4712 GNDA_2.n2744 GNDA_2.n2743 185
R4713 GNDA_2.n2746 GNDA_2.n2711 185
R4714 GNDA_2.n2749 GNDA_2.n2748 185
R4715 GNDA_2.n2750 GNDA_2.n2710 185
R4716 GNDA_2.n2807 GNDA_2.n2806 185
R4717 GNDA_2.n2719 GNDA_2.n2675 185
R4718 GNDA_2.n2721 GNDA_2.n2720 185
R4719 GNDA_2.n2723 GNDA_2.n2717 185
R4720 GNDA_2.n2725 GNDA_2.n2724 185
R4721 GNDA_2.n2726 GNDA_2.n2716 185
R4722 GNDA_2.n2728 GNDA_2.n2727 185
R4723 GNDA_2.n2730 GNDA_2.n2715 185
R4724 GNDA_2.n2733 GNDA_2.n2732 185
R4725 GNDA_2.n2805 GNDA_2.n2674 185
R4726 GNDA_2.n2803 GNDA_2.n2802 185
R4727 GNDA_2.n2678 GNDA_2.n2677 185
R4728 GNDA_2.n2792 GNDA_2.n2791 185
R4729 GNDA_2.n2789 GNDA_2.n2682 185
R4730 GNDA_2.n2787 GNDA_2.n2786 185
R4731 GNDA_2.n2684 GNDA_2.n2683 185
R4732 GNDA_2.n2776 GNDA_2.n2775 185
R4733 GNDA_2.n2773 GNDA_2.n2704 185
R4734 GNDA_2.n2085 GNDA_2.n2084 185
R4735 GNDA_2.n2087 GNDA_2.n2086 185
R4736 GNDA_2.n2089 GNDA_2.n2088 185
R4737 GNDA_2.n2091 GNDA_2.n2090 185
R4738 GNDA_2.n2093 GNDA_2.n2092 185
R4739 GNDA_2.n2095 GNDA_2.n2094 185
R4740 GNDA_2.n2097 GNDA_2.n2096 185
R4741 GNDA_2.n2099 GNDA_2.n2098 185
R4742 GNDA_2.n2100 GNDA_2.n2048 185
R4743 GNDA_2.n2067 GNDA_2.n2066 185
R4744 GNDA_2.n2069 GNDA_2.n2068 185
R4745 GNDA_2.n2071 GNDA_2.n2070 185
R4746 GNDA_2.n2073 GNDA_2.n2072 185
R4747 GNDA_2.n2075 GNDA_2.n2074 185
R4748 GNDA_2.n2077 GNDA_2.n2076 185
R4749 GNDA_2.n2079 GNDA_2.n2078 185
R4750 GNDA_2.n2081 GNDA_2.n2080 185
R4751 GNDA_2.n2083 GNDA_2.n2082 185
R4752 GNDA_2.n2040 GNDA_2.n2026 185
R4753 GNDA_2.n2051 GNDA_2.n2050 185
R4754 GNDA_2.n2053 GNDA_2.n2052 185
R4755 GNDA_2.n2055 GNDA_2.n2054 185
R4756 GNDA_2.n2057 GNDA_2.n2056 185
R4757 GNDA_2.n2059 GNDA_2.n2058 185
R4758 GNDA_2.n2061 GNDA_2.n2060 185
R4759 GNDA_2.n2063 GNDA_2.n2062 185
R4760 GNDA_2.n2065 GNDA_2.n2064 185
R4761 GNDA_2.n2030 GNDA_2.n2027 185
R4762 GNDA_2.n2137 GNDA_2.n2136 185
R4763 GNDA_2.n2110 GNDA_2.n2029 185
R4764 GNDA_2.n2116 GNDA_2.n2115 185
R4765 GNDA_2.n2114 GNDA_2.n2109 185
R4766 GNDA_2.n2123 GNDA_2.n2122 185
R4767 GNDA_2.n2121 GNDA_2.n2108 185
R4768 GNDA_2.n2128 GNDA_2.n2049 185
R4769 GNDA_2.n2133 GNDA_2.n2132 185
R4770 GNDA_2.n5428 GNDA_2.n5427 185
R4771 GNDA_2.n5430 GNDA_2.n5429 185
R4772 GNDA_2.n5432 GNDA_2.n5431 185
R4773 GNDA_2.n5434 GNDA_2.n5433 185
R4774 GNDA_2.n5436 GNDA_2.n5435 185
R4775 GNDA_2.n5438 GNDA_2.n5437 185
R4776 GNDA_2.n5440 GNDA_2.n5439 185
R4777 GNDA_2.n5442 GNDA_2.n5441 185
R4778 GNDA_2.n5443 GNDA_2.n89 185
R4779 GNDA_2.n5410 GNDA_2.n5409 185
R4780 GNDA_2.n5412 GNDA_2.n5411 185
R4781 GNDA_2.n5414 GNDA_2.n5413 185
R4782 GNDA_2.n5416 GNDA_2.n5415 185
R4783 GNDA_2.n5418 GNDA_2.n5417 185
R4784 GNDA_2.n5420 GNDA_2.n5419 185
R4785 GNDA_2.n5422 GNDA_2.n5421 185
R4786 GNDA_2.n5424 GNDA_2.n5423 185
R4787 GNDA_2.n5426 GNDA_2.n5425 185
R4788 GNDA_2.n5392 GNDA_2.n5391 185
R4789 GNDA_2.n5394 GNDA_2.n5393 185
R4790 GNDA_2.n5396 GNDA_2.n5395 185
R4791 GNDA_2.n5398 GNDA_2.n5397 185
R4792 GNDA_2.n5400 GNDA_2.n5399 185
R4793 GNDA_2.n5402 GNDA_2.n5401 185
R4794 GNDA_2.n5404 GNDA_2.n5403 185
R4795 GNDA_2.n5406 GNDA_2.n5405 185
R4796 GNDA_2.n5408 GNDA_2.n5407 185
R4797 GNDA_2.n5390 GNDA_2.n5389 185
R4798 GNDA_2.n5384 GNDA_2.n5383 185
R4799 GNDA_2.n5382 GNDA_2.n5381 185
R4800 GNDA_2.n5377 GNDA_2.n5376 185
R4801 GNDA_2.n5375 GNDA_2.n5374 185
R4802 GNDA_2.n5369 GNDA_2.n5368 185
R4803 GNDA_2.n5364 GNDA_2.n93 185
R4804 GNDA_2.n5447 GNDA_2.n5446 185
R4805 GNDA_2.n92 GNDA_2.n90 185
R4806 GNDA_2.n2301 GNDA_2.n2300 185
R4807 GNDA_2.n2303 GNDA_2.n2302 185
R4808 GNDA_2.n2305 GNDA_2.n2304 185
R4809 GNDA_2.n2307 GNDA_2.n2306 185
R4810 GNDA_2.n2309 GNDA_2.n2308 185
R4811 GNDA_2.n2311 GNDA_2.n2310 185
R4812 GNDA_2.n2313 GNDA_2.n2312 185
R4813 GNDA_2.n2315 GNDA_2.n2314 185
R4814 GNDA_2.n2316 GNDA_2.n2144 185
R4815 GNDA_2.n2283 GNDA_2.n2282 185
R4816 GNDA_2.n2285 GNDA_2.n2284 185
R4817 GNDA_2.n2287 GNDA_2.n2286 185
R4818 GNDA_2.n2289 GNDA_2.n2288 185
R4819 GNDA_2.n2291 GNDA_2.n2290 185
R4820 GNDA_2.n2293 GNDA_2.n2292 185
R4821 GNDA_2.n2295 GNDA_2.n2294 185
R4822 GNDA_2.n2297 GNDA_2.n2296 185
R4823 GNDA_2.n2299 GNDA_2.n2298 185
R4824 GNDA_2.n2265 GNDA_2.n2264 185
R4825 GNDA_2.n2267 GNDA_2.n2266 185
R4826 GNDA_2.n2269 GNDA_2.n2268 185
R4827 GNDA_2.n2271 GNDA_2.n2270 185
R4828 GNDA_2.n2273 GNDA_2.n2272 185
R4829 GNDA_2.n2275 GNDA_2.n2274 185
R4830 GNDA_2.n2277 GNDA_2.n2276 185
R4831 GNDA_2.n2279 GNDA_2.n2278 185
R4832 GNDA_2.n2281 GNDA_2.n2280 185
R4833 GNDA_2.n2263 GNDA_2.n2262 185
R4834 GNDA_2.n2257 GNDA_2.n2256 185
R4835 GNDA_2.n2255 GNDA_2.n2254 185
R4836 GNDA_2.n2250 GNDA_2.n2249 185
R4837 GNDA_2.n2248 GNDA_2.n2247 185
R4838 GNDA_2.n2242 GNDA_2.n2241 185
R4839 GNDA_2.n2237 GNDA_2.n2148 185
R4840 GNDA_2.n2320 GNDA_2.n2319 185
R4841 GNDA_2.n2147 GNDA_2.n2145 185
R4842 GNDA_2.n1764 GNDA_2.n1763 185
R4843 GNDA_2.n1766 GNDA_2.n1765 185
R4844 GNDA_2.n1768 GNDA_2.n1767 185
R4845 GNDA_2.n1770 GNDA_2.n1769 185
R4846 GNDA_2.n1772 GNDA_2.n1771 185
R4847 GNDA_2.n1774 GNDA_2.n1773 185
R4848 GNDA_2.n1776 GNDA_2.n1775 185
R4849 GNDA_2.n1778 GNDA_2.n1777 185
R4850 GNDA_2.n1779 GNDA_2.n1723 185
R4851 GNDA_2.n1746 GNDA_2.n1745 185
R4852 GNDA_2.n1748 GNDA_2.n1747 185
R4853 GNDA_2.n1750 GNDA_2.n1749 185
R4854 GNDA_2.n1752 GNDA_2.n1751 185
R4855 GNDA_2.n1754 GNDA_2.n1753 185
R4856 GNDA_2.n1756 GNDA_2.n1755 185
R4857 GNDA_2.n1758 GNDA_2.n1757 185
R4858 GNDA_2.n1760 GNDA_2.n1759 185
R4859 GNDA_2.n1762 GNDA_2.n1761 185
R4860 GNDA_2.n1715 GNDA_2.n1672 185
R4861 GNDA_2.n1730 GNDA_2.n1729 185
R4862 GNDA_2.n1732 GNDA_2.n1731 185
R4863 GNDA_2.n1734 GNDA_2.n1733 185
R4864 GNDA_2.n1736 GNDA_2.n1735 185
R4865 GNDA_2.n1738 GNDA_2.n1737 185
R4866 GNDA_2.n1740 GNDA_2.n1739 185
R4867 GNDA_2.n1742 GNDA_2.n1741 185
R4868 GNDA_2.n1744 GNDA_2.n1743 185
R4869 GNDA_2.n1714 GNDA_2.n1671 185
R4870 GNDA_2.n1708 GNDA_2.n1707 185
R4871 GNDA_2.n1701 GNDA_2.n1696 185
R4872 GNDA_2.n3365 GNDA_2.n3364 185
R4873 GNDA_2.n3348 GNDA_2.n1695 185
R4874 GNDA_2.n3352 GNDA_2.n3351 185
R4875 GNDA_2.n3350 GNDA_2.n3347 185
R4876 GNDA_2.n1726 GNDA_2.n1724 185
R4877 GNDA_2.n3361 GNDA_2.n3360 185
R4878 GNDA_2.n3381 GNDA_2.n1685 185
R4879 GNDA_2.n3373 GNDA_2.n3372 185
R4880 GNDA_2.n2838 GNDA_2.n2837 185
R4881 GNDA_2.n2837 GNDA_2.n2836 185
R4882 GNDA_2.n2838 GNDA_2.n2828 185
R4883 GNDA_2.n2831 GNDA_2.n2828 185
R4884 GNDA_2.n5336 GNDA_2.n5335 185
R4885 GNDA_2.n5338 GNDA_2.n5337 185
R4886 GNDA_2.n5340 GNDA_2.n5339 185
R4887 GNDA_2.n5342 GNDA_2.n5341 185
R4888 GNDA_2.n5344 GNDA_2.n5343 185
R4889 GNDA_2.n5346 GNDA_2.n5345 185
R4890 GNDA_2.n5348 GNDA_2.n5347 185
R4891 GNDA_2.n5350 GNDA_2.n5349 185
R4892 GNDA_2.n5351 GNDA_2.n20 185
R4893 GNDA_2.n5318 GNDA_2.n5317 185
R4894 GNDA_2.n5320 GNDA_2.n5319 185
R4895 GNDA_2.n5322 GNDA_2.n5321 185
R4896 GNDA_2.n5324 GNDA_2.n5323 185
R4897 GNDA_2.n5326 GNDA_2.n5325 185
R4898 GNDA_2.n5328 GNDA_2.n5327 185
R4899 GNDA_2.n5330 GNDA_2.n5329 185
R4900 GNDA_2.n5332 GNDA_2.n5331 185
R4901 GNDA_2.n5334 GNDA_2.n5333 185
R4902 GNDA_2.n5300 GNDA_2.n5299 185
R4903 GNDA_2.n5302 GNDA_2.n5301 185
R4904 GNDA_2.n5304 GNDA_2.n5303 185
R4905 GNDA_2.n5306 GNDA_2.n5305 185
R4906 GNDA_2.n5308 GNDA_2.n5307 185
R4907 GNDA_2.n5310 GNDA_2.n5309 185
R4908 GNDA_2.n5312 GNDA_2.n5311 185
R4909 GNDA_2.n5314 GNDA_2.n5313 185
R4910 GNDA_2.n5316 GNDA_2.n5315 185
R4911 GNDA_2.n5298 GNDA_2.n5297 185
R4912 GNDA_2.n5292 GNDA_2.n5291 185
R4913 GNDA_2.n5287 GNDA_2.n3 185
R4914 GNDA_2.n5560 GNDA_2.n5559 185
R4915 GNDA_2.n34 GNDA_2.n2 185
R4916 GNDA_2.n38 GNDA_2.n37 185
R4917 GNDA_2.n36 GNDA_2.n33 185
R4918 GNDA_2.n23 GNDA_2.n21 185
R4919 GNDA_2.n5556 GNDA_2.n5555 185
R4920 GNDA_2.n2947 GNDA_2.n2946 175.546
R4921 GNDA_2.n3259 GNDA_2.n2946 175.546
R4922 GNDA_2.n3257 GNDA_2.n3256 175.546
R4923 GNDA_2.n3253 GNDA_2.n3252 175.546
R4924 GNDA_2.n3249 GNDA_2.n3248 175.546
R4925 GNDA_2.n3245 GNDA_2.n3244 175.546
R4926 GNDA_2.n3241 GNDA_2.n2948 175.546
R4927 GNDA_2.n3241 GNDA_2.n2950 175.546
R4928 GNDA_2.n3237 GNDA_2.n2950 175.546
R4929 GNDA_2.n3237 GNDA_2.n2953 175.546
R4930 GNDA_2.n3233 GNDA_2.n2953 175.546
R4931 GNDA_2.n3233 GNDA_2.n2955 175.546
R4932 GNDA_2.n3229 GNDA_2.n2955 175.546
R4933 GNDA_2.n3229 GNDA_2.n2957 175.546
R4934 GNDA_2.n3225 GNDA_2.n2957 175.546
R4935 GNDA_2.n3225 GNDA_2.n2959 175.546
R4936 GNDA_2.n3221 GNDA_2.n2959 175.546
R4937 GNDA_2.n58 GNDA_2.n54 175.546
R4938 GNDA_2.n5540 GNDA_2.n5539 175.546
R4939 GNDA_2.n5466 GNDA_2.n5465 175.546
R4940 GNDA_2.n5471 GNDA_2.n5470 175.546
R4941 GNDA_2.n5479 GNDA_2.n5478 175.546
R4942 GNDA_2.n3181 GNDA_2.n2961 175.546
R4943 GNDA_2.n3182 GNDA_2.n3181 175.546
R4944 GNDA_2.n3185 GNDA_2.n3182 175.546
R4945 GNDA_2.n3186 GNDA_2.n3185 175.546
R4946 GNDA_2.n3206 GNDA_2.n3186 175.546
R4947 GNDA_2.n3206 GNDA_2.n3205 175.546
R4948 GNDA_2.n3205 GNDA_2.n3189 175.546
R4949 GNDA_2.n3193 GNDA_2.n3189 175.546
R4950 GNDA_2.n3194 GNDA_2.n3193 175.546
R4951 GNDA_2.n3194 GNDA_2.n85 175.546
R4952 GNDA_2.n5458 GNDA_2.n85 175.546
R4953 GNDA_2.n1961 GNDA_2.n1960 175.546
R4954 GNDA_2.n1957 GNDA_2.n1956 175.546
R4955 GNDA_2.n1953 GNDA_2.n1952 175.546
R4956 GNDA_2.n1949 GNDA_2.n1948 175.546
R4957 GNDA_2.n1945 GNDA_2.n1944 175.546
R4958 GNDA_2.n1969 GNDA_2.n1968 175.546
R4959 GNDA_2.n1973 GNDA_2.n1972 175.546
R4960 GNDA_2.n1977 GNDA_2.n1976 175.546
R4961 GNDA_2.n1981 GNDA_2.n1980 175.546
R4962 GNDA_2.n1983 GNDA_2.n1943 175.546
R4963 GNDA_2.n2600 GNDA_2.n1849 175.546
R4964 GNDA_2.n2596 GNDA_2.n1867 175.546
R4965 GNDA_2.n1897 GNDA_2.n1896 175.546
R4966 GNDA_2.n1900 GNDA_2.n1899 175.546
R4967 GNDA_2.n1911 GNDA_2.n1910 175.546
R4968 GNDA_2.n2510 GNDA_2.n2509 175.546
R4969 GNDA_2.n1933 GNDA_2.n1932 175.546
R4970 GNDA_2.n2520 GNDA_2.n2519 175.546
R4971 GNDA_2.n1928 GNDA_2.n1923 175.546
R4972 GNDA_2.n2529 GNDA_2.n1917 175.546
R4973 GNDA_2.n3268 GNDA_2.n1830 175.546
R4974 GNDA_2.n2944 GNDA_2.n2612 175.546
R4975 GNDA_2.n2940 GNDA_2.n2939 175.546
R4976 GNDA_2.n2936 GNDA_2.n2935 175.546
R4977 GNDA_2.n2932 GNDA_2.n2931 175.546
R4978 GNDA_2.n3276 GNDA_2.n3274 175.546
R4979 GNDA_2.n3280 GNDA_2.n1826 175.546
R4980 GNDA_2.n3284 GNDA_2.n3282 175.546
R4981 GNDA_2.n3288 GNDA_2.n1824 175.546
R4982 GNDA_2.n3291 GNDA_2.n3290 175.546
R4983 GNDA_2.n2927 GNDA_2.n2615 175.546
R4984 GNDA_2.n2921 GNDA_2.n2615 175.546
R4985 GNDA_2.n2921 GNDA_2.n2618 175.546
R4986 GNDA_2.n2652 GNDA_2.n2618 175.546
R4987 GNDA_2.n2656 GNDA_2.n2652 175.546
R4988 GNDA_2.n2842 GNDA_2.n2656 175.546
R4989 GNDA_2.n2842 GNDA_2.n2646 175.546
R4990 GNDA_2.n2854 GNDA_2.n2646 175.546
R4991 GNDA_2.n2854 GNDA_2.n2644 175.546
R4992 GNDA_2.n2859 GNDA_2.n2644 175.546
R4993 GNDA_2.n2859 GNDA_2.n1807 175.546
R4994 GNDA_2.n3304 GNDA_2.n1818 175.546
R4995 GNDA_2.n3308 GNDA_2.n3306 175.546
R4996 GNDA_2.n3316 GNDA_2.n1814 175.546
R4997 GNDA_2.n3320 GNDA_2.n3318 175.546
R4998 GNDA_2.n3328 GNDA_2.n1810 175.546
R4999 GNDA_2.n3302 GNDA_2.n3300 175.546
R5000 GNDA_2.n3310 GNDA_2.n1816 175.546
R5001 GNDA_2.n3314 GNDA_2.n3312 175.546
R5002 GNDA_2.n3322 GNDA_2.n1812 175.546
R5003 GNDA_2.n3326 GNDA_2.n3324 175.546
R5004 GNDA_2.n2436 GNDA_2.n2432 175.546
R5005 GNDA_2.n2440 GNDA_2.n2438 175.546
R5006 GNDA_2.n2444 GNDA_2.n2429 175.546
R5007 GNDA_2.n2447 GNDA_2.n2446 175.546
R5008 GNDA_2.n2451 GNDA_2.n2450 175.546
R5009 GNDA_2.n2703 GNDA_2.n1805 175.546
R5010 GNDA_2.n2778 GNDA_2.n2703 175.546
R5011 GNDA_2.n2778 GNDA_2.n2685 175.546
R5012 GNDA_2.n2783 GNDA_2.n2685 175.546
R5013 GNDA_2.n2783 GNDA_2.n2680 175.546
R5014 GNDA_2.n2794 GNDA_2.n2680 175.546
R5015 GNDA_2.n2794 GNDA_2.n2679 175.546
R5016 GNDA_2.n2799 GNDA_2.n2679 175.546
R5017 GNDA_2.n2799 GNDA_2.n2673 175.546
R5018 GNDA_2.n2811 GNDA_2.n2673 175.546
R5019 GNDA_2.n2811 GNDA_2.n1783 175.546
R5020 GNDA_2.n2392 GNDA_2.n2391 175.546
R5021 GNDA_2.n2394 GNDA_2.n2393 175.546
R5022 GNDA_2.n2398 GNDA_2.n2397 175.546
R5023 GNDA_2.n2400 GNDA_2.n2399 175.546
R5024 GNDA_2.n2404 GNDA_2.n1786 175.546
R5025 GNDA_2.n2512 GNDA_2.n1934 175.546
R5026 GNDA_2.n2516 GNDA_2.n2514 175.546
R5027 GNDA_2.n2522 GNDA_2.n1930 175.546
R5028 GNDA_2.n2525 GNDA_2.n2524 175.546
R5029 GNDA_2.n2527 GNDA_2.n1926 175.546
R5030 GNDA_2.n2502 GNDA_2.n1990 175.546
R5031 GNDA_2.n2498 GNDA_2.n2497 175.546
R5032 GNDA_2.n2495 GNDA_2.n1993 175.546
R5033 GNDA_2.n2491 GNDA_2.n2490 175.546
R5034 GNDA_2.n2488 GNDA_2.n1996 175.546
R5035 GNDA_2.n2130 GNDA_2.n2129 175.546
R5036 GNDA_2.n2126 GNDA_2.n2125 175.546
R5037 GNDA_2.n2119 GNDA_2.n2118 175.546
R5038 GNDA_2.n2112 GNDA_2.n2111 175.546
R5039 GNDA_2.n2140 GNDA_2.n2139 175.546
R5040 GNDA_2.n2010 GNDA_2.n2009 175.546
R5041 GNDA_2.n2012 GNDA_2.n2011 175.546
R5042 GNDA_2.n2014 GNDA_2.n2013 175.546
R5043 GNDA_2.n2016 GNDA_2.n2015 175.546
R5044 GNDA_2.n2018 GNDA_2.n2017 175.546
R5045 GNDA_2.n3217 GNDA_2.n3180 175.546
R5046 GNDA_2.n3213 GNDA_2.n3180 175.546
R5047 GNDA_2.n3213 GNDA_2.n3184 175.546
R5048 GNDA_2.n3209 GNDA_2.n3184 175.546
R5049 GNDA_2.n3209 GNDA_2.n3188 175.546
R5050 GNDA_2.n3203 GNDA_2.n3188 175.546
R5051 GNDA_2.n3203 GNDA_2.n3202 175.546
R5052 GNDA_2.n3202 GNDA_2.n3192 175.546
R5053 GNDA_2.n3198 GNDA_2.n3192 175.546
R5054 GNDA_2.n3198 GNDA_2.n88 175.546
R5055 GNDA_2.n5456 GNDA_2.n88 175.546
R5056 GNDA_2.n3179 GNDA_2.n2964 175.546
R5057 GNDA_2.n3175 GNDA_2.n2964 175.546
R5058 GNDA_2.n3175 GNDA_2.n2966 175.546
R5059 GNDA_2.n3171 GNDA_2.n2966 175.546
R5060 GNDA_2.n3171 GNDA_2.n2969 175.546
R5061 GNDA_2.n3164 GNDA_2.n2969 175.546
R5062 GNDA_2.n3164 GNDA_2.n3163 175.546
R5063 GNDA_2.n3163 GNDA_2.n3071 175.546
R5064 GNDA_2.n3159 GNDA_2.n3071 175.546
R5065 GNDA_2.n3159 GNDA_2.n3073 175.546
R5066 GNDA_2.n3155 GNDA_2.n3073 175.546
R5067 GNDA_2.n5450 GNDA_2.n5449 175.546
R5068 GNDA_2.n5366 GNDA_2.n5365 175.546
R5069 GNDA_2.n5372 GNDA_2.n5371 175.546
R5070 GNDA_2.n5379 GNDA_2.n5378 175.546
R5071 GNDA_2.n5387 GNDA_2.n5386 175.546
R5072 GNDA_2.n3080 GNDA_2.n3076 175.546
R5073 GNDA_2.n3081 GNDA_2.n3080 175.546
R5074 GNDA_2.n3085 GNDA_2.n3081 175.546
R5075 GNDA_2.n3086 GNDA_2.n3085 175.546
R5076 GNDA_2.n3089 GNDA_2.n3086 175.546
R5077 GNDA_2.n3090 GNDA_2.n3089 175.546
R5078 GNDA_2.n3093 GNDA_2.n3090 175.546
R5079 GNDA_2.n3094 GNDA_2.n3093 175.546
R5080 GNDA_2.n3097 GNDA_2.n3094 175.546
R5081 GNDA_2.n3097 GNDA_2.n112 175.546
R5082 GNDA_2.n5358 GNDA_2.n112 175.546
R5083 GNDA_2.n2478 GNDA_2.n2002 175.546
R5084 GNDA_2.n2478 GNDA_2.n2008 175.546
R5085 GNDA_2.n2474 GNDA_2.n2473 175.546
R5086 GNDA_2.n2470 GNDA_2.n2469 175.546
R5087 GNDA_2.n2466 GNDA_2.n2465 175.546
R5088 GNDA_2.n2462 GNDA_2.n2007 175.546
R5089 GNDA_2.n2186 GNDA_2.n2184 175.546
R5090 GNDA_2.n2190 GNDA_2.n2180 175.546
R5091 GNDA_2.n2194 GNDA_2.n2192 175.546
R5092 GNDA_2.n2198 GNDA_2.n2178 175.546
R5093 GNDA_2.n2201 GNDA_2.n2200 175.546
R5094 GNDA_2.n2323 GNDA_2.n2322 175.546
R5095 GNDA_2.n2239 GNDA_2.n2238 175.546
R5096 GNDA_2.n2245 GNDA_2.n2244 175.546
R5097 GNDA_2.n2252 GNDA_2.n2251 175.546
R5098 GNDA_2.n2260 GNDA_2.n2259 175.546
R5099 GNDA_2.n2208 GNDA_2.n2205 175.546
R5100 GNDA_2.n2208 GNDA_2.n2174 175.546
R5101 GNDA_2.n2213 GNDA_2.n2174 175.546
R5102 GNDA_2.n2213 GNDA_2.n2171 175.546
R5103 GNDA_2.n2217 GNDA_2.n2171 175.546
R5104 GNDA_2.n2218 GNDA_2.n2217 175.546
R5105 GNDA_2.n2221 GNDA_2.n2218 175.546
R5106 GNDA_2.n2221 GNDA_2.n2169 175.546
R5107 GNDA_2.n2226 GNDA_2.n2169 175.546
R5108 GNDA_2.n2226 GNDA_2.n2167 175.546
R5109 GNDA_2.n2230 GNDA_2.n2167 175.546
R5110 GNDA_2.n2422 GNDA_2.n2421 175.546
R5111 GNDA_2.n2418 GNDA_2.n2417 175.546
R5112 GNDA_2.n2415 GNDA_2.n2396 175.546
R5113 GNDA_2.n2411 GNDA_2.n2409 175.546
R5114 GNDA_2.n2407 GNDA_2.n2403 175.546
R5115 GNDA_2.n2387 GNDA_2.n2331 175.546
R5116 GNDA_2.n2383 GNDA_2.n2382 175.546
R5117 GNDA_2.n2380 GNDA_2.n2334 175.546
R5118 GNDA_2.n2376 GNDA_2.n2375 175.546
R5119 GNDA_2.n2373 GNDA_2.n2337 175.546
R5120 GNDA_2.n3344 GNDA_2.n1727 175.546
R5121 GNDA_2.n3358 GNDA_2.n3344 175.546
R5122 GNDA_2.n3358 GNDA_2.n3345 175.546
R5123 GNDA_2.n3354 GNDA_2.n3345 175.546
R5124 GNDA_2.n3354 GNDA_2.n1692 175.546
R5125 GNDA_2.n3367 GNDA_2.n1692 175.546
R5126 GNDA_2.n3367 GNDA_2.n1693 175.546
R5127 GNDA_2.n1704 GNDA_2.n1693 175.546
R5128 GNDA_2.n1704 GNDA_2.n1669 175.546
R5129 GNDA_2.n3401 GNDA_2.n1669 175.546
R5130 GNDA_2.n3401 GNDA_2.n1670 175.546
R5131 GNDA_2.n2368 GNDA_2.n2340 175.546
R5132 GNDA_2.n2364 GNDA_2.n2340 175.546
R5133 GNDA_2.n2364 GNDA_2.n2342 175.546
R5134 GNDA_2.n2360 GNDA_2.n2342 175.546
R5135 GNDA_2.n2360 GNDA_2.n2358 175.546
R5136 GNDA_2.n2358 GNDA_2.n2357 175.546
R5137 GNDA_2.n2357 GNDA_2.n2345 175.546
R5138 GNDA_2.n2353 GNDA_2.n2345 175.546
R5139 GNDA_2.n2353 GNDA_2.n2347 175.546
R5140 GNDA_2.n2349 GNDA_2.n2347 175.546
R5141 GNDA_2.n2349 GNDA_2.n1674 175.546
R5142 GNDA_2.n3117 GNDA_2.n3079 175.546
R5143 GNDA_2.n3113 GNDA_2.n3079 175.546
R5144 GNDA_2.n3113 GNDA_2.n3083 175.546
R5145 GNDA_2.n3109 GNDA_2.n3083 175.546
R5146 GNDA_2.n3109 GNDA_2.n3088 175.546
R5147 GNDA_2.n3105 GNDA_2.n3088 175.546
R5148 GNDA_2.n3105 GNDA_2.n3092 175.546
R5149 GNDA_2.n3101 GNDA_2.n3092 175.546
R5150 GNDA_2.n3101 GNDA_2.n3096 175.546
R5151 GNDA_2.n3096 GNDA_2.n115 175.546
R5152 GNDA_2.n5356 GNDA_2.n115 175.546
R5153 GNDA_2.n3151 GNDA_2.n3118 175.546
R5154 GNDA_2.n3147 GNDA_2.n3118 175.546
R5155 GNDA_2.n3147 GNDA_2.n3120 175.546
R5156 GNDA_2.n3143 GNDA_2.n3120 175.546
R5157 GNDA_2.n3143 GNDA_2.n3122 175.546
R5158 GNDA_2.n3139 GNDA_2.n3122 175.546
R5159 GNDA_2.n3139 GNDA_2.n3124 175.546
R5160 GNDA_2.n3135 GNDA_2.n3124 175.546
R5161 GNDA_2.n3135 GNDA_2.n3126 175.546
R5162 GNDA_2.n3131 GNDA_2.n3126 175.546
R5163 GNDA_2.n3131 GNDA_2.n3128 175.546
R5164 GNDA_2.n5553 GNDA_2.n24 175.546
R5165 GNDA_2.n40 GNDA_2.n25 175.546
R5166 GNDA_2.n31 GNDA_2.n30 175.546
R5167 GNDA_2.n5289 GNDA_2.n5288 175.546
R5168 GNDA_2.n5295 GNDA_2.n5294 175.546
R5169 GNDA_2.n5259 GNDA_2.n127 175.546
R5170 GNDA_2.n5259 GNDA_2.n125 175.546
R5171 GNDA_2.n5264 GNDA_2.n125 175.546
R5172 GNDA_2.n5264 GNDA_2.n122 175.546
R5173 GNDA_2.n5268 GNDA_2.n122 175.546
R5174 GNDA_2.n5269 GNDA_2.n5268 175.546
R5175 GNDA_2.n5272 GNDA_2.n5269 175.546
R5176 GNDA_2.n5272 GNDA_2.n120 175.546
R5177 GNDA_2.n5277 GNDA_2.n120 175.546
R5178 GNDA_2.n5277 GNDA_2.n118 175.546
R5179 GNDA_2.n5281 GNDA_2.n118 175.546
R5180 GNDA_2.n2531 GNDA_2.n1918 173.881
R5181 GNDA_2.n2023 GNDA_2.t73 172.876
R5182 GNDA_2.n2479 GNDA_2.t73 172.615
R5183 GNDA_2.n1927 GNDA_2.n1918 171.624
R5184 GNDA_2.n4372 GNDA_2.n4371 166.4
R5185 GNDA_2.n4367 GNDA_2.n4366 166.4
R5186 GNDA_2.n5483 GNDA_2.n5482 163.333
R5187 GNDA_2.n2539 GNDA_2.n1887 163.333
R5188 GNDA_2.n2863 GNDA_2.n2862 163.333
R5189 GNDA_2.n2806 GNDA_2.n2805 163.333
R5190 GNDA_2.n2040 GNDA_2.n2030 163.333
R5191 GNDA_2.n5391 GNDA_2.n5390 163.333
R5192 GNDA_2.n2264 GNDA_2.n2263 163.333
R5193 GNDA_2.n1715 GNDA_2.n1714 163.333
R5194 GNDA_2.n5299 GNDA_2.n5298 163.333
R5195 GNDA_2.n3168 GNDA_2.n2972 157.601
R5196 GNDA_2.n5515 GNDA_2.n5514 150
R5197 GNDA_2.n5511 GNDA_2.n5510 150
R5198 GNDA_2.n5507 GNDA_2.n5506 150
R5199 GNDA_2.n5503 GNDA_2.n5502 150
R5200 GNDA_2.n5499 GNDA_2.n5498 150
R5201 GNDA_2.n5495 GNDA_2.n5494 150
R5202 GNDA_2.n5491 GNDA_2.n5490 150
R5203 GNDA_2.n5487 GNDA_2.n5486 150
R5204 GNDA_2.n5544 GNDA_2.n5543 150
R5205 GNDA_2.n5536 GNDA_2.n64 150
R5206 GNDA_2.n5468 GNDA_2.n65 150
R5207 GNDA_2.n5475 GNDA_2.n5474 150
R5208 GNDA_2.n5533 GNDA_2.n81 150
R5209 GNDA_2.n5529 GNDA_2.n5528 150
R5210 GNDA_2.n5525 GNDA_2.n5524 150
R5211 GNDA_2.n5521 GNDA_2.n5520 150
R5212 GNDA_2.n2569 GNDA_2.n1877 150
R5213 GNDA_2.n2565 GNDA_2.n2563 150
R5214 GNDA_2.n2561 GNDA_2.n1879 150
R5215 GNDA_2.n2557 GNDA_2.n2555 150
R5216 GNDA_2.n2553 GNDA_2.n1881 150
R5217 GNDA_2.n2549 GNDA_2.n2548 150
R5218 GNDA_2.n2546 GNDA_2.n1884 150
R5219 GNDA_2.n2542 GNDA_2.n2541 150
R5220 GNDA_2.n2591 GNDA_2.n2590 150
R5221 GNDA_2.n2593 GNDA_2.n1871 150
R5222 GNDA_2.n1903 GNDA_2.n1892 150
R5223 GNDA_2.n1907 GNDA_2.n1905 150
R5224 GNDA_2.n2577 GNDA_2.n1875 150
R5225 GNDA_2.n2581 GNDA_2.n2579 150
R5226 GNDA_2.n2585 GNDA_2.n1873 150
R5227 GNDA_2.n2588 GNDA_2.n2587 150
R5228 GNDA_2.n2895 GNDA_2.n2894 150
R5229 GNDA_2.n2891 GNDA_2.n2890 150
R5230 GNDA_2.n2887 GNDA_2.n2886 150
R5231 GNDA_2.n2883 GNDA_2.n2882 150
R5232 GNDA_2.n2879 GNDA_2.n2878 150
R5233 GNDA_2.n2875 GNDA_2.n2874 150
R5234 GNDA_2.n2871 GNDA_2.n2870 150
R5235 GNDA_2.n2867 GNDA_2.n2866 150
R5236 GNDA_2.n2918 GNDA_2.n2622 150
R5237 GNDA_2.n2649 GNDA_2.n2623 150
R5238 GNDA_2.n2846 GNDA_2.n2845 150
R5239 GNDA_2.n2851 GNDA_2.n2850 150
R5240 GNDA_2.n2903 GNDA_2.n2902 150
R5241 GNDA_2.n2907 GNDA_2.n2906 150
R5242 GNDA_2.n2911 GNDA_2.n2910 150
R5243 GNDA_2.n2915 GNDA_2.n2640 150
R5244 GNDA_2.n2748 GNDA_2.n2746 150
R5245 GNDA_2.n2744 GNDA_2.n2712 150
R5246 GNDA_2.n2740 GNDA_2.n2738 150
R5247 GNDA_2.n2736 GNDA_2.n2714 150
R5248 GNDA_2.n2732 GNDA_2.n2730 150
R5249 GNDA_2.n2728 GNDA_2.n2716 150
R5250 GNDA_2.n2724 GNDA_2.n2723 150
R5251 GNDA_2.n2721 GNDA_2.n2719 150
R5252 GNDA_2.n2775 GNDA_2.n2773 150
R5253 GNDA_2.n2787 GNDA_2.n2683 150
R5254 GNDA_2.n2791 GNDA_2.n2789 150
R5255 GNDA_2.n2803 GNDA_2.n2677 150
R5256 GNDA_2.n2756 GNDA_2.n2754 150
R5257 GNDA_2.n2760 GNDA_2.n2708 150
R5258 GNDA_2.n2764 GNDA_2.n2762 150
R5259 GNDA_2.n2771 GNDA_2.n2706 150
R5260 GNDA_2.n2080 GNDA_2.n2079 150
R5261 GNDA_2.n2076 GNDA_2.n2075 150
R5262 GNDA_2.n2072 GNDA_2.n2071 150
R5263 GNDA_2.n2068 GNDA_2.n2067 150
R5264 GNDA_2.n2064 GNDA_2.n2063 150
R5265 GNDA_2.n2060 GNDA_2.n2059 150
R5266 GNDA_2.n2056 GNDA_2.n2055 150
R5267 GNDA_2.n2052 GNDA_2.n2051 150
R5268 GNDA_2.n2133 GNDA_2.n2049 150
R5269 GNDA_2.n2122 GNDA_2.n2121 150
R5270 GNDA_2.n2115 GNDA_2.n2114 150
R5271 GNDA_2.n2136 GNDA_2.n2029 150
R5272 GNDA_2.n2088 GNDA_2.n2087 150
R5273 GNDA_2.n2092 GNDA_2.n2091 150
R5274 GNDA_2.n2096 GNDA_2.n2095 150
R5275 GNDA_2.n2098 GNDA_2.n2048 150
R5276 GNDA_2.n5423 GNDA_2.n5422 150
R5277 GNDA_2.n5419 GNDA_2.n5418 150
R5278 GNDA_2.n5415 GNDA_2.n5414 150
R5279 GNDA_2.n5411 GNDA_2.n5410 150
R5280 GNDA_2.n5407 GNDA_2.n5406 150
R5281 GNDA_2.n5403 GNDA_2.n5402 150
R5282 GNDA_2.n5399 GNDA_2.n5398 150
R5283 GNDA_2.n5395 GNDA_2.n5394 150
R5284 GNDA_2.n5446 GNDA_2.n92 150
R5285 GNDA_2.n5368 GNDA_2.n93 150
R5286 GNDA_2.n5376 GNDA_2.n5375 150
R5287 GNDA_2.n5383 GNDA_2.n5382 150
R5288 GNDA_2.n5431 GNDA_2.n5430 150
R5289 GNDA_2.n5435 GNDA_2.n5434 150
R5290 GNDA_2.n5439 GNDA_2.n5438 150
R5291 GNDA_2.n5443 GNDA_2.n5442 150
R5292 GNDA_2.n2296 GNDA_2.n2295 150
R5293 GNDA_2.n2292 GNDA_2.n2291 150
R5294 GNDA_2.n2288 GNDA_2.n2287 150
R5295 GNDA_2.n2284 GNDA_2.n2283 150
R5296 GNDA_2.n2280 GNDA_2.n2279 150
R5297 GNDA_2.n2276 GNDA_2.n2275 150
R5298 GNDA_2.n2272 GNDA_2.n2271 150
R5299 GNDA_2.n2268 GNDA_2.n2267 150
R5300 GNDA_2.n2319 GNDA_2.n2147 150
R5301 GNDA_2.n2241 GNDA_2.n2148 150
R5302 GNDA_2.n2249 GNDA_2.n2248 150
R5303 GNDA_2.n2256 GNDA_2.n2255 150
R5304 GNDA_2.n2304 GNDA_2.n2303 150
R5305 GNDA_2.n2308 GNDA_2.n2307 150
R5306 GNDA_2.n2312 GNDA_2.n2311 150
R5307 GNDA_2.n2316 GNDA_2.n2315 150
R5308 GNDA_2.n1759 GNDA_2.n1758 150
R5309 GNDA_2.n1755 GNDA_2.n1754 150
R5310 GNDA_2.n1751 GNDA_2.n1750 150
R5311 GNDA_2.n1747 GNDA_2.n1746 150
R5312 GNDA_2.n1743 GNDA_2.n1742 150
R5313 GNDA_2.n1739 GNDA_2.n1738 150
R5314 GNDA_2.n1735 GNDA_2.n1734 150
R5315 GNDA_2.n1731 GNDA_2.n1730 150
R5316 GNDA_2.n3361 GNDA_2.n1724 150
R5317 GNDA_2.n3351 GNDA_2.n3350 150
R5318 GNDA_2.n3364 GNDA_2.n1695 150
R5319 GNDA_2.n1708 GNDA_2.n1696 150
R5320 GNDA_2.n1767 GNDA_2.n1766 150
R5321 GNDA_2.n1771 GNDA_2.n1770 150
R5322 GNDA_2.n1775 GNDA_2.n1774 150
R5323 GNDA_2.n1777 GNDA_2.n1723 150
R5324 GNDA_2.n5331 GNDA_2.n5330 150
R5325 GNDA_2.n5327 GNDA_2.n5326 150
R5326 GNDA_2.n5323 GNDA_2.n5322 150
R5327 GNDA_2.n5319 GNDA_2.n5318 150
R5328 GNDA_2.n5315 GNDA_2.n5314 150
R5329 GNDA_2.n5311 GNDA_2.n5310 150
R5330 GNDA_2.n5307 GNDA_2.n5306 150
R5331 GNDA_2.n5303 GNDA_2.n5302 150
R5332 GNDA_2.n5556 GNDA_2.n21 150
R5333 GNDA_2.n37 GNDA_2.n36 150
R5334 GNDA_2.n5559 GNDA_2.n2 150
R5335 GNDA_2.n5291 GNDA_2.n3 150
R5336 GNDA_2.n5339 GNDA_2.n5338 150
R5337 GNDA_2.n5343 GNDA_2.n5342 150
R5338 GNDA_2.n5347 GNDA_2.n5346 150
R5339 GNDA_2.n5349 GNDA_2.n20 150
R5340 GNDA_2.n5255 GNDA_2.n5254 148.017
R5341 GNDA_2.n4469 GNDA_2.n4468 148.017
R5342 GNDA_2.n4408 GNDA_2.n4407 148.017
R5343 GNDA_2.n4317 GNDA_2.n4316 148.017
R5344 GNDA_2.n3406 GNDA_2.n1666 136.145
R5345 GNDA_2.n3407 GNDA_2.n1665 136.145
R5346 GNDA_2.n3408 GNDA_2.n1664 136.145
R5347 GNDA_2.n3411 GNDA_2.n1661 136.145
R5348 GNDA_2.n3412 GNDA_2.n1660 136.145
R5349 GNDA_2.n3413 GNDA_2.n1659 136.145
R5350 GNDA_2.n3416 GNDA_2.n1656 136.145
R5351 GNDA_2.n3417 GNDA_2.n1655 136.145
R5352 GNDA_2.n3418 GNDA_2.n1654 136.145
R5353 GNDA_2.n3421 GNDA_2.n1651 136.145
R5354 GNDA_2.n3422 GNDA_2.n1650 136.145
R5355 GNDA_2.n2837 GNDA_2.n2830 134.268
R5356 GNDA_2.n2830 GNDA_2.n2828 134.268
R5357 GNDA_2.n2605 GNDA_2.n1844 132.721
R5358 GNDA_2.n2613 GNDA_2.n2608 132.721
R5359 GNDA_2.n1831 GNDA_2.t67 130.001
R5360 GNDA_2.n3404 GNDA_2.t140 130.001
R5361 GNDA_2.n1798 GNDA_2.t82 130.001
R5362 GNDA_2.n2813 GNDA_2.t148 130.001
R5363 GNDA_2.n2700 GNDA_2.t118 130.001
R5364 GNDA_2.n1802 GNDA_2.t79 130.001
R5365 GNDA_2.n2616 GNDA_2.t163 130.001
R5366 GNDA_2.n2923 GNDA_2.t132 130.001
R5367 GNDA_2.n5270 GNDA_2.t73 127.219
R5368 GNDA_2.n2219 GNDA_2.t73 127.219
R5369 GNDA_2.t73 GNDA_2.n1691 127.219
R5370 GNDA_2.n5459 GNDA_2.n5458 124.832
R5371 GNDA_2.n2534 GNDA_2.n2533 124.832
R5372 GNDA_2.n3331 GNDA_2.n3330 124.832
R5373 GNDA_2.n3333 GNDA_2.n1804 124.832
R5374 GNDA_2.n3338 GNDA_2.n3337 124.832
R5375 GNDA_2.n2103 GNDA_2.n2102 124.832
R5376 GNDA_2.n2328 GNDA_2.n2025 124.832
R5377 GNDA_2.n5456 GNDA_2.n5455 124.832
R5378 GNDA_2.n5359 GNDA_2.n5358 124.832
R5379 GNDA_2.n2458 GNDA_2.n2007 124.832
R5380 GNDA_2.n3340 GNDA_2.n1728 124.832
R5381 GNDA_2.n5356 GNDA_2.n5355 124.832
R5382 GNDA_2.n5231 GNDA_2.n5229 121.251
R5383 GNDA_2.n3984 GNDA_2.n3982 121.251
R5384 GNDA_2.n5239 GNDA_2.n5238 121.136
R5385 GNDA_2.n5237 GNDA_2.n5236 121.136
R5386 GNDA_2.n5235 GNDA_2.n5234 121.136
R5387 GNDA_2.n5233 GNDA_2.n5232 121.136
R5388 GNDA_2.n5231 GNDA_2.n5230 121.136
R5389 GNDA_2.n3984 GNDA_2.n3983 121.136
R5390 GNDA_2.n3986 GNDA_2.n3985 121.136
R5391 GNDA_2.n3988 GNDA_2.n3987 121.136
R5392 GNDA_2.n3990 GNDA_2.n3989 121.136
R5393 GNDA_2.n3992 GNDA_2.n3991 121.136
R5394 GNDA_2.n3064 GNDA_2.t175 111.799
R5395 GNDA_2.n3065 GNDA_2.t17 111.331
R5396 GNDA_2.n3430 GNDA_2.t195 111.206
R5397 GNDA_2.n3430 GNDA_2.t281 111.076
R5398 GNDA_2.n3222 GNDA_2.n2960 105.719
R5399 GNDA_2.n3154 GNDA_2.n3153 105.719
R5400 GNDA_2.n3178 GNDA_2.n2960 103.457
R5401 GNDA_2.n3153 GNDA_2.n3152 103.457
R5402 GNDA_2.n3369 GNDA_2.n1688 101.718
R5403 GNDA_2.n2833 GNDA_2.n2657 101.718
R5404 GNDA_2.n2839 GNDA_2.n2659 101.718
R5405 GNDA_2.n3380 GNDA_2.n1686 101.718
R5406 GNDA_2.n1800 GNDA_2.t73 47.6748
R5407 GNDA_2.n4369 GNDA_2.t52 97.7783
R5408 GNDA_2.n4342 GNDA_2.n4341 92.8005
R5409 GNDA_2.n597 GNDA_2.n384 92.8005
R5410 GNDA_2.n3376 GNDA_2.n1685 91.069
R5411 GNDA_2.n3371 GNDA_2.n1685 91.069
R5412 GNDA_2.n3373 GNDA_2.n1684 91.069
R5413 GNDA_2.n3374 GNDA_2.n3373 91.069
R5414 GNDA_2.n2837 GNDA_2.n2832 91.069
R5415 GNDA_2.n2835 GNDA_2.n2828 91.069
R5416 GNDA_2.n2926 GNDA_2.n2925 90.1439
R5417 GNDA_2.n2855 GNDA_2.n2645 90.1439
R5418 GNDA_2.n2779 GNDA_2.n2702 90.1439
R5419 GNDA_2.n3356 GNDA_2.n3355 90.1439
R5420 GNDA_2.n1703 GNDA_2.n1667 90.1439
R5421 GNDA_2.n3402 GNDA_2.n1668 90.1439
R5422 GNDA_2.n4348 GNDA_2.n381 89.6005
R5423 GNDA_2.n4354 GNDA_2.n4348 89.6005
R5424 GNDA_2.n2922 GNDA_2.n2617 87.1391
R5425 GNDA_2.t73 GNDA_2.n3334 87.1391
R5426 GNDA_2.n2698 GNDA_2.n2688 84.306
R5427 GNDA_2.n2817 GNDA_2.n2672 84.306
R5428 GNDA_2.n2654 GNDA_2.t201 83.1328
R5429 GNDA_2.n2841 GNDA_2.t254 82.1312
R5430 GNDA_2.n2782 GNDA_2.t221 82.1312
R5431 GNDA_2.n3357 GNDA_2.t231 82.1312
R5432 GNDA_2.n3153 GNDA_2.n3077 80.9821
R5433 GNDA_2.n3216 GNDA_2.n2960 80.9821
R5434 GNDA_2.n1676 GNDA_2.t258 78.5658
R5435 GNDA_2.n2856 GNDA_2.t11 78.1248
R5436 GNDA_2.n2796 GNDA_2.t44 78.1248
R5437 GNDA_2.t272 GNDA_2.n1687 78.1248
R5438 GNDA_2.n1918 GNDA_2.t73 76.3879
R5439 GNDA_2.n3265 GNDA_2.n3264 76.3222
R5440 GNDA_2.n3259 GNDA_2.n1834 76.3222
R5441 GNDA_2.n3256 GNDA_2.n1835 76.3222
R5442 GNDA_2.n3252 GNDA_2.n1836 76.3222
R5443 GNDA_2.n3248 GNDA_2.n1837 76.3222
R5444 GNDA_2.n5550 GNDA_2.n5549 76.3222
R5445 GNDA_2.n58 GNDA_2.n53 76.3222
R5446 GNDA_2.n5539 GNDA_2.n52 76.3222
R5447 GNDA_2.n5466 GNDA_2.n51 76.3222
R5448 GNDA_2.n5470 GNDA_2.n50 76.3222
R5449 GNDA_2.n5479 GNDA_2.n49 76.3222
R5450 GNDA_2.n1964 GNDA_2.n1839 76.3222
R5451 GNDA_2.n1960 GNDA_2.n1840 76.3222
R5452 GNDA_2.n1956 GNDA_2.n1841 76.3222
R5453 GNDA_2.n1952 GNDA_2.n1842 76.3222
R5454 GNDA_2.n1948 GNDA_2.n1843 76.3222
R5455 GNDA_2.n1944 GNDA_2.n1844 76.3222
R5456 GNDA_2.n1968 GNDA_2.n1938 76.3222
R5457 GNDA_2.n1972 GNDA_2.n1939 76.3222
R5458 GNDA_2.n1976 GNDA_2.n1940 76.3222
R5459 GNDA_2.n1980 GNDA_2.n1941 76.3222
R5460 GNDA_2.n1983 GNDA_2.n1942 76.3222
R5461 GNDA_2.n1988 GNDA_2.n1987 76.3222
R5462 GNDA_2.n2599 GNDA_2.n1845 76.3222
R5463 GNDA_2.n2597 GNDA_2.n1849 76.3222
R5464 GNDA_2.n1867 GNDA_2.n1866 76.3222
R5465 GNDA_2.n1897 GNDA_2.n1865 76.3222
R5466 GNDA_2.n1899 GNDA_2.n1864 76.3222
R5467 GNDA_2.n1911 GNDA_2.n1863 76.3222
R5468 GNDA_2.n1936 GNDA_2.n1919 76.3222
R5469 GNDA_2.n2510 GNDA_2.n1920 76.3222
R5470 GNDA_2.n1933 GNDA_2.n1921 76.3222
R5471 GNDA_2.n2520 GNDA_2.n1922 76.3222
R5472 GNDA_2.n2530 GNDA_2.n1923 76.3222
R5473 GNDA_2.n2532 GNDA_2.n1917 76.3222
R5474 GNDA_2.n3267 GNDA_2.n1828 76.3222
R5475 GNDA_2.n2945 GNDA_2.n1830 76.3222
R5476 GNDA_2.n2612 GNDA_2.n2611 76.3222
R5477 GNDA_2.n2939 GNDA_2.n2610 76.3222
R5478 GNDA_2.n2935 GNDA_2.n2609 76.3222
R5479 GNDA_2.n2931 GNDA_2.n2608 76.3222
R5480 GNDA_2.n3274 GNDA_2.n3273 76.3222
R5481 GNDA_2.n3275 GNDA_2.n1826 76.3222
R5482 GNDA_2.n3282 GNDA_2.n3281 76.3222
R5483 GNDA_2.n3283 GNDA_2.n1824 76.3222
R5484 GNDA_2.n3290 GNDA_2.n3289 76.3222
R5485 GNDA_2.n3294 GNDA_2.n1822 76.3222
R5486 GNDA_2.n3296 GNDA_2.n3295 76.3222
R5487 GNDA_2.n3305 GNDA_2.n3304 76.3222
R5488 GNDA_2.n3308 GNDA_2.n3307 76.3222
R5489 GNDA_2.n3317 GNDA_2.n3316 76.3222
R5490 GNDA_2.n3320 GNDA_2.n3319 76.3222
R5491 GNDA_2.n3329 GNDA_2.n3328 76.3222
R5492 GNDA_2.n3299 GNDA_2.n3298 76.3222
R5493 GNDA_2.n3302 GNDA_2.n3301 76.3222
R5494 GNDA_2.n3311 GNDA_2.n3310 76.3222
R5495 GNDA_2.n3314 GNDA_2.n3313 76.3222
R5496 GNDA_2.n3323 GNDA_2.n3322 76.3222
R5497 GNDA_2.n3326 GNDA_2.n3325 76.3222
R5498 GNDA_2.n2432 GNDA_2.n2431 76.3222
R5499 GNDA_2.n2438 GNDA_2.n2437 76.3222
R5500 GNDA_2.n2439 GNDA_2.n2429 76.3222
R5501 GNDA_2.n2446 GNDA_2.n2445 76.3222
R5502 GNDA_2.n2450 GNDA_2.n2427 76.3222
R5503 GNDA_2.n2454 GNDA_2.n2452 76.3222
R5504 GNDA_2.n2453 GNDA_2.n1792 76.3222
R5505 GNDA_2.n2392 GNDA_2.n1793 76.3222
R5506 GNDA_2.n2394 GNDA_2.n1794 76.3222
R5507 GNDA_2.n2398 GNDA_2.n1795 76.3222
R5508 GNDA_2.n2400 GNDA_2.n1796 76.3222
R5509 GNDA_2.n3336 GNDA_2.n1786 76.3222
R5510 GNDA_2.n2506 GNDA_2.n2505 76.3222
R5511 GNDA_2.n2513 GNDA_2.n2512 76.3222
R5512 GNDA_2.n2516 GNDA_2.n2515 76.3222
R5513 GNDA_2.n2523 GNDA_2.n2522 76.3222
R5514 GNDA_2.n2526 GNDA_2.n2525 76.3222
R5515 GNDA_2.n2101 GNDA_2.n1926 76.3222
R5516 GNDA_2.n2503 GNDA_2.n2502 76.3222
R5517 GNDA_2.n2498 GNDA_2.n1992 76.3222
R5518 GNDA_2.n2496 GNDA_2.n2495 76.3222
R5519 GNDA_2.n2491 GNDA_2.n1995 76.3222
R5520 GNDA_2.n2489 GNDA_2.n2488 76.3222
R5521 GNDA_2.n2484 GNDA_2.n1998 76.3222
R5522 GNDA_2.n2104 GNDA_2.n1862 76.3222
R5523 GNDA_2.n2130 GNDA_2.n1861 76.3222
R5524 GNDA_2.n2125 GNDA_2.n1860 76.3222
R5525 GNDA_2.n2118 GNDA_2.n1859 76.3222
R5526 GNDA_2.n2111 GNDA_2.n1858 76.3222
R5527 GNDA_2.n2140 GNDA_2.n1857 76.3222
R5528 GNDA_2.n2483 GNDA_2.n1999 76.3222
R5529 GNDA_2.n2019 GNDA_2.n2010 76.3222
R5530 GNDA_2.n2020 GNDA_2.n2012 76.3222
R5531 GNDA_2.n2021 GNDA_2.n2014 76.3222
R5532 GNDA_2.n2022 GNDA_2.n2016 76.3222
R5533 GNDA_2.n2024 GNDA_2.n2018 76.3222
R5534 GNDA_2.n5454 GNDA_2.n48 76.3222
R5535 GNDA_2.n5449 GNDA_2.n47 76.3222
R5536 GNDA_2.n5366 GNDA_2.n46 76.3222
R5537 GNDA_2.n5372 GNDA_2.n45 76.3222
R5538 GNDA_2.n5378 GNDA_2.n44 76.3222
R5539 GNDA_2.n5387 GNDA_2.n43 76.3222
R5540 GNDA_2.n2481 GNDA_2.n2480 76.3222
R5541 GNDA_2.n2008 GNDA_2.n2003 76.3222
R5542 GNDA_2.n2473 GNDA_2.n2004 76.3222
R5543 GNDA_2.n2469 GNDA_2.n2005 76.3222
R5544 GNDA_2.n2465 GNDA_2.n2006 76.3222
R5545 GNDA_2.n2184 GNDA_2.n2183 76.3222
R5546 GNDA_2.n2185 GNDA_2.n2180 76.3222
R5547 GNDA_2.n2192 GNDA_2.n2191 76.3222
R5548 GNDA_2.n2193 GNDA_2.n2178 76.3222
R5549 GNDA_2.n2200 GNDA_2.n2199 76.3222
R5550 GNDA_2.n2204 GNDA_2.n2176 76.3222
R5551 GNDA_2.n2457 GNDA_2.n1856 76.3222
R5552 GNDA_2.n2322 GNDA_2.n1855 76.3222
R5553 GNDA_2.n2239 GNDA_2.n1854 76.3222
R5554 GNDA_2.n2245 GNDA_2.n1853 76.3222
R5555 GNDA_2.n2251 GNDA_2.n1852 76.3222
R5556 GNDA_2.n2260 GNDA_2.n1851 76.3222
R5557 GNDA_2.n2424 GNDA_2.n2423 76.3222
R5558 GNDA_2.n2421 GNDA_2.n2390 76.3222
R5559 GNDA_2.n2417 GNDA_2.n2416 76.3222
R5560 GNDA_2.n2410 GNDA_2.n2396 76.3222
R5561 GNDA_2.n2409 GNDA_2.n2408 76.3222
R5562 GNDA_2.n2403 GNDA_2.n2402 76.3222
R5563 GNDA_2.n2388 GNDA_2.n2387 76.3222
R5564 GNDA_2.n2383 GNDA_2.n2333 76.3222
R5565 GNDA_2.n2381 GNDA_2.n2380 76.3222
R5566 GNDA_2.n2376 GNDA_2.n2336 76.3222
R5567 GNDA_2.n2374 GNDA_2.n2373 76.3222
R5568 GNDA_2.n2369 GNDA_2.n2339 76.3222
R5569 GNDA_2.n5354 GNDA_2.n42 76.3222
R5570 GNDA_2.n5553 GNDA_2.n5552 76.3222
R5571 GNDA_2.n41 GNDA_2.n40 76.3222
R5572 GNDA_2.n30 GNDA_2.n29 76.3222
R5573 GNDA_2.n5289 GNDA_2.n28 76.3222
R5574 GNDA_2.n5295 GNDA_2.n27 76.3222
R5575 GNDA_2.n2025 GNDA_2.n2024 76.3222
R5576 GNDA_2.n2022 GNDA_2.n2017 76.3222
R5577 GNDA_2.n2021 GNDA_2.n2015 76.3222
R5578 GNDA_2.n2020 GNDA_2.n2013 76.3222
R5579 GNDA_2.n2019 GNDA_2.n2011 76.3222
R5580 GNDA_2.n2009 GNDA_2.n1999 76.3222
R5581 GNDA_2.n2480 GNDA_2.n2002 76.3222
R5582 GNDA_2.n2474 GNDA_2.n2003 76.3222
R5583 GNDA_2.n2470 GNDA_2.n2004 76.3222
R5584 GNDA_2.n2466 GNDA_2.n2005 76.3222
R5585 GNDA_2.n2462 GNDA_2.n2006 76.3222
R5586 GNDA_2.n3337 GNDA_2.n3336 76.3222
R5587 GNDA_2.n2404 GNDA_2.n1796 76.3222
R5588 GNDA_2.n2399 GNDA_2.n1795 76.3222
R5589 GNDA_2.n2397 GNDA_2.n1794 76.3222
R5590 GNDA_2.n2393 GNDA_2.n1793 76.3222
R5591 GNDA_2.n2391 GNDA_2.n1792 76.3222
R5592 GNDA_2.n2423 GNDA_2.n2422 76.3222
R5593 GNDA_2.n2418 GNDA_2.n2390 76.3222
R5594 GNDA_2.n2416 GNDA_2.n2415 76.3222
R5595 GNDA_2.n2411 GNDA_2.n2410 76.3222
R5596 GNDA_2.n2408 GNDA_2.n2407 76.3222
R5597 GNDA_2.n2402 GNDA_2.n1728 76.3222
R5598 GNDA_2.n3330 GNDA_2.n3329 76.3222
R5599 GNDA_2.n3319 GNDA_2.n1810 76.3222
R5600 GNDA_2.n3318 GNDA_2.n3317 76.3222
R5601 GNDA_2.n3307 GNDA_2.n1814 76.3222
R5602 GNDA_2.n3306 GNDA_2.n3305 76.3222
R5603 GNDA_2.n3295 GNDA_2.n1818 76.3222
R5604 GNDA_2.n3300 GNDA_2.n3299 76.3222
R5605 GNDA_2.n3301 GNDA_2.n1816 76.3222
R5606 GNDA_2.n3312 GNDA_2.n3311 76.3222
R5607 GNDA_2.n3313 GNDA_2.n1812 76.3222
R5608 GNDA_2.n3324 GNDA_2.n3323 76.3222
R5609 GNDA_2.n3325 GNDA_2.n1804 76.3222
R5610 GNDA_2.n2533 GNDA_2.n2532 76.3222
R5611 GNDA_2.n2530 GNDA_2.n2529 76.3222
R5612 GNDA_2.n1928 GNDA_2.n1922 76.3222
R5613 GNDA_2.n2519 GNDA_2.n1921 76.3222
R5614 GNDA_2.n1932 GNDA_2.n1920 76.3222
R5615 GNDA_2.n2509 GNDA_2.n1919 76.3222
R5616 GNDA_2.n2505 GNDA_2.n1934 76.3222
R5617 GNDA_2.n2514 GNDA_2.n2513 76.3222
R5618 GNDA_2.n2515 GNDA_2.n1930 76.3222
R5619 GNDA_2.n2524 GNDA_2.n2523 76.3222
R5620 GNDA_2.n2527 GNDA_2.n2526 76.3222
R5621 GNDA_2.n2102 GNDA_2.n2101 76.3222
R5622 GNDA_2.n1988 GNDA_2.n1943 76.3222
R5623 GNDA_2.n1981 GNDA_2.n1942 76.3222
R5624 GNDA_2.n1977 GNDA_2.n1941 76.3222
R5625 GNDA_2.n1973 GNDA_2.n1940 76.3222
R5626 GNDA_2.n1969 GNDA_2.n1939 76.3222
R5627 GNDA_2.n1965 GNDA_2.n1938 76.3222
R5628 GNDA_2.n1998 GNDA_2.n1996 76.3222
R5629 GNDA_2.n2490 GNDA_2.n2489 76.3222
R5630 GNDA_2.n1995 GNDA_2.n1993 76.3222
R5631 GNDA_2.n2497 GNDA_2.n2496 76.3222
R5632 GNDA_2.n1992 GNDA_2.n1990 76.3222
R5633 GNDA_2.n2504 GNDA_2.n2503 76.3222
R5634 GNDA_2.n2201 GNDA_2.n2176 76.3222
R5635 GNDA_2.n2199 GNDA_2.n2198 76.3222
R5636 GNDA_2.n2194 GNDA_2.n2193 76.3222
R5637 GNDA_2.n2191 GNDA_2.n2190 76.3222
R5638 GNDA_2.n2186 GNDA_2.n2185 76.3222
R5639 GNDA_2.n2183 GNDA_2.n2001 76.3222
R5640 GNDA_2.n5550 GNDA_2.n54 76.3222
R5641 GNDA_2.n5540 GNDA_2.n53 76.3222
R5642 GNDA_2.n5465 GNDA_2.n52 76.3222
R5643 GNDA_2.n5471 GNDA_2.n51 76.3222
R5644 GNDA_2.n5478 GNDA_2.n50 76.3222
R5645 GNDA_2.n5460 GNDA_2.n49 76.3222
R5646 GNDA_2.n5450 GNDA_2.n48 76.3222
R5647 GNDA_2.n5365 GNDA_2.n47 76.3222
R5648 GNDA_2.n5371 GNDA_2.n46 76.3222
R5649 GNDA_2.n5379 GNDA_2.n45 76.3222
R5650 GNDA_2.n5386 GNDA_2.n44 76.3222
R5651 GNDA_2.n5360 GNDA_2.n43 76.3222
R5652 GNDA_2.n42 GNDA_2.n24 76.3222
R5653 GNDA_2.n5552 GNDA_2.n25 76.3222
R5654 GNDA_2.n41 GNDA_2.n31 76.3222
R5655 GNDA_2.n5288 GNDA_2.n29 76.3222
R5656 GNDA_2.n5294 GNDA_2.n28 76.3222
R5657 GNDA_2.n5284 GNDA_2.n27 76.3222
R5658 GNDA_2.n3291 GNDA_2.n1822 76.3222
R5659 GNDA_2.n3289 GNDA_2.n3288 76.3222
R5660 GNDA_2.n3284 GNDA_2.n3283 76.3222
R5661 GNDA_2.n3281 GNDA_2.n3280 76.3222
R5662 GNDA_2.n3276 GNDA_2.n3275 76.3222
R5663 GNDA_2.n3273 GNDA_2.n3272 76.3222
R5664 GNDA_2.n2452 GNDA_2.n2451 76.3222
R5665 GNDA_2.n2447 GNDA_2.n2427 76.3222
R5666 GNDA_2.n2445 GNDA_2.n2444 76.3222
R5667 GNDA_2.n2440 GNDA_2.n2439 76.3222
R5668 GNDA_2.n2437 GNDA_2.n2436 76.3222
R5669 GNDA_2.n2431 GNDA_2.n1820 76.3222
R5670 GNDA_2.n2339 GNDA_2.n2337 76.3222
R5671 GNDA_2.n2375 GNDA_2.n2374 76.3222
R5672 GNDA_2.n2336 GNDA_2.n2334 76.3222
R5673 GNDA_2.n2382 GNDA_2.n2381 76.3222
R5674 GNDA_2.n2333 GNDA_2.n2331 76.3222
R5675 GNDA_2.n2389 GNDA_2.n2388 76.3222
R5676 GNDA_2.n2600 GNDA_2.n2599 76.3222
R5677 GNDA_2.n2597 GNDA_2.n2596 76.3222
R5678 GNDA_2.n1896 GNDA_2.n1866 76.3222
R5679 GNDA_2.n1900 GNDA_2.n1865 76.3222
R5680 GNDA_2.n1910 GNDA_2.n1864 76.3222
R5681 GNDA_2.n2535 GNDA_2.n1863 76.3222
R5682 GNDA_2.n2129 GNDA_2.n1862 76.3222
R5683 GNDA_2.n2126 GNDA_2.n1861 76.3222
R5684 GNDA_2.n2119 GNDA_2.n1860 76.3222
R5685 GNDA_2.n2112 GNDA_2.n1859 76.3222
R5686 GNDA_2.n2139 GNDA_2.n1858 76.3222
R5687 GNDA_2.n2327 GNDA_2.n1857 76.3222
R5688 GNDA_2.n2323 GNDA_2.n1856 76.3222
R5689 GNDA_2.n2238 GNDA_2.n1855 76.3222
R5690 GNDA_2.n2244 GNDA_2.n1854 76.3222
R5691 GNDA_2.n2252 GNDA_2.n1853 76.3222
R5692 GNDA_2.n2259 GNDA_2.n1852 76.3222
R5693 GNDA_2.n2233 GNDA_2.n1851 76.3222
R5694 GNDA_2.n3268 GNDA_2.n3267 76.3222
R5695 GNDA_2.n2945 GNDA_2.n2944 76.3222
R5696 GNDA_2.n2940 GNDA_2.n2611 76.3222
R5697 GNDA_2.n2936 GNDA_2.n2610 76.3222
R5698 GNDA_2.n2932 GNDA_2.n2609 76.3222
R5699 GNDA_2.n1961 GNDA_2.n1839 76.3222
R5700 GNDA_2.n1957 GNDA_2.n1840 76.3222
R5701 GNDA_2.n1953 GNDA_2.n1841 76.3222
R5702 GNDA_2.n1949 GNDA_2.n1842 76.3222
R5703 GNDA_2.n1945 GNDA_2.n1843 76.3222
R5704 GNDA_2.n3265 GNDA_2.n2947 76.3222
R5705 GNDA_2.n3257 GNDA_2.n1834 76.3222
R5706 GNDA_2.n3253 GNDA_2.n1835 76.3222
R5707 GNDA_2.n3249 GNDA_2.n1836 76.3222
R5708 GNDA_2.n3245 GNDA_2.n1837 76.3222
R5709 GNDA_2.n5502 GNDA_2.n70 74.5978
R5710 GNDA_2.n5499 GNDA_2.n70 74.5978
R5711 GNDA_2.n2555 GNDA_2.n2554 74.5978
R5712 GNDA_2.n2554 GNDA_2.n2553 74.5978
R5713 GNDA_2.n2882 GNDA_2.n2629 74.5978
R5714 GNDA_2.n2879 GNDA_2.n2629 74.5978
R5715 GNDA_2.n2731 GNDA_2.n2714 74.5978
R5716 GNDA_2.n2732 GNDA_2.n2731 74.5978
R5717 GNDA_2.n2067 GNDA_2.n2036 74.5978
R5718 GNDA_2.n2064 GNDA_2.n2036 74.5978
R5719 GNDA_2.n5410 GNDA_2.n99 74.5978
R5720 GNDA_2.n5407 GNDA_2.n99 74.5978
R5721 GNDA_2.n2283 GNDA_2.n2154 74.5978
R5722 GNDA_2.n2280 GNDA_2.n2154 74.5978
R5723 GNDA_2.n1746 GNDA_2.n1710 74.5978
R5724 GNDA_2.n1743 GNDA_2.n1710 74.5978
R5725 GNDA_2.n5318 GNDA_2.n9 74.5978
R5726 GNDA_2.n5315 GNDA_2.n9 74.5978
R5727 GNDA_2.n2814 GNDA_2.n1784 74.1184
R5728 GNDA_2.n2857 GNDA_2.t27 72.1152
R5729 GNDA_2.n2797 GNDA_2.t146 72.1152
R5730 GNDA_2.t139 GNDA_2.n1702 72.1152
R5731 GNDA_2.n4469 GNDA_2.n4466 71.0215
R5732 GNDA_2.n2972 GNDA_2.n2970 69.4466
R5733 GNDA_2.n5544 GNDA_2.n60 69.3109
R5734 GNDA_2.n5520 GNDA_2.n60 69.3109
R5735 GNDA_2.n2590 GNDA_2.n2589 69.3109
R5736 GNDA_2.n2589 GNDA_2.n2588 69.3109
R5737 GNDA_2.n2916 GNDA_2.n2622 69.3109
R5738 GNDA_2.n2916 GNDA_2.n2915 69.3109
R5739 GNDA_2.n2773 GNDA_2.n2772 69.3109
R5740 GNDA_2.n2772 GNDA_2.n2771 69.3109
R5741 GNDA_2.n2134 GNDA_2.n2133 69.3109
R5742 GNDA_2.n2134 GNDA_2.n2048 69.3109
R5743 GNDA_2.n5444 GNDA_2.n92 69.3109
R5744 GNDA_2.n5444 GNDA_2.n5443 69.3109
R5745 GNDA_2.n2317 GNDA_2.n2147 69.3109
R5746 GNDA_2.n2317 GNDA_2.n2316 69.3109
R5747 GNDA_2.n3362 GNDA_2.n3361 69.3109
R5748 GNDA_2.n3362 GNDA_2.n1723 69.3109
R5749 GNDA_2.n5557 GNDA_2.n5556 69.3109
R5750 GNDA_2.n5557 GNDA_2.n20 69.3109
R5751 GNDA_2.n3342 GNDA_2.t81 68.1089
R5752 GNDA_2.n1799 GNDA_2.n1784 66.1057
R5753 GNDA_2.t72 GNDA_2.n5534 65.8183
R5754 GNDA_2.t72 GNDA_2.n79 65.8183
R5755 GNDA_2.t72 GNDA_2.n78 65.8183
R5756 GNDA_2.t72 GNDA_2.n77 65.8183
R5757 GNDA_2.t72 GNDA_2.n68 65.8183
R5758 GNDA_2.t72 GNDA_2.n75 65.8183
R5759 GNDA_2.t72 GNDA_2.n66 65.8183
R5760 GNDA_2.t72 GNDA_2.n76 65.8183
R5761 GNDA_2.t72 GNDA_2.n74 65.8183
R5762 GNDA_2.t72 GNDA_2.n73 65.8183
R5763 GNDA_2.t72 GNDA_2.n72 65.8183
R5764 GNDA_2.t72 GNDA_2.n71 65.8183
R5765 GNDA_2.t72 GNDA_2.n69 65.8183
R5766 GNDA_2.t72 GNDA_2.n67 65.8183
R5767 GNDA_2.n5535 GNDA_2.t72 65.8183
R5768 GNDA_2.t72 GNDA_2.n61 65.8183
R5769 GNDA_2.n2572 GNDA_2.t152 65.8183
R5770 GNDA_2.n2578 GNDA_2.t152 65.8183
R5771 GNDA_2.n2580 GNDA_2.t152 65.8183
R5772 GNDA_2.n2586 GNDA_2.t152 65.8183
R5773 GNDA_2.n2556 GNDA_2.t152 65.8183
R5774 GNDA_2.n2562 GNDA_2.t152 65.8183
R5775 GNDA_2.n2564 GNDA_2.t152 65.8183
R5776 GNDA_2.n2570 GNDA_2.t152 65.8183
R5777 GNDA_2.n2540 GNDA_2.t152 65.8183
R5778 GNDA_2.n1886 GNDA_2.t152 65.8183
R5779 GNDA_2.n2547 GNDA_2.t152 65.8183
R5780 GNDA_2.n1883 GNDA_2.t152 65.8183
R5781 GNDA_2.n1906 GNDA_2.t152 65.8183
R5782 GNDA_2.n1904 GNDA_2.t152 65.8183
R5783 GNDA_2.n1891 GNDA_2.t152 65.8183
R5784 GNDA_2.n2592 GNDA_2.t152 65.8183
R5785 GNDA_2.t160 GNDA_2.n2639 65.8183
R5786 GNDA_2.t160 GNDA_2.n2638 65.8183
R5787 GNDA_2.t160 GNDA_2.n2637 65.8183
R5788 GNDA_2.t160 GNDA_2.n2636 65.8183
R5789 GNDA_2.t160 GNDA_2.n2627 65.8183
R5790 GNDA_2.t160 GNDA_2.n2634 65.8183
R5791 GNDA_2.t160 GNDA_2.n2624 65.8183
R5792 GNDA_2.t160 GNDA_2.n2635 65.8183
R5793 GNDA_2.t160 GNDA_2.n2633 65.8183
R5794 GNDA_2.t160 GNDA_2.n2632 65.8183
R5795 GNDA_2.t160 GNDA_2.n2631 65.8183
R5796 GNDA_2.t160 GNDA_2.n2630 65.8183
R5797 GNDA_2.t160 GNDA_2.n2628 65.8183
R5798 GNDA_2.t160 GNDA_2.n2626 65.8183
R5799 GNDA_2.t160 GNDA_2.n2625 65.8183
R5800 GNDA_2.n2917 GNDA_2.t160 65.8183
R5801 GNDA_2.n2753 GNDA_2.t119 65.8183
R5802 GNDA_2.n2755 GNDA_2.t119 65.8183
R5803 GNDA_2.n2761 GNDA_2.t119 65.8183
R5804 GNDA_2.n2763 GNDA_2.t119 65.8183
R5805 GNDA_2.n2737 GNDA_2.t119 65.8183
R5806 GNDA_2.n2739 GNDA_2.t119 65.8183
R5807 GNDA_2.n2745 GNDA_2.t119 65.8183
R5808 GNDA_2.n2747 GNDA_2.t119 65.8183
R5809 GNDA_2.t119 GNDA_2.n2676 65.8183
R5810 GNDA_2.n2722 GNDA_2.t119 65.8183
R5811 GNDA_2.n2718 GNDA_2.t119 65.8183
R5812 GNDA_2.n2729 GNDA_2.t119 65.8183
R5813 GNDA_2.n2804 GNDA_2.t119 65.8183
R5814 GNDA_2.n2790 GNDA_2.t119 65.8183
R5815 GNDA_2.n2788 GNDA_2.t119 65.8183
R5816 GNDA_2.n2774 GNDA_2.t119 65.8183
R5817 GNDA_2.t99 GNDA_2.n2047 65.8183
R5818 GNDA_2.t99 GNDA_2.n2046 65.8183
R5819 GNDA_2.t99 GNDA_2.n2045 65.8183
R5820 GNDA_2.t99 GNDA_2.n2044 65.8183
R5821 GNDA_2.t99 GNDA_2.n2035 65.8183
R5822 GNDA_2.t99 GNDA_2.n2042 65.8183
R5823 GNDA_2.t99 GNDA_2.n2032 65.8183
R5824 GNDA_2.t99 GNDA_2.n2043 65.8183
R5825 GNDA_2.t99 GNDA_2.n2041 65.8183
R5826 GNDA_2.t99 GNDA_2.n2039 65.8183
R5827 GNDA_2.t99 GNDA_2.n2038 65.8183
R5828 GNDA_2.t99 GNDA_2.n2037 65.8183
R5829 GNDA_2.n2135 GNDA_2.t99 65.8183
R5830 GNDA_2.t99 GNDA_2.n2034 65.8183
R5831 GNDA_2.t99 GNDA_2.n2033 65.8183
R5832 GNDA_2.t99 GNDA_2.n2031 65.8183
R5833 GNDA_2.t98 GNDA_2.n109 65.8183
R5834 GNDA_2.t98 GNDA_2.n108 65.8183
R5835 GNDA_2.t98 GNDA_2.n107 65.8183
R5836 GNDA_2.t98 GNDA_2.n106 65.8183
R5837 GNDA_2.t98 GNDA_2.n97 65.8183
R5838 GNDA_2.t98 GNDA_2.n104 65.8183
R5839 GNDA_2.t98 GNDA_2.n94 65.8183
R5840 GNDA_2.t98 GNDA_2.n105 65.8183
R5841 GNDA_2.t98 GNDA_2.n103 65.8183
R5842 GNDA_2.t98 GNDA_2.n102 65.8183
R5843 GNDA_2.t98 GNDA_2.n101 65.8183
R5844 GNDA_2.t98 GNDA_2.n100 65.8183
R5845 GNDA_2.t98 GNDA_2.n98 65.8183
R5846 GNDA_2.t98 GNDA_2.n96 65.8183
R5847 GNDA_2.t98 GNDA_2.n95 65.8183
R5848 GNDA_2.n5445 GNDA_2.t98 65.8183
R5849 GNDA_2.t85 GNDA_2.n2164 65.8183
R5850 GNDA_2.t85 GNDA_2.n2163 65.8183
R5851 GNDA_2.t85 GNDA_2.n2162 65.8183
R5852 GNDA_2.t85 GNDA_2.n2161 65.8183
R5853 GNDA_2.t85 GNDA_2.n2152 65.8183
R5854 GNDA_2.t85 GNDA_2.n2159 65.8183
R5855 GNDA_2.t85 GNDA_2.n2149 65.8183
R5856 GNDA_2.t85 GNDA_2.n2160 65.8183
R5857 GNDA_2.t85 GNDA_2.n2158 65.8183
R5858 GNDA_2.t85 GNDA_2.n2157 65.8183
R5859 GNDA_2.t85 GNDA_2.n2156 65.8183
R5860 GNDA_2.t85 GNDA_2.n2155 65.8183
R5861 GNDA_2.t85 GNDA_2.n2153 65.8183
R5862 GNDA_2.t85 GNDA_2.n2151 65.8183
R5863 GNDA_2.t85 GNDA_2.n2150 65.8183
R5864 GNDA_2.n2318 GNDA_2.t85 65.8183
R5865 GNDA_2.t75 GNDA_2.n1722 65.8183
R5866 GNDA_2.t75 GNDA_2.n1721 65.8183
R5867 GNDA_2.t75 GNDA_2.n1720 65.8183
R5868 GNDA_2.t75 GNDA_2.n1719 65.8183
R5869 GNDA_2.t75 GNDA_2.n1700 65.8183
R5870 GNDA_2.t75 GNDA_2.n1717 65.8183
R5871 GNDA_2.t75 GNDA_2.n1698 65.8183
R5872 GNDA_2.t75 GNDA_2.n1718 65.8183
R5873 GNDA_2.t75 GNDA_2.n1716 65.8183
R5874 GNDA_2.t75 GNDA_2.n1713 65.8183
R5875 GNDA_2.t75 GNDA_2.n1712 65.8183
R5876 GNDA_2.t75 GNDA_2.n1711 65.8183
R5877 GNDA_2.t75 GNDA_2.n1709 65.8183
R5878 GNDA_2.n3363 GNDA_2.t75 65.8183
R5879 GNDA_2.t75 GNDA_2.n1699 65.8183
R5880 GNDA_2.t75 GNDA_2.n1697 65.8183
R5881 GNDA_2.t74 GNDA_2.n19 65.8183
R5882 GNDA_2.t74 GNDA_2.n18 65.8183
R5883 GNDA_2.t74 GNDA_2.n17 65.8183
R5884 GNDA_2.t74 GNDA_2.n16 65.8183
R5885 GNDA_2.t74 GNDA_2.n7 65.8183
R5886 GNDA_2.t74 GNDA_2.n14 65.8183
R5887 GNDA_2.t74 GNDA_2.n5 65.8183
R5888 GNDA_2.t74 GNDA_2.n15 65.8183
R5889 GNDA_2.t74 GNDA_2.n13 65.8183
R5890 GNDA_2.t74 GNDA_2.n12 65.8183
R5891 GNDA_2.t74 GNDA_2.n11 65.8183
R5892 GNDA_2.t74 GNDA_2.n10 65.8183
R5893 GNDA_2.t74 GNDA_2.n8 65.8183
R5894 GNDA_2.n5558 GNDA_2.t74 65.8183
R5895 GNDA_2.t74 GNDA_2.n6 65.8183
R5896 GNDA_2.t74 GNDA_2.n4 65.8183
R5897 GNDA_2.n4351 GNDA_2.t137 65.3505
R5898 GNDA_2.n4350 GNDA_2.t115 65.3505
R5899 GNDA_2.n378 GNDA_2.t154 65.3505
R5900 GNDA_2.n377 GNDA_2.t128 65.3505
R5901 GNDA_2.n4431 GNDA_2.t84 65.3505
R5902 GNDA_2.n4429 GNDA_2.t69 65.3505
R5903 GNDA_2.t14 GNDA_2.t284 64.5256
R5904 GNDA_2.n4366 GNDA_2.n345 64.0005
R5905 GNDA_2.n4372 GNDA_2.n345 64.0005
R5906 GNDA_2.n388 GNDA_2.t107 63.4011
R5907 GNDA_2.n1076 GNDA_2.t144 63.4011
R5908 GNDA_2.n3403 GNDA_2.n3402 63.1009
R5909 GNDA_2.t166 GNDA_2.t188 62.9893
R5910 GNDA_2.n372 GNDA_2.t142 62.2505
R5911 GNDA_2.n351 GNDA_2.t156 62.2505
R5912 GNDA_2.n4399 GNDA_2.t88 62.2505
R5913 GNDA_2.n307 GNDA_2.t97 62.2505
R5914 GNDA_2.t4 GNDA_2.n2780 62.0993
R5915 GNDA_2.n3343 GNDA_2.t9 62.0993
R5916 GNDA_2.n4620 GNDA_2.n132 59.2425
R5917 GNDA_2.n4208 GNDA_2.n332 59.2425
R5918 GNDA_2.n4314 GNDA_2.n4313 59.2425
R5919 GNDA_2.n4471 GNDA_2.n4470 59.2425
R5920 GNDA_2.n2858 GNDA_2.t172 58.0929
R5921 GNDA_2.n2798 GNDA_2.t1 58.0929
R5922 GNDA_2.t72 GNDA_2.n60 57.8461
R5923 GNDA_2.n2589 GNDA_2.t152 57.8461
R5924 GNDA_2.t160 GNDA_2.n2916 57.8461
R5925 GNDA_2.n2772 GNDA_2.t119 57.8461
R5926 GNDA_2.t99 GNDA_2.n2134 57.8461
R5927 GNDA_2.t98 GNDA_2.n5444 57.8461
R5928 GNDA_2.t85 GNDA_2.n2317 57.8461
R5929 GNDA_2.t75 GNDA_2.n3362 57.8461
R5930 GNDA_2.t74 GNDA_2.n5557 57.8461
R5931 GNDA_2.n2699 GNDA_2.n2686 57.0913
R5932 GNDA_2.n3244 GNDA_2.n1838 56.3995
R5933 GNDA_2.n1838 GNDA_2.n55 56.3995
R5934 GNDA_2.n2231 GNDA_2.n2230 56.3995
R5935 GNDA_2.n3396 GNDA_2.n1674 56.3995
R5936 GNDA_2.n3396 GNDA_2.n3395 56.3995
R5937 GNDA_2.n2232 GNDA_2.n2231 56.3995
R5938 GNDA_2.n5282 GNDA_2.n5281 56.3995
R5939 GNDA_2.n5283 GNDA_2.n5282 56.3995
R5940 GNDA_2.n2613 GNDA_2.n2607 56.3995
R5941 GNDA_2.n2606 GNDA_2.n2605 56.3995
R5942 GNDA_2.t72 GNDA_2.n70 55.2026
R5943 GNDA_2.n2554 GNDA_2.t152 55.2026
R5944 GNDA_2.t160 GNDA_2.n2629 55.2026
R5945 GNDA_2.n2731 GNDA_2.t119 55.2026
R5946 GNDA_2.t99 GNDA_2.n2036 55.2026
R5947 GNDA_2.t98 GNDA_2.n99 55.2026
R5948 GNDA_2.t85 GNDA_2.n2154 55.2026
R5949 GNDA_2.t75 GNDA_2.n1710 55.2026
R5950 GNDA_2.t74 GNDA_2.n9 55.2026
R5951 GNDA_2.n5517 GNDA_2.n76 53.3664
R5952 GNDA_2.n5514 GNDA_2.n66 53.3664
R5953 GNDA_2.n5510 GNDA_2.n75 53.3664
R5954 GNDA_2.n5506 GNDA_2.n68 53.3664
R5955 GNDA_2.n5495 GNDA_2.n71 53.3664
R5956 GNDA_2.n5491 GNDA_2.n72 53.3664
R5957 GNDA_2.n5487 GNDA_2.n73 53.3664
R5958 GNDA_2.n5483 GNDA_2.n74 53.3664
R5959 GNDA_2.n5543 GNDA_2.n61 53.3664
R5960 GNDA_2.n5536 GNDA_2.n5535 53.3664
R5961 GNDA_2.n5468 GNDA_2.n67 53.3664
R5962 GNDA_2.n5475 GNDA_2.n69 53.3664
R5963 GNDA_2.n5534 GNDA_2.n5533 53.3664
R5964 GNDA_2.n81 GNDA_2.n79 53.3664
R5965 GNDA_2.n5528 GNDA_2.n78 53.3664
R5966 GNDA_2.n5524 GNDA_2.n77 53.3664
R5967 GNDA_2.n5534 GNDA_2.n80 53.3664
R5968 GNDA_2.n5529 GNDA_2.n79 53.3664
R5969 GNDA_2.n5525 GNDA_2.n78 53.3664
R5970 GNDA_2.n5521 GNDA_2.n77 53.3664
R5971 GNDA_2.n5503 GNDA_2.n68 53.3664
R5972 GNDA_2.n5507 GNDA_2.n75 53.3664
R5973 GNDA_2.n5511 GNDA_2.n66 53.3664
R5974 GNDA_2.n5515 GNDA_2.n76 53.3664
R5975 GNDA_2.n5486 GNDA_2.n74 53.3664
R5976 GNDA_2.n5490 GNDA_2.n73 53.3664
R5977 GNDA_2.n5494 GNDA_2.n72 53.3664
R5978 GNDA_2.n5498 GNDA_2.n71 53.3664
R5979 GNDA_2.n5482 GNDA_2.n69 53.3664
R5980 GNDA_2.n5474 GNDA_2.n67 53.3664
R5981 GNDA_2.n5535 GNDA_2.n65 53.3664
R5982 GNDA_2.n64 GNDA_2.n61 53.3664
R5983 GNDA_2.n2571 GNDA_2.n2570 53.3664
R5984 GNDA_2.n2564 GNDA_2.n1877 53.3664
R5985 GNDA_2.n2563 GNDA_2.n2562 53.3664
R5986 GNDA_2.n2556 GNDA_2.n1879 53.3664
R5987 GNDA_2.n2549 GNDA_2.n1883 53.3664
R5988 GNDA_2.n2547 GNDA_2.n2546 53.3664
R5989 GNDA_2.n2542 GNDA_2.n1886 53.3664
R5990 GNDA_2.n2540 GNDA_2.n2539 53.3664
R5991 GNDA_2.n2592 GNDA_2.n2591 53.3664
R5992 GNDA_2.n1891 GNDA_2.n1871 53.3664
R5993 GNDA_2.n1904 GNDA_2.n1903 53.3664
R5994 GNDA_2.n1907 GNDA_2.n1906 53.3664
R5995 GNDA_2.n2572 GNDA_2.n1875 53.3664
R5996 GNDA_2.n2578 GNDA_2.n2577 53.3664
R5997 GNDA_2.n2581 GNDA_2.n2580 53.3664
R5998 GNDA_2.n2586 GNDA_2.n2585 53.3664
R5999 GNDA_2.n2573 GNDA_2.n2572 53.3664
R6000 GNDA_2.n2579 GNDA_2.n2578 53.3664
R6001 GNDA_2.n2580 GNDA_2.n1873 53.3664
R6002 GNDA_2.n2587 GNDA_2.n2586 53.3664
R6003 GNDA_2.n2557 GNDA_2.n2556 53.3664
R6004 GNDA_2.n2562 GNDA_2.n2561 53.3664
R6005 GNDA_2.n2565 GNDA_2.n2564 53.3664
R6006 GNDA_2.n2570 GNDA_2.n2569 53.3664
R6007 GNDA_2.n2541 GNDA_2.n2540 53.3664
R6008 GNDA_2.n1886 GNDA_2.n1884 53.3664
R6009 GNDA_2.n2548 GNDA_2.n2547 53.3664
R6010 GNDA_2.n1883 GNDA_2.n1881 53.3664
R6011 GNDA_2.n1906 GNDA_2.n1887 53.3664
R6012 GNDA_2.n1905 GNDA_2.n1904 53.3664
R6013 GNDA_2.n1892 GNDA_2.n1891 53.3664
R6014 GNDA_2.n2593 GNDA_2.n2592 53.3664
R6015 GNDA_2.n2898 GNDA_2.n2635 53.3664
R6016 GNDA_2.n2894 GNDA_2.n2624 53.3664
R6017 GNDA_2.n2890 GNDA_2.n2634 53.3664
R6018 GNDA_2.n2886 GNDA_2.n2627 53.3664
R6019 GNDA_2.n2875 GNDA_2.n2630 53.3664
R6020 GNDA_2.n2871 GNDA_2.n2631 53.3664
R6021 GNDA_2.n2867 GNDA_2.n2632 53.3664
R6022 GNDA_2.n2863 GNDA_2.n2633 53.3664
R6023 GNDA_2.n2918 GNDA_2.n2917 53.3664
R6024 GNDA_2.n2649 GNDA_2.n2625 53.3664
R6025 GNDA_2.n2846 GNDA_2.n2626 53.3664
R6026 GNDA_2.n2851 GNDA_2.n2628 53.3664
R6027 GNDA_2.n2902 GNDA_2.n2639 53.3664
R6028 GNDA_2.n2903 GNDA_2.n2638 53.3664
R6029 GNDA_2.n2907 GNDA_2.n2637 53.3664
R6030 GNDA_2.n2911 GNDA_2.n2636 53.3664
R6031 GNDA_2.n2899 GNDA_2.n2639 53.3664
R6032 GNDA_2.n2906 GNDA_2.n2638 53.3664
R6033 GNDA_2.n2910 GNDA_2.n2637 53.3664
R6034 GNDA_2.n2640 GNDA_2.n2636 53.3664
R6035 GNDA_2.n2883 GNDA_2.n2627 53.3664
R6036 GNDA_2.n2887 GNDA_2.n2634 53.3664
R6037 GNDA_2.n2891 GNDA_2.n2624 53.3664
R6038 GNDA_2.n2895 GNDA_2.n2635 53.3664
R6039 GNDA_2.n2866 GNDA_2.n2633 53.3664
R6040 GNDA_2.n2870 GNDA_2.n2632 53.3664
R6041 GNDA_2.n2874 GNDA_2.n2631 53.3664
R6042 GNDA_2.n2878 GNDA_2.n2630 53.3664
R6043 GNDA_2.n2862 GNDA_2.n2628 53.3664
R6044 GNDA_2.n2850 GNDA_2.n2626 53.3664
R6045 GNDA_2.n2845 GNDA_2.n2625 53.3664
R6046 GNDA_2.n2917 GNDA_2.n2623 53.3664
R6047 GNDA_2.n2747 GNDA_2.n2710 53.3664
R6048 GNDA_2.n2746 GNDA_2.n2745 53.3664
R6049 GNDA_2.n2739 GNDA_2.n2712 53.3664
R6050 GNDA_2.n2738 GNDA_2.n2737 53.3664
R6051 GNDA_2.n2729 GNDA_2.n2728 53.3664
R6052 GNDA_2.n2724 GNDA_2.n2718 53.3664
R6053 GNDA_2.n2722 GNDA_2.n2721 53.3664
R6054 GNDA_2.n2806 GNDA_2.n2676 53.3664
R6055 GNDA_2.n2775 GNDA_2.n2774 53.3664
R6056 GNDA_2.n2788 GNDA_2.n2787 53.3664
R6057 GNDA_2.n2791 GNDA_2.n2790 53.3664
R6058 GNDA_2.n2804 GNDA_2.n2803 53.3664
R6059 GNDA_2.n2754 GNDA_2.n2753 53.3664
R6060 GNDA_2.n2756 GNDA_2.n2755 53.3664
R6061 GNDA_2.n2761 GNDA_2.n2760 53.3664
R6062 GNDA_2.n2764 GNDA_2.n2763 53.3664
R6063 GNDA_2.n2753 GNDA_2.n2752 53.3664
R6064 GNDA_2.n2755 GNDA_2.n2708 53.3664
R6065 GNDA_2.n2762 GNDA_2.n2761 53.3664
R6066 GNDA_2.n2763 GNDA_2.n2706 53.3664
R6067 GNDA_2.n2737 GNDA_2.n2736 53.3664
R6068 GNDA_2.n2740 GNDA_2.n2739 53.3664
R6069 GNDA_2.n2745 GNDA_2.n2744 53.3664
R6070 GNDA_2.n2748 GNDA_2.n2747 53.3664
R6071 GNDA_2.n2719 GNDA_2.n2676 53.3664
R6072 GNDA_2.n2723 GNDA_2.n2722 53.3664
R6073 GNDA_2.n2718 GNDA_2.n2716 53.3664
R6074 GNDA_2.n2730 GNDA_2.n2729 53.3664
R6075 GNDA_2.n2805 GNDA_2.n2804 53.3664
R6076 GNDA_2.n2790 GNDA_2.n2677 53.3664
R6077 GNDA_2.n2789 GNDA_2.n2788 53.3664
R6078 GNDA_2.n2774 GNDA_2.n2683 53.3664
R6079 GNDA_2.n2083 GNDA_2.n2043 53.3664
R6080 GNDA_2.n2079 GNDA_2.n2032 53.3664
R6081 GNDA_2.n2075 GNDA_2.n2042 53.3664
R6082 GNDA_2.n2071 GNDA_2.n2035 53.3664
R6083 GNDA_2.n2060 GNDA_2.n2037 53.3664
R6084 GNDA_2.n2056 GNDA_2.n2038 53.3664
R6085 GNDA_2.n2052 GNDA_2.n2039 53.3664
R6086 GNDA_2.n2041 GNDA_2.n2040 53.3664
R6087 GNDA_2.n2049 GNDA_2.n2031 53.3664
R6088 GNDA_2.n2122 GNDA_2.n2033 53.3664
R6089 GNDA_2.n2115 GNDA_2.n2034 53.3664
R6090 GNDA_2.n2136 GNDA_2.n2135 53.3664
R6091 GNDA_2.n2087 GNDA_2.n2047 53.3664
R6092 GNDA_2.n2088 GNDA_2.n2046 53.3664
R6093 GNDA_2.n2092 GNDA_2.n2045 53.3664
R6094 GNDA_2.n2096 GNDA_2.n2044 53.3664
R6095 GNDA_2.n2084 GNDA_2.n2047 53.3664
R6096 GNDA_2.n2091 GNDA_2.n2046 53.3664
R6097 GNDA_2.n2095 GNDA_2.n2045 53.3664
R6098 GNDA_2.n2098 GNDA_2.n2044 53.3664
R6099 GNDA_2.n2068 GNDA_2.n2035 53.3664
R6100 GNDA_2.n2072 GNDA_2.n2042 53.3664
R6101 GNDA_2.n2076 GNDA_2.n2032 53.3664
R6102 GNDA_2.n2080 GNDA_2.n2043 53.3664
R6103 GNDA_2.n2051 GNDA_2.n2041 53.3664
R6104 GNDA_2.n2055 GNDA_2.n2039 53.3664
R6105 GNDA_2.n2059 GNDA_2.n2038 53.3664
R6106 GNDA_2.n2063 GNDA_2.n2037 53.3664
R6107 GNDA_2.n2135 GNDA_2.n2030 53.3664
R6108 GNDA_2.n2034 GNDA_2.n2029 53.3664
R6109 GNDA_2.n2114 GNDA_2.n2033 53.3664
R6110 GNDA_2.n2121 GNDA_2.n2031 53.3664
R6111 GNDA_2.n5426 GNDA_2.n105 53.3664
R6112 GNDA_2.n5422 GNDA_2.n94 53.3664
R6113 GNDA_2.n5418 GNDA_2.n104 53.3664
R6114 GNDA_2.n5414 GNDA_2.n97 53.3664
R6115 GNDA_2.n5403 GNDA_2.n100 53.3664
R6116 GNDA_2.n5399 GNDA_2.n101 53.3664
R6117 GNDA_2.n5395 GNDA_2.n102 53.3664
R6118 GNDA_2.n5391 GNDA_2.n103 53.3664
R6119 GNDA_2.n5446 GNDA_2.n5445 53.3664
R6120 GNDA_2.n5368 GNDA_2.n95 53.3664
R6121 GNDA_2.n5376 GNDA_2.n96 53.3664
R6122 GNDA_2.n5383 GNDA_2.n98 53.3664
R6123 GNDA_2.n5430 GNDA_2.n109 53.3664
R6124 GNDA_2.n5431 GNDA_2.n108 53.3664
R6125 GNDA_2.n5435 GNDA_2.n107 53.3664
R6126 GNDA_2.n5439 GNDA_2.n106 53.3664
R6127 GNDA_2.n5427 GNDA_2.n109 53.3664
R6128 GNDA_2.n5434 GNDA_2.n108 53.3664
R6129 GNDA_2.n5438 GNDA_2.n107 53.3664
R6130 GNDA_2.n5442 GNDA_2.n106 53.3664
R6131 GNDA_2.n5411 GNDA_2.n97 53.3664
R6132 GNDA_2.n5415 GNDA_2.n104 53.3664
R6133 GNDA_2.n5419 GNDA_2.n94 53.3664
R6134 GNDA_2.n5423 GNDA_2.n105 53.3664
R6135 GNDA_2.n5394 GNDA_2.n103 53.3664
R6136 GNDA_2.n5398 GNDA_2.n102 53.3664
R6137 GNDA_2.n5402 GNDA_2.n101 53.3664
R6138 GNDA_2.n5406 GNDA_2.n100 53.3664
R6139 GNDA_2.n5390 GNDA_2.n98 53.3664
R6140 GNDA_2.n5382 GNDA_2.n96 53.3664
R6141 GNDA_2.n5375 GNDA_2.n95 53.3664
R6142 GNDA_2.n5445 GNDA_2.n93 53.3664
R6143 GNDA_2.n2299 GNDA_2.n2160 53.3664
R6144 GNDA_2.n2295 GNDA_2.n2149 53.3664
R6145 GNDA_2.n2291 GNDA_2.n2159 53.3664
R6146 GNDA_2.n2287 GNDA_2.n2152 53.3664
R6147 GNDA_2.n2276 GNDA_2.n2155 53.3664
R6148 GNDA_2.n2272 GNDA_2.n2156 53.3664
R6149 GNDA_2.n2268 GNDA_2.n2157 53.3664
R6150 GNDA_2.n2264 GNDA_2.n2158 53.3664
R6151 GNDA_2.n2319 GNDA_2.n2318 53.3664
R6152 GNDA_2.n2241 GNDA_2.n2150 53.3664
R6153 GNDA_2.n2249 GNDA_2.n2151 53.3664
R6154 GNDA_2.n2256 GNDA_2.n2153 53.3664
R6155 GNDA_2.n2303 GNDA_2.n2164 53.3664
R6156 GNDA_2.n2304 GNDA_2.n2163 53.3664
R6157 GNDA_2.n2308 GNDA_2.n2162 53.3664
R6158 GNDA_2.n2312 GNDA_2.n2161 53.3664
R6159 GNDA_2.n2300 GNDA_2.n2164 53.3664
R6160 GNDA_2.n2307 GNDA_2.n2163 53.3664
R6161 GNDA_2.n2311 GNDA_2.n2162 53.3664
R6162 GNDA_2.n2315 GNDA_2.n2161 53.3664
R6163 GNDA_2.n2284 GNDA_2.n2152 53.3664
R6164 GNDA_2.n2288 GNDA_2.n2159 53.3664
R6165 GNDA_2.n2292 GNDA_2.n2149 53.3664
R6166 GNDA_2.n2296 GNDA_2.n2160 53.3664
R6167 GNDA_2.n2267 GNDA_2.n2158 53.3664
R6168 GNDA_2.n2271 GNDA_2.n2157 53.3664
R6169 GNDA_2.n2275 GNDA_2.n2156 53.3664
R6170 GNDA_2.n2279 GNDA_2.n2155 53.3664
R6171 GNDA_2.n2263 GNDA_2.n2153 53.3664
R6172 GNDA_2.n2255 GNDA_2.n2151 53.3664
R6173 GNDA_2.n2248 GNDA_2.n2150 53.3664
R6174 GNDA_2.n2318 GNDA_2.n2148 53.3664
R6175 GNDA_2.n1762 GNDA_2.n1718 53.3664
R6176 GNDA_2.n1758 GNDA_2.n1698 53.3664
R6177 GNDA_2.n1754 GNDA_2.n1717 53.3664
R6178 GNDA_2.n1750 GNDA_2.n1700 53.3664
R6179 GNDA_2.n1739 GNDA_2.n1711 53.3664
R6180 GNDA_2.n1735 GNDA_2.n1712 53.3664
R6181 GNDA_2.n1731 GNDA_2.n1713 53.3664
R6182 GNDA_2.n1716 GNDA_2.n1715 53.3664
R6183 GNDA_2.n1724 GNDA_2.n1697 53.3664
R6184 GNDA_2.n3351 GNDA_2.n1699 53.3664
R6185 GNDA_2.n3364 GNDA_2.n3363 53.3664
R6186 GNDA_2.n1709 GNDA_2.n1708 53.3664
R6187 GNDA_2.n1766 GNDA_2.n1722 53.3664
R6188 GNDA_2.n1767 GNDA_2.n1721 53.3664
R6189 GNDA_2.n1771 GNDA_2.n1720 53.3664
R6190 GNDA_2.n1775 GNDA_2.n1719 53.3664
R6191 GNDA_2.n1763 GNDA_2.n1722 53.3664
R6192 GNDA_2.n1770 GNDA_2.n1721 53.3664
R6193 GNDA_2.n1774 GNDA_2.n1720 53.3664
R6194 GNDA_2.n1777 GNDA_2.n1719 53.3664
R6195 GNDA_2.n1747 GNDA_2.n1700 53.3664
R6196 GNDA_2.n1751 GNDA_2.n1717 53.3664
R6197 GNDA_2.n1755 GNDA_2.n1698 53.3664
R6198 GNDA_2.n1759 GNDA_2.n1718 53.3664
R6199 GNDA_2.n1730 GNDA_2.n1716 53.3664
R6200 GNDA_2.n1734 GNDA_2.n1713 53.3664
R6201 GNDA_2.n1738 GNDA_2.n1712 53.3664
R6202 GNDA_2.n1742 GNDA_2.n1711 53.3664
R6203 GNDA_2.n1714 GNDA_2.n1709 53.3664
R6204 GNDA_2.n3363 GNDA_2.n1696 53.3664
R6205 GNDA_2.n1699 GNDA_2.n1695 53.3664
R6206 GNDA_2.n3350 GNDA_2.n1697 53.3664
R6207 GNDA_2.n5334 GNDA_2.n15 53.3664
R6208 GNDA_2.n5330 GNDA_2.n5 53.3664
R6209 GNDA_2.n5326 GNDA_2.n14 53.3664
R6210 GNDA_2.n5322 GNDA_2.n7 53.3664
R6211 GNDA_2.n5311 GNDA_2.n10 53.3664
R6212 GNDA_2.n5307 GNDA_2.n11 53.3664
R6213 GNDA_2.n5303 GNDA_2.n12 53.3664
R6214 GNDA_2.n5299 GNDA_2.n13 53.3664
R6215 GNDA_2.n21 GNDA_2.n4 53.3664
R6216 GNDA_2.n37 GNDA_2.n6 53.3664
R6217 GNDA_2.n5559 GNDA_2.n5558 53.3664
R6218 GNDA_2.n5291 GNDA_2.n8 53.3664
R6219 GNDA_2.n5338 GNDA_2.n19 53.3664
R6220 GNDA_2.n5339 GNDA_2.n18 53.3664
R6221 GNDA_2.n5343 GNDA_2.n17 53.3664
R6222 GNDA_2.n5347 GNDA_2.n16 53.3664
R6223 GNDA_2.n5335 GNDA_2.n19 53.3664
R6224 GNDA_2.n5342 GNDA_2.n18 53.3664
R6225 GNDA_2.n5346 GNDA_2.n17 53.3664
R6226 GNDA_2.n5349 GNDA_2.n16 53.3664
R6227 GNDA_2.n5319 GNDA_2.n7 53.3664
R6228 GNDA_2.n5323 GNDA_2.n14 53.3664
R6229 GNDA_2.n5327 GNDA_2.n5 53.3664
R6230 GNDA_2.n5331 GNDA_2.n15 53.3664
R6231 GNDA_2.n5302 GNDA_2.n13 53.3664
R6232 GNDA_2.n5306 GNDA_2.n12 53.3664
R6233 GNDA_2.n5310 GNDA_2.n11 53.3664
R6234 GNDA_2.n5314 GNDA_2.n10 53.3664
R6235 GNDA_2.n5298 GNDA_2.n8 53.3664
R6236 GNDA_2.n5558 GNDA_2.n3 53.3664
R6237 GNDA_2.n6 GNDA_2.n2 53.3664
R6238 GNDA_2.n36 GNDA_2.n4 53.3664
R6239 GNDA_2.n2924 GNDA_2.n2922 53.085
R6240 GNDA_2.n2686 GNDA_2.n1803 53.085
R6241 GNDA_2.n2818 GNDA_2.n2815 53.085
R6242 GNDA_2.n2858 GNDA_2.t241 52.0834
R6243 GNDA_2.n2798 GNDA_2.t245 52.0834
R6244 GNDA_2.n3368 GNDA_2.t35 52.0834
R6245 GNDA_2.n3240 GNDA_2.n2951 50.8806
R6246 GNDA_2.n3240 GNDA_2.n3239 50.8806
R6247 GNDA_2.n3239 GNDA_2.n3238 50.8806
R6248 GNDA_2.n3238 GNDA_2.n2952 50.8806
R6249 GNDA_2.n3232 GNDA_2.n2952 50.8806
R6250 GNDA_2.n3231 GNDA_2.n3230 50.8806
R6251 GNDA_2.n3230 GNDA_2.n2956 50.8806
R6252 GNDA_2.n3224 GNDA_2.n2956 50.8806
R6253 GNDA_2.n3224 GNDA_2.n3223 50.8806
R6254 GNDA_2.n3223 GNDA_2.n3222 50.8806
R6255 GNDA_2.n3178 GNDA_2.n3177 50.8806
R6256 GNDA_2.n3177 GNDA_2.n3176 50.8806
R6257 GNDA_2.n3176 GNDA_2.n2965 50.8806
R6258 GNDA_2.n3170 GNDA_2.n2965 50.8806
R6259 GNDA_2.n3170 GNDA_2.n3169 50.8806
R6260 GNDA_2.n3162 GNDA_2.n2971 50.8806
R6261 GNDA_2.n3162 GNDA_2.n3161 50.8806
R6262 GNDA_2.n3161 GNDA_2.n3160 50.8806
R6263 GNDA_2.n3160 GNDA_2.n3072 50.8806
R6264 GNDA_2.n3154 GNDA_2.n3072 50.8806
R6265 GNDA_2.n3152 GNDA_2.n3078 50.8806
R6266 GNDA_2.n3146 GNDA_2.n3078 50.8806
R6267 GNDA_2.n3146 GNDA_2.n3145 50.8806
R6268 GNDA_2.n3145 GNDA_2.n3144 50.8806
R6269 GNDA_2.n3144 GNDA_2.n3121 50.8806
R6270 GNDA_2.n3138 GNDA_2.n3137 50.8806
R6271 GNDA_2.n3137 GNDA_2.n3136 50.8806
R6272 GNDA_2.n3136 GNDA_2.n3125 50.8806
R6273 GNDA_2.n3130 GNDA_2.n3125 50.8806
R6274 GNDA_2.n3130 GNDA_2.n3129 50.8806
R6275 GNDA_2.n2655 GNDA_2.t162 48.077
R6276 GNDA_2.n2780 GNDA_2.t117 48.077
R6277 GNDA_2.n3343 GNDA_2.t55 48.077
R6278 GNDA_2.n1989 GNDA_2.t73 47.6748
R6279 GNDA_2.n2655 GNDA_2.t73 47.0754
R6280 GNDA_2.n3341 GNDA_2.t261 47.0754
R6281 GNDA_2.n1808 GNDA_2.t267 46.0738
R6282 GNDA_2.n3334 GNDA_2.n1803 43.069
R6283 GNDA_2.n2795 GNDA_2.t73 43.069
R6284 GNDA_2.t73 GNDA_2.n3368 43.069
R6285 GNDA_2.n569 GNDA_2.t123 42.6297
R6286 GNDA_2.t151 GNDA_2.n568 42.6297
R6287 GNDA_2.n4373 GNDA_2.t71 42.6297
R6288 GNDA_2.n343 GNDA_2.t104 42.6297
R6289 GNDA_2.n4405 GNDA_2.t87 42.4481
R6290 GNDA_2.n4461 GNDA_2.t96 42.4481
R6291 GNDA_2.t117 GNDA_2.n2779 42.0674
R6292 GNDA_2.t55 GNDA_2.n3342 42.0674
R6293 GNDA_2.n2781 GNDA_2.t276 41.0658
R6294 GNDA_2.t73 GNDA_2.t261 40.0642
R6295 GNDA_2.t241 GNDA_2.n2857 38.0611
R6296 GNDA_2.t245 GNDA_2.n2797 38.0611
R6297 GNDA_2.n2925 GNDA_2.n2924 37.0595
R6298 GNDA_2.t176 GNDA_2.n2654 37.0595
R6299 GNDA_2.n2818 GNDA_2.n2812 37.0595
R6300 GNDA_2.t288 GNDA_2.t226 36.3368
R6301 GNDA_2.t23 GNDA_2.t26 36.3368
R6302 GNDA_2.t208 GNDA_2.t228 36.3368
R6303 GNDA_2.t225 GNDA_2.t237 36.3368
R6304 GNDA_2.t22 GNDA_2.t21 36.3368
R6305 GNDA_2.t199 GNDA_2.t244 36.3368
R6306 GNDA_2.t62 GNDA_2.t248 36.3368
R6307 GNDA_2.t202 GNDA_2.t192 36.3368
R6308 GNDA_2.t198 GNDA_2.t178 36.3368
R6309 GNDA_2.t271 GNDA_2.t220 36.3368
R6310 GNDA_2.t267 GNDA_2.t78 35.0563
R6311 GNDA_2.t109 GNDA_2.t158 34.6852
R6312 GNDA_2.t134 GNDA_2.t125 34.6852
R6313 GNDA_2.t93 GNDA_2.t112 34.6852
R6314 GNDA_2.t90 GNDA_2.t101 34.6852
R6315 GNDA_2.n572 GNDA_2.n571 34.5991
R6316 GNDA_2.n574 GNDA_2.n573 34.5991
R6317 GNDA_2.n576 GNDA_2.n575 34.5991
R6318 GNDA_2.n578 GNDA_2.n577 34.5991
R6319 GNDA_2.n580 GNDA_2.n579 34.5991
R6320 GNDA_2.n582 GNDA_2.n581 34.5991
R6321 GNDA_2.n584 GNDA_2.n583 34.5991
R6322 GNDA_2.n586 GNDA_2.n585 34.5991
R6323 GNDA_2.n588 GNDA_2.n587 34.5991
R6324 GNDA_2.n590 GNDA_2.n589 34.5991
R6325 GNDA_2.n592 GNDA_2.n591 34.5991
R6326 GNDA_2.n594 GNDA_2.n593 34.5991
R6327 GNDA_2.n4384 GNDA_2.n4383 34.5991
R6328 GNDA_2.t34 GNDA_2.t196 33.1455
R6329 GNDA_2.n2838 GNDA_2.n2827 33.0531
R6330 GNDA_2.n1702 GNDA_2.t270 33.0531
R6331 GNDA_2.t73 GNDA_2.n26 32.9056
R6332 GNDA_2.n1850 GNDA_2.t73 32.9056
R6333 GNDA_2.n3382 GNDA_2.n3381 32.3969
R6334 GNDA_2.t1 GNDA_2.n2796 32.0515
R6335 GNDA_2.n4406 GNDA_2.n4405 31.533
R6336 GNDA_2.n3167 GNDA_2.n3166 31.3605
R6337 GNDA_2.n5254 GNDA_2.t126 31.1255
R6338 GNDA_2.n4468 GNDA_2.t110 31.1255
R6339 GNDA_2.n4408 GNDA_2.t102 31.1255
R6340 GNDA_2.n4316 GNDA_2.t94 31.1255
R6341 GNDA_2.t37 GNDA_2.t66 30.3834
R6342 GNDA_2.t250 GNDA_2.t37 30.3834
R6343 GNDA_2.t290 GNDA_2.t250 30.3834
R6344 GNDA_2.n2701 GNDA_2.n2699 30.0483
R6345 GNDA_2.t27 GNDA_2.n1808 29.0467
R6346 GNDA_2.t226 GNDA_2.t59 28.0786
R6347 GNDA_2.t216 GNDA_2.t22 28.0786
R6348 GNDA_2.t244 GNDA_2.t282 28.0786
R6349 GNDA_2.t190 GNDA_2.t271 28.0786
R6350 GNDA_2.n2782 GNDA_2.t4 28.0451
R6351 GNDA_2.t81 GNDA_2.n3341 28.0451
R6352 GNDA_2.n5519 GNDA_2.n5518 27.5561
R6353 GNDA_2.n2574 GNDA_2.n1876 27.5561
R6354 GNDA_2.n2900 GNDA_2.n2897 27.5561
R6355 GNDA_2.n2751 GNDA_2.n2750 27.5561
R6356 GNDA_2.n2085 GNDA_2.n2082 27.5561
R6357 GNDA_2.n5428 GNDA_2.n5425 27.5561
R6358 GNDA_2.n2301 GNDA_2.n2298 27.5561
R6359 GNDA_2.n1764 GNDA_2.n1761 27.5561
R6360 GNDA_2.n5336 GNDA_2.n5333 27.5561
R6361 GNDA_2.n2815 GNDA_2.n2814 27.0435
R6362 GNDA_2.n3379 GNDA_2.n1687 27.0435
R6363 GNDA_2.n3403 GNDA_2.n1667 27.0435
R6364 GNDA_2.t177 GNDA_2.t87 26.6819
R6365 GNDA_2.t15 GNDA_2.t235 26.6819
R6366 GNDA_2.t43 GNDA_2.t183 26.6819
R6367 GNDA_2.t50 GNDA_2.t96 26.6819
R6368 GNDA_2.n5501 GNDA_2.n5500 26.6672
R6369 GNDA_2.n2552 GNDA_2.n1880 26.6672
R6370 GNDA_2.n2881 GNDA_2.n2880 26.6672
R6371 GNDA_2.n2734 GNDA_2.n2733 26.6672
R6372 GNDA_2.n2066 GNDA_2.n2065 26.6672
R6373 GNDA_2.n5409 GNDA_2.n5408 26.6672
R6374 GNDA_2.n2282 GNDA_2.n2281 26.6672
R6375 GNDA_2.n1745 GNDA_2.n1744 26.6672
R6376 GNDA_2.n5317 GNDA_2.n5316 26.6672
R6377 GNDA_2.n3232 GNDA_2.t73 26.5712
R6378 GNDA_2.n3169 GNDA_2.t73 26.5712
R6379 GNDA_2.t73 GNDA_2.n3121 26.5712
R6380 GNDA_2.n2830 GNDA_2.n2829 25.3679
R6381 GNDA_2.t172 GNDA_2.t29 25.0403
R6382 GNDA_2.t9 GNDA_2.t48 25.0403
R6383 GNDA_2.n4470 GNDA_2.t109 24.7753
R6384 GNDA_2.t125 GNDA_2.n132 24.7753
R6385 GNDA_2.n4314 GNDA_2.t93 24.7753
R6386 GNDA_2.t101 GNDA_2.n332 24.7753
R6387 GNDA_2.t73 GNDA_2.n3231 24.3099
R6388 GNDA_2.t73 GNDA_2.n2971 24.3099
R6389 GNDA_2.n3138 GNDA_2.t73 24.3099
R6390 GNDA_2.n1676 GNDA_2.n1668 24.0387
R6391 GNDA_2.n1666 GNDA_2.t31 24.0005
R6392 GNDA_2.n1666 GNDA_2.t36 24.0005
R6393 GNDA_2.n1665 GNDA_2.t232 24.0005
R6394 GNDA_2.n1665 GNDA_2.t273 24.0005
R6395 GNDA_2.n1664 GNDA_2.t56 24.0005
R6396 GNDA_2.n1664 GNDA_2.t10 24.0005
R6397 GNDA_2.n1661 GNDA_2.t246 24.0005
R6398 GNDA_2.n1661 GNDA_2.t147 24.0005
R6399 GNDA_2.n1660 GNDA_2.t45 24.0005
R6400 GNDA_2.n1660 GNDA_2.t2 24.0005
R6401 GNDA_2.n1659 GNDA_2.t5 24.0005
R6402 GNDA_2.n1659 GNDA_2.t222 24.0005
R6403 GNDA_2.n1656 GNDA_2.t242 24.0005
R6404 GNDA_2.n1656 GNDA_2.t28 24.0005
R6405 GNDA_2.n1655 GNDA_2.t12 24.0005
R6406 GNDA_2.n1655 GNDA_2.t173 24.0005
R6407 GNDA_2.n1654 GNDA_2.t253 24.0005
R6408 GNDA_2.n1654 GNDA_2.t255 24.0005
R6409 GNDA_2.n1651 GNDA_2.t291 24.0005
R6410 GNDA_2.n1651 GNDA_2.t131 24.0005
R6411 GNDA_2.n1650 GNDA_2.t38 24.0005
R6412 GNDA_2.n1650 GNDA_2.t251 24.0005
R6413 GNDA_2.t280 GNDA_2.n1832 23.4782
R6414 GNDA_2.n5256 GNDA_2.t171 23.4439
R6415 GNDA_2.n4318 GNDA_2.t209 23.4439
R6416 GNDA_2.n4322 GNDA_2.t177 23.0435
R6417 GNDA_2.n4324 GNDA_2.t50 23.0435
R6418 GNDA_2.n2841 GNDA_2.n2840 23.0371
R6419 GNDA_2.n2813 GNDA_2.n1662 22.53
R6420 GNDA_2.t26 GNDA_2.t274 21.472
R6421 GNDA_2.t185 GNDA_2.t225 21.472
R6422 GNDA_2.t248 GNDA_2.t277 21.472
R6423 GNDA_2.t18 GNDA_2.t198 21.472
R6424 GNDA_2.n3405 GNDA_2.n3404 20.8233
R6425 GNDA_2.n1798 GNDA_2.n1663 20.8233
R6426 GNDA_2.n2700 GNDA_2.n1658 20.8233
R6427 GNDA_2.n1802 GNDA_2.n1657 20.8233
R6428 GNDA_2.n2616 GNDA_2.n1653 20.8233
R6429 GNDA_2.n2923 GNDA_2.n1652 20.8233
R6430 GNDA_2.n1831 GNDA_2.n1649 20.8233
R6431 GNDA_2.t54 GNDA_2.t168 20.5939
R6432 GNDA_2.t184 GNDA_2.t279 20.5939
R6433 GNDA_2.t73 GNDA_2.n1799 20.0324
R6434 GNDA_2.n4470 GNDA_2.n4469 19.8203
R6435 GNDA_2.n5255 GNDA_2.n132 19.8203
R6436 GNDA_2.n4317 GNDA_2.n4314 19.8203
R6437 GNDA_2.n4407 GNDA_2.n332 19.8203
R6438 GNDA_2.n5238 GNDA_2.t227 19.7005
R6439 GNDA_2.n5238 GNDA_2.t269 19.7005
R6440 GNDA_2.n5236 GNDA_2.t20 19.7005
R6441 GNDA_2.n5236 GNDA_2.t240 19.7005
R6442 GNDA_2.n5234 GNDA_2.t58 19.7005
R6443 GNDA_2.n5234 GNDA_2.t0 19.7005
R6444 GNDA_2.n5232 GNDA_2.t236 19.7005
R6445 GNDA_2.n5232 GNDA_2.t285 19.7005
R6446 GNDA_2.n5230 GNDA_2.t204 19.7005
R6447 GNDA_2.n5230 GNDA_2.t218 19.7005
R6448 GNDA_2.n5229 GNDA_2.t266 19.7005
R6449 GNDA_2.n5229 GNDA_2.t210 19.7005
R6450 GNDA_2.n3982 GNDA_2.t33 19.7005
R6451 GNDA_2.n3982 GNDA_2.t265 19.7005
R6452 GNDA_2.n3983 GNDA_2.t211 19.7005
R6453 GNDA_2.n3983 GNDA_2.t42 19.7005
R6454 GNDA_2.n3985 GNDA_2.t180 19.7005
R6455 GNDA_2.n3985 GNDA_2.t249 19.7005
R6456 GNDA_2.n3987 GNDA_2.t203 19.7005
R6457 GNDA_2.n3987 GNDA_2.t219 19.7005
R6458 GNDA_2.n3989 GNDA_2.t213 19.7005
R6459 GNDA_2.n3989 GNDA_2.t179 19.7005
R6460 GNDA_2.n3991 GNDA_2.t260 19.7005
R6461 GNDA_2.n3991 GNDA_2.t181 19.7005
R6462 GNDA_2.n5257 GNDA_2.t174 19.2044
R6463 GNDA_2.t174 GNDA_2.t189 18.4363
R6464 GNDA_2.t189 GNDA_2.t166 18.4363
R6465 GNDA_2.t230 GNDA_2.t14 18.4363
R6466 GNDA_2.t194 GNDA_2.t230 18.4363
R6467 GNDA_2.n2812 GNDA_2.t146 18.0292
R6468 GNDA_2.n2203 GNDA_2.n2175 17.5843
R6469 GNDA_2.n2370 GNDA_2.n2338 17.5843
R6470 GNDA_2.n3127 GNDA_2.n126 17.5843
R6471 GNDA_2.n5257 GNDA_2.n124 17.5479
R6472 GNDA_2.n3263 GNDA_2.n3243 16.9379
R6473 GNDA_2.n1966 GNDA_2.n1963 16.9379
R6474 GNDA_2.n3271 GNDA_2.n3270 16.9379
R6475 GNDA_2.n1997 GNDA_2.n111 16.7709
R6476 GNDA_2.n2459 GNDA_2.n2456 16.7709
R6477 GNDA_2.n1915 GNDA_2.n1821 16.7709
R6478 GNDA_2.n1935 GNDA_2.n84 16.7709
R6479 GNDA_2.n1833 GNDA_2.t73 16.4553
R6480 GNDA_2.n5532 GNDA_2.n5519 16.0005
R6481 GNDA_2.n5532 GNDA_2.n5531 16.0005
R6482 GNDA_2.n5531 GNDA_2.n5530 16.0005
R6483 GNDA_2.n5530 GNDA_2.n5527 16.0005
R6484 GNDA_2.n5527 GNDA_2.n5526 16.0005
R6485 GNDA_2.n5526 GNDA_2.n5523 16.0005
R6486 GNDA_2.n5523 GNDA_2.n5522 16.0005
R6487 GNDA_2.n5522 GNDA_2.n57 16.0005
R6488 GNDA_2.n5518 GNDA_2.n5516 16.0005
R6489 GNDA_2.n5516 GNDA_2.n5513 16.0005
R6490 GNDA_2.n5513 GNDA_2.n5512 16.0005
R6491 GNDA_2.n5512 GNDA_2.n5509 16.0005
R6492 GNDA_2.n5509 GNDA_2.n5508 16.0005
R6493 GNDA_2.n5508 GNDA_2.n5505 16.0005
R6494 GNDA_2.n5505 GNDA_2.n5504 16.0005
R6495 GNDA_2.n5504 GNDA_2.n5501 16.0005
R6496 GNDA_2.n5500 GNDA_2.n5497 16.0005
R6497 GNDA_2.n5497 GNDA_2.n5496 16.0005
R6498 GNDA_2.n5496 GNDA_2.n5493 16.0005
R6499 GNDA_2.n5493 GNDA_2.n5492 16.0005
R6500 GNDA_2.n5492 GNDA_2.n5489 16.0005
R6501 GNDA_2.n5489 GNDA_2.n5488 16.0005
R6502 GNDA_2.n5488 GNDA_2.n5485 16.0005
R6503 GNDA_2.n5485 GNDA_2.n5484 16.0005
R6504 GNDA_2.n2575 GNDA_2.n2574 16.0005
R6505 GNDA_2.n2576 GNDA_2.n2575 16.0005
R6506 GNDA_2.n2576 GNDA_2.n1874 16.0005
R6507 GNDA_2.n2582 GNDA_2.n1874 16.0005
R6508 GNDA_2.n2583 GNDA_2.n2582 16.0005
R6509 GNDA_2.n2584 GNDA_2.n2583 16.0005
R6510 GNDA_2.n2584 GNDA_2.n1872 16.0005
R6511 GNDA_2.n1872 GNDA_2.n1847 16.0005
R6512 GNDA_2.n2568 GNDA_2.n1876 16.0005
R6513 GNDA_2.n2568 GNDA_2.n2567 16.0005
R6514 GNDA_2.n2567 GNDA_2.n2566 16.0005
R6515 GNDA_2.n2566 GNDA_2.n1878 16.0005
R6516 GNDA_2.n2560 GNDA_2.n1878 16.0005
R6517 GNDA_2.n2560 GNDA_2.n2559 16.0005
R6518 GNDA_2.n2559 GNDA_2.n2558 16.0005
R6519 GNDA_2.n2558 GNDA_2.n1880 16.0005
R6520 GNDA_2.n2552 GNDA_2.n2551 16.0005
R6521 GNDA_2.n2551 GNDA_2.n2550 16.0005
R6522 GNDA_2.n2550 GNDA_2.n1882 16.0005
R6523 GNDA_2.n2545 GNDA_2.n1882 16.0005
R6524 GNDA_2.n2545 GNDA_2.n2544 16.0005
R6525 GNDA_2.n2544 GNDA_2.n2543 16.0005
R6526 GNDA_2.n2543 GNDA_2.n1885 16.0005
R6527 GNDA_2.n2538 GNDA_2.n1885 16.0005
R6528 GNDA_2.n2901 GNDA_2.n2900 16.0005
R6529 GNDA_2.n2904 GNDA_2.n2901 16.0005
R6530 GNDA_2.n2905 GNDA_2.n2904 16.0005
R6531 GNDA_2.n2908 GNDA_2.n2905 16.0005
R6532 GNDA_2.n2909 GNDA_2.n2908 16.0005
R6533 GNDA_2.n2912 GNDA_2.n2909 16.0005
R6534 GNDA_2.n2913 GNDA_2.n2912 16.0005
R6535 GNDA_2.n2914 GNDA_2.n2913 16.0005
R6536 GNDA_2.n2897 GNDA_2.n2896 16.0005
R6537 GNDA_2.n2896 GNDA_2.n2893 16.0005
R6538 GNDA_2.n2893 GNDA_2.n2892 16.0005
R6539 GNDA_2.n2892 GNDA_2.n2889 16.0005
R6540 GNDA_2.n2889 GNDA_2.n2888 16.0005
R6541 GNDA_2.n2888 GNDA_2.n2885 16.0005
R6542 GNDA_2.n2885 GNDA_2.n2884 16.0005
R6543 GNDA_2.n2884 GNDA_2.n2881 16.0005
R6544 GNDA_2.n2880 GNDA_2.n2877 16.0005
R6545 GNDA_2.n2877 GNDA_2.n2876 16.0005
R6546 GNDA_2.n2876 GNDA_2.n2873 16.0005
R6547 GNDA_2.n2873 GNDA_2.n2872 16.0005
R6548 GNDA_2.n2872 GNDA_2.n2869 16.0005
R6549 GNDA_2.n2869 GNDA_2.n2868 16.0005
R6550 GNDA_2.n2868 GNDA_2.n2865 16.0005
R6551 GNDA_2.n2865 GNDA_2.n2864 16.0005
R6552 GNDA_2.n2751 GNDA_2.n2709 16.0005
R6553 GNDA_2.n2757 GNDA_2.n2709 16.0005
R6554 GNDA_2.n2758 GNDA_2.n2757 16.0005
R6555 GNDA_2.n2759 GNDA_2.n2758 16.0005
R6556 GNDA_2.n2759 GNDA_2.n2707 16.0005
R6557 GNDA_2.n2765 GNDA_2.n2707 16.0005
R6558 GNDA_2.n2766 GNDA_2.n2765 16.0005
R6559 GNDA_2.n2770 GNDA_2.n2766 16.0005
R6560 GNDA_2.n2750 GNDA_2.n2749 16.0005
R6561 GNDA_2.n2749 GNDA_2.n2711 16.0005
R6562 GNDA_2.n2743 GNDA_2.n2711 16.0005
R6563 GNDA_2.n2743 GNDA_2.n2742 16.0005
R6564 GNDA_2.n2742 GNDA_2.n2741 16.0005
R6565 GNDA_2.n2741 GNDA_2.n2713 16.0005
R6566 GNDA_2.n2735 GNDA_2.n2713 16.0005
R6567 GNDA_2.n2735 GNDA_2.n2734 16.0005
R6568 GNDA_2.n2733 GNDA_2.n2715 16.0005
R6569 GNDA_2.n2727 GNDA_2.n2715 16.0005
R6570 GNDA_2.n2727 GNDA_2.n2726 16.0005
R6571 GNDA_2.n2726 GNDA_2.n2725 16.0005
R6572 GNDA_2.n2725 GNDA_2.n2717 16.0005
R6573 GNDA_2.n2720 GNDA_2.n2717 16.0005
R6574 GNDA_2.n2720 GNDA_2.n2675 16.0005
R6575 GNDA_2.n2807 GNDA_2.n2675 16.0005
R6576 GNDA_2.n2086 GNDA_2.n2085 16.0005
R6577 GNDA_2.n2089 GNDA_2.n2086 16.0005
R6578 GNDA_2.n2090 GNDA_2.n2089 16.0005
R6579 GNDA_2.n2093 GNDA_2.n2090 16.0005
R6580 GNDA_2.n2094 GNDA_2.n2093 16.0005
R6581 GNDA_2.n2097 GNDA_2.n2094 16.0005
R6582 GNDA_2.n2099 GNDA_2.n2097 16.0005
R6583 GNDA_2.n2100 GNDA_2.n2099 16.0005
R6584 GNDA_2.n2082 GNDA_2.n2081 16.0005
R6585 GNDA_2.n2081 GNDA_2.n2078 16.0005
R6586 GNDA_2.n2078 GNDA_2.n2077 16.0005
R6587 GNDA_2.n2077 GNDA_2.n2074 16.0005
R6588 GNDA_2.n2074 GNDA_2.n2073 16.0005
R6589 GNDA_2.n2073 GNDA_2.n2070 16.0005
R6590 GNDA_2.n2070 GNDA_2.n2069 16.0005
R6591 GNDA_2.n2069 GNDA_2.n2066 16.0005
R6592 GNDA_2.n2065 GNDA_2.n2062 16.0005
R6593 GNDA_2.n2062 GNDA_2.n2061 16.0005
R6594 GNDA_2.n2061 GNDA_2.n2058 16.0005
R6595 GNDA_2.n2058 GNDA_2.n2057 16.0005
R6596 GNDA_2.n2057 GNDA_2.n2054 16.0005
R6597 GNDA_2.n2054 GNDA_2.n2053 16.0005
R6598 GNDA_2.n2053 GNDA_2.n2050 16.0005
R6599 GNDA_2.n2050 GNDA_2.n2026 16.0005
R6600 GNDA_2.n5429 GNDA_2.n5428 16.0005
R6601 GNDA_2.n5432 GNDA_2.n5429 16.0005
R6602 GNDA_2.n5433 GNDA_2.n5432 16.0005
R6603 GNDA_2.n5436 GNDA_2.n5433 16.0005
R6604 GNDA_2.n5437 GNDA_2.n5436 16.0005
R6605 GNDA_2.n5440 GNDA_2.n5437 16.0005
R6606 GNDA_2.n5441 GNDA_2.n5440 16.0005
R6607 GNDA_2.n5441 GNDA_2.n89 16.0005
R6608 GNDA_2.n5425 GNDA_2.n5424 16.0005
R6609 GNDA_2.n5424 GNDA_2.n5421 16.0005
R6610 GNDA_2.n5421 GNDA_2.n5420 16.0005
R6611 GNDA_2.n5420 GNDA_2.n5417 16.0005
R6612 GNDA_2.n5417 GNDA_2.n5416 16.0005
R6613 GNDA_2.n5416 GNDA_2.n5413 16.0005
R6614 GNDA_2.n5413 GNDA_2.n5412 16.0005
R6615 GNDA_2.n5412 GNDA_2.n5409 16.0005
R6616 GNDA_2.n5408 GNDA_2.n5405 16.0005
R6617 GNDA_2.n5405 GNDA_2.n5404 16.0005
R6618 GNDA_2.n5404 GNDA_2.n5401 16.0005
R6619 GNDA_2.n5401 GNDA_2.n5400 16.0005
R6620 GNDA_2.n5400 GNDA_2.n5397 16.0005
R6621 GNDA_2.n5397 GNDA_2.n5396 16.0005
R6622 GNDA_2.n5396 GNDA_2.n5393 16.0005
R6623 GNDA_2.n5393 GNDA_2.n5392 16.0005
R6624 GNDA_2.n2302 GNDA_2.n2301 16.0005
R6625 GNDA_2.n2305 GNDA_2.n2302 16.0005
R6626 GNDA_2.n2306 GNDA_2.n2305 16.0005
R6627 GNDA_2.n2309 GNDA_2.n2306 16.0005
R6628 GNDA_2.n2310 GNDA_2.n2309 16.0005
R6629 GNDA_2.n2313 GNDA_2.n2310 16.0005
R6630 GNDA_2.n2314 GNDA_2.n2313 16.0005
R6631 GNDA_2.n2314 GNDA_2.n2144 16.0005
R6632 GNDA_2.n2298 GNDA_2.n2297 16.0005
R6633 GNDA_2.n2297 GNDA_2.n2294 16.0005
R6634 GNDA_2.n2294 GNDA_2.n2293 16.0005
R6635 GNDA_2.n2293 GNDA_2.n2290 16.0005
R6636 GNDA_2.n2290 GNDA_2.n2289 16.0005
R6637 GNDA_2.n2289 GNDA_2.n2286 16.0005
R6638 GNDA_2.n2286 GNDA_2.n2285 16.0005
R6639 GNDA_2.n2285 GNDA_2.n2282 16.0005
R6640 GNDA_2.n2281 GNDA_2.n2278 16.0005
R6641 GNDA_2.n2278 GNDA_2.n2277 16.0005
R6642 GNDA_2.n2277 GNDA_2.n2274 16.0005
R6643 GNDA_2.n2274 GNDA_2.n2273 16.0005
R6644 GNDA_2.n2273 GNDA_2.n2270 16.0005
R6645 GNDA_2.n2270 GNDA_2.n2269 16.0005
R6646 GNDA_2.n2269 GNDA_2.n2266 16.0005
R6647 GNDA_2.n2266 GNDA_2.n2265 16.0005
R6648 GNDA_2.n1765 GNDA_2.n1764 16.0005
R6649 GNDA_2.n1768 GNDA_2.n1765 16.0005
R6650 GNDA_2.n1769 GNDA_2.n1768 16.0005
R6651 GNDA_2.n1772 GNDA_2.n1769 16.0005
R6652 GNDA_2.n1773 GNDA_2.n1772 16.0005
R6653 GNDA_2.n1776 GNDA_2.n1773 16.0005
R6654 GNDA_2.n1778 GNDA_2.n1776 16.0005
R6655 GNDA_2.n1779 GNDA_2.n1778 16.0005
R6656 GNDA_2.n1761 GNDA_2.n1760 16.0005
R6657 GNDA_2.n1760 GNDA_2.n1757 16.0005
R6658 GNDA_2.n1757 GNDA_2.n1756 16.0005
R6659 GNDA_2.n1756 GNDA_2.n1753 16.0005
R6660 GNDA_2.n1753 GNDA_2.n1752 16.0005
R6661 GNDA_2.n1752 GNDA_2.n1749 16.0005
R6662 GNDA_2.n1749 GNDA_2.n1748 16.0005
R6663 GNDA_2.n1748 GNDA_2.n1745 16.0005
R6664 GNDA_2.n1744 GNDA_2.n1741 16.0005
R6665 GNDA_2.n1741 GNDA_2.n1740 16.0005
R6666 GNDA_2.n1740 GNDA_2.n1737 16.0005
R6667 GNDA_2.n1737 GNDA_2.n1736 16.0005
R6668 GNDA_2.n1736 GNDA_2.n1733 16.0005
R6669 GNDA_2.n1733 GNDA_2.n1732 16.0005
R6670 GNDA_2.n1732 GNDA_2.n1729 16.0005
R6671 GNDA_2.n1729 GNDA_2.n1672 16.0005
R6672 GNDA_2.n5337 GNDA_2.n5336 16.0005
R6673 GNDA_2.n5340 GNDA_2.n5337 16.0005
R6674 GNDA_2.n5341 GNDA_2.n5340 16.0005
R6675 GNDA_2.n5344 GNDA_2.n5341 16.0005
R6676 GNDA_2.n5345 GNDA_2.n5344 16.0005
R6677 GNDA_2.n5348 GNDA_2.n5345 16.0005
R6678 GNDA_2.n5350 GNDA_2.n5348 16.0005
R6679 GNDA_2.n5351 GNDA_2.n5350 16.0005
R6680 GNDA_2.n5333 GNDA_2.n5332 16.0005
R6681 GNDA_2.n5332 GNDA_2.n5329 16.0005
R6682 GNDA_2.n5329 GNDA_2.n5328 16.0005
R6683 GNDA_2.n5328 GNDA_2.n5325 16.0005
R6684 GNDA_2.n5325 GNDA_2.n5324 16.0005
R6685 GNDA_2.n5324 GNDA_2.n5321 16.0005
R6686 GNDA_2.n5321 GNDA_2.n5320 16.0005
R6687 GNDA_2.n5320 GNDA_2.n5317 16.0005
R6688 GNDA_2.n5316 GNDA_2.n5313 16.0005
R6689 GNDA_2.n5313 GNDA_2.n5312 16.0005
R6690 GNDA_2.n5312 GNDA_2.n5309 16.0005
R6691 GNDA_2.n5309 GNDA_2.n5308 16.0005
R6692 GNDA_2.n5308 GNDA_2.n5305 16.0005
R6693 GNDA_2.n5305 GNDA_2.n5304 16.0005
R6694 GNDA_2.n5304 GNDA_2.n5301 16.0005
R6695 GNDA_2.n5301 GNDA_2.n5300 16.0005
R6696 GNDA_2.t252 GNDA_2.t73 15.0244
R6697 GNDA_2.t30 GNDA_2.t73 15.0244
R6698 GNDA_2.t165 GNDA_2.t139 15.0244
R6699 GNDA_2.t274 GNDA_2.t208 14.8654
R6700 GNDA_2.t228 GNDA_2.t185 14.8654
R6701 GNDA_2.t277 GNDA_2.t202 14.8654
R6702 GNDA_2.t192 GNDA_2.t18 14.8654
R6703 GNDA_2.n5551 GNDA_2.n26 14.555
R6704 GNDA_2.n2598 GNDA_2.n1850 14.555
R6705 GNDA_2.t164 GNDA_2.t150 14.554
R6706 GNDA_2.t61 GNDA_2.t223 14.554
R6707 GNDA_2.t170 GNDA_2.t46 14.554
R6708 GNDA_2.t25 GNDA_2.t121 14.554
R6709 GNDA_2.n4354 GNDA_2.n4353 14.238
R6710 GNDA_2.n381 GNDA_2.n380 14.238
R6711 GNDA_2.t66 GNDA_2.t280 13.8109
R6712 GNDA_2.n4476 GNDA_2.n4475 13.5941
R6713 GNDA_2.n4303 GNDA_2.n1092 13.5941
R6714 GNDA_2.n4618 GNDA_2.n180 13.5697
R6715 GNDA_2.n4306 GNDA_2.n4305 13.5697
R6716 GNDA_2.n4341 GNDA_2.n385 12.8005
R6717 GNDA_2.n4337 GNDA_2.n385 12.8005
R6718 GNDA_2.n598 GNDA_2.n597 12.8005
R6719 GNDA_2.n598 GNDA_2.n387 12.8005
R6720 GNDA_2.n369 GNDA_2.n349 12.8005
R6721 GNDA_2.n375 GNDA_2.n369 12.8005
R6722 GNDA_2.n4359 GNDA_2.n350 12.8005
R6723 GNDA_2.n4355 GNDA_2.n350 12.8005
R6724 GNDA_2.n4403 GNDA_2.n336 12.8005
R6725 GNDA_2.n4403 GNDA_2.n4402 12.8005
R6726 GNDA_2.n4459 GNDA_2.n304 12.8005
R6727 GNDA_2.n4459 GNDA_2.n305 12.8005
R6728 GNDA_2.n2816 GNDA_2.n2671 12.8005
R6729 GNDA_2.n2820 GNDA_2.n2671 12.8005
R6730 GNDA_2.n2697 GNDA_2.n2696 12.8005
R6731 GNDA_2.n2696 GNDA_2.n2690 12.8005
R6732 GNDA_2.n3066 GNDA_2.n2973 12.8005
R6733 GNDA_2.n3167 GNDA_2.n2973 12.8005
R6734 GNDA_2.n4471 GNDA_2.t159 12.6791
R6735 GNDA_2.n4620 GNDA_2.t135 12.6791
R6736 GNDA_2.n4208 GNDA_2.t91 12.6791
R6737 GNDA_2.n4313 GNDA_2.t113 12.6791
R6738 GNDA_2.t51 GNDA_2.t54 12.5036
R6739 GNDA_2.t215 GNDA_2.t184 12.5036
R6740 GNDA_2.t150 GNDA_2.t15 12.1284
R6741 GNDA_2.t286 GNDA_2.t164 12.1284
R6742 GNDA_2.t223 GNDA_2.t41 12.1284
R6743 GNDA_2.t205 GNDA_2.t61 12.1284
R6744 GNDA_2.t238 GNDA_2.t170 12.1284
R6745 GNDA_2.t46 GNDA_2.t229 12.1284
R6746 GNDA_2.t233 GNDA_2.t25 12.1284
R6747 GNDA_2.t121 GNDA_2.t43 12.1284
R6748 GNDA_2.t11 GNDA_2.n2855 12.0196
R6749 GNDA_2.t44 GNDA_2.n2795 12.0196
R6750 GNDA_2.n3355 GNDA_2.t272 12.0196
R6751 GNDA_2.n3263 GNDA_2.n3262 11.6369
R6752 GNDA_2.n3262 GNDA_2.n3261 11.6369
R6753 GNDA_2.n3261 GNDA_2.n3260 11.6369
R6754 GNDA_2.n3260 GNDA_2.n3258 11.6369
R6755 GNDA_2.n3258 GNDA_2.n3255 11.6369
R6756 GNDA_2.n3255 GNDA_2.n3254 11.6369
R6757 GNDA_2.n3254 GNDA_2.n3251 11.6369
R6758 GNDA_2.n3251 GNDA_2.n3250 11.6369
R6759 GNDA_2.n3250 GNDA_2.n3247 11.6369
R6760 GNDA_2.n3247 GNDA_2.n3246 11.6369
R6761 GNDA_2.n3243 GNDA_2.n3242 11.6369
R6762 GNDA_2.n3242 GNDA_2.n2949 11.6369
R6763 GNDA_2.n3236 GNDA_2.n2949 11.6369
R6764 GNDA_2.n3236 GNDA_2.n3235 11.6369
R6765 GNDA_2.n3235 GNDA_2.n3234 11.6369
R6766 GNDA_2.n3234 GNDA_2.n2954 11.6369
R6767 GNDA_2.n3228 GNDA_2.n2954 11.6369
R6768 GNDA_2.n3228 GNDA_2.n3227 11.6369
R6769 GNDA_2.n3227 GNDA_2.n3226 11.6369
R6770 GNDA_2.n3226 GNDA_2.n2958 11.6369
R6771 GNDA_2.n3220 GNDA_2.n2958 11.6369
R6772 GNDA_2.n1963 GNDA_2.n1962 11.6369
R6773 GNDA_2.n1962 GNDA_2.n1959 11.6369
R6774 GNDA_2.n1959 GNDA_2.n1958 11.6369
R6775 GNDA_2.n1958 GNDA_2.n1955 11.6369
R6776 GNDA_2.n1955 GNDA_2.n1954 11.6369
R6777 GNDA_2.n1954 GNDA_2.n1951 11.6369
R6778 GNDA_2.n1951 GNDA_2.n1950 11.6369
R6779 GNDA_2.n1950 GNDA_2.n1947 11.6369
R6780 GNDA_2.n1947 GNDA_2.n1946 11.6369
R6781 GNDA_2.n1946 GNDA_2.n1846 11.6369
R6782 GNDA_2.n1967 GNDA_2.n1966 11.6369
R6783 GNDA_2.n1970 GNDA_2.n1967 11.6369
R6784 GNDA_2.n1971 GNDA_2.n1970 11.6369
R6785 GNDA_2.n1974 GNDA_2.n1971 11.6369
R6786 GNDA_2.n1975 GNDA_2.n1974 11.6369
R6787 GNDA_2.n1978 GNDA_2.n1975 11.6369
R6788 GNDA_2.n1979 GNDA_2.n1978 11.6369
R6789 GNDA_2.n1982 GNDA_2.n1979 11.6369
R6790 GNDA_2.n1984 GNDA_2.n1982 11.6369
R6791 GNDA_2.n1985 GNDA_2.n1984 11.6369
R6792 GNDA_2.n1986 GNDA_2.n1985 11.6369
R6793 GNDA_2.n3270 GNDA_2.n3269 11.6369
R6794 GNDA_2.n3269 GNDA_2.n1829 11.6369
R6795 GNDA_2.n2943 GNDA_2.n1829 11.6369
R6796 GNDA_2.n2943 GNDA_2.n2942 11.6369
R6797 GNDA_2.n2942 GNDA_2.n2941 11.6369
R6798 GNDA_2.n2941 GNDA_2.n2938 11.6369
R6799 GNDA_2.n2938 GNDA_2.n2937 11.6369
R6800 GNDA_2.n2937 GNDA_2.n2934 11.6369
R6801 GNDA_2.n2934 GNDA_2.n2933 11.6369
R6802 GNDA_2.n2933 GNDA_2.n2930 11.6369
R6803 GNDA_2.n2501 GNDA_2.n1937 11.6369
R6804 GNDA_2.n2501 GNDA_2.n2500 11.6369
R6805 GNDA_2.n2500 GNDA_2.n2499 11.6369
R6806 GNDA_2.n2499 GNDA_2.n1991 11.6369
R6807 GNDA_2.n2494 GNDA_2.n1991 11.6369
R6808 GNDA_2.n2494 GNDA_2.n2493 11.6369
R6809 GNDA_2.n2493 GNDA_2.n2492 11.6369
R6810 GNDA_2.n2492 GNDA_2.n1994 11.6369
R6811 GNDA_2.n2487 GNDA_2.n1994 11.6369
R6812 GNDA_2.n2487 GNDA_2.n2486 11.6369
R6813 GNDA_2.n2486 GNDA_2.n2485 11.6369
R6814 GNDA_2.n2182 GNDA_2.n2181 11.6369
R6815 GNDA_2.n2187 GNDA_2.n2182 11.6369
R6816 GNDA_2.n2188 GNDA_2.n2187 11.6369
R6817 GNDA_2.n2189 GNDA_2.n2188 11.6369
R6818 GNDA_2.n2189 GNDA_2.n2179 11.6369
R6819 GNDA_2.n2195 GNDA_2.n2179 11.6369
R6820 GNDA_2.n2196 GNDA_2.n2195 11.6369
R6821 GNDA_2.n2197 GNDA_2.n2196 11.6369
R6822 GNDA_2.n2197 GNDA_2.n2177 11.6369
R6823 GNDA_2.n2202 GNDA_2.n2177 11.6369
R6824 GNDA_2.n2203 GNDA_2.n2202 11.6369
R6825 GNDA_2.n2209 GNDA_2.n2175 11.6369
R6826 GNDA_2.n2210 GNDA_2.n2209 11.6369
R6827 GNDA_2.n2212 GNDA_2.n2210 11.6369
R6828 GNDA_2.n2212 GNDA_2.n2211 11.6369
R6829 GNDA_2.n2211 GNDA_2.n2172 11.6369
R6830 GNDA_2.n2172 GNDA_2.n2170 11.6369
R6831 GNDA_2.n2222 GNDA_2.n2170 11.6369
R6832 GNDA_2.n2223 GNDA_2.n2222 11.6369
R6833 GNDA_2.n2225 GNDA_2.n2223 11.6369
R6834 GNDA_2.n2225 GNDA_2.n2224 11.6369
R6835 GNDA_2.n2386 GNDA_2.n2329 11.6369
R6836 GNDA_2.n2386 GNDA_2.n2385 11.6369
R6837 GNDA_2.n2385 GNDA_2.n2384 11.6369
R6838 GNDA_2.n2384 GNDA_2.n2332 11.6369
R6839 GNDA_2.n2379 GNDA_2.n2332 11.6369
R6840 GNDA_2.n2379 GNDA_2.n2378 11.6369
R6841 GNDA_2.n2378 GNDA_2.n2377 11.6369
R6842 GNDA_2.n2377 GNDA_2.n2335 11.6369
R6843 GNDA_2.n2372 GNDA_2.n2335 11.6369
R6844 GNDA_2.n2372 GNDA_2.n2371 11.6369
R6845 GNDA_2.n2371 GNDA_2.n2370 11.6369
R6846 GNDA_2.n2343 GNDA_2.n2338 11.6369
R6847 GNDA_2.n2363 GNDA_2.n2343 11.6369
R6848 GNDA_2.n2363 GNDA_2.n2362 11.6369
R6849 GNDA_2.n2362 GNDA_2.n2361 11.6369
R6850 GNDA_2.n2361 GNDA_2.n2344 11.6369
R6851 GNDA_2.n2356 GNDA_2.n2344 11.6369
R6852 GNDA_2.n2356 GNDA_2.n2355 11.6369
R6853 GNDA_2.n2355 GNDA_2.n2354 11.6369
R6854 GNDA_2.n2354 GNDA_2.n2346 11.6369
R6855 GNDA_2.n2346 GNDA_2.n1673 11.6369
R6856 GNDA_2.n5260 GNDA_2.n126 11.6369
R6857 GNDA_2.n5261 GNDA_2.n5260 11.6369
R6858 GNDA_2.n5263 GNDA_2.n5261 11.6369
R6859 GNDA_2.n5263 GNDA_2.n5262 11.6369
R6860 GNDA_2.n5262 GNDA_2.n123 11.6369
R6861 GNDA_2.n123 GNDA_2.n121 11.6369
R6862 GNDA_2.n5273 GNDA_2.n121 11.6369
R6863 GNDA_2.n5274 GNDA_2.n5273 11.6369
R6864 GNDA_2.n5276 GNDA_2.n5274 11.6369
R6865 GNDA_2.n5276 GNDA_2.n5275 11.6369
R6866 GNDA_2.n3150 GNDA_2.n3149 11.6369
R6867 GNDA_2.n3149 GNDA_2.n3148 11.6369
R6868 GNDA_2.n3148 GNDA_2.n3119 11.6369
R6869 GNDA_2.n3142 GNDA_2.n3119 11.6369
R6870 GNDA_2.n3142 GNDA_2.n3141 11.6369
R6871 GNDA_2.n3141 GNDA_2.n3140 11.6369
R6872 GNDA_2.n3140 GNDA_2.n3123 11.6369
R6873 GNDA_2.n3134 GNDA_2.n3123 11.6369
R6874 GNDA_2.n3134 GNDA_2.n3133 11.6369
R6875 GNDA_2.n3133 GNDA_2.n3132 11.6369
R6876 GNDA_2.n3132 GNDA_2.n3127 11.6369
R6877 GNDA_2.n2967 GNDA_2.n2962 11.6369
R6878 GNDA_2.n3174 GNDA_2.n2967 11.6369
R6879 GNDA_2.n3174 GNDA_2.n3173 11.6369
R6880 GNDA_2.n3173 GNDA_2.n3172 11.6369
R6881 GNDA_2.n3172 GNDA_2.n2968 11.6369
R6882 GNDA_2.n3165 GNDA_2.n3070 11.6369
R6883 GNDA_2.n3074 GNDA_2.n3070 11.6369
R6884 GNDA_2.n3158 GNDA_2.n3074 11.6369
R6885 GNDA_2.n3158 GNDA_2.n3157 11.6369
R6886 GNDA_2.n3157 GNDA_2.n3156 11.6369
R6887 GNDA_2.n2434 GNDA_2.n2433 11.6369
R6888 GNDA_2.n2435 GNDA_2.n2434 11.6369
R6889 GNDA_2.n2435 GNDA_2.n2430 11.6369
R6890 GNDA_2.n2441 GNDA_2.n2430 11.6369
R6891 GNDA_2.n2442 GNDA_2.n2441 11.6369
R6892 GNDA_2.n2443 GNDA_2.n2442 11.6369
R6893 GNDA_2.n2443 GNDA_2.n2428 11.6369
R6894 GNDA_2.n2448 GNDA_2.n2428 11.6369
R6895 GNDA_2.n2449 GNDA_2.n2448 11.6369
R6896 GNDA_2.n2449 GNDA_2.n2426 11.6369
R6897 GNDA_2.n2455 GNDA_2.n2426 11.6369
R6898 GNDA_2.n3271 GNDA_2.n1827 11.6369
R6899 GNDA_2.n3277 GNDA_2.n1827 11.6369
R6900 GNDA_2.n3278 GNDA_2.n3277 11.6369
R6901 GNDA_2.n3279 GNDA_2.n3278 11.6369
R6902 GNDA_2.n3279 GNDA_2.n1825 11.6369
R6903 GNDA_2.n3285 GNDA_2.n1825 11.6369
R6904 GNDA_2.n3286 GNDA_2.n3285 11.6369
R6905 GNDA_2.n3287 GNDA_2.n3286 11.6369
R6906 GNDA_2.n3287 GNDA_2.n1823 11.6369
R6907 GNDA_2.n3292 GNDA_2.n1823 11.6369
R6908 GNDA_2.n3293 GNDA_2.n3292 11.6369
R6909 GNDA_2.n2951 GNDA_2.t73 11.3072
R6910 GNDA_2.t171 GNDA_2.t51 11.0327
R6911 GNDA_2.t168 GNDA_2.t169 11.0327
R6912 GNDA_2.t169 GNDA_2.t214 11.0327
R6913 GNDA_2.t214 GNDA_2.t182 11.0327
R6914 GNDA_2.t193 GNDA_2.t289 11.0327
R6915 GNDA_2.t167 GNDA_2.t193 11.0327
R6916 GNDA_2.t279 GNDA_2.t167 11.0327
R6917 GNDA_2.t209 GNDA_2.t215 11.0327
R6918 GNDA_2.n3406 GNDA_2.n3405 10.9846
R6919 GNDA_2.t41 GNDA_2.n4323 10.9156
R6920 GNDA_2.t229 GNDA_2.n4325 10.9156
R6921 GNDA_2.n3409 GNDA_2.n1663 10.87
R6922 GNDA_2.n3410 GNDA_2.n1662 10.87
R6923 GNDA_2.n3414 GNDA_2.n1658 10.87
R6924 GNDA_2.n3415 GNDA_2.n1657 10.87
R6925 GNDA_2.n3419 GNDA_2.n1653 10.87
R6926 GNDA_2.n3420 GNDA_2.n1652 10.87
R6927 GNDA_2.n3423 GNDA_2.n1649 10.87
R6928 GNDA_2.n1832 GNDA_2.t34 9.66779
R6929 GNDA_2.n571 GNDA_2.t234 9.6005
R6930 GNDA_2.n571 GNDA_2.t122 9.6005
R6931 GNDA_2.n573 GNDA_2.t239 9.6005
R6932 GNDA_2.n573 GNDA_2.t47 9.6005
R6933 GNDA_2.n575 GNDA_2.t63 9.6005
R6934 GNDA_2.n575 GNDA_2.t197 9.6005
R6935 GNDA_2.n577 GNDA_2.t257 9.6005
R6936 GNDA_2.n577 GNDA_2.t200 9.6005
R6937 GNDA_2.n579 GNDA_2.t8 9.6005
R6938 GNDA_2.n579 GNDA_2.t40 9.6005
R6939 GNDA_2.n581 GNDA_2.t243 9.6005
R6940 GNDA_2.n581 GNDA_2.t64 9.6005
R6941 GNDA_2.n583 GNDA_2.t7 9.6005
R6942 GNDA_2.n583 GNDA_2.t39 9.6005
R6943 GNDA_2.n585 GNDA_2.t247 9.6005
R6944 GNDA_2.n585 GNDA_2.t32 9.6005
R6945 GNDA_2.n587 GNDA_2.t207 9.6005
R6946 GNDA_2.n587 GNDA_2.t212 9.6005
R6947 GNDA_2.n589 GNDA_2.t13 9.6005
R6948 GNDA_2.n589 GNDA_2.t57 9.6005
R6949 GNDA_2.n591 GNDA_2.t224 9.6005
R6950 GNDA_2.n591 GNDA_2.t206 9.6005
R6951 GNDA_2.n593 GNDA_2.t151 9.6005
R6952 GNDA_2.n593 GNDA_2.t287 9.6005
R6953 GNDA_2.n4383 GNDA_2.t187 9.6005
R6954 GNDA_2.n4383 GNDA_2.t53 9.6005
R6955 GNDA_2.n3373 GNDA_2.t259 9.6005
R6956 GNDA_2.n1685 GNDA_2.t262 9.6005
R6957 GNDA_2.n2828 GNDA_2.t264 9.6005
R6958 GNDA_2.n2837 GNDA_2.t268 9.6005
R6959 GNDA_2.n4374 GNDA_2.n4372 9.42329
R6960 GNDA_2.n4366 GNDA_2.n344 9.42293
R6961 GNDA_2.n375 GNDA_2.n374 9.36264
R6962 GNDA_2.n4359 GNDA_2.n4358 9.36264
R6963 GNDA_2.n4402 GNDA_2.n4401 9.36264
R6964 GNDA_2.n306 GNDA_2.n304 9.36264
R6965 GNDA_2.n2816 GNDA_2.n2669 9.36264
R6966 GNDA_2.n2697 GNDA_2.n2689 9.36264
R6967 GNDA_2.n3067 GNDA_2.n3066 9.36264
R6968 GNDA_2.n597 GNDA_2.n596 9.36264
R6969 GNDA_2.n4341 GNDA_2.n4340 9.36264
R6970 GNDA_2.n4339 GNDA_2.n385 9.3005
R6971 GNDA_2.n4338 GNDA_2.n4337 9.3005
R6972 GNDA_2.n599 GNDA_2.n598 9.3005
R6973 GNDA_2.n600 GNDA_2.n387 9.3005
R6974 GNDA_2.n370 GNDA_2.n369 9.3005
R6975 GNDA_2.n371 GNDA_2.n349 9.3005
R6976 GNDA_2.n4357 GNDA_2.n350 9.3005
R6977 GNDA_2.n4356 GNDA_2.n4355 9.3005
R6978 GNDA_2.n4403 GNDA_2.n337 9.3005
R6979 GNDA_2.n4398 GNDA_2.n336 9.3005
R6980 GNDA_2.n4459 GNDA_2.n4458 9.3005
R6981 GNDA_2.n4457 GNDA_2.n305 9.3005
R6982 GNDA_2.n2671 GNDA_2.n2670 9.3005
R6983 GNDA_2.n2821 GNDA_2.n2820 9.3005
R6984 GNDA_2.n2696 GNDA_2.n2695 9.3005
R6985 GNDA_2.n2694 GNDA_2.n2690 9.3005
R6986 GNDA_2.n2974 GNDA_2.n2973 9.3005
R6987 GNDA_2.n3167 GNDA_2.n3069 9.3005
R6988 GNDA_2.n3390 GNDA_2.n3388 8.62751
R6989 GNDA_2.n83 GNDA_2.n26 8.60107
R6990 GNDA_2.n1914 GNDA_2.n1850 8.60107
R6991 GNDA_2.n4326 GNDA_2.t205 8.49003
R6992 GNDA_2.n4326 GNDA_2.t238 8.49003
R6993 GNDA_2.t59 GNDA_2.t23 8.25876
R6994 GNDA_2.t237 GNDA_2.t216 8.25876
R6995 GNDA_2.t282 GNDA_2.t62 8.25876
R6996 GNDA_2.t178 GNDA_2.t190 8.25876
R6997 GNDA_2.n2926 GNDA_2.t130 8.01325
R6998 GNDA_2.t254 GNDA_2.n2645 8.01325
R6999 GNDA_2.t221 GNDA_2.n2781 8.01325
R7000 GNDA_2.t231 GNDA_2.n3356 8.01325
R7001 GNDA_2.t201 GNDA_2.n2653 7.01165
R7002 GNDA_2.t29 GNDA_2.n2856 7.01165
R7003 GNDA_2.n3220 GNDA_2.n3219 6.72373
R7004 GNDA_2.n1986 GNDA_2.n1935 6.72373
R7005 GNDA_2.n2485 GNDA_2.n1997 6.72373
R7006 GNDA_2.n3156 GNDA_2.n3075 6.72373
R7007 GNDA_2.n2456 GNDA_2.n2455 6.72373
R7008 GNDA_2.n3293 GNDA_2.n1821 6.72373
R7009 GNDA_2.n1937 GNDA_2.n1935 6.20656
R7010 GNDA_2.n2181 GNDA_2.n1997 6.20656
R7011 GNDA_2.n2456 GNDA_2.n2329 6.20656
R7012 GNDA_2.n3150 GNDA_2.n3075 6.20656
R7013 GNDA_2.n3219 GNDA_2.n2962 6.20656
R7014 GNDA_2.n2433 GNDA_2.n1821 6.20656
R7015 GNDA_2.n3166 GNDA_2.n2968 6.07727
R7016 GNDA_2.t276 GNDA_2.t73 6.01006
R7017 GNDA_2.n2838 GNDA_2.n2829 5.81868
R7018 GNDA_2.n2836 GNDA_2.n2829 5.81868
R7019 GNDA_2.n3166 GNDA_2.n3165 5.5601
R7020 GNDA_2.n5484 GNDA_2.n5462 5.51161
R7021 GNDA_2.n2538 GNDA_2.n2537 5.51161
R7022 GNDA_2.n2864 GNDA_2.n2642 5.51161
R7023 GNDA_2.n2809 GNDA_2.n2807 5.51161
R7024 GNDA_2.n2142 GNDA_2.n2026 5.51161
R7025 GNDA_2.n5392 GNDA_2.n5362 5.51161
R7026 GNDA_2.n2265 GNDA_2.n2235 5.51161
R7027 GNDA_2.n3399 GNDA_2.n1672 5.51161
R7028 GNDA_2.n5300 GNDA_2.n5286 5.51161
R7029 GNDA_2.n4319 GNDA_2.t194 5.3776
R7030 GNDA_2.n2234 GNDA_2.n2165 5.1717
R7031 GNDA_2.n3398 GNDA_2.n3397 5.1717
R7032 GNDA_2.n5285 GNDA_2.n116 5.1717
R7033 GNDA_2.t162 GNDA_2.t176 5.00847
R7034 GNDA_2.n2840 GNDA_2.t252 5.00847
R7035 GNDA_2.t73 GNDA_2.t78 5.00847
R7036 GNDA_2.n3379 GNDA_2.t30 5.00847
R7037 GNDA_2.t270 GNDA_2.t35 5.00847
R7038 GNDA_2.n5548 GNDA_2.n56 4.9157
R7039 GNDA_2.n2604 GNDA_2.n2603 4.9157
R7040 GNDA_2.n2929 GNDA_2.n2928 4.9157
R7041 GNDA_2.n373 GNDA_2.n372 4.663
R7042 GNDA_2.n368 GNDA_2.n351 4.663
R7043 GNDA_2.n4400 GNDA_2.n4399 4.663
R7044 GNDA_2.n4456 GNDA_2.n307 4.663
R7045 GNDA_2.n4353 GNDA_2.n4349 4.64112
R7046 GNDA_2.n4353 GNDA_2.n4352 4.64112
R7047 GNDA_2.n380 GNDA_2.n376 4.64112
R7048 GNDA_2.n380 GNDA_2.n379 4.64112
R7049 GNDA_2.n1067 GNDA_2.n1066 4.5005
R7050 GNDA_2.n1065 GNDA_2.n401 4.5005
R7051 GNDA_2.n1064 GNDA_2.n1063 4.5005
R7052 GNDA_2.n1062 GNDA_2.n405 4.5005
R7053 GNDA_2.n1061 GNDA_2.n1060 4.5005
R7054 GNDA_2.n1059 GNDA_2.n406 4.5005
R7055 GNDA_2.n1058 GNDA_2.n1057 4.5005
R7056 GNDA_2.n1056 GNDA_2.n410 4.5005
R7057 GNDA_2.n1055 GNDA_2.n1054 4.5005
R7058 GNDA_2.n1053 GNDA_2.n411 4.5005
R7059 GNDA_2.n1052 GNDA_2.n1051 4.5005
R7060 GNDA_2.n1050 GNDA_2.n415 4.5005
R7061 GNDA_2.n1049 GNDA_2.n1048 4.5005
R7062 GNDA_2.n1047 GNDA_2.n416 4.5005
R7063 GNDA_2.n1046 GNDA_2.n1045 4.5005
R7064 GNDA_2.n1044 GNDA_2.n420 4.5005
R7065 GNDA_2.n1043 GNDA_2.n1042 4.5005
R7066 GNDA_2.n1041 GNDA_2.n421 4.5005
R7067 GNDA_2.n1040 GNDA_2.n1039 4.5005
R7068 GNDA_2.n1038 GNDA_2.n425 4.5005
R7069 GNDA_2.n1037 GNDA_2.n1036 4.5005
R7070 GNDA_2.n1035 GNDA_2.n426 4.5005
R7071 GNDA_2.n5066 GNDA_2.n5065 4.5005
R7072 GNDA_2.n4904 GNDA_2.n4903 4.5005
R7073 GNDA_2.n5011 GNDA_2.n5010 4.5005
R7074 GNDA_2.n5015 GNDA_2.n5012 4.5005
R7075 GNDA_2.n5016 GNDA_2.n5009 4.5005
R7076 GNDA_2.n5020 GNDA_2.n5019 4.5005
R7077 GNDA_2.n5021 GNDA_2.n5008 4.5005
R7078 GNDA_2.n5025 GNDA_2.n5022 4.5005
R7079 GNDA_2.n5026 GNDA_2.n5007 4.5005
R7080 GNDA_2.n5030 GNDA_2.n5029 4.5005
R7081 GNDA_2.n5031 GNDA_2.n5006 4.5005
R7082 GNDA_2.n5035 GNDA_2.n5032 4.5005
R7083 GNDA_2.n5036 GNDA_2.n5005 4.5005
R7084 GNDA_2.n5040 GNDA_2.n5039 4.5005
R7085 GNDA_2.n5041 GNDA_2.n5004 4.5005
R7086 GNDA_2.n5045 GNDA_2.n5042 4.5005
R7087 GNDA_2.n5046 GNDA_2.n5003 4.5005
R7088 GNDA_2.n5050 GNDA_2.n5049 4.5005
R7089 GNDA_2.n5051 GNDA_2.n5002 4.5005
R7090 GNDA_2.n5055 GNDA_2.n5052 4.5005
R7091 GNDA_2.n5056 GNDA_2.n5001 4.5005
R7092 GNDA_2.n5060 GNDA_2.n5059 4.5005
R7093 GNDA_2.n4931 GNDA_2.n4930 4.5005
R7094 GNDA_2.n4934 GNDA_2.n4933 4.5005
R7095 GNDA_2.n4935 GNDA_2.n4929 4.5005
R7096 GNDA_2.n4939 GNDA_2.n4936 4.5005
R7097 GNDA_2.n4940 GNDA_2.n4928 4.5005
R7098 GNDA_2.n4944 GNDA_2.n4943 4.5005
R7099 GNDA_2.n4945 GNDA_2.n4927 4.5005
R7100 GNDA_2.n4949 GNDA_2.n4946 4.5005
R7101 GNDA_2.n4950 GNDA_2.n4926 4.5005
R7102 GNDA_2.n4954 GNDA_2.n4953 4.5005
R7103 GNDA_2.n4955 GNDA_2.n4925 4.5005
R7104 GNDA_2.n4959 GNDA_2.n4956 4.5005
R7105 GNDA_2.n4960 GNDA_2.n4924 4.5005
R7106 GNDA_2.n4964 GNDA_2.n4963 4.5005
R7107 GNDA_2.n4965 GNDA_2.n4923 4.5005
R7108 GNDA_2.n4969 GNDA_2.n4966 4.5005
R7109 GNDA_2.n4970 GNDA_2.n4922 4.5005
R7110 GNDA_2.n4974 GNDA_2.n4973 4.5005
R7111 GNDA_2.n4975 GNDA_2.n4921 4.5005
R7112 GNDA_2.n4979 GNDA_2.n4976 4.5005
R7113 GNDA_2.n4980 GNDA_2.n4920 4.5005
R7114 GNDA_2.n4984 GNDA_2.n4983 4.5005
R7115 GNDA_2.n4892 GNDA_2.n4891 4.5005
R7116 GNDA_2.n4813 GNDA_2.n4812 4.5005
R7117 GNDA_2.n4835 GNDA_2.n4814 4.5005
R7118 GNDA_2.n4836 GNDA_2.n4815 4.5005
R7119 GNDA_2.n4837 GNDA_2.n4816 4.5005
R7120 GNDA_2.n4838 GNDA_2.n4817 4.5005
R7121 GNDA_2.n4839 GNDA_2.n4818 4.5005
R7122 GNDA_2.n4840 GNDA_2.n4819 4.5005
R7123 GNDA_2.n4841 GNDA_2.n4820 4.5005
R7124 GNDA_2.n4842 GNDA_2.n4821 4.5005
R7125 GNDA_2.n4843 GNDA_2.n4822 4.5005
R7126 GNDA_2.n4844 GNDA_2.n4823 4.5005
R7127 GNDA_2.n4845 GNDA_2.n4824 4.5005
R7128 GNDA_2.n4846 GNDA_2.n4825 4.5005
R7129 GNDA_2.n4847 GNDA_2.n4826 4.5005
R7130 GNDA_2.n4848 GNDA_2.n4827 4.5005
R7131 GNDA_2.n4849 GNDA_2.n4828 4.5005
R7132 GNDA_2.n4850 GNDA_2.n4829 4.5005
R7133 GNDA_2.n4851 GNDA_2.n4830 4.5005
R7134 GNDA_2.n4852 GNDA_2.n4831 4.5005
R7135 GNDA_2.n4853 GNDA_2.n4832 4.5005
R7136 GNDA_2.n4854 GNDA_2.n4833 4.5005
R7137 GNDA_2.n5091 GNDA_2.n5090 4.5005
R7138 GNDA_2.n5094 GNDA_2.n5093 4.5005
R7139 GNDA_2.n5095 GNDA_2.n4808 4.5005
R7140 GNDA_2.n5099 GNDA_2.n5096 4.5005
R7141 GNDA_2.n5100 GNDA_2.n4807 4.5005
R7142 GNDA_2.n5104 GNDA_2.n5103 4.5005
R7143 GNDA_2.n5105 GNDA_2.n4806 4.5005
R7144 GNDA_2.n5109 GNDA_2.n5106 4.5005
R7145 GNDA_2.n5110 GNDA_2.n4805 4.5005
R7146 GNDA_2.n5114 GNDA_2.n5113 4.5005
R7147 GNDA_2.n5115 GNDA_2.n4804 4.5005
R7148 GNDA_2.n5119 GNDA_2.n5116 4.5005
R7149 GNDA_2.n5120 GNDA_2.n4803 4.5005
R7150 GNDA_2.n5124 GNDA_2.n5123 4.5005
R7151 GNDA_2.n5125 GNDA_2.n4802 4.5005
R7152 GNDA_2.n5129 GNDA_2.n5126 4.5005
R7153 GNDA_2.n5130 GNDA_2.n4801 4.5005
R7154 GNDA_2.n5134 GNDA_2.n5133 4.5005
R7155 GNDA_2.n5135 GNDA_2.n4800 4.5005
R7156 GNDA_2.n5139 GNDA_2.n5136 4.5005
R7157 GNDA_2.n5140 GNDA_2.n4799 4.5005
R7158 GNDA_2.n5144 GNDA_2.n5143 4.5005
R7159 GNDA_2.n4614 GNDA_2.n4613 4.5005
R7160 GNDA_2.n185 GNDA_2.n184 4.5005
R7161 GNDA_2.n4559 GNDA_2.n4558 4.5005
R7162 GNDA_2.n4563 GNDA_2.n4560 4.5005
R7163 GNDA_2.n4564 GNDA_2.n4557 4.5005
R7164 GNDA_2.n4568 GNDA_2.n4567 4.5005
R7165 GNDA_2.n4569 GNDA_2.n4556 4.5005
R7166 GNDA_2.n4573 GNDA_2.n4570 4.5005
R7167 GNDA_2.n4574 GNDA_2.n4555 4.5005
R7168 GNDA_2.n4578 GNDA_2.n4577 4.5005
R7169 GNDA_2.n4579 GNDA_2.n4554 4.5005
R7170 GNDA_2.n4583 GNDA_2.n4580 4.5005
R7171 GNDA_2.n4584 GNDA_2.n4553 4.5005
R7172 GNDA_2.n4588 GNDA_2.n4587 4.5005
R7173 GNDA_2.n4589 GNDA_2.n4552 4.5005
R7174 GNDA_2.n4593 GNDA_2.n4590 4.5005
R7175 GNDA_2.n4594 GNDA_2.n4551 4.5005
R7176 GNDA_2.n4598 GNDA_2.n4597 4.5005
R7177 GNDA_2.n4599 GNDA_2.n4550 4.5005
R7178 GNDA_2.n4603 GNDA_2.n4600 4.5005
R7179 GNDA_2.n4604 GNDA_2.n4549 4.5005
R7180 GNDA_2.n4608 GNDA_2.n4607 4.5005
R7181 GNDA_2.n5215 GNDA_2.n5214 4.5005
R7182 GNDA_2.n145 GNDA_2.n144 4.5005
R7183 GNDA_2.n5160 GNDA_2.n5159 4.5005
R7184 GNDA_2.n5164 GNDA_2.n5161 4.5005
R7185 GNDA_2.n5165 GNDA_2.n5158 4.5005
R7186 GNDA_2.n5169 GNDA_2.n5168 4.5005
R7187 GNDA_2.n5170 GNDA_2.n5157 4.5005
R7188 GNDA_2.n5174 GNDA_2.n5171 4.5005
R7189 GNDA_2.n5175 GNDA_2.n5156 4.5005
R7190 GNDA_2.n5179 GNDA_2.n5178 4.5005
R7191 GNDA_2.n5180 GNDA_2.n5155 4.5005
R7192 GNDA_2.n5184 GNDA_2.n5181 4.5005
R7193 GNDA_2.n5185 GNDA_2.n5154 4.5005
R7194 GNDA_2.n5189 GNDA_2.n5188 4.5005
R7195 GNDA_2.n5190 GNDA_2.n5153 4.5005
R7196 GNDA_2.n5194 GNDA_2.n5191 4.5005
R7197 GNDA_2.n5195 GNDA_2.n5152 4.5005
R7198 GNDA_2.n5199 GNDA_2.n5198 4.5005
R7199 GNDA_2.n5200 GNDA_2.n5151 4.5005
R7200 GNDA_2.n5204 GNDA_2.n5201 4.5005
R7201 GNDA_2.n5205 GNDA_2.n5150 4.5005
R7202 GNDA_2.n5209 GNDA_2.n5208 4.5005
R7203 GNDA_2.n4716 GNDA_2.n4715 4.5005
R7204 GNDA_2.n4719 GNDA_2.n4718 4.5005
R7205 GNDA_2.n4720 GNDA_2.n171 4.5005
R7206 GNDA_2.n4724 GNDA_2.n4721 4.5005
R7207 GNDA_2.n4725 GNDA_2.n170 4.5005
R7208 GNDA_2.n4729 GNDA_2.n4728 4.5005
R7209 GNDA_2.n4730 GNDA_2.n169 4.5005
R7210 GNDA_2.n4734 GNDA_2.n4731 4.5005
R7211 GNDA_2.n4735 GNDA_2.n168 4.5005
R7212 GNDA_2.n4739 GNDA_2.n4738 4.5005
R7213 GNDA_2.n4740 GNDA_2.n167 4.5005
R7214 GNDA_2.n4744 GNDA_2.n4741 4.5005
R7215 GNDA_2.n4745 GNDA_2.n166 4.5005
R7216 GNDA_2.n4749 GNDA_2.n4748 4.5005
R7217 GNDA_2.n4750 GNDA_2.n165 4.5005
R7218 GNDA_2.n4754 GNDA_2.n4751 4.5005
R7219 GNDA_2.n4755 GNDA_2.n164 4.5005
R7220 GNDA_2.n4759 GNDA_2.n4758 4.5005
R7221 GNDA_2.n4760 GNDA_2.n163 4.5005
R7222 GNDA_2.n4764 GNDA_2.n4761 4.5005
R7223 GNDA_2.n4765 GNDA_2.n162 4.5005
R7224 GNDA_2.n4769 GNDA_2.n4768 4.5005
R7225 GNDA_2.n4704 GNDA_2.n4703 4.5005
R7226 GNDA_2.n4625 GNDA_2.n4624 4.5005
R7227 GNDA_2.n4647 GNDA_2.n4626 4.5005
R7228 GNDA_2.n4648 GNDA_2.n4627 4.5005
R7229 GNDA_2.n4649 GNDA_2.n4628 4.5005
R7230 GNDA_2.n4650 GNDA_2.n4629 4.5005
R7231 GNDA_2.n4651 GNDA_2.n4630 4.5005
R7232 GNDA_2.n4652 GNDA_2.n4631 4.5005
R7233 GNDA_2.n4653 GNDA_2.n4632 4.5005
R7234 GNDA_2.n4654 GNDA_2.n4633 4.5005
R7235 GNDA_2.n4655 GNDA_2.n4634 4.5005
R7236 GNDA_2.n4656 GNDA_2.n4635 4.5005
R7237 GNDA_2.n4657 GNDA_2.n4636 4.5005
R7238 GNDA_2.n4658 GNDA_2.n4637 4.5005
R7239 GNDA_2.n4659 GNDA_2.n4638 4.5005
R7240 GNDA_2.n4660 GNDA_2.n4639 4.5005
R7241 GNDA_2.n4661 GNDA_2.n4640 4.5005
R7242 GNDA_2.n4662 GNDA_2.n4641 4.5005
R7243 GNDA_2.n4663 GNDA_2.n4642 4.5005
R7244 GNDA_2.n4664 GNDA_2.n4643 4.5005
R7245 GNDA_2.n4665 GNDA_2.n4644 4.5005
R7246 GNDA_2.n4666 GNDA_2.n4645 4.5005
R7247 GNDA_2.n4479 GNDA_2.n4478 4.5005
R7248 GNDA_2.n4482 GNDA_2.n4481 4.5005
R7249 GNDA_2.n4483 GNDA_2.n211 4.5005
R7250 GNDA_2.n4487 GNDA_2.n4484 4.5005
R7251 GNDA_2.n4488 GNDA_2.n210 4.5005
R7252 GNDA_2.n4492 GNDA_2.n4491 4.5005
R7253 GNDA_2.n4493 GNDA_2.n209 4.5005
R7254 GNDA_2.n4497 GNDA_2.n4494 4.5005
R7255 GNDA_2.n4498 GNDA_2.n208 4.5005
R7256 GNDA_2.n4502 GNDA_2.n4501 4.5005
R7257 GNDA_2.n4503 GNDA_2.n207 4.5005
R7258 GNDA_2.n4507 GNDA_2.n4504 4.5005
R7259 GNDA_2.n4508 GNDA_2.n206 4.5005
R7260 GNDA_2.n4512 GNDA_2.n4511 4.5005
R7261 GNDA_2.n4513 GNDA_2.n205 4.5005
R7262 GNDA_2.n4517 GNDA_2.n4514 4.5005
R7263 GNDA_2.n4518 GNDA_2.n204 4.5005
R7264 GNDA_2.n4522 GNDA_2.n4521 4.5005
R7265 GNDA_2.n4523 GNDA_2.n203 4.5005
R7266 GNDA_2.n4527 GNDA_2.n4524 4.5005
R7267 GNDA_2.n4528 GNDA_2.n202 4.5005
R7268 GNDA_2.n4532 GNDA_2.n4531 4.5005
R7269 GNDA_2.n5244 GNDA_2.n5243 4.5005
R7270 GNDA_2.n5251 GNDA_2.n134 4.5005
R7271 GNDA_2.n5250 GNDA_2.n5249 4.5005
R7272 GNDA_2.n5251 GNDA_2.n5250 4.5005
R7273 GNDA_2.n373 GNDA_2.n371 4.5005
R7274 GNDA_2.n4356 GNDA_2.n368 4.5005
R7275 GNDA_2.n4436 GNDA_2.n4435 4.5005
R7276 GNDA_2.n4441 GNDA_2.n4427 4.5005
R7277 GNDA_2.n4443 GNDA_2.n4442 4.5005
R7278 GNDA_2.n4442 GNDA_2.n4441 4.5005
R7279 GNDA_2.n4400 GNDA_2.n4398 4.5005
R7280 GNDA_2.n4457 GNDA_2.n4456 4.5005
R7281 GNDA_2.n311 GNDA_2.n309 4.5005
R7282 GNDA_2.n314 GNDA_2.n313 4.5005
R7283 GNDA_2.n365 GNDA_2.n353 4.5005
R7284 GNDA_2.n356 GNDA_2.n355 4.5005
R7285 GNDA_2.n4381 GNDA_2.n4375 4.5005
R7286 GNDA_2.n4378 GNDA_2.n310 4.5005
R7287 GNDA_2.n4381 GNDA_2.n310 4.5005
R7288 GNDA_2.n4389 GNDA_2.n4388 4.5005
R7289 GNDA_2.n4397 GNDA_2.n4396 4.5005
R7290 GNDA_2.n4396 GNDA_2.n4395 4.5005
R7291 GNDA_2.n4395 GNDA_2.n4393 4.5005
R7292 GNDA_2.n4426 GNDA_2.n4425 4.5005
R7293 GNDA_2.n4425 GNDA_2.n4424 4.5005
R7294 GNDA_2.n4424 GNDA_2.n323 4.5005
R7295 GNDA_2.n4421 GNDA_2.n325 4.5005
R7296 GNDA_2.n4421 GNDA_2.n4420 4.5005
R7297 GNDA_2.n4420 GNDA_2.n326 4.5005
R7298 GNDA_2.n4411 GNDA_2.n328 4.5005
R7299 GNDA_2.n4413 GNDA_2.n4412 4.5005
R7300 GNDA_2.n4412 GNDA_2.n4411 4.5005
R7301 GNDA_2.n3996 GNDA_2.n3995 4.5005
R7302 GNDA_2.n4003 GNDA_2.n4002 4.5005
R7303 GNDA_2.n4301 GNDA_2.n4300 4.5005
R7304 GNDA_2.n4299 GNDA_2.n1093 4.5005
R7305 GNDA_2.n4298 GNDA_2.n4297 4.5005
R7306 GNDA_2.n4296 GNDA_2.n1097 4.5005
R7307 GNDA_2.n4295 GNDA_2.n4294 4.5005
R7308 GNDA_2.n4293 GNDA_2.n1098 4.5005
R7309 GNDA_2.n4292 GNDA_2.n4291 4.5005
R7310 GNDA_2.n4290 GNDA_2.n1102 4.5005
R7311 GNDA_2.n4289 GNDA_2.n4288 4.5005
R7312 GNDA_2.n4287 GNDA_2.n1103 4.5005
R7313 GNDA_2.n4286 GNDA_2.n4285 4.5005
R7314 GNDA_2.n4284 GNDA_2.n1107 4.5005
R7315 GNDA_2.n4283 GNDA_2.n4282 4.5005
R7316 GNDA_2.n4281 GNDA_2.n1108 4.5005
R7317 GNDA_2.n4280 GNDA_2.n4279 4.5005
R7318 GNDA_2.n4278 GNDA_2.n1112 4.5005
R7319 GNDA_2.n4277 GNDA_2.n4276 4.5005
R7320 GNDA_2.n4275 GNDA_2.n1113 4.5005
R7321 GNDA_2.n4274 GNDA_2.n4273 4.5005
R7322 GNDA_2.n4272 GNDA_2.n1117 4.5005
R7323 GNDA_2.n4271 GNDA_2.n4270 4.5005
R7324 GNDA_2.n4269 GNDA_2.n1118 4.5005
R7325 GNDA_2.n4218 GNDA_2.n4217 4.5005
R7326 GNDA_2.n4221 GNDA_2.n4220 4.5005
R7327 GNDA_2.n4222 GNDA_2.n4203 4.5005
R7328 GNDA_2.n4224 GNDA_2.n4223 4.5005
R7329 GNDA_2.n4225 GNDA_2.n4202 4.5005
R7330 GNDA_2.n4229 GNDA_2.n4228 4.5005
R7331 GNDA_2.n4230 GNDA_2.n4199 4.5005
R7332 GNDA_2.n4232 GNDA_2.n4231 4.5005
R7333 GNDA_2.n4233 GNDA_2.n4198 4.5005
R7334 GNDA_2.n4237 GNDA_2.n4236 4.5005
R7335 GNDA_2.n4238 GNDA_2.n4195 4.5005
R7336 GNDA_2.n4240 GNDA_2.n4239 4.5005
R7337 GNDA_2.n4241 GNDA_2.n4194 4.5005
R7338 GNDA_2.n4245 GNDA_2.n4244 4.5005
R7339 GNDA_2.n4246 GNDA_2.n4191 4.5005
R7340 GNDA_2.n4248 GNDA_2.n4247 4.5005
R7341 GNDA_2.n4249 GNDA_2.n4190 4.5005
R7342 GNDA_2.n4253 GNDA_2.n4252 4.5005
R7343 GNDA_2.n4254 GNDA_2.n4187 4.5005
R7344 GNDA_2.n4256 GNDA_2.n4255 4.5005
R7345 GNDA_2.n4257 GNDA_2.n4186 4.5005
R7346 GNDA_2.n4261 GNDA_2.n4260 4.5005
R7347 GNDA_2.n4109 GNDA_2.n1089 4.5005
R7348 GNDA_2.n4112 GNDA_2.n4111 4.5005
R7349 GNDA_2.n4113 GNDA_2.n4106 4.5005
R7350 GNDA_2.n4115 GNDA_2.n4114 4.5005
R7351 GNDA_2.n4116 GNDA_2.n4105 4.5005
R7352 GNDA_2.n4120 GNDA_2.n4119 4.5005
R7353 GNDA_2.n4121 GNDA_2.n4102 4.5005
R7354 GNDA_2.n4123 GNDA_2.n4122 4.5005
R7355 GNDA_2.n4124 GNDA_2.n4101 4.5005
R7356 GNDA_2.n4128 GNDA_2.n4127 4.5005
R7357 GNDA_2.n4129 GNDA_2.n4098 4.5005
R7358 GNDA_2.n4131 GNDA_2.n4130 4.5005
R7359 GNDA_2.n4132 GNDA_2.n4097 4.5005
R7360 GNDA_2.n4136 GNDA_2.n4135 4.5005
R7361 GNDA_2.n4137 GNDA_2.n4094 4.5005
R7362 GNDA_2.n4139 GNDA_2.n4138 4.5005
R7363 GNDA_2.n4140 GNDA_2.n4093 4.5005
R7364 GNDA_2.n4144 GNDA_2.n4143 4.5005
R7365 GNDA_2.n4145 GNDA_2.n4090 4.5005
R7366 GNDA_2.n4147 GNDA_2.n4146 4.5005
R7367 GNDA_2.n4148 GNDA_2.n4089 4.5005
R7368 GNDA_2.n4152 GNDA_2.n4151 4.5005
R7369 GNDA_2.n4028 GNDA_2.n4027 4.5005
R7370 GNDA_2.n4031 GNDA_2.n4030 4.5005
R7371 GNDA_2.n4032 GNDA_2.n1154 4.5005
R7372 GNDA_2.n4034 GNDA_2.n4033 4.5005
R7373 GNDA_2.n4035 GNDA_2.n1153 4.5005
R7374 GNDA_2.n4039 GNDA_2.n4038 4.5005
R7375 GNDA_2.n4040 GNDA_2.n1150 4.5005
R7376 GNDA_2.n4042 GNDA_2.n4041 4.5005
R7377 GNDA_2.n4043 GNDA_2.n1149 4.5005
R7378 GNDA_2.n4047 GNDA_2.n4046 4.5005
R7379 GNDA_2.n4048 GNDA_2.n1146 4.5005
R7380 GNDA_2.n4050 GNDA_2.n4049 4.5005
R7381 GNDA_2.n4051 GNDA_2.n1145 4.5005
R7382 GNDA_2.n4055 GNDA_2.n4054 4.5005
R7383 GNDA_2.n4056 GNDA_2.n1142 4.5005
R7384 GNDA_2.n4058 GNDA_2.n4057 4.5005
R7385 GNDA_2.n4059 GNDA_2.n1141 4.5005
R7386 GNDA_2.n4063 GNDA_2.n4062 4.5005
R7387 GNDA_2.n4064 GNDA_2.n1138 4.5005
R7388 GNDA_2.n4066 GNDA_2.n4065 4.5005
R7389 GNDA_2.n4067 GNDA_2.n1137 4.5005
R7390 GNDA_2.n4071 GNDA_2.n4070 4.5005
R7391 GNDA_2.n1241 GNDA_2.n1240 4.5005
R7392 GNDA_2.n1239 GNDA_2.n1161 4.5005
R7393 GNDA_2.n1238 GNDA_2.n1237 4.5005
R7394 GNDA_2.n1236 GNDA_2.n1166 4.5005
R7395 GNDA_2.n1235 GNDA_2.n1234 4.5005
R7396 GNDA_2.n1233 GNDA_2.n1167 4.5005
R7397 GNDA_2.n1232 GNDA_2.n1231 4.5005
R7398 GNDA_2.n1230 GNDA_2.n1174 4.5005
R7399 GNDA_2.n1229 GNDA_2.n1228 4.5005
R7400 GNDA_2.n1227 GNDA_2.n1175 4.5005
R7401 GNDA_2.n1226 GNDA_2.n1225 4.5005
R7402 GNDA_2.n1224 GNDA_2.n1182 4.5005
R7403 GNDA_2.n1223 GNDA_2.n1222 4.5005
R7404 GNDA_2.n1221 GNDA_2.n1183 4.5005
R7405 GNDA_2.n1220 GNDA_2.n1219 4.5005
R7406 GNDA_2.n1218 GNDA_2.n1190 4.5005
R7407 GNDA_2.n1217 GNDA_2.n1216 4.5005
R7408 GNDA_2.n1215 GNDA_2.n1191 4.5005
R7409 GNDA_2.n1214 GNDA_2.n1213 4.5005
R7410 GNDA_2.n1212 GNDA_2.n1198 4.5005
R7411 GNDA_2.n1211 GNDA_2.n1210 4.5005
R7412 GNDA_2.n1209 GNDA_2.n1199 4.5005
R7413 GNDA_2.n3635 GNDA_2.n1245 4.5005
R7414 GNDA_2.n3638 GNDA_2.n3637 4.5005
R7415 GNDA_2.n3639 GNDA_2.n3632 4.5005
R7416 GNDA_2.n3641 GNDA_2.n3640 4.5005
R7417 GNDA_2.n3642 GNDA_2.n3631 4.5005
R7418 GNDA_2.n3646 GNDA_2.n3645 4.5005
R7419 GNDA_2.n3647 GNDA_2.n3628 4.5005
R7420 GNDA_2.n3649 GNDA_2.n3648 4.5005
R7421 GNDA_2.n3650 GNDA_2.n3627 4.5005
R7422 GNDA_2.n3654 GNDA_2.n3653 4.5005
R7423 GNDA_2.n3655 GNDA_2.n3624 4.5005
R7424 GNDA_2.n3657 GNDA_2.n3656 4.5005
R7425 GNDA_2.n3658 GNDA_2.n3623 4.5005
R7426 GNDA_2.n3662 GNDA_2.n3661 4.5005
R7427 GNDA_2.n3663 GNDA_2.n3620 4.5005
R7428 GNDA_2.n3665 GNDA_2.n3664 4.5005
R7429 GNDA_2.n3666 GNDA_2.n3619 4.5005
R7430 GNDA_2.n3670 GNDA_2.n3669 4.5005
R7431 GNDA_2.n3671 GNDA_2.n3616 4.5005
R7432 GNDA_2.n3673 GNDA_2.n3672 4.5005
R7433 GNDA_2.n3674 GNDA_2.n3615 4.5005
R7434 GNDA_2.n3678 GNDA_2.n3677 4.5005
R7435 GNDA_2.n3704 GNDA_2.n1252 4.5005
R7436 GNDA_2.n3707 GNDA_2.n3706 4.5005
R7437 GNDA_2.n3708 GNDA_2.n3701 4.5005
R7438 GNDA_2.n3710 GNDA_2.n3709 4.5005
R7439 GNDA_2.n3711 GNDA_2.n3700 4.5005
R7440 GNDA_2.n3715 GNDA_2.n3714 4.5005
R7441 GNDA_2.n3716 GNDA_2.n3697 4.5005
R7442 GNDA_2.n3718 GNDA_2.n3717 4.5005
R7443 GNDA_2.n3719 GNDA_2.n3696 4.5005
R7444 GNDA_2.n3723 GNDA_2.n3722 4.5005
R7445 GNDA_2.n3724 GNDA_2.n3693 4.5005
R7446 GNDA_2.n3726 GNDA_2.n3725 4.5005
R7447 GNDA_2.n3727 GNDA_2.n3692 4.5005
R7448 GNDA_2.n3731 GNDA_2.n3730 4.5005
R7449 GNDA_2.n3732 GNDA_2.n3689 4.5005
R7450 GNDA_2.n3734 GNDA_2.n3733 4.5005
R7451 GNDA_2.n3735 GNDA_2.n3688 4.5005
R7452 GNDA_2.n3739 GNDA_2.n3738 4.5005
R7453 GNDA_2.n3740 GNDA_2.n3685 4.5005
R7454 GNDA_2.n3742 GNDA_2.n3741 4.5005
R7455 GNDA_2.n3743 GNDA_2.n3684 4.5005
R7456 GNDA_2.n3747 GNDA_2.n3746 4.5005
R7457 GNDA_2.n3773 GNDA_2.n1256 4.5005
R7458 GNDA_2.n3776 GNDA_2.n3775 4.5005
R7459 GNDA_2.n3777 GNDA_2.n3770 4.5005
R7460 GNDA_2.n3779 GNDA_2.n3778 4.5005
R7461 GNDA_2.n3780 GNDA_2.n3769 4.5005
R7462 GNDA_2.n3784 GNDA_2.n3783 4.5005
R7463 GNDA_2.n3785 GNDA_2.n3766 4.5005
R7464 GNDA_2.n3787 GNDA_2.n3786 4.5005
R7465 GNDA_2.n3788 GNDA_2.n3765 4.5005
R7466 GNDA_2.n3792 GNDA_2.n3791 4.5005
R7467 GNDA_2.n3793 GNDA_2.n3762 4.5005
R7468 GNDA_2.n3795 GNDA_2.n3794 4.5005
R7469 GNDA_2.n3796 GNDA_2.n3761 4.5005
R7470 GNDA_2.n3800 GNDA_2.n3799 4.5005
R7471 GNDA_2.n3801 GNDA_2.n3758 4.5005
R7472 GNDA_2.n3803 GNDA_2.n3802 4.5005
R7473 GNDA_2.n3804 GNDA_2.n3757 4.5005
R7474 GNDA_2.n3808 GNDA_2.n3807 4.5005
R7475 GNDA_2.n3809 GNDA_2.n3754 4.5005
R7476 GNDA_2.n3811 GNDA_2.n3810 4.5005
R7477 GNDA_2.n3812 GNDA_2.n3753 4.5005
R7478 GNDA_2.n3816 GNDA_2.n3815 4.5005
R7479 GNDA_2.n3842 GNDA_2.n1260 4.5005
R7480 GNDA_2.n3845 GNDA_2.n3844 4.5005
R7481 GNDA_2.n3846 GNDA_2.n3839 4.5005
R7482 GNDA_2.n3848 GNDA_2.n3847 4.5005
R7483 GNDA_2.n3849 GNDA_2.n3838 4.5005
R7484 GNDA_2.n3853 GNDA_2.n3852 4.5005
R7485 GNDA_2.n3854 GNDA_2.n3835 4.5005
R7486 GNDA_2.n3856 GNDA_2.n3855 4.5005
R7487 GNDA_2.n3857 GNDA_2.n3834 4.5005
R7488 GNDA_2.n3861 GNDA_2.n3860 4.5005
R7489 GNDA_2.n3862 GNDA_2.n3831 4.5005
R7490 GNDA_2.n3864 GNDA_2.n3863 4.5005
R7491 GNDA_2.n3865 GNDA_2.n3830 4.5005
R7492 GNDA_2.n3869 GNDA_2.n3868 4.5005
R7493 GNDA_2.n3870 GNDA_2.n3827 4.5005
R7494 GNDA_2.n3872 GNDA_2.n3871 4.5005
R7495 GNDA_2.n3873 GNDA_2.n3826 4.5005
R7496 GNDA_2.n3877 GNDA_2.n3876 4.5005
R7497 GNDA_2.n3878 GNDA_2.n3823 4.5005
R7498 GNDA_2.n3880 GNDA_2.n3879 4.5005
R7499 GNDA_2.n3881 GNDA_2.n3822 4.5005
R7500 GNDA_2.n3885 GNDA_2.n3884 4.5005
R7501 GNDA_2.n3964 GNDA_2.n3962 4.5005
R7502 GNDA_2.n3966 GNDA_2.n3965 4.5005
R7503 GNDA_2.n3965 GNDA_2.n3964 4.5005
R7504 GNDA_2.n3969 GNDA_2.n3967 4.5005
R7505 GNDA_2.n3971 GNDA_2.n3970 4.5005
R7506 GNDA_2.n3970 GNDA_2.n3969 4.5005
R7507 GNDA_2.n3974 GNDA_2.n3972 4.5005
R7508 GNDA_2.n3976 GNDA_2.n3975 4.5005
R7509 GNDA_2.n3975 GNDA_2.n3974 4.5005
R7510 GNDA_2.n4013 GNDA_2.n4011 4.5005
R7511 GNDA_2.n4015 GNDA_2.n4014 4.5005
R7512 GNDA_2.n4014 GNDA_2.n4013 4.5005
R7513 GNDA_2.n4018 GNDA_2.n4016 4.5005
R7514 GNDA_2.n4020 GNDA_2.n4019 4.5005
R7515 GNDA_2.n4019 GNDA_2.n4018 4.5005
R7516 GNDA_2.n4025 GNDA_2.n4021 4.5005
R7517 GNDA_2.n4026 GNDA_2.n1085 4.5005
R7518 GNDA_2.n4026 GNDA_2.n4025 4.5005
R7519 GNDA_2.n4310 GNDA_2.n1086 4.5005
R7520 GNDA_2.n4309 GNDA_2.n4308 4.5005
R7521 GNDA_2.n4310 GNDA_2.n4309 4.5005
R7522 GNDA_2.n4215 GNDA_2.n4211 4.5005
R7523 GNDA_2.n4216 GNDA_2.n4207 4.5005
R7524 GNDA_2.n4216 GNDA_2.n4215 4.5005
R7525 GNDA_2.n4008 GNDA_2.n3977 4.5005
R7526 GNDA_2.n4010 GNDA_2.n4009 4.5005
R7527 GNDA_2.n4009 GNDA_2.n4008 4.5005
R7528 GNDA_2.n1263 GNDA_2.n1262 4.5005
R7529 GNDA_2.n3956 GNDA_2.n3955 4.5005
R7530 GNDA_2.n1265 GNDA_2.n1264 4.5005
R7531 GNDA_2.n3901 GNDA_2.n3900 4.5005
R7532 GNDA_2.n3905 GNDA_2.n3902 4.5005
R7533 GNDA_2.n3906 GNDA_2.n3899 4.5005
R7534 GNDA_2.n3910 GNDA_2.n3909 4.5005
R7535 GNDA_2.n3911 GNDA_2.n3898 4.5005
R7536 GNDA_2.n3915 GNDA_2.n3912 4.5005
R7537 GNDA_2.n3916 GNDA_2.n3897 4.5005
R7538 GNDA_2.n3920 GNDA_2.n3919 4.5005
R7539 GNDA_2.n3921 GNDA_2.n3896 4.5005
R7540 GNDA_2.n3925 GNDA_2.n3922 4.5005
R7541 GNDA_2.n3926 GNDA_2.n3895 4.5005
R7542 GNDA_2.n3930 GNDA_2.n3929 4.5005
R7543 GNDA_2.n3931 GNDA_2.n3894 4.5005
R7544 GNDA_2.n3935 GNDA_2.n3932 4.5005
R7545 GNDA_2.n3936 GNDA_2.n3893 4.5005
R7546 GNDA_2.n3940 GNDA_2.n3939 4.5005
R7547 GNDA_2.n3941 GNDA_2.n3892 4.5005
R7548 GNDA_2.n3945 GNDA_2.n3942 4.5005
R7549 GNDA_2.n3946 GNDA_2.n3891 4.5005
R7550 GNDA_2.n3950 GNDA_2.n3949 4.5005
R7551 GNDA_2.n2694 GNDA_2.n2693 4.5005
R7552 GNDA_2.n2822 GNDA_2.n2821 4.5005
R7553 GNDA_2.n2667 GNDA_2.n2666 4.5005
R7554 GNDA_2.n2827 GNDA_2.n2660 4.5005
R7555 GNDA_2.n2826 GNDA_2.n1683 4.5005
R7556 GNDA_2.n2827 GNDA_2.n2826 4.5005
R7557 GNDA_2.n3069 GNDA_2.n3068 4.5005
R7558 GNDA_2.n3058 GNDA_2.n2976 4.5005
R7559 GNDA_2.n1682 GNDA_2.n1681 4.5005
R7560 GNDA_2.n2998 GNDA_2.n2997 4.5005
R7561 GNDA_2.n3008 GNDA_2.n3007 4.5005
R7562 GNDA_2.n3009 GNDA_2.n2996 4.5005
R7563 GNDA_2.n3011 GNDA_2.n3010 4.5005
R7564 GNDA_2.n2994 GNDA_2.n2993 4.5005
R7565 GNDA_2.n3018 GNDA_2.n3017 4.5005
R7566 GNDA_2.n3019 GNDA_2.n2992 4.5005
R7567 GNDA_2.n3021 GNDA_2.n3020 4.5005
R7568 GNDA_2.n2990 GNDA_2.n2989 4.5005
R7569 GNDA_2.n3028 GNDA_2.n3027 4.5005
R7570 GNDA_2.n3029 GNDA_2.n2988 4.5005
R7571 GNDA_2.n3031 GNDA_2.n3030 4.5005
R7572 GNDA_2.n2986 GNDA_2.n2985 4.5005
R7573 GNDA_2.n3038 GNDA_2.n3037 4.5005
R7574 GNDA_2.n3039 GNDA_2.n2984 4.5005
R7575 GNDA_2.n3041 GNDA_2.n3040 4.5005
R7576 GNDA_2.n2982 GNDA_2.n2981 4.5005
R7577 GNDA_2.n3048 GNDA_2.n3047 4.5005
R7578 GNDA_2.n3049 GNDA_2.n2980 4.5005
R7579 GNDA_2.n3051 GNDA_2.n3050 4.5005
R7580 GNDA_2.n2978 GNDA_2.n2977 4.5005
R7581 GNDA_2.n3057 GNDA_2.n3056 4.5005
R7582 GNDA_2.n1643 GNDA_2.n1642 4.5005
R7583 GNDA_2.n1646 GNDA_2.n1645 4.5005
R7584 GNDA_2.n1590 GNDA_2.n1586 4.5005
R7585 GNDA_2.n1594 GNDA_2.n1591 4.5005
R7586 GNDA_2.n1595 GNDA_2.n1585 4.5005
R7587 GNDA_2.n1599 GNDA_2.n1598 4.5005
R7588 GNDA_2.n1600 GNDA_2.n1584 4.5005
R7589 GNDA_2.n1604 GNDA_2.n1601 4.5005
R7590 GNDA_2.n1605 GNDA_2.n1583 4.5005
R7591 GNDA_2.n1609 GNDA_2.n1608 4.5005
R7592 GNDA_2.n1610 GNDA_2.n1582 4.5005
R7593 GNDA_2.n1614 GNDA_2.n1611 4.5005
R7594 GNDA_2.n1615 GNDA_2.n1581 4.5005
R7595 GNDA_2.n1619 GNDA_2.n1618 4.5005
R7596 GNDA_2.n1620 GNDA_2.n1580 4.5005
R7597 GNDA_2.n1624 GNDA_2.n1621 4.5005
R7598 GNDA_2.n1625 GNDA_2.n1579 4.5005
R7599 GNDA_2.n1629 GNDA_2.n1628 4.5005
R7600 GNDA_2.n1630 GNDA_2.n1578 4.5005
R7601 GNDA_2.n1634 GNDA_2.n1631 4.5005
R7602 GNDA_2.n1635 GNDA_2.n1577 4.5005
R7603 GNDA_2.n1639 GNDA_2.n1638 4.5005
R7604 GNDA_2.n1640 GNDA_2.n1576 4.5005
R7605 GNDA_2.n3435 GNDA_2.n3434 4.5005
R7606 GNDA_2.n294 GNDA_2.n293 4.5005
R7607 GNDA_2.n292 GNDA_2.n215 4.5005
R7608 GNDA_2.n291 GNDA_2.n290 4.5005
R7609 GNDA_2.n289 GNDA_2.n219 4.5005
R7610 GNDA_2.n288 GNDA_2.n287 4.5005
R7611 GNDA_2.n286 GNDA_2.n220 4.5005
R7612 GNDA_2.n285 GNDA_2.n284 4.5005
R7613 GNDA_2.n283 GNDA_2.n227 4.5005
R7614 GNDA_2.n282 GNDA_2.n281 4.5005
R7615 GNDA_2.n280 GNDA_2.n228 4.5005
R7616 GNDA_2.n279 GNDA_2.n278 4.5005
R7617 GNDA_2.n277 GNDA_2.n235 4.5005
R7618 GNDA_2.n276 GNDA_2.n275 4.5005
R7619 GNDA_2.n274 GNDA_2.n236 4.5005
R7620 GNDA_2.n273 GNDA_2.n272 4.5005
R7621 GNDA_2.n271 GNDA_2.n243 4.5005
R7622 GNDA_2.n270 GNDA_2.n269 4.5005
R7623 GNDA_2.n268 GNDA_2.n244 4.5005
R7624 GNDA_2.n267 GNDA_2.n266 4.5005
R7625 GNDA_2.n265 GNDA_2.n251 4.5005
R7626 GNDA_2.n264 GNDA_2.n263 4.5005
R7627 GNDA_2.n262 GNDA_2.n252 4.5005
R7628 GNDA_2.n297 GNDA_2.n295 4.5005
R7629 GNDA_2.n299 GNDA_2.n298 4.5005
R7630 GNDA_2.n298 GNDA_2.n297 4.5005
R7631 GNDA_2.n4709 GNDA_2.n4708 4.5005
R7632 GNDA_2.n4708 GNDA_2.n4707 4.5005
R7633 GNDA_2.n4707 GNDA_2.n4623 4.5005
R7634 GNDA_2.n4710 GNDA_2.n142 4.5005
R7635 GNDA_2.n4711 GNDA_2.n4710 4.5005
R7636 GNDA_2.n4712 GNDA_2.n4711 4.5005
R7637 GNDA_2.n5220 GNDA_2.n5219 4.5005
R7638 GNDA_2.n5219 GNDA_2.n5218 4.5005
R7639 GNDA_2.n5218 GNDA_2.n143 4.5005
R7640 GNDA_2.n4619 GNDA_2.n4618 4.5005
R7641 GNDA_2.n4618 GNDA_2.n4617 4.5005
R7642 GNDA_2.n4617 GNDA_2.n183 4.5005
R7643 GNDA_2.n5085 GNDA_2.n5082 4.5005
R7644 GNDA_2.n5086 GNDA_2.n5085 4.5005
R7645 GNDA_2.n5087 GNDA_2.n5086 4.5005
R7646 GNDA_2.n5078 GNDA_2.n4811 4.5005
R7647 GNDA_2.n5081 GNDA_2.n4811 4.5005
R7648 GNDA_2.n5081 GNDA_2.n4810 4.5005
R7649 GNDA_2.n5074 GNDA_2.n4897 4.5005
R7650 GNDA_2.n5077 GNDA_2.n4897 4.5005
R7651 GNDA_2.n5077 GNDA_2.n4896 4.5005
R7652 GNDA_2.n5070 GNDA_2.n4902 4.5005
R7653 GNDA_2.n5073 GNDA_2.n4902 4.5005
R7654 GNDA_2.n5073 GNDA_2.n4901 4.5005
R7655 GNDA_2.n5226 GNDA_2.n138 4.5005
R7656 GNDA_2.n5226 GNDA_2.n5225 4.5005
R7657 GNDA_2.n5225 GNDA_2.n5221 4.5005
R7658 GNDA_2.n399 GNDA_2.n390 4.5005
R7659 GNDA_2.n397 GNDA_2.n393 4.5005
R7660 GNDA_2.n398 GNDA_2.n392 4.5005
R7661 GNDA_2.n398 GNDA_2.n397 4.5005
R7662 GNDA_2.n601 GNDA_2.n600 4.5005
R7663 GNDA_2.n4338 GNDA_2.n386 4.5005
R7664 GNDA_2.n605 GNDA_2.n604 4.5005
R7665 GNDA_2.n608 GNDA_2.n563 4.5005
R7666 GNDA_2.n609 GNDA_2.n608 4.5005
R7667 GNDA_2.n610 GNDA_2.n609 4.5005
R7668 GNDA_2.n652 GNDA_2.n651 4.5005
R7669 GNDA_2.n655 GNDA_2.n654 4.5005
R7670 GNDA_2.n656 GNDA_2.n648 4.5005
R7671 GNDA_2.n658 GNDA_2.n657 4.5005
R7672 GNDA_2.n659 GNDA_2.n647 4.5005
R7673 GNDA_2.n663 GNDA_2.n662 4.5005
R7674 GNDA_2.n664 GNDA_2.n644 4.5005
R7675 GNDA_2.n666 GNDA_2.n665 4.5005
R7676 GNDA_2.n667 GNDA_2.n643 4.5005
R7677 GNDA_2.n671 GNDA_2.n670 4.5005
R7678 GNDA_2.n672 GNDA_2.n640 4.5005
R7679 GNDA_2.n674 GNDA_2.n673 4.5005
R7680 GNDA_2.n675 GNDA_2.n639 4.5005
R7681 GNDA_2.n679 GNDA_2.n678 4.5005
R7682 GNDA_2.n680 GNDA_2.n636 4.5005
R7683 GNDA_2.n682 GNDA_2.n681 4.5005
R7684 GNDA_2.n683 GNDA_2.n635 4.5005
R7685 GNDA_2.n687 GNDA_2.n686 4.5005
R7686 GNDA_2.n688 GNDA_2.n632 4.5005
R7687 GNDA_2.n690 GNDA_2.n689 4.5005
R7688 GNDA_2.n691 GNDA_2.n631 4.5005
R7689 GNDA_2.n695 GNDA_2.n694 4.5005
R7690 GNDA_2.n968 GNDA_2.n967 4.5005
R7691 GNDA_2.n971 GNDA_2.n970 4.5005
R7692 GNDA_2.n972 GNDA_2.n462 4.5005
R7693 GNDA_2.n974 GNDA_2.n973 4.5005
R7694 GNDA_2.n975 GNDA_2.n461 4.5005
R7695 GNDA_2.n979 GNDA_2.n978 4.5005
R7696 GNDA_2.n980 GNDA_2.n458 4.5005
R7697 GNDA_2.n982 GNDA_2.n981 4.5005
R7698 GNDA_2.n983 GNDA_2.n457 4.5005
R7699 GNDA_2.n987 GNDA_2.n986 4.5005
R7700 GNDA_2.n988 GNDA_2.n454 4.5005
R7701 GNDA_2.n990 GNDA_2.n989 4.5005
R7702 GNDA_2.n991 GNDA_2.n453 4.5005
R7703 GNDA_2.n995 GNDA_2.n994 4.5005
R7704 GNDA_2.n996 GNDA_2.n450 4.5005
R7705 GNDA_2.n998 GNDA_2.n997 4.5005
R7706 GNDA_2.n999 GNDA_2.n449 4.5005
R7707 GNDA_2.n1003 GNDA_2.n1002 4.5005
R7708 GNDA_2.n1004 GNDA_2.n446 4.5005
R7709 GNDA_2.n1006 GNDA_2.n1005 4.5005
R7710 GNDA_2.n1007 GNDA_2.n445 4.5005
R7711 GNDA_2.n1011 GNDA_2.n1010 4.5005
R7712 GNDA_2.n549 GNDA_2.n548 4.5005
R7713 GNDA_2.n547 GNDA_2.n469 4.5005
R7714 GNDA_2.n546 GNDA_2.n545 4.5005
R7715 GNDA_2.n544 GNDA_2.n474 4.5005
R7716 GNDA_2.n543 GNDA_2.n542 4.5005
R7717 GNDA_2.n541 GNDA_2.n475 4.5005
R7718 GNDA_2.n540 GNDA_2.n539 4.5005
R7719 GNDA_2.n538 GNDA_2.n482 4.5005
R7720 GNDA_2.n537 GNDA_2.n536 4.5005
R7721 GNDA_2.n535 GNDA_2.n483 4.5005
R7722 GNDA_2.n534 GNDA_2.n533 4.5005
R7723 GNDA_2.n532 GNDA_2.n490 4.5005
R7724 GNDA_2.n531 GNDA_2.n530 4.5005
R7725 GNDA_2.n529 GNDA_2.n491 4.5005
R7726 GNDA_2.n528 GNDA_2.n527 4.5005
R7727 GNDA_2.n526 GNDA_2.n498 4.5005
R7728 GNDA_2.n525 GNDA_2.n524 4.5005
R7729 GNDA_2.n523 GNDA_2.n499 4.5005
R7730 GNDA_2.n522 GNDA_2.n521 4.5005
R7731 GNDA_2.n520 GNDA_2.n506 4.5005
R7732 GNDA_2.n519 GNDA_2.n518 4.5005
R7733 GNDA_2.n517 GNDA_2.n507 4.5005
R7734 GNDA_2.n756 GNDA_2.n553 4.5005
R7735 GNDA_2.n759 GNDA_2.n758 4.5005
R7736 GNDA_2.n760 GNDA_2.n753 4.5005
R7737 GNDA_2.n762 GNDA_2.n761 4.5005
R7738 GNDA_2.n763 GNDA_2.n752 4.5005
R7739 GNDA_2.n767 GNDA_2.n766 4.5005
R7740 GNDA_2.n768 GNDA_2.n749 4.5005
R7741 GNDA_2.n770 GNDA_2.n769 4.5005
R7742 GNDA_2.n771 GNDA_2.n748 4.5005
R7743 GNDA_2.n775 GNDA_2.n774 4.5005
R7744 GNDA_2.n776 GNDA_2.n745 4.5005
R7745 GNDA_2.n778 GNDA_2.n777 4.5005
R7746 GNDA_2.n779 GNDA_2.n744 4.5005
R7747 GNDA_2.n783 GNDA_2.n782 4.5005
R7748 GNDA_2.n784 GNDA_2.n741 4.5005
R7749 GNDA_2.n786 GNDA_2.n785 4.5005
R7750 GNDA_2.n787 GNDA_2.n740 4.5005
R7751 GNDA_2.n791 GNDA_2.n790 4.5005
R7752 GNDA_2.n792 GNDA_2.n737 4.5005
R7753 GNDA_2.n794 GNDA_2.n793 4.5005
R7754 GNDA_2.n795 GNDA_2.n736 4.5005
R7755 GNDA_2.n799 GNDA_2.n798 4.5005
R7756 GNDA_2.n825 GNDA_2.n557 4.5005
R7757 GNDA_2.n828 GNDA_2.n827 4.5005
R7758 GNDA_2.n829 GNDA_2.n822 4.5005
R7759 GNDA_2.n831 GNDA_2.n830 4.5005
R7760 GNDA_2.n832 GNDA_2.n821 4.5005
R7761 GNDA_2.n836 GNDA_2.n835 4.5005
R7762 GNDA_2.n837 GNDA_2.n818 4.5005
R7763 GNDA_2.n839 GNDA_2.n838 4.5005
R7764 GNDA_2.n840 GNDA_2.n817 4.5005
R7765 GNDA_2.n844 GNDA_2.n843 4.5005
R7766 GNDA_2.n845 GNDA_2.n814 4.5005
R7767 GNDA_2.n847 GNDA_2.n846 4.5005
R7768 GNDA_2.n848 GNDA_2.n813 4.5005
R7769 GNDA_2.n852 GNDA_2.n851 4.5005
R7770 GNDA_2.n853 GNDA_2.n810 4.5005
R7771 GNDA_2.n855 GNDA_2.n854 4.5005
R7772 GNDA_2.n856 GNDA_2.n809 4.5005
R7773 GNDA_2.n860 GNDA_2.n859 4.5005
R7774 GNDA_2.n861 GNDA_2.n806 4.5005
R7775 GNDA_2.n863 GNDA_2.n862 4.5005
R7776 GNDA_2.n864 GNDA_2.n805 4.5005
R7777 GNDA_2.n868 GNDA_2.n867 4.5005
R7778 GNDA_2.n948 GNDA_2.n946 4.5005
R7779 GNDA_2.n950 GNDA_2.n949 4.5005
R7780 GNDA_2.n949 GNDA_2.n948 4.5005
R7781 GNDA_2.n953 GNDA_2.n951 4.5005
R7782 GNDA_2.n955 GNDA_2.n954 4.5005
R7783 GNDA_2.n954 GNDA_2.n953 4.5005
R7784 GNDA_2.n958 GNDA_2.n956 4.5005
R7785 GNDA_2.n960 GNDA_2.n959 4.5005
R7786 GNDA_2.n959 GNDA_2.n958 4.5005
R7787 GNDA_2.n965 GNDA_2.n961 4.5005
R7788 GNDA_2.n966 GNDA_2.n400 4.5005
R7789 GNDA_2.n966 GNDA_2.n965 4.5005
R7790 GNDA_2.n560 GNDA_2.n559 4.5005
R7791 GNDA_2.n939 GNDA_2.n938 4.5005
R7792 GNDA_2.n615 GNDA_2.n614 4.5005
R7793 GNDA_2.n884 GNDA_2.n883 4.5005
R7794 GNDA_2.n888 GNDA_2.n885 4.5005
R7795 GNDA_2.n889 GNDA_2.n882 4.5005
R7796 GNDA_2.n893 GNDA_2.n892 4.5005
R7797 GNDA_2.n894 GNDA_2.n881 4.5005
R7798 GNDA_2.n898 GNDA_2.n895 4.5005
R7799 GNDA_2.n899 GNDA_2.n880 4.5005
R7800 GNDA_2.n903 GNDA_2.n902 4.5005
R7801 GNDA_2.n904 GNDA_2.n879 4.5005
R7802 GNDA_2.n908 GNDA_2.n905 4.5005
R7803 GNDA_2.n909 GNDA_2.n878 4.5005
R7804 GNDA_2.n913 GNDA_2.n912 4.5005
R7805 GNDA_2.n914 GNDA_2.n877 4.5005
R7806 GNDA_2.n918 GNDA_2.n915 4.5005
R7807 GNDA_2.n919 GNDA_2.n876 4.5005
R7808 GNDA_2.n923 GNDA_2.n922 4.5005
R7809 GNDA_2.n924 GNDA_2.n875 4.5005
R7810 GNDA_2.n928 GNDA_2.n925 4.5005
R7811 GNDA_2.n929 GNDA_2.n874 4.5005
R7812 GNDA_2.n933 GNDA_2.n932 4.5005
R7813 GNDA_2.n3116 GNDA_2.n3115 4.26717
R7814 GNDA_2.n3115 GNDA_2.n3114 4.26717
R7815 GNDA_2.n3114 GNDA_2.n3082 4.26717
R7816 GNDA_2.n3108 GNDA_2.n3082 4.26717
R7817 GNDA_2.n3108 GNDA_2.n3107 4.26717
R7818 GNDA_2.n3107 GNDA_2.n3106 4.26717
R7819 GNDA_2.n3106 GNDA_2.n3091 4.26717
R7820 GNDA_2.n3100 GNDA_2.n3091 4.26717
R7821 GNDA_2.n3100 GNDA_2.n3099 4.26717
R7822 GNDA_2.n3099 GNDA_2.n3098 4.26717
R7823 GNDA_2.n3098 GNDA_2.n113 4.26717
R7824 GNDA_2.n2482 GNDA_2.n2000 4.26717
R7825 GNDA_2.n2477 GNDA_2.n2000 4.26717
R7826 GNDA_2.n2477 GNDA_2.n2476 4.26717
R7827 GNDA_2.n2476 GNDA_2.n2475 4.26717
R7828 GNDA_2.n2475 GNDA_2.n2472 4.26717
R7829 GNDA_2.n2472 GNDA_2.n2471 4.26717
R7830 GNDA_2.n2471 GNDA_2.n2468 4.26717
R7831 GNDA_2.n2468 GNDA_2.n2467 4.26717
R7832 GNDA_2.n2467 GNDA_2.n2464 4.26717
R7833 GNDA_2.n2464 GNDA_2.n2463 4.26717
R7834 GNDA_2.n2463 GNDA_2.n2461 4.26717
R7835 GNDA_2.n2425 GNDA_2.n2330 4.26717
R7836 GNDA_2.n2420 GNDA_2.n2330 4.26717
R7837 GNDA_2.n2420 GNDA_2.n2419 4.26717
R7838 GNDA_2.n2419 GNDA_2.n2395 4.26717
R7839 GNDA_2.n2414 GNDA_2.n2395 4.26717
R7840 GNDA_2.n2414 GNDA_2.n2413 4.26717
R7841 GNDA_2.n2413 GNDA_2.n2412 4.26717
R7842 GNDA_2.n2412 GNDA_2.n2401 4.26717
R7843 GNDA_2.n2406 GNDA_2.n2401 4.26717
R7844 GNDA_2.n2406 GNDA_2.n2405 4.26717
R7845 GNDA_2.n2405 GNDA_2.n1785 4.26717
R7846 GNDA_2.n3297 GNDA_2.n1819 4.26717
R7847 GNDA_2.n3303 GNDA_2.n1819 4.26717
R7848 GNDA_2.n3303 GNDA_2.n1817 4.26717
R7849 GNDA_2.n3309 GNDA_2.n1817 4.26717
R7850 GNDA_2.n3309 GNDA_2.n1815 4.26717
R7851 GNDA_2.n3315 GNDA_2.n1815 4.26717
R7852 GNDA_2.n3315 GNDA_2.n1813 4.26717
R7853 GNDA_2.n3321 GNDA_2.n1813 4.26717
R7854 GNDA_2.n3321 GNDA_2.n1811 4.26717
R7855 GNDA_2.n3327 GNDA_2.n1811 4.26717
R7856 GNDA_2.n3327 GNDA_2.n1809 4.26717
R7857 GNDA_2.n2508 GNDA_2.n2507 4.26717
R7858 GNDA_2.n2511 GNDA_2.n2508 4.26717
R7859 GNDA_2.n2511 GNDA_2.n1931 4.26717
R7860 GNDA_2.n2517 GNDA_2.n1931 4.26717
R7861 GNDA_2.n2518 GNDA_2.n2517 4.26717
R7862 GNDA_2.n2521 GNDA_2.n2518 4.26717
R7863 GNDA_2.n2521 GNDA_2.n1929 4.26717
R7864 GNDA_2.n1929 GNDA_2.n1924 4.26717
R7865 GNDA_2.n2528 GNDA_2.n1924 4.26717
R7866 GNDA_2.n2528 GNDA_2.n1925 4.26717
R7867 GNDA_2.n1925 GNDA_2.n1916 4.26717
R7868 GNDA_2.n3218 GNDA_2.n2963 4.26717
R7869 GNDA_2.n3212 GNDA_2.n2963 4.26717
R7870 GNDA_2.n3212 GNDA_2.n3211 4.26717
R7871 GNDA_2.n3211 GNDA_2.n3210 4.26717
R7872 GNDA_2.n3210 GNDA_2.n3187 4.26717
R7873 GNDA_2.n3190 GNDA_2.n3187 4.26717
R7874 GNDA_2.n3201 GNDA_2.n3190 4.26717
R7875 GNDA_2.n3201 GNDA_2.n3200 4.26717
R7876 GNDA_2.n3200 GNDA_2.n3199 4.26717
R7877 GNDA_2.n3199 GNDA_2.n3195 4.26717
R7878 GNDA_2.n3195 GNDA_2.n86 4.26717
R7879 GNDA_2.t263 GNDA_2.t290 4.14363
R7880 GNDA_2.n3116 GNDA_2.n3075 3.93531
R7881 GNDA_2.n2482 GNDA_2.n1997 3.93531
R7882 GNDA_2.n2456 GNDA_2.n2425 3.93531
R7883 GNDA_2.n3297 GNDA_2.n1821 3.93531
R7884 GNDA_2.n2507 GNDA_2.n1935 3.93531
R7885 GNDA_2.n3219 GNDA_2.n3218 3.93531
R7886 GNDA_2.n4622 GNDA_2.n4621 3.84081
R7887 GNDA_2.n4210 GNDA_2.n4209 3.84081
R7888 GNDA_2.n4312 GNDA_2.n4311 3.84081
R7889 GNDA_2.n4473 GNDA_2.n4472 3.84045
R7890 GNDA_2.n5546 GNDA_2.n5545 3.7893
R7891 GNDA_2.n5542 GNDA_2.n59 3.7893
R7892 GNDA_2.n5541 GNDA_2.n62 3.7893
R7893 GNDA_2.n5538 GNDA_2.n5537 3.7893
R7894 GNDA_2.n5464 GNDA_2.n63 3.7893
R7895 GNDA_2.n5473 GNDA_2.n5472 3.7893
R7896 GNDA_2.n5476 GNDA_2.n5463 3.7893
R7897 GNDA_2.n5481 GNDA_2.n5477 3.7893
R7898 GNDA_2.n2601 GNDA_2.n1848 3.7893
R7899 GNDA_2.n1869 GNDA_2.n1868 3.7893
R7900 GNDA_2.n2595 GNDA_2.n2594 3.7893
R7901 GNDA_2.n1893 GNDA_2.n1870 3.7893
R7902 GNDA_2.n1895 GNDA_2.n1894 3.7893
R7903 GNDA_2.n1901 GNDA_2.n1890 3.7893
R7904 GNDA_2.n1908 GNDA_2.n1889 3.7893
R7905 GNDA_2.n1909 GNDA_2.n1888 3.7893
R7906 GNDA_2.n2620 GNDA_2.n2619 3.7893
R7907 GNDA_2.n2920 GNDA_2.n2919 3.7893
R7908 GNDA_2.n2648 GNDA_2.n2621 3.7893
R7909 GNDA_2.n2651 GNDA_2.n2650 3.7893
R7910 GNDA_2.n2844 GNDA_2.n2647 3.7893
R7911 GNDA_2.n2849 GNDA_2.n2848 3.7893
R7912 GNDA_2.n2853 GNDA_2.n2852 3.7893
R7913 GNDA_2.n2861 GNDA_2.n2643 3.7893
R7914 GNDA_2.n2768 GNDA_2.n2704 3.7893
R7915 GNDA_2.n2777 GNDA_2.n2776 3.7893
R7916 GNDA_2.n2705 GNDA_2.n2684 3.7893
R7917 GNDA_2.n2786 GNDA_2.n2784 3.7893
R7918 GNDA_2.n2785 GNDA_2.n2682 3.7893
R7919 GNDA_2.n2681 GNDA_2.n2678 3.7893
R7920 GNDA_2.n2802 GNDA_2.n2800 3.7893
R7921 GNDA_2.n2801 GNDA_2.n2674 3.7893
R7922 GNDA_2.n2132 GNDA_2.n2107 3.7893
R7923 GNDA_2.n2131 GNDA_2.n2128 3.7893
R7924 GNDA_2.n2127 GNDA_2.n2108 3.7893
R7925 GNDA_2.n2124 GNDA_2.n2123 3.7893
R7926 GNDA_2.n2120 GNDA_2.n2109 3.7893
R7927 GNDA_2.n2113 GNDA_2.n2110 3.7893
R7928 GNDA_2.n2137 GNDA_2.n2028 3.7893
R7929 GNDA_2.n2138 GNDA_2.n2027 3.7893
R7930 GNDA_2.n5451 GNDA_2.n90 3.7893
R7931 GNDA_2.n5448 GNDA_2.n5447 3.7893
R7932 GNDA_2.n5364 GNDA_2.n91 3.7893
R7933 GNDA_2.n5369 GNDA_2.n5367 3.7893
R7934 GNDA_2.n5374 GNDA_2.n5370 3.7893
R7935 GNDA_2.n5381 GNDA_2.n5380 3.7893
R7936 GNDA_2.n5384 GNDA_2.n5363 3.7893
R7937 GNDA_2.n5389 GNDA_2.n5385 3.7893
R7938 GNDA_2.n2324 GNDA_2.n2145 3.7893
R7939 GNDA_2.n2321 GNDA_2.n2320 3.7893
R7940 GNDA_2.n2237 GNDA_2.n2146 3.7893
R7941 GNDA_2.n2242 GNDA_2.n2240 3.7893
R7942 GNDA_2.n2247 GNDA_2.n2243 3.7893
R7943 GNDA_2.n2254 GNDA_2.n2253 3.7893
R7944 GNDA_2.n2257 GNDA_2.n2236 3.7893
R7945 GNDA_2.n2262 GNDA_2.n2258 3.7893
R7946 GNDA_2.n3360 GNDA_2.n1725 3.7893
R7947 GNDA_2.n3359 GNDA_2.n1726 3.7893
R7948 GNDA_2.n3347 GNDA_2.n3346 3.7893
R7949 GNDA_2.n3353 GNDA_2.n3352 3.7893
R7950 GNDA_2.n3349 GNDA_2.n3348 3.7893
R7951 GNDA_2.n1701 GNDA_2.n1694 3.7893
R7952 GNDA_2.n1707 GNDA_2.n1705 3.7893
R7953 GNDA_2.n1706 GNDA_2.n1671 3.7893
R7954 GNDA_2.n5555 GNDA_2.n22 3.7893
R7955 GNDA_2.n5554 GNDA_2.n23 3.7893
R7956 GNDA_2.n33 GNDA_2.n32 3.7893
R7957 GNDA_2.n39 GNDA_2.n38 3.7893
R7958 GNDA_2.n35 GNDA_2.n34 3.7893
R7959 GNDA_2.n5287 GNDA_2.n1 3.7893
R7960 GNDA_2.n5292 GNDA_2.n5290 3.7893
R7961 GNDA_2.n5297 GNDA_2.n5293 3.7893
R7962 GNDA_2.n5469 GNDA_2 3.7381
R7963 GNDA_2.n1902 GNDA_2 3.7381
R7964 GNDA_2.n2847 GNDA_2 3.7381
R7965 GNDA_2 GNDA_2.n2792 3.7381
R7966 GNDA_2 GNDA_2.n2116 3.7381
R7967 GNDA_2.n5377 GNDA_2 3.7381
R7968 GNDA_2.n2250 GNDA_2 3.7381
R7969 GNDA_2 GNDA_2.n3365 3.7381
R7970 GNDA_2 GNDA_2.n5560 3.7381
R7971 GNDA_2.t235 GNDA_2.n4322 3.63887
R7972 GNDA_2.n4323 GNDA_2.t286 3.63887
R7973 GNDA_2.n4325 GNDA_2.t233 3.63887
R7974 GNDA_2.t183 GNDA_2.n4324 3.63887
R7975 GNDA_2.n260 GNDA_2.n259 3.50398
R7976 GNDA_2.n1589 GNDA_2.n1562 3.47871
R7977 GNDA_2.n1033 GNDA_2.n1032 3.47821
R7978 GNDA_2.n5062 GNDA_2.n5061 3.47821
R7979 GNDA_2.n4986 GNDA_2.n4985 3.47821
R7980 GNDA_2.n4856 GNDA_2.n4855 3.47821
R7981 GNDA_2.n5146 GNDA_2.n5145 3.47821
R7982 GNDA_2.n4610 GNDA_2.n4609 3.47821
R7983 GNDA_2.n5211 GNDA_2.n5210 3.47821
R7984 GNDA_2.n4771 GNDA_2.n4770 3.47821
R7985 GNDA_2.n4668 GNDA_2.n4667 3.47821
R7986 GNDA_2.n4534 GNDA_2.n4533 3.47821
R7987 GNDA_2.n4267 GNDA_2.n4266 3.47821
R7988 GNDA_2.n4263 GNDA_2.n4262 3.47821
R7989 GNDA_2.n4154 GNDA_2.n4153 3.47821
R7990 GNDA_2.n4073 GNDA_2.n4072 3.47821
R7991 GNDA_2.n1207 GNDA_2.n1206 3.47821
R7992 GNDA_2.n3680 GNDA_2.n3679 3.47821
R7993 GNDA_2.n3749 GNDA_2.n3748 3.47821
R7994 GNDA_2.n3818 GNDA_2.n3817 3.47821
R7995 GNDA_2.n3887 GNDA_2.n3886 3.47821
R7996 GNDA_2.n3952 GNDA_2.n3951 3.47821
R7997 GNDA_2.n3000 GNDA_2.n2999 3.47821
R7998 GNDA_2.n697 GNDA_2.n696 3.47821
R7999 GNDA_2.n1013 GNDA_2.n1012 3.47821
R8000 GNDA_2.n515 GNDA_2.n514 3.47821
R8001 GNDA_2.n801 GNDA_2.n800 3.47821
R8002 GNDA_2.n870 GNDA_2.n869 3.47821
R8003 GNDA_2.n935 GNDA_2.n934 3.47821
R8004 GNDA_2.n293 GNDA_2.n216 3.43627
R8005 GNDA_2.n180 GNDA_2.t186 3.42907
R8006 GNDA_2.n180 GNDA_2.t217 3.42907
R8007 GNDA_2.n4475 GNDA_2.t60 3.42907
R8008 GNDA_2.n4475 GNDA_2.t275 3.42907
R8009 GNDA_2.n1092 GNDA_2.t19 3.42907
R8010 GNDA_2.n1092 GNDA_2.t191 3.42907
R8011 GNDA_2.n4305 GNDA_2.t283 3.42907
R8012 GNDA_2.n4305 GNDA_2.t278 3.42907
R8013 GNDA_2.n1034 GNDA_2.n429 3.4105
R8014 GNDA_2.n1035 GNDA_2.n428 3.4105
R8015 GNDA_2.n1036 GNDA_2.n427 3.4105
R8016 GNDA_2.n1028 GNDA_2.n425 3.4105
R8017 GNDA_2.n1040 GNDA_2.n424 3.4105
R8018 GNDA_2.n1041 GNDA_2.n423 3.4105
R8019 GNDA_2.n1042 GNDA_2.n422 3.4105
R8020 GNDA_2.n1025 GNDA_2.n420 3.4105
R8021 GNDA_2.n1046 GNDA_2.n419 3.4105
R8022 GNDA_2.n1047 GNDA_2.n418 3.4105
R8023 GNDA_2.n1048 GNDA_2.n417 3.4105
R8024 GNDA_2.n1022 GNDA_2.n415 3.4105
R8025 GNDA_2.n1052 GNDA_2.n414 3.4105
R8026 GNDA_2.n1053 GNDA_2.n413 3.4105
R8027 GNDA_2.n1054 GNDA_2.n412 3.4105
R8028 GNDA_2.n1019 GNDA_2.n410 3.4105
R8029 GNDA_2.n1058 GNDA_2.n409 3.4105
R8030 GNDA_2.n1059 GNDA_2.n408 3.4105
R8031 GNDA_2.n1060 GNDA_2.n407 3.4105
R8032 GNDA_2.n1016 GNDA_2.n405 3.4105
R8033 GNDA_2.n1064 GNDA_2.n404 3.4105
R8034 GNDA_2.n1065 GNDA_2.n403 3.4105
R8035 GNDA_2.n1066 GNDA_2.n402 3.4105
R8036 GNDA_2.n5000 GNDA_2.n4999 3.4105
R8037 GNDA_2.n5059 GNDA_2.n5058 3.4105
R8038 GNDA_2.n5057 GNDA_2.n5056 3.4105
R8039 GNDA_2.n5055 GNDA_2.n5054 3.4105
R8040 GNDA_2.n5053 GNDA_2.n5002 3.4105
R8041 GNDA_2.n5049 GNDA_2.n5048 3.4105
R8042 GNDA_2.n5047 GNDA_2.n5046 3.4105
R8043 GNDA_2.n5045 GNDA_2.n5044 3.4105
R8044 GNDA_2.n5043 GNDA_2.n5004 3.4105
R8045 GNDA_2.n5039 GNDA_2.n5038 3.4105
R8046 GNDA_2.n5037 GNDA_2.n5036 3.4105
R8047 GNDA_2.n5035 GNDA_2.n5034 3.4105
R8048 GNDA_2.n5033 GNDA_2.n5006 3.4105
R8049 GNDA_2.n5029 GNDA_2.n5028 3.4105
R8050 GNDA_2.n5027 GNDA_2.n5026 3.4105
R8051 GNDA_2.n5025 GNDA_2.n5024 3.4105
R8052 GNDA_2.n5023 GNDA_2.n5008 3.4105
R8053 GNDA_2.n5019 GNDA_2.n5018 3.4105
R8054 GNDA_2.n5017 GNDA_2.n5016 3.4105
R8055 GNDA_2.n5015 GNDA_2.n5014 3.4105
R8056 GNDA_2.n5013 GNDA_2.n5010 3.4105
R8057 GNDA_2.n4905 GNDA_2.n4904 3.4105
R8058 GNDA_2.n5065 GNDA_2.n5064 3.4105
R8059 GNDA_2.n4919 GNDA_2.n4918 3.4105
R8060 GNDA_2.n4983 GNDA_2.n4982 3.4105
R8061 GNDA_2.n4981 GNDA_2.n4980 3.4105
R8062 GNDA_2.n4979 GNDA_2.n4978 3.4105
R8063 GNDA_2.n4977 GNDA_2.n4921 3.4105
R8064 GNDA_2.n4973 GNDA_2.n4972 3.4105
R8065 GNDA_2.n4971 GNDA_2.n4970 3.4105
R8066 GNDA_2.n4969 GNDA_2.n4968 3.4105
R8067 GNDA_2.n4967 GNDA_2.n4923 3.4105
R8068 GNDA_2.n4963 GNDA_2.n4962 3.4105
R8069 GNDA_2.n4961 GNDA_2.n4960 3.4105
R8070 GNDA_2.n4959 GNDA_2.n4958 3.4105
R8071 GNDA_2.n4957 GNDA_2.n4925 3.4105
R8072 GNDA_2.n4953 GNDA_2.n4952 3.4105
R8073 GNDA_2.n4951 GNDA_2.n4950 3.4105
R8074 GNDA_2.n4949 GNDA_2.n4948 3.4105
R8075 GNDA_2.n4947 GNDA_2.n4927 3.4105
R8076 GNDA_2.n4943 GNDA_2.n4942 3.4105
R8077 GNDA_2.n4941 GNDA_2.n4940 3.4105
R8078 GNDA_2.n4939 GNDA_2.n4938 3.4105
R8079 GNDA_2.n4937 GNDA_2.n4929 3.4105
R8080 GNDA_2.n4933 GNDA_2.n4932 3.4105
R8081 GNDA_2.n4931 GNDA_2.n4906 3.4105
R8082 GNDA_2.n4857 GNDA_2.n4834 3.4105
R8083 GNDA_2.n4859 GNDA_2.n4833 3.4105
R8084 GNDA_2.n4860 GNDA_2.n4832 3.4105
R8085 GNDA_2.n4862 GNDA_2.n4831 3.4105
R8086 GNDA_2.n4863 GNDA_2.n4830 3.4105
R8087 GNDA_2.n4865 GNDA_2.n4829 3.4105
R8088 GNDA_2.n4866 GNDA_2.n4828 3.4105
R8089 GNDA_2.n4868 GNDA_2.n4827 3.4105
R8090 GNDA_2.n4869 GNDA_2.n4826 3.4105
R8091 GNDA_2.n4871 GNDA_2.n4825 3.4105
R8092 GNDA_2.n4872 GNDA_2.n4824 3.4105
R8093 GNDA_2.n4874 GNDA_2.n4823 3.4105
R8094 GNDA_2.n4875 GNDA_2.n4822 3.4105
R8095 GNDA_2.n4877 GNDA_2.n4821 3.4105
R8096 GNDA_2.n4878 GNDA_2.n4820 3.4105
R8097 GNDA_2.n4880 GNDA_2.n4819 3.4105
R8098 GNDA_2.n4881 GNDA_2.n4818 3.4105
R8099 GNDA_2.n4883 GNDA_2.n4817 3.4105
R8100 GNDA_2.n4884 GNDA_2.n4816 3.4105
R8101 GNDA_2.n4886 GNDA_2.n4815 3.4105
R8102 GNDA_2.n4887 GNDA_2.n4814 3.4105
R8103 GNDA_2.n4889 GNDA_2.n4813 3.4105
R8104 GNDA_2.n4891 GNDA_2.n4890 3.4105
R8105 GNDA_2.n4798 GNDA_2.n4797 3.4105
R8106 GNDA_2.n5143 GNDA_2.n5142 3.4105
R8107 GNDA_2.n5141 GNDA_2.n5140 3.4105
R8108 GNDA_2.n5139 GNDA_2.n5138 3.4105
R8109 GNDA_2.n5137 GNDA_2.n4800 3.4105
R8110 GNDA_2.n5133 GNDA_2.n5132 3.4105
R8111 GNDA_2.n5131 GNDA_2.n5130 3.4105
R8112 GNDA_2.n5129 GNDA_2.n5128 3.4105
R8113 GNDA_2.n5127 GNDA_2.n4802 3.4105
R8114 GNDA_2.n5123 GNDA_2.n5122 3.4105
R8115 GNDA_2.n5121 GNDA_2.n5120 3.4105
R8116 GNDA_2.n5119 GNDA_2.n5118 3.4105
R8117 GNDA_2.n5117 GNDA_2.n4804 3.4105
R8118 GNDA_2.n5113 GNDA_2.n5112 3.4105
R8119 GNDA_2.n5111 GNDA_2.n5110 3.4105
R8120 GNDA_2.n5109 GNDA_2.n5108 3.4105
R8121 GNDA_2.n5107 GNDA_2.n4806 3.4105
R8122 GNDA_2.n5103 GNDA_2.n5102 3.4105
R8123 GNDA_2.n5101 GNDA_2.n5100 3.4105
R8124 GNDA_2.n5099 GNDA_2.n5098 3.4105
R8125 GNDA_2.n5097 GNDA_2.n4808 3.4105
R8126 GNDA_2.n5093 GNDA_2.n5092 3.4105
R8127 GNDA_2.n5091 GNDA_2.n4784 3.4105
R8128 GNDA_2.n4548 GNDA_2.n4547 3.4105
R8129 GNDA_2.n4607 GNDA_2.n4606 3.4105
R8130 GNDA_2.n4605 GNDA_2.n4604 3.4105
R8131 GNDA_2.n4603 GNDA_2.n4602 3.4105
R8132 GNDA_2.n4601 GNDA_2.n4550 3.4105
R8133 GNDA_2.n4597 GNDA_2.n4596 3.4105
R8134 GNDA_2.n4595 GNDA_2.n4594 3.4105
R8135 GNDA_2.n4593 GNDA_2.n4592 3.4105
R8136 GNDA_2.n4591 GNDA_2.n4552 3.4105
R8137 GNDA_2.n4587 GNDA_2.n4586 3.4105
R8138 GNDA_2.n4585 GNDA_2.n4584 3.4105
R8139 GNDA_2.n4583 GNDA_2.n4582 3.4105
R8140 GNDA_2.n4581 GNDA_2.n4554 3.4105
R8141 GNDA_2.n4577 GNDA_2.n4576 3.4105
R8142 GNDA_2.n4575 GNDA_2.n4574 3.4105
R8143 GNDA_2.n4573 GNDA_2.n4572 3.4105
R8144 GNDA_2.n4571 GNDA_2.n4556 3.4105
R8145 GNDA_2.n4567 GNDA_2.n4566 3.4105
R8146 GNDA_2.n4565 GNDA_2.n4564 3.4105
R8147 GNDA_2.n4563 GNDA_2.n4562 3.4105
R8148 GNDA_2.n4561 GNDA_2.n4558 3.4105
R8149 GNDA_2.n186 GNDA_2.n185 3.4105
R8150 GNDA_2.n4613 GNDA_2.n4612 3.4105
R8151 GNDA_2.n5149 GNDA_2.n5148 3.4105
R8152 GNDA_2.n5208 GNDA_2.n5207 3.4105
R8153 GNDA_2.n5206 GNDA_2.n5205 3.4105
R8154 GNDA_2.n5204 GNDA_2.n5203 3.4105
R8155 GNDA_2.n5202 GNDA_2.n5151 3.4105
R8156 GNDA_2.n5198 GNDA_2.n5197 3.4105
R8157 GNDA_2.n5196 GNDA_2.n5195 3.4105
R8158 GNDA_2.n5194 GNDA_2.n5193 3.4105
R8159 GNDA_2.n5192 GNDA_2.n5153 3.4105
R8160 GNDA_2.n5188 GNDA_2.n5187 3.4105
R8161 GNDA_2.n5186 GNDA_2.n5185 3.4105
R8162 GNDA_2.n5184 GNDA_2.n5183 3.4105
R8163 GNDA_2.n5182 GNDA_2.n5155 3.4105
R8164 GNDA_2.n5178 GNDA_2.n5177 3.4105
R8165 GNDA_2.n5176 GNDA_2.n5175 3.4105
R8166 GNDA_2.n5174 GNDA_2.n5173 3.4105
R8167 GNDA_2.n5172 GNDA_2.n5157 3.4105
R8168 GNDA_2.n5168 GNDA_2.n5167 3.4105
R8169 GNDA_2.n5166 GNDA_2.n5165 3.4105
R8170 GNDA_2.n5164 GNDA_2.n5163 3.4105
R8171 GNDA_2.n5162 GNDA_2.n5159 3.4105
R8172 GNDA_2.n146 GNDA_2.n145 3.4105
R8173 GNDA_2.n5214 GNDA_2.n5213 3.4105
R8174 GNDA_2.n161 GNDA_2.n160 3.4105
R8175 GNDA_2.n4768 GNDA_2.n4767 3.4105
R8176 GNDA_2.n4766 GNDA_2.n4765 3.4105
R8177 GNDA_2.n4764 GNDA_2.n4763 3.4105
R8178 GNDA_2.n4762 GNDA_2.n163 3.4105
R8179 GNDA_2.n4758 GNDA_2.n4757 3.4105
R8180 GNDA_2.n4756 GNDA_2.n4755 3.4105
R8181 GNDA_2.n4754 GNDA_2.n4753 3.4105
R8182 GNDA_2.n4752 GNDA_2.n165 3.4105
R8183 GNDA_2.n4748 GNDA_2.n4747 3.4105
R8184 GNDA_2.n4746 GNDA_2.n4745 3.4105
R8185 GNDA_2.n4744 GNDA_2.n4743 3.4105
R8186 GNDA_2.n4742 GNDA_2.n167 3.4105
R8187 GNDA_2.n4738 GNDA_2.n4737 3.4105
R8188 GNDA_2.n4736 GNDA_2.n4735 3.4105
R8189 GNDA_2.n4734 GNDA_2.n4733 3.4105
R8190 GNDA_2.n4732 GNDA_2.n169 3.4105
R8191 GNDA_2.n4728 GNDA_2.n4727 3.4105
R8192 GNDA_2.n4726 GNDA_2.n4725 3.4105
R8193 GNDA_2.n4724 GNDA_2.n4723 3.4105
R8194 GNDA_2.n4722 GNDA_2.n171 3.4105
R8195 GNDA_2.n4718 GNDA_2.n4717 3.4105
R8196 GNDA_2.n4716 GNDA_2.n148 3.4105
R8197 GNDA_2.n4669 GNDA_2.n4646 3.4105
R8198 GNDA_2.n4671 GNDA_2.n4645 3.4105
R8199 GNDA_2.n4672 GNDA_2.n4644 3.4105
R8200 GNDA_2.n4674 GNDA_2.n4643 3.4105
R8201 GNDA_2.n4675 GNDA_2.n4642 3.4105
R8202 GNDA_2.n4677 GNDA_2.n4641 3.4105
R8203 GNDA_2.n4678 GNDA_2.n4640 3.4105
R8204 GNDA_2.n4680 GNDA_2.n4639 3.4105
R8205 GNDA_2.n4681 GNDA_2.n4638 3.4105
R8206 GNDA_2.n4683 GNDA_2.n4637 3.4105
R8207 GNDA_2.n4684 GNDA_2.n4636 3.4105
R8208 GNDA_2.n4686 GNDA_2.n4635 3.4105
R8209 GNDA_2.n4687 GNDA_2.n4634 3.4105
R8210 GNDA_2.n4689 GNDA_2.n4633 3.4105
R8211 GNDA_2.n4690 GNDA_2.n4632 3.4105
R8212 GNDA_2.n4692 GNDA_2.n4631 3.4105
R8213 GNDA_2.n4693 GNDA_2.n4630 3.4105
R8214 GNDA_2.n4695 GNDA_2.n4629 3.4105
R8215 GNDA_2.n4696 GNDA_2.n4628 3.4105
R8216 GNDA_2.n4698 GNDA_2.n4627 3.4105
R8217 GNDA_2.n4699 GNDA_2.n4626 3.4105
R8218 GNDA_2.n4701 GNDA_2.n4625 3.4105
R8219 GNDA_2.n4703 GNDA_2.n4702 3.4105
R8220 GNDA_2.n201 GNDA_2.n200 3.4105
R8221 GNDA_2.n4531 GNDA_2.n4530 3.4105
R8222 GNDA_2.n4529 GNDA_2.n4528 3.4105
R8223 GNDA_2.n4527 GNDA_2.n4526 3.4105
R8224 GNDA_2.n4525 GNDA_2.n203 3.4105
R8225 GNDA_2.n4521 GNDA_2.n4520 3.4105
R8226 GNDA_2.n4519 GNDA_2.n4518 3.4105
R8227 GNDA_2.n4517 GNDA_2.n4516 3.4105
R8228 GNDA_2.n4515 GNDA_2.n205 3.4105
R8229 GNDA_2.n4511 GNDA_2.n4510 3.4105
R8230 GNDA_2.n4509 GNDA_2.n4508 3.4105
R8231 GNDA_2.n4507 GNDA_2.n4506 3.4105
R8232 GNDA_2.n4505 GNDA_2.n207 3.4105
R8233 GNDA_2.n4501 GNDA_2.n4500 3.4105
R8234 GNDA_2.n4499 GNDA_2.n4498 3.4105
R8235 GNDA_2.n4497 GNDA_2.n4496 3.4105
R8236 GNDA_2.n4495 GNDA_2.n209 3.4105
R8237 GNDA_2.n4491 GNDA_2.n4490 3.4105
R8238 GNDA_2.n4489 GNDA_2.n4488 3.4105
R8239 GNDA_2.n4487 GNDA_2.n4486 3.4105
R8240 GNDA_2.n4485 GNDA_2.n211 3.4105
R8241 GNDA_2.n4481 GNDA_2.n4480 3.4105
R8242 GNDA_2.n4479 GNDA_2.n188 3.4105
R8243 GNDA_2.n4268 GNDA_2.n1121 3.4105
R8244 GNDA_2.n4269 GNDA_2.n1120 3.4105
R8245 GNDA_2.n4270 GNDA_2.n1119 3.4105
R8246 GNDA_2.n4169 GNDA_2.n1117 3.4105
R8247 GNDA_2.n4274 GNDA_2.n1116 3.4105
R8248 GNDA_2.n4275 GNDA_2.n1115 3.4105
R8249 GNDA_2.n4276 GNDA_2.n1114 3.4105
R8250 GNDA_2.n4166 GNDA_2.n1112 3.4105
R8251 GNDA_2.n4280 GNDA_2.n1111 3.4105
R8252 GNDA_2.n4281 GNDA_2.n1110 3.4105
R8253 GNDA_2.n4282 GNDA_2.n1109 3.4105
R8254 GNDA_2.n4163 GNDA_2.n1107 3.4105
R8255 GNDA_2.n4286 GNDA_2.n1106 3.4105
R8256 GNDA_2.n4287 GNDA_2.n1105 3.4105
R8257 GNDA_2.n4288 GNDA_2.n1104 3.4105
R8258 GNDA_2.n4160 GNDA_2.n1102 3.4105
R8259 GNDA_2.n4292 GNDA_2.n1101 3.4105
R8260 GNDA_2.n4293 GNDA_2.n1100 3.4105
R8261 GNDA_2.n4294 GNDA_2.n1099 3.4105
R8262 GNDA_2.n4157 GNDA_2.n1097 3.4105
R8263 GNDA_2.n4298 GNDA_2.n1096 3.4105
R8264 GNDA_2.n4299 GNDA_2.n1095 3.4105
R8265 GNDA_2.n4300 GNDA_2.n1094 3.4105
R8266 GNDA_2.n4185 GNDA_2.n4184 3.4105
R8267 GNDA_2.n4260 GNDA_2.n4259 3.4105
R8268 GNDA_2.n4258 GNDA_2.n4257 3.4105
R8269 GNDA_2.n4256 GNDA_2.n4189 3.4105
R8270 GNDA_2.n4188 GNDA_2.n4187 3.4105
R8271 GNDA_2.n4252 GNDA_2.n4251 3.4105
R8272 GNDA_2.n4250 GNDA_2.n4249 3.4105
R8273 GNDA_2.n4248 GNDA_2.n4193 3.4105
R8274 GNDA_2.n4192 GNDA_2.n4191 3.4105
R8275 GNDA_2.n4244 GNDA_2.n4243 3.4105
R8276 GNDA_2.n4242 GNDA_2.n4241 3.4105
R8277 GNDA_2.n4240 GNDA_2.n4197 3.4105
R8278 GNDA_2.n4196 GNDA_2.n4195 3.4105
R8279 GNDA_2.n4236 GNDA_2.n4235 3.4105
R8280 GNDA_2.n4234 GNDA_2.n4233 3.4105
R8281 GNDA_2.n4232 GNDA_2.n4201 3.4105
R8282 GNDA_2.n4200 GNDA_2.n4199 3.4105
R8283 GNDA_2.n4228 GNDA_2.n4227 3.4105
R8284 GNDA_2.n4226 GNDA_2.n4225 3.4105
R8285 GNDA_2.n4224 GNDA_2.n4205 3.4105
R8286 GNDA_2.n4204 GNDA_2.n4203 3.4105
R8287 GNDA_2.n4220 GNDA_2.n4219 3.4105
R8288 GNDA_2.n4218 GNDA_2.n4172 3.4105
R8289 GNDA_2.n4088 GNDA_2.n4087 3.4105
R8290 GNDA_2.n4151 GNDA_2.n4150 3.4105
R8291 GNDA_2.n4149 GNDA_2.n4148 3.4105
R8292 GNDA_2.n4147 GNDA_2.n4092 3.4105
R8293 GNDA_2.n4091 GNDA_2.n4090 3.4105
R8294 GNDA_2.n4143 GNDA_2.n4142 3.4105
R8295 GNDA_2.n4141 GNDA_2.n4140 3.4105
R8296 GNDA_2.n4139 GNDA_2.n4096 3.4105
R8297 GNDA_2.n4095 GNDA_2.n4094 3.4105
R8298 GNDA_2.n4135 GNDA_2.n4134 3.4105
R8299 GNDA_2.n4133 GNDA_2.n4132 3.4105
R8300 GNDA_2.n4131 GNDA_2.n4100 3.4105
R8301 GNDA_2.n4099 GNDA_2.n4098 3.4105
R8302 GNDA_2.n4127 GNDA_2.n4126 3.4105
R8303 GNDA_2.n4125 GNDA_2.n4124 3.4105
R8304 GNDA_2.n4123 GNDA_2.n4104 3.4105
R8305 GNDA_2.n4103 GNDA_2.n4102 3.4105
R8306 GNDA_2.n4119 GNDA_2.n4118 3.4105
R8307 GNDA_2.n4117 GNDA_2.n4116 3.4105
R8308 GNDA_2.n4115 GNDA_2.n4108 3.4105
R8309 GNDA_2.n4107 GNDA_2.n4106 3.4105
R8310 GNDA_2.n4111 GNDA_2.n4110 3.4105
R8311 GNDA_2.n4109 GNDA_2.n4075 3.4105
R8312 GNDA_2.n1136 GNDA_2.n1135 3.4105
R8313 GNDA_2.n4070 GNDA_2.n4069 3.4105
R8314 GNDA_2.n4068 GNDA_2.n4067 3.4105
R8315 GNDA_2.n4066 GNDA_2.n1140 3.4105
R8316 GNDA_2.n1139 GNDA_2.n1138 3.4105
R8317 GNDA_2.n4062 GNDA_2.n4061 3.4105
R8318 GNDA_2.n4060 GNDA_2.n4059 3.4105
R8319 GNDA_2.n4058 GNDA_2.n1144 3.4105
R8320 GNDA_2.n1143 GNDA_2.n1142 3.4105
R8321 GNDA_2.n4054 GNDA_2.n4053 3.4105
R8322 GNDA_2.n4052 GNDA_2.n4051 3.4105
R8323 GNDA_2.n4050 GNDA_2.n1148 3.4105
R8324 GNDA_2.n1147 GNDA_2.n1146 3.4105
R8325 GNDA_2.n4046 GNDA_2.n4045 3.4105
R8326 GNDA_2.n4044 GNDA_2.n4043 3.4105
R8327 GNDA_2.n4042 GNDA_2.n1152 3.4105
R8328 GNDA_2.n1151 GNDA_2.n1150 3.4105
R8329 GNDA_2.n4038 GNDA_2.n4037 3.4105
R8330 GNDA_2.n4036 GNDA_2.n4035 3.4105
R8331 GNDA_2.n4034 GNDA_2.n1156 3.4105
R8332 GNDA_2.n1155 GNDA_2.n1154 3.4105
R8333 GNDA_2.n4030 GNDA_2.n4029 3.4105
R8334 GNDA_2.n4028 GNDA_2.n1123 3.4105
R8335 GNDA_2.n1208 GNDA_2.n1205 3.4105
R8336 GNDA_2.n1209 GNDA_2.n1203 3.4105
R8337 GNDA_2.n1210 GNDA_2.n1202 3.4105
R8338 GNDA_2.n1200 GNDA_2.n1198 3.4105
R8339 GNDA_2.n1214 GNDA_2.n1197 3.4105
R8340 GNDA_2.n1215 GNDA_2.n1195 3.4105
R8341 GNDA_2.n1216 GNDA_2.n1194 3.4105
R8342 GNDA_2.n1192 GNDA_2.n1190 3.4105
R8343 GNDA_2.n1220 GNDA_2.n1189 3.4105
R8344 GNDA_2.n1221 GNDA_2.n1187 3.4105
R8345 GNDA_2.n1222 GNDA_2.n1186 3.4105
R8346 GNDA_2.n1184 GNDA_2.n1182 3.4105
R8347 GNDA_2.n1226 GNDA_2.n1181 3.4105
R8348 GNDA_2.n1227 GNDA_2.n1179 3.4105
R8349 GNDA_2.n1228 GNDA_2.n1178 3.4105
R8350 GNDA_2.n1176 GNDA_2.n1174 3.4105
R8351 GNDA_2.n1232 GNDA_2.n1173 3.4105
R8352 GNDA_2.n1233 GNDA_2.n1171 3.4105
R8353 GNDA_2.n1234 GNDA_2.n1170 3.4105
R8354 GNDA_2.n1168 GNDA_2.n1166 3.4105
R8355 GNDA_2.n1238 GNDA_2.n1165 3.4105
R8356 GNDA_2.n1239 GNDA_2.n1163 3.4105
R8357 GNDA_2.n1240 GNDA_2.n1162 3.4105
R8358 GNDA_2.n3614 GNDA_2.n3613 3.4105
R8359 GNDA_2.n3677 GNDA_2.n3676 3.4105
R8360 GNDA_2.n3675 GNDA_2.n3674 3.4105
R8361 GNDA_2.n3673 GNDA_2.n3618 3.4105
R8362 GNDA_2.n3617 GNDA_2.n3616 3.4105
R8363 GNDA_2.n3669 GNDA_2.n3668 3.4105
R8364 GNDA_2.n3667 GNDA_2.n3666 3.4105
R8365 GNDA_2.n3665 GNDA_2.n3622 3.4105
R8366 GNDA_2.n3621 GNDA_2.n3620 3.4105
R8367 GNDA_2.n3661 GNDA_2.n3660 3.4105
R8368 GNDA_2.n3659 GNDA_2.n3658 3.4105
R8369 GNDA_2.n3657 GNDA_2.n3626 3.4105
R8370 GNDA_2.n3625 GNDA_2.n3624 3.4105
R8371 GNDA_2.n3653 GNDA_2.n3652 3.4105
R8372 GNDA_2.n3651 GNDA_2.n3650 3.4105
R8373 GNDA_2.n3649 GNDA_2.n3630 3.4105
R8374 GNDA_2.n3629 GNDA_2.n3628 3.4105
R8375 GNDA_2.n3645 GNDA_2.n3644 3.4105
R8376 GNDA_2.n3643 GNDA_2.n3642 3.4105
R8377 GNDA_2.n3641 GNDA_2.n3634 3.4105
R8378 GNDA_2.n3633 GNDA_2.n3632 3.4105
R8379 GNDA_2.n3637 GNDA_2.n3636 3.4105
R8380 GNDA_2.n3635 GNDA_2.n3601 3.4105
R8381 GNDA_2.n3683 GNDA_2.n3682 3.4105
R8382 GNDA_2.n3746 GNDA_2.n3745 3.4105
R8383 GNDA_2.n3744 GNDA_2.n3743 3.4105
R8384 GNDA_2.n3742 GNDA_2.n3687 3.4105
R8385 GNDA_2.n3686 GNDA_2.n3685 3.4105
R8386 GNDA_2.n3738 GNDA_2.n3737 3.4105
R8387 GNDA_2.n3736 GNDA_2.n3735 3.4105
R8388 GNDA_2.n3734 GNDA_2.n3691 3.4105
R8389 GNDA_2.n3690 GNDA_2.n3689 3.4105
R8390 GNDA_2.n3730 GNDA_2.n3729 3.4105
R8391 GNDA_2.n3728 GNDA_2.n3727 3.4105
R8392 GNDA_2.n3726 GNDA_2.n3695 3.4105
R8393 GNDA_2.n3694 GNDA_2.n3693 3.4105
R8394 GNDA_2.n3722 GNDA_2.n3721 3.4105
R8395 GNDA_2.n3720 GNDA_2.n3719 3.4105
R8396 GNDA_2.n3718 GNDA_2.n3699 3.4105
R8397 GNDA_2.n3698 GNDA_2.n3697 3.4105
R8398 GNDA_2.n3714 GNDA_2.n3713 3.4105
R8399 GNDA_2.n3712 GNDA_2.n3711 3.4105
R8400 GNDA_2.n3710 GNDA_2.n3703 3.4105
R8401 GNDA_2.n3702 GNDA_2.n3701 3.4105
R8402 GNDA_2.n3706 GNDA_2.n3705 3.4105
R8403 GNDA_2.n3704 GNDA_2.n3589 3.4105
R8404 GNDA_2.n3752 GNDA_2.n3751 3.4105
R8405 GNDA_2.n3815 GNDA_2.n3814 3.4105
R8406 GNDA_2.n3813 GNDA_2.n3812 3.4105
R8407 GNDA_2.n3811 GNDA_2.n3756 3.4105
R8408 GNDA_2.n3755 GNDA_2.n3754 3.4105
R8409 GNDA_2.n3807 GNDA_2.n3806 3.4105
R8410 GNDA_2.n3805 GNDA_2.n3804 3.4105
R8411 GNDA_2.n3803 GNDA_2.n3760 3.4105
R8412 GNDA_2.n3759 GNDA_2.n3758 3.4105
R8413 GNDA_2.n3799 GNDA_2.n3798 3.4105
R8414 GNDA_2.n3797 GNDA_2.n3796 3.4105
R8415 GNDA_2.n3795 GNDA_2.n3764 3.4105
R8416 GNDA_2.n3763 GNDA_2.n3762 3.4105
R8417 GNDA_2.n3791 GNDA_2.n3790 3.4105
R8418 GNDA_2.n3789 GNDA_2.n3788 3.4105
R8419 GNDA_2.n3787 GNDA_2.n3768 3.4105
R8420 GNDA_2.n3767 GNDA_2.n3766 3.4105
R8421 GNDA_2.n3783 GNDA_2.n3782 3.4105
R8422 GNDA_2.n3781 GNDA_2.n3780 3.4105
R8423 GNDA_2.n3779 GNDA_2.n3772 3.4105
R8424 GNDA_2.n3771 GNDA_2.n3770 3.4105
R8425 GNDA_2.n3775 GNDA_2.n3774 3.4105
R8426 GNDA_2.n3773 GNDA_2.n3577 3.4105
R8427 GNDA_2.n3821 GNDA_2.n3820 3.4105
R8428 GNDA_2.n3884 GNDA_2.n3883 3.4105
R8429 GNDA_2.n3882 GNDA_2.n3881 3.4105
R8430 GNDA_2.n3880 GNDA_2.n3825 3.4105
R8431 GNDA_2.n3824 GNDA_2.n3823 3.4105
R8432 GNDA_2.n3876 GNDA_2.n3875 3.4105
R8433 GNDA_2.n3874 GNDA_2.n3873 3.4105
R8434 GNDA_2.n3872 GNDA_2.n3829 3.4105
R8435 GNDA_2.n3828 GNDA_2.n3827 3.4105
R8436 GNDA_2.n3868 GNDA_2.n3867 3.4105
R8437 GNDA_2.n3866 GNDA_2.n3865 3.4105
R8438 GNDA_2.n3864 GNDA_2.n3833 3.4105
R8439 GNDA_2.n3832 GNDA_2.n3831 3.4105
R8440 GNDA_2.n3860 GNDA_2.n3859 3.4105
R8441 GNDA_2.n3858 GNDA_2.n3857 3.4105
R8442 GNDA_2.n3856 GNDA_2.n3837 3.4105
R8443 GNDA_2.n3836 GNDA_2.n3835 3.4105
R8444 GNDA_2.n3852 GNDA_2.n3851 3.4105
R8445 GNDA_2.n3850 GNDA_2.n3849 3.4105
R8446 GNDA_2.n3848 GNDA_2.n3841 3.4105
R8447 GNDA_2.n3840 GNDA_2.n3839 3.4105
R8448 GNDA_2.n3844 GNDA_2.n3843 3.4105
R8449 GNDA_2.n3842 GNDA_2.n3565 3.4105
R8450 GNDA_2.n3890 GNDA_2.n3889 3.4105
R8451 GNDA_2.n3949 GNDA_2.n3948 3.4105
R8452 GNDA_2.n3947 GNDA_2.n3946 3.4105
R8453 GNDA_2.n3945 GNDA_2.n3944 3.4105
R8454 GNDA_2.n3943 GNDA_2.n3892 3.4105
R8455 GNDA_2.n3939 GNDA_2.n3938 3.4105
R8456 GNDA_2.n3937 GNDA_2.n3936 3.4105
R8457 GNDA_2.n3935 GNDA_2.n3934 3.4105
R8458 GNDA_2.n3933 GNDA_2.n3894 3.4105
R8459 GNDA_2.n3929 GNDA_2.n3928 3.4105
R8460 GNDA_2.n3927 GNDA_2.n3926 3.4105
R8461 GNDA_2.n3925 GNDA_2.n3924 3.4105
R8462 GNDA_2.n3923 GNDA_2.n3896 3.4105
R8463 GNDA_2.n3919 GNDA_2.n3918 3.4105
R8464 GNDA_2.n3917 GNDA_2.n3916 3.4105
R8465 GNDA_2.n3915 GNDA_2.n3914 3.4105
R8466 GNDA_2.n3913 GNDA_2.n3898 3.4105
R8467 GNDA_2.n3909 GNDA_2.n3908 3.4105
R8468 GNDA_2.n3907 GNDA_2.n3906 3.4105
R8469 GNDA_2.n3905 GNDA_2.n3904 3.4105
R8470 GNDA_2.n3903 GNDA_2.n3900 3.4105
R8471 GNDA_2.n1266 GNDA_2.n1265 3.4105
R8472 GNDA_2.n3955 GNDA_2.n3954 3.4105
R8473 GNDA_2.n3054 GNDA_2.n2978 3.4105
R8474 GNDA_2.n3052 GNDA_2.n3051 3.4105
R8475 GNDA_2.n2980 GNDA_2.n2979 3.4105
R8476 GNDA_2.n3047 GNDA_2.n3046 3.4105
R8477 GNDA_2.n3044 GNDA_2.n2982 3.4105
R8478 GNDA_2.n3042 GNDA_2.n3041 3.4105
R8479 GNDA_2.n2984 GNDA_2.n2983 3.4105
R8480 GNDA_2.n3037 GNDA_2.n3036 3.4105
R8481 GNDA_2.n3034 GNDA_2.n2986 3.4105
R8482 GNDA_2.n3032 GNDA_2.n3031 3.4105
R8483 GNDA_2.n2988 GNDA_2.n2987 3.4105
R8484 GNDA_2.n3027 GNDA_2.n3026 3.4105
R8485 GNDA_2.n3024 GNDA_2.n2990 3.4105
R8486 GNDA_2.n3022 GNDA_2.n3021 3.4105
R8487 GNDA_2.n2992 GNDA_2.n2991 3.4105
R8488 GNDA_2.n3017 GNDA_2.n3016 3.4105
R8489 GNDA_2.n3014 GNDA_2.n2994 3.4105
R8490 GNDA_2.n3012 GNDA_2.n3011 3.4105
R8491 GNDA_2.n2996 GNDA_2.n2995 3.4105
R8492 GNDA_2.n3007 GNDA_2.n3006 3.4105
R8493 GNDA_2.n3004 GNDA_2.n2998 3.4105
R8494 GNDA_2.n3002 GNDA_2.n3001 3.4105
R8495 GNDA_2.n3056 GNDA_2.n3055 3.4105
R8496 GNDA_2.n1576 GNDA_2.n1575 3.4105
R8497 GNDA_2.n1638 GNDA_2.n1637 3.4105
R8498 GNDA_2.n1636 GNDA_2.n1635 3.4105
R8499 GNDA_2.n1634 GNDA_2.n1633 3.4105
R8500 GNDA_2.n1632 GNDA_2.n1578 3.4105
R8501 GNDA_2.n1628 GNDA_2.n1627 3.4105
R8502 GNDA_2.n1626 GNDA_2.n1625 3.4105
R8503 GNDA_2.n1624 GNDA_2.n1623 3.4105
R8504 GNDA_2.n1622 GNDA_2.n1580 3.4105
R8505 GNDA_2.n1618 GNDA_2.n1617 3.4105
R8506 GNDA_2.n1616 GNDA_2.n1615 3.4105
R8507 GNDA_2.n1614 GNDA_2.n1613 3.4105
R8508 GNDA_2.n1612 GNDA_2.n1582 3.4105
R8509 GNDA_2.n1608 GNDA_2.n1607 3.4105
R8510 GNDA_2.n1606 GNDA_2.n1605 3.4105
R8511 GNDA_2.n1604 GNDA_2.n1603 3.4105
R8512 GNDA_2.n1602 GNDA_2.n1584 3.4105
R8513 GNDA_2.n1598 GNDA_2.n1597 3.4105
R8514 GNDA_2.n1596 GNDA_2.n1595 3.4105
R8515 GNDA_2.n1594 GNDA_2.n1593 3.4105
R8516 GNDA_2.n1592 GNDA_2.n1586 3.4105
R8517 GNDA_2.n1588 GNDA_2.n1587 3.4105
R8518 GNDA_2.n3436 GNDA_2.n3435 3.4105
R8519 GNDA_2.n3437 GNDA_2.n1562 3.4105
R8520 GNDA_2.n3437 GNDA_2.n3436 3.4105
R8521 GNDA_2.n2999 GNDA_2.n1574 3.4105
R8522 GNDA_2.n3055 GNDA_2.n1574 3.4105
R8523 GNDA_2.n1545 GNDA_2.n1512 3.4105
R8524 GNDA_2.n3441 GNDA_2.n1512 3.4105
R8525 GNDA_2.n3441 GNDA_2.n1494 3.4105
R8526 GNDA_2.n1545 GNDA_2.n1514 3.4105
R8527 GNDA_2.n1514 GNDA_2.n1447 3.4105
R8528 GNDA_2.n1514 GNDA_2.n1445 3.4105
R8529 GNDA_2.n1514 GNDA_2.n1448 3.4105
R8530 GNDA_2.n1514 GNDA_2.n1444 3.4105
R8531 GNDA_2.n1514 GNDA_2.n1449 3.4105
R8532 GNDA_2.n1514 GNDA_2.n1443 3.4105
R8533 GNDA_2.n1514 GNDA_2.n1450 3.4105
R8534 GNDA_2.n1514 GNDA_2.n1442 3.4105
R8535 GNDA_2.n1514 GNDA_2.n1451 3.4105
R8536 GNDA_2.n1514 GNDA_2.n1441 3.4105
R8537 GNDA_2.n1514 GNDA_2.n1452 3.4105
R8538 GNDA_2.n1514 GNDA_2.n1440 3.4105
R8539 GNDA_2.n1514 GNDA_2.n1453 3.4105
R8540 GNDA_2.n1514 GNDA_2.n1439 3.4105
R8541 GNDA_2.n1514 GNDA_2.n1454 3.4105
R8542 GNDA_2.n1514 GNDA_2.n1438 3.4105
R8543 GNDA_2.n1514 GNDA_2.n1455 3.4105
R8544 GNDA_2.n1514 GNDA_2.n1437 3.4105
R8545 GNDA_2.n1514 GNDA_2.n1456 3.4105
R8546 GNDA_2.n1514 GNDA_2.n1436 3.4105
R8547 GNDA_2.n1514 GNDA_2.n1457 3.4105
R8548 GNDA_2.n1514 GNDA_2.n1435 3.4105
R8549 GNDA_2.n1514 GNDA_2.n1458 3.4105
R8550 GNDA_2.n1514 GNDA_2.n1434 3.4105
R8551 GNDA_2.n1514 GNDA_2.n1459 3.4105
R8552 GNDA_2.n1514 GNDA_2.n1433 3.4105
R8553 GNDA_2.n1514 GNDA_2.n1460 3.4105
R8554 GNDA_2.n1514 GNDA_2.n1432 3.4105
R8555 GNDA_2.n1514 GNDA_2.n1461 3.4105
R8556 GNDA_2.n1514 GNDA_2.n1431 3.4105
R8557 GNDA_2.n1514 GNDA_2.n1462 3.4105
R8558 GNDA_2.n3441 GNDA_2.n1514 3.4105
R8559 GNDA_2.n1545 GNDA_2.n1478 3.4105
R8560 GNDA_2.n1478 GNDA_2.n1447 3.4105
R8561 GNDA_2.n1478 GNDA_2.n1445 3.4105
R8562 GNDA_2.n1478 GNDA_2.n1448 3.4105
R8563 GNDA_2.n1478 GNDA_2.n1444 3.4105
R8564 GNDA_2.n1478 GNDA_2.n1449 3.4105
R8565 GNDA_2.n1478 GNDA_2.n1443 3.4105
R8566 GNDA_2.n1478 GNDA_2.n1450 3.4105
R8567 GNDA_2.n1478 GNDA_2.n1442 3.4105
R8568 GNDA_2.n1478 GNDA_2.n1451 3.4105
R8569 GNDA_2.n1478 GNDA_2.n1441 3.4105
R8570 GNDA_2.n1478 GNDA_2.n1452 3.4105
R8571 GNDA_2.n1478 GNDA_2.n1440 3.4105
R8572 GNDA_2.n1478 GNDA_2.n1453 3.4105
R8573 GNDA_2.n1478 GNDA_2.n1439 3.4105
R8574 GNDA_2.n1478 GNDA_2.n1454 3.4105
R8575 GNDA_2.n1478 GNDA_2.n1438 3.4105
R8576 GNDA_2.n1478 GNDA_2.n1455 3.4105
R8577 GNDA_2.n1478 GNDA_2.n1437 3.4105
R8578 GNDA_2.n1478 GNDA_2.n1456 3.4105
R8579 GNDA_2.n1478 GNDA_2.n1436 3.4105
R8580 GNDA_2.n1478 GNDA_2.n1457 3.4105
R8581 GNDA_2.n1478 GNDA_2.n1435 3.4105
R8582 GNDA_2.n1478 GNDA_2.n1458 3.4105
R8583 GNDA_2.n1478 GNDA_2.n1434 3.4105
R8584 GNDA_2.n1478 GNDA_2.n1459 3.4105
R8585 GNDA_2.n1478 GNDA_2.n1433 3.4105
R8586 GNDA_2.n1478 GNDA_2.n1460 3.4105
R8587 GNDA_2.n1478 GNDA_2.n1432 3.4105
R8588 GNDA_2.n1478 GNDA_2.n1461 3.4105
R8589 GNDA_2.n1478 GNDA_2.n1431 3.4105
R8590 GNDA_2.n1478 GNDA_2.n1462 3.4105
R8591 GNDA_2.n3441 GNDA_2.n1478 3.4105
R8592 GNDA_2.n1545 GNDA_2.n1516 3.4105
R8593 GNDA_2.n1516 GNDA_2.n1447 3.4105
R8594 GNDA_2.n1516 GNDA_2.n1445 3.4105
R8595 GNDA_2.n1516 GNDA_2.n1448 3.4105
R8596 GNDA_2.n1516 GNDA_2.n1444 3.4105
R8597 GNDA_2.n1516 GNDA_2.n1449 3.4105
R8598 GNDA_2.n1516 GNDA_2.n1443 3.4105
R8599 GNDA_2.n1516 GNDA_2.n1450 3.4105
R8600 GNDA_2.n1516 GNDA_2.n1442 3.4105
R8601 GNDA_2.n1516 GNDA_2.n1451 3.4105
R8602 GNDA_2.n1516 GNDA_2.n1441 3.4105
R8603 GNDA_2.n1516 GNDA_2.n1452 3.4105
R8604 GNDA_2.n1516 GNDA_2.n1440 3.4105
R8605 GNDA_2.n1516 GNDA_2.n1453 3.4105
R8606 GNDA_2.n1516 GNDA_2.n1439 3.4105
R8607 GNDA_2.n1516 GNDA_2.n1454 3.4105
R8608 GNDA_2.n1516 GNDA_2.n1438 3.4105
R8609 GNDA_2.n1516 GNDA_2.n1455 3.4105
R8610 GNDA_2.n1516 GNDA_2.n1437 3.4105
R8611 GNDA_2.n1516 GNDA_2.n1456 3.4105
R8612 GNDA_2.n1516 GNDA_2.n1436 3.4105
R8613 GNDA_2.n1516 GNDA_2.n1457 3.4105
R8614 GNDA_2.n1516 GNDA_2.n1435 3.4105
R8615 GNDA_2.n1516 GNDA_2.n1458 3.4105
R8616 GNDA_2.n1516 GNDA_2.n1434 3.4105
R8617 GNDA_2.n1516 GNDA_2.n1459 3.4105
R8618 GNDA_2.n1516 GNDA_2.n1433 3.4105
R8619 GNDA_2.n1516 GNDA_2.n1460 3.4105
R8620 GNDA_2.n1516 GNDA_2.n1432 3.4105
R8621 GNDA_2.n1516 GNDA_2.n1461 3.4105
R8622 GNDA_2.n1516 GNDA_2.n1431 3.4105
R8623 GNDA_2.n1516 GNDA_2.n1462 3.4105
R8624 GNDA_2.n3441 GNDA_2.n1516 3.4105
R8625 GNDA_2.n1545 GNDA_2.n1477 3.4105
R8626 GNDA_2.n1477 GNDA_2.n1447 3.4105
R8627 GNDA_2.n1477 GNDA_2.n1445 3.4105
R8628 GNDA_2.n1477 GNDA_2.n1448 3.4105
R8629 GNDA_2.n1477 GNDA_2.n1444 3.4105
R8630 GNDA_2.n1477 GNDA_2.n1449 3.4105
R8631 GNDA_2.n1477 GNDA_2.n1443 3.4105
R8632 GNDA_2.n1477 GNDA_2.n1450 3.4105
R8633 GNDA_2.n1477 GNDA_2.n1442 3.4105
R8634 GNDA_2.n1477 GNDA_2.n1451 3.4105
R8635 GNDA_2.n1477 GNDA_2.n1441 3.4105
R8636 GNDA_2.n1477 GNDA_2.n1452 3.4105
R8637 GNDA_2.n1477 GNDA_2.n1440 3.4105
R8638 GNDA_2.n1477 GNDA_2.n1453 3.4105
R8639 GNDA_2.n1477 GNDA_2.n1439 3.4105
R8640 GNDA_2.n1477 GNDA_2.n1454 3.4105
R8641 GNDA_2.n1477 GNDA_2.n1438 3.4105
R8642 GNDA_2.n1477 GNDA_2.n1455 3.4105
R8643 GNDA_2.n1477 GNDA_2.n1437 3.4105
R8644 GNDA_2.n1477 GNDA_2.n1456 3.4105
R8645 GNDA_2.n1477 GNDA_2.n1436 3.4105
R8646 GNDA_2.n1477 GNDA_2.n1457 3.4105
R8647 GNDA_2.n1477 GNDA_2.n1435 3.4105
R8648 GNDA_2.n1477 GNDA_2.n1458 3.4105
R8649 GNDA_2.n1477 GNDA_2.n1434 3.4105
R8650 GNDA_2.n1477 GNDA_2.n1459 3.4105
R8651 GNDA_2.n1477 GNDA_2.n1433 3.4105
R8652 GNDA_2.n1477 GNDA_2.n1460 3.4105
R8653 GNDA_2.n1477 GNDA_2.n1432 3.4105
R8654 GNDA_2.n1477 GNDA_2.n1461 3.4105
R8655 GNDA_2.n1477 GNDA_2.n1431 3.4105
R8656 GNDA_2.n1477 GNDA_2.n1462 3.4105
R8657 GNDA_2.n3441 GNDA_2.n1477 3.4105
R8658 GNDA_2.n1545 GNDA_2.n1518 3.4105
R8659 GNDA_2.n1518 GNDA_2.n1447 3.4105
R8660 GNDA_2.n1518 GNDA_2.n1445 3.4105
R8661 GNDA_2.n1518 GNDA_2.n1448 3.4105
R8662 GNDA_2.n1518 GNDA_2.n1444 3.4105
R8663 GNDA_2.n1518 GNDA_2.n1449 3.4105
R8664 GNDA_2.n1518 GNDA_2.n1443 3.4105
R8665 GNDA_2.n1518 GNDA_2.n1450 3.4105
R8666 GNDA_2.n1518 GNDA_2.n1442 3.4105
R8667 GNDA_2.n1518 GNDA_2.n1451 3.4105
R8668 GNDA_2.n1518 GNDA_2.n1441 3.4105
R8669 GNDA_2.n1518 GNDA_2.n1452 3.4105
R8670 GNDA_2.n1518 GNDA_2.n1440 3.4105
R8671 GNDA_2.n1518 GNDA_2.n1453 3.4105
R8672 GNDA_2.n1518 GNDA_2.n1439 3.4105
R8673 GNDA_2.n1518 GNDA_2.n1454 3.4105
R8674 GNDA_2.n1518 GNDA_2.n1438 3.4105
R8675 GNDA_2.n1518 GNDA_2.n1455 3.4105
R8676 GNDA_2.n1518 GNDA_2.n1437 3.4105
R8677 GNDA_2.n1518 GNDA_2.n1456 3.4105
R8678 GNDA_2.n1518 GNDA_2.n1436 3.4105
R8679 GNDA_2.n1518 GNDA_2.n1457 3.4105
R8680 GNDA_2.n1518 GNDA_2.n1435 3.4105
R8681 GNDA_2.n1518 GNDA_2.n1458 3.4105
R8682 GNDA_2.n1518 GNDA_2.n1434 3.4105
R8683 GNDA_2.n1518 GNDA_2.n1459 3.4105
R8684 GNDA_2.n1518 GNDA_2.n1433 3.4105
R8685 GNDA_2.n1518 GNDA_2.n1460 3.4105
R8686 GNDA_2.n1518 GNDA_2.n1432 3.4105
R8687 GNDA_2.n1518 GNDA_2.n1461 3.4105
R8688 GNDA_2.n1518 GNDA_2.n1431 3.4105
R8689 GNDA_2.n1518 GNDA_2.n1462 3.4105
R8690 GNDA_2.n3441 GNDA_2.n1518 3.4105
R8691 GNDA_2.n1545 GNDA_2.n1476 3.4105
R8692 GNDA_2.n1476 GNDA_2.n1447 3.4105
R8693 GNDA_2.n1476 GNDA_2.n1445 3.4105
R8694 GNDA_2.n1476 GNDA_2.n1448 3.4105
R8695 GNDA_2.n1476 GNDA_2.n1444 3.4105
R8696 GNDA_2.n1476 GNDA_2.n1449 3.4105
R8697 GNDA_2.n1476 GNDA_2.n1443 3.4105
R8698 GNDA_2.n1476 GNDA_2.n1450 3.4105
R8699 GNDA_2.n1476 GNDA_2.n1442 3.4105
R8700 GNDA_2.n1476 GNDA_2.n1451 3.4105
R8701 GNDA_2.n1476 GNDA_2.n1441 3.4105
R8702 GNDA_2.n1476 GNDA_2.n1452 3.4105
R8703 GNDA_2.n1476 GNDA_2.n1440 3.4105
R8704 GNDA_2.n1476 GNDA_2.n1453 3.4105
R8705 GNDA_2.n1476 GNDA_2.n1439 3.4105
R8706 GNDA_2.n1476 GNDA_2.n1454 3.4105
R8707 GNDA_2.n1476 GNDA_2.n1438 3.4105
R8708 GNDA_2.n1476 GNDA_2.n1455 3.4105
R8709 GNDA_2.n1476 GNDA_2.n1437 3.4105
R8710 GNDA_2.n1476 GNDA_2.n1456 3.4105
R8711 GNDA_2.n1476 GNDA_2.n1436 3.4105
R8712 GNDA_2.n1476 GNDA_2.n1457 3.4105
R8713 GNDA_2.n1476 GNDA_2.n1435 3.4105
R8714 GNDA_2.n1476 GNDA_2.n1458 3.4105
R8715 GNDA_2.n1476 GNDA_2.n1434 3.4105
R8716 GNDA_2.n1476 GNDA_2.n1459 3.4105
R8717 GNDA_2.n1476 GNDA_2.n1433 3.4105
R8718 GNDA_2.n1476 GNDA_2.n1460 3.4105
R8719 GNDA_2.n1476 GNDA_2.n1432 3.4105
R8720 GNDA_2.n1476 GNDA_2.n1461 3.4105
R8721 GNDA_2.n1476 GNDA_2.n1431 3.4105
R8722 GNDA_2.n1476 GNDA_2.n1462 3.4105
R8723 GNDA_2.n3441 GNDA_2.n1476 3.4105
R8724 GNDA_2.n1545 GNDA_2.n1520 3.4105
R8725 GNDA_2.n1520 GNDA_2.n1447 3.4105
R8726 GNDA_2.n1520 GNDA_2.n1445 3.4105
R8727 GNDA_2.n1520 GNDA_2.n1448 3.4105
R8728 GNDA_2.n1520 GNDA_2.n1444 3.4105
R8729 GNDA_2.n1520 GNDA_2.n1449 3.4105
R8730 GNDA_2.n1520 GNDA_2.n1443 3.4105
R8731 GNDA_2.n1520 GNDA_2.n1450 3.4105
R8732 GNDA_2.n1520 GNDA_2.n1442 3.4105
R8733 GNDA_2.n1520 GNDA_2.n1451 3.4105
R8734 GNDA_2.n1520 GNDA_2.n1441 3.4105
R8735 GNDA_2.n1520 GNDA_2.n1452 3.4105
R8736 GNDA_2.n1520 GNDA_2.n1440 3.4105
R8737 GNDA_2.n1520 GNDA_2.n1453 3.4105
R8738 GNDA_2.n1520 GNDA_2.n1439 3.4105
R8739 GNDA_2.n1520 GNDA_2.n1454 3.4105
R8740 GNDA_2.n1520 GNDA_2.n1438 3.4105
R8741 GNDA_2.n1520 GNDA_2.n1455 3.4105
R8742 GNDA_2.n1520 GNDA_2.n1437 3.4105
R8743 GNDA_2.n1520 GNDA_2.n1456 3.4105
R8744 GNDA_2.n1520 GNDA_2.n1436 3.4105
R8745 GNDA_2.n1520 GNDA_2.n1457 3.4105
R8746 GNDA_2.n1520 GNDA_2.n1435 3.4105
R8747 GNDA_2.n1520 GNDA_2.n1458 3.4105
R8748 GNDA_2.n1520 GNDA_2.n1434 3.4105
R8749 GNDA_2.n1520 GNDA_2.n1459 3.4105
R8750 GNDA_2.n1520 GNDA_2.n1433 3.4105
R8751 GNDA_2.n1520 GNDA_2.n1460 3.4105
R8752 GNDA_2.n1520 GNDA_2.n1432 3.4105
R8753 GNDA_2.n1520 GNDA_2.n1461 3.4105
R8754 GNDA_2.n1520 GNDA_2.n1431 3.4105
R8755 GNDA_2.n1520 GNDA_2.n1462 3.4105
R8756 GNDA_2.n3441 GNDA_2.n1520 3.4105
R8757 GNDA_2.n1545 GNDA_2.n1475 3.4105
R8758 GNDA_2.n1475 GNDA_2.n1447 3.4105
R8759 GNDA_2.n1475 GNDA_2.n1445 3.4105
R8760 GNDA_2.n1475 GNDA_2.n1448 3.4105
R8761 GNDA_2.n1475 GNDA_2.n1444 3.4105
R8762 GNDA_2.n1475 GNDA_2.n1449 3.4105
R8763 GNDA_2.n1475 GNDA_2.n1443 3.4105
R8764 GNDA_2.n1475 GNDA_2.n1450 3.4105
R8765 GNDA_2.n1475 GNDA_2.n1442 3.4105
R8766 GNDA_2.n1475 GNDA_2.n1451 3.4105
R8767 GNDA_2.n1475 GNDA_2.n1441 3.4105
R8768 GNDA_2.n1475 GNDA_2.n1452 3.4105
R8769 GNDA_2.n1475 GNDA_2.n1440 3.4105
R8770 GNDA_2.n1475 GNDA_2.n1453 3.4105
R8771 GNDA_2.n1475 GNDA_2.n1439 3.4105
R8772 GNDA_2.n1475 GNDA_2.n1454 3.4105
R8773 GNDA_2.n1475 GNDA_2.n1438 3.4105
R8774 GNDA_2.n1475 GNDA_2.n1455 3.4105
R8775 GNDA_2.n1475 GNDA_2.n1437 3.4105
R8776 GNDA_2.n1475 GNDA_2.n1456 3.4105
R8777 GNDA_2.n1475 GNDA_2.n1436 3.4105
R8778 GNDA_2.n1475 GNDA_2.n1457 3.4105
R8779 GNDA_2.n1475 GNDA_2.n1435 3.4105
R8780 GNDA_2.n1475 GNDA_2.n1458 3.4105
R8781 GNDA_2.n1475 GNDA_2.n1434 3.4105
R8782 GNDA_2.n1475 GNDA_2.n1459 3.4105
R8783 GNDA_2.n1475 GNDA_2.n1433 3.4105
R8784 GNDA_2.n1475 GNDA_2.n1460 3.4105
R8785 GNDA_2.n1475 GNDA_2.n1432 3.4105
R8786 GNDA_2.n1475 GNDA_2.n1461 3.4105
R8787 GNDA_2.n1475 GNDA_2.n1431 3.4105
R8788 GNDA_2.n1475 GNDA_2.n1462 3.4105
R8789 GNDA_2.n3441 GNDA_2.n1475 3.4105
R8790 GNDA_2.n1545 GNDA_2.n1522 3.4105
R8791 GNDA_2.n1522 GNDA_2.n1447 3.4105
R8792 GNDA_2.n1522 GNDA_2.n1445 3.4105
R8793 GNDA_2.n1522 GNDA_2.n1448 3.4105
R8794 GNDA_2.n1522 GNDA_2.n1444 3.4105
R8795 GNDA_2.n1522 GNDA_2.n1449 3.4105
R8796 GNDA_2.n1522 GNDA_2.n1443 3.4105
R8797 GNDA_2.n1522 GNDA_2.n1450 3.4105
R8798 GNDA_2.n1522 GNDA_2.n1442 3.4105
R8799 GNDA_2.n1522 GNDA_2.n1451 3.4105
R8800 GNDA_2.n1522 GNDA_2.n1441 3.4105
R8801 GNDA_2.n1522 GNDA_2.n1452 3.4105
R8802 GNDA_2.n1522 GNDA_2.n1440 3.4105
R8803 GNDA_2.n1522 GNDA_2.n1453 3.4105
R8804 GNDA_2.n1522 GNDA_2.n1439 3.4105
R8805 GNDA_2.n1522 GNDA_2.n1454 3.4105
R8806 GNDA_2.n1522 GNDA_2.n1438 3.4105
R8807 GNDA_2.n1522 GNDA_2.n1455 3.4105
R8808 GNDA_2.n1522 GNDA_2.n1437 3.4105
R8809 GNDA_2.n1522 GNDA_2.n1456 3.4105
R8810 GNDA_2.n1522 GNDA_2.n1436 3.4105
R8811 GNDA_2.n1522 GNDA_2.n1457 3.4105
R8812 GNDA_2.n1522 GNDA_2.n1435 3.4105
R8813 GNDA_2.n1522 GNDA_2.n1458 3.4105
R8814 GNDA_2.n1522 GNDA_2.n1434 3.4105
R8815 GNDA_2.n1522 GNDA_2.n1459 3.4105
R8816 GNDA_2.n1522 GNDA_2.n1433 3.4105
R8817 GNDA_2.n1522 GNDA_2.n1460 3.4105
R8818 GNDA_2.n1522 GNDA_2.n1432 3.4105
R8819 GNDA_2.n1522 GNDA_2.n1461 3.4105
R8820 GNDA_2.n1522 GNDA_2.n1431 3.4105
R8821 GNDA_2.n1522 GNDA_2.n1462 3.4105
R8822 GNDA_2.n3441 GNDA_2.n1522 3.4105
R8823 GNDA_2.n1545 GNDA_2.n1474 3.4105
R8824 GNDA_2.n1474 GNDA_2.n1447 3.4105
R8825 GNDA_2.n1474 GNDA_2.n1445 3.4105
R8826 GNDA_2.n1474 GNDA_2.n1448 3.4105
R8827 GNDA_2.n1474 GNDA_2.n1444 3.4105
R8828 GNDA_2.n1474 GNDA_2.n1449 3.4105
R8829 GNDA_2.n1474 GNDA_2.n1443 3.4105
R8830 GNDA_2.n1474 GNDA_2.n1450 3.4105
R8831 GNDA_2.n1474 GNDA_2.n1442 3.4105
R8832 GNDA_2.n1474 GNDA_2.n1451 3.4105
R8833 GNDA_2.n1474 GNDA_2.n1441 3.4105
R8834 GNDA_2.n1474 GNDA_2.n1452 3.4105
R8835 GNDA_2.n1474 GNDA_2.n1440 3.4105
R8836 GNDA_2.n1474 GNDA_2.n1453 3.4105
R8837 GNDA_2.n1474 GNDA_2.n1439 3.4105
R8838 GNDA_2.n1474 GNDA_2.n1454 3.4105
R8839 GNDA_2.n1474 GNDA_2.n1438 3.4105
R8840 GNDA_2.n1474 GNDA_2.n1455 3.4105
R8841 GNDA_2.n1474 GNDA_2.n1437 3.4105
R8842 GNDA_2.n1474 GNDA_2.n1456 3.4105
R8843 GNDA_2.n1474 GNDA_2.n1436 3.4105
R8844 GNDA_2.n1474 GNDA_2.n1457 3.4105
R8845 GNDA_2.n1474 GNDA_2.n1435 3.4105
R8846 GNDA_2.n1474 GNDA_2.n1458 3.4105
R8847 GNDA_2.n1474 GNDA_2.n1434 3.4105
R8848 GNDA_2.n1474 GNDA_2.n1459 3.4105
R8849 GNDA_2.n1474 GNDA_2.n1433 3.4105
R8850 GNDA_2.n1474 GNDA_2.n1460 3.4105
R8851 GNDA_2.n1474 GNDA_2.n1432 3.4105
R8852 GNDA_2.n1474 GNDA_2.n1461 3.4105
R8853 GNDA_2.n1474 GNDA_2.n1431 3.4105
R8854 GNDA_2.n1474 GNDA_2.n1462 3.4105
R8855 GNDA_2.n3441 GNDA_2.n1474 3.4105
R8856 GNDA_2.n1545 GNDA_2.n1524 3.4105
R8857 GNDA_2.n1524 GNDA_2.n1447 3.4105
R8858 GNDA_2.n1524 GNDA_2.n1445 3.4105
R8859 GNDA_2.n1524 GNDA_2.n1448 3.4105
R8860 GNDA_2.n1524 GNDA_2.n1444 3.4105
R8861 GNDA_2.n1524 GNDA_2.n1449 3.4105
R8862 GNDA_2.n1524 GNDA_2.n1443 3.4105
R8863 GNDA_2.n1524 GNDA_2.n1450 3.4105
R8864 GNDA_2.n1524 GNDA_2.n1442 3.4105
R8865 GNDA_2.n1524 GNDA_2.n1451 3.4105
R8866 GNDA_2.n1524 GNDA_2.n1441 3.4105
R8867 GNDA_2.n1524 GNDA_2.n1452 3.4105
R8868 GNDA_2.n1524 GNDA_2.n1440 3.4105
R8869 GNDA_2.n1524 GNDA_2.n1453 3.4105
R8870 GNDA_2.n1524 GNDA_2.n1439 3.4105
R8871 GNDA_2.n1524 GNDA_2.n1454 3.4105
R8872 GNDA_2.n1524 GNDA_2.n1438 3.4105
R8873 GNDA_2.n1524 GNDA_2.n1455 3.4105
R8874 GNDA_2.n1524 GNDA_2.n1437 3.4105
R8875 GNDA_2.n1524 GNDA_2.n1456 3.4105
R8876 GNDA_2.n1524 GNDA_2.n1436 3.4105
R8877 GNDA_2.n1524 GNDA_2.n1457 3.4105
R8878 GNDA_2.n1524 GNDA_2.n1435 3.4105
R8879 GNDA_2.n1524 GNDA_2.n1458 3.4105
R8880 GNDA_2.n1524 GNDA_2.n1434 3.4105
R8881 GNDA_2.n1524 GNDA_2.n1459 3.4105
R8882 GNDA_2.n1524 GNDA_2.n1433 3.4105
R8883 GNDA_2.n1524 GNDA_2.n1460 3.4105
R8884 GNDA_2.n1524 GNDA_2.n1432 3.4105
R8885 GNDA_2.n1524 GNDA_2.n1461 3.4105
R8886 GNDA_2.n1524 GNDA_2.n1431 3.4105
R8887 GNDA_2.n1524 GNDA_2.n1462 3.4105
R8888 GNDA_2.n3441 GNDA_2.n1524 3.4105
R8889 GNDA_2.n1545 GNDA_2.n1473 3.4105
R8890 GNDA_2.n1473 GNDA_2.n1447 3.4105
R8891 GNDA_2.n1473 GNDA_2.n1445 3.4105
R8892 GNDA_2.n1473 GNDA_2.n1448 3.4105
R8893 GNDA_2.n1473 GNDA_2.n1444 3.4105
R8894 GNDA_2.n1473 GNDA_2.n1449 3.4105
R8895 GNDA_2.n1473 GNDA_2.n1443 3.4105
R8896 GNDA_2.n1473 GNDA_2.n1450 3.4105
R8897 GNDA_2.n1473 GNDA_2.n1442 3.4105
R8898 GNDA_2.n1473 GNDA_2.n1451 3.4105
R8899 GNDA_2.n1473 GNDA_2.n1441 3.4105
R8900 GNDA_2.n1473 GNDA_2.n1452 3.4105
R8901 GNDA_2.n1473 GNDA_2.n1440 3.4105
R8902 GNDA_2.n1473 GNDA_2.n1453 3.4105
R8903 GNDA_2.n1473 GNDA_2.n1439 3.4105
R8904 GNDA_2.n1473 GNDA_2.n1454 3.4105
R8905 GNDA_2.n1473 GNDA_2.n1438 3.4105
R8906 GNDA_2.n1473 GNDA_2.n1455 3.4105
R8907 GNDA_2.n1473 GNDA_2.n1437 3.4105
R8908 GNDA_2.n1473 GNDA_2.n1456 3.4105
R8909 GNDA_2.n1473 GNDA_2.n1436 3.4105
R8910 GNDA_2.n1473 GNDA_2.n1457 3.4105
R8911 GNDA_2.n1473 GNDA_2.n1435 3.4105
R8912 GNDA_2.n1473 GNDA_2.n1458 3.4105
R8913 GNDA_2.n1473 GNDA_2.n1434 3.4105
R8914 GNDA_2.n1473 GNDA_2.n1459 3.4105
R8915 GNDA_2.n1473 GNDA_2.n1433 3.4105
R8916 GNDA_2.n1473 GNDA_2.n1460 3.4105
R8917 GNDA_2.n1473 GNDA_2.n1432 3.4105
R8918 GNDA_2.n1473 GNDA_2.n1461 3.4105
R8919 GNDA_2.n1473 GNDA_2.n1431 3.4105
R8920 GNDA_2.n1473 GNDA_2.n1462 3.4105
R8921 GNDA_2.n3441 GNDA_2.n1473 3.4105
R8922 GNDA_2.n1545 GNDA_2.n1526 3.4105
R8923 GNDA_2.n1526 GNDA_2.n1447 3.4105
R8924 GNDA_2.n1526 GNDA_2.n1445 3.4105
R8925 GNDA_2.n1526 GNDA_2.n1448 3.4105
R8926 GNDA_2.n1526 GNDA_2.n1444 3.4105
R8927 GNDA_2.n1526 GNDA_2.n1449 3.4105
R8928 GNDA_2.n1526 GNDA_2.n1443 3.4105
R8929 GNDA_2.n1526 GNDA_2.n1450 3.4105
R8930 GNDA_2.n1526 GNDA_2.n1442 3.4105
R8931 GNDA_2.n1526 GNDA_2.n1451 3.4105
R8932 GNDA_2.n1526 GNDA_2.n1441 3.4105
R8933 GNDA_2.n1526 GNDA_2.n1452 3.4105
R8934 GNDA_2.n1526 GNDA_2.n1440 3.4105
R8935 GNDA_2.n1526 GNDA_2.n1453 3.4105
R8936 GNDA_2.n1526 GNDA_2.n1439 3.4105
R8937 GNDA_2.n1526 GNDA_2.n1454 3.4105
R8938 GNDA_2.n1526 GNDA_2.n1438 3.4105
R8939 GNDA_2.n1526 GNDA_2.n1455 3.4105
R8940 GNDA_2.n1526 GNDA_2.n1437 3.4105
R8941 GNDA_2.n1526 GNDA_2.n1456 3.4105
R8942 GNDA_2.n1526 GNDA_2.n1436 3.4105
R8943 GNDA_2.n1526 GNDA_2.n1457 3.4105
R8944 GNDA_2.n1526 GNDA_2.n1435 3.4105
R8945 GNDA_2.n1526 GNDA_2.n1458 3.4105
R8946 GNDA_2.n1526 GNDA_2.n1434 3.4105
R8947 GNDA_2.n1526 GNDA_2.n1459 3.4105
R8948 GNDA_2.n1526 GNDA_2.n1433 3.4105
R8949 GNDA_2.n1526 GNDA_2.n1460 3.4105
R8950 GNDA_2.n1526 GNDA_2.n1432 3.4105
R8951 GNDA_2.n1526 GNDA_2.n1461 3.4105
R8952 GNDA_2.n1526 GNDA_2.n1431 3.4105
R8953 GNDA_2.n1526 GNDA_2.n1462 3.4105
R8954 GNDA_2.n3441 GNDA_2.n1526 3.4105
R8955 GNDA_2.n1545 GNDA_2.n1472 3.4105
R8956 GNDA_2.n1472 GNDA_2.n1447 3.4105
R8957 GNDA_2.n1472 GNDA_2.n1445 3.4105
R8958 GNDA_2.n1472 GNDA_2.n1448 3.4105
R8959 GNDA_2.n1472 GNDA_2.n1444 3.4105
R8960 GNDA_2.n1472 GNDA_2.n1449 3.4105
R8961 GNDA_2.n1472 GNDA_2.n1443 3.4105
R8962 GNDA_2.n1472 GNDA_2.n1450 3.4105
R8963 GNDA_2.n1472 GNDA_2.n1442 3.4105
R8964 GNDA_2.n1472 GNDA_2.n1451 3.4105
R8965 GNDA_2.n1472 GNDA_2.n1441 3.4105
R8966 GNDA_2.n1472 GNDA_2.n1452 3.4105
R8967 GNDA_2.n1472 GNDA_2.n1440 3.4105
R8968 GNDA_2.n1472 GNDA_2.n1453 3.4105
R8969 GNDA_2.n1472 GNDA_2.n1439 3.4105
R8970 GNDA_2.n1472 GNDA_2.n1454 3.4105
R8971 GNDA_2.n1472 GNDA_2.n1438 3.4105
R8972 GNDA_2.n1472 GNDA_2.n1455 3.4105
R8973 GNDA_2.n1472 GNDA_2.n1437 3.4105
R8974 GNDA_2.n1472 GNDA_2.n1456 3.4105
R8975 GNDA_2.n1472 GNDA_2.n1436 3.4105
R8976 GNDA_2.n1472 GNDA_2.n1457 3.4105
R8977 GNDA_2.n1472 GNDA_2.n1435 3.4105
R8978 GNDA_2.n1472 GNDA_2.n1458 3.4105
R8979 GNDA_2.n1472 GNDA_2.n1434 3.4105
R8980 GNDA_2.n1472 GNDA_2.n1459 3.4105
R8981 GNDA_2.n1472 GNDA_2.n1433 3.4105
R8982 GNDA_2.n1472 GNDA_2.n1460 3.4105
R8983 GNDA_2.n1472 GNDA_2.n1432 3.4105
R8984 GNDA_2.n1472 GNDA_2.n1461 3.4105
R8985 GNDA_2.n1472 GNDA_2.n1431 3.4105
R8986 GNDA_2.n1472 GNDA_2.n1462 3.4105
R8987 GNDA_2.n3441 GNDA_2.n1472 3.4105
R8988 GNDA_2.n1545 GNDA_2.n1528 3.4105
R8989 GNDA_2.n1528 GNDA_2.n1447 3.4105
R8990 GNDA_2.n1528 GNDA_2.n1445 3.4105
R8991 GNDA_2.n1528 GNDA_2.n1448 3.4105
R8992 GNDA_2.n1528 GNDA_2.n1444 3.4105
R8993 GNDA_2.n1528 GNDA_2.n1449 3.4105
R8994 GNDA_2.n1528 GNDA_2.n1443 3.4105
R8995 GNDA_2.n1528 GNDA_2.n1450 3.4105
R8996 GNDA_2.n1528 GNDA_2.n1442 3.4105
R8997 GNDA_2.n1528 GNDA_2.n1451 3.4105
R8998 GNDA_2.n1528 GNDA_2.n1441 3.4105
R8999 GNDA_2.n1528 GNDA_2.n1452 3.4105
R9000 GNDA_2.n1528 GNDA_2.n1440 3.4105
R9001 GNDA_2.n1528 GNDA_2.n1453 3.4105
R9002 GNDA_2.n1528 GNDA_2.n1439 3.4105
R9003 GNDA_2.n1528 GNDA_2.n1454 3.4105
R9004 GNDA_2.n1528 GNDA_2.n1438 3.4105
R9005 GNDA_2.n1528 GNDA_2.n1455 3.4105
R9006 GNDA_2.n1528 GNDA_2.n1437 3.4105
R9007 GNDA_2.n1528 GNDA_2.n1456 3.4105
R9008 GNDA_2.n1528 GNDA_2.n1436 3.4105
R9009 GNDA_2.n1528 GNDA_2.n1457 3.4105
R9010 GNDA_2.n1528 GNDA_2.n1435 3.4105
R9011 GNDA_2.n1528 GNDA_2.n1458 3.4105
R9012 GNDA_2.n1528 GNDA_2.n1434 3.4105
R9013 GNDA_2.n1528 GNDA_2.n1459 3.4105
R9014 GNDA_2.n1528 GNDA_2.n1433 3.4105
R9015 GNDA_2.n1528 GNDA_2.n1460 3.4105
R9016 GNDA_2.n1528 GNDA_2.n1432 3.4105
R9017 GNDA_2.n1528 GNDA_2.n1461 3.4105
R9018 GNDA_2.n1528 GNDA_2.n1431 3.4105
R9019 GNDA_2.n1528 GNDA_2.n1462 3.4105
R9020 GNDA_2.n3441 GNDA_2.n1528 3.4105
R9021 GNDA_2.n1545 GNDA_2.n1471 3.4105
R9022 GNDA_2.n1471 GNDA_2.n1447 3.4105
R9023 GNDA_2.n1471 GNDA_2.n1445 3.4105
R9024 GNDA_2.n1471 GNDA_2.n1448 3.4105
R9025 GNDA_2.n1471 GNDA_2.n1444 3.4105
R9026 GNDA_2.n1471 GNDA_2.n1449 3.4105
R9027 GNDA_2.n1471 GNDA_2.n1443 3.4105
R9028 GNDA_2.n1471 GNDA_2.n1450 3.4105
R9029 GNDA_2.n1471 GNDA_2.n1442 3.4105
R9030 GNDA_2.n1471 GNDA_2.n1451 3.4105
R9031 GNDA_2.n1471 GNDA_2.n1441 3.4105
R9032 GNDA_2.n1471 GNDA_2.n1452 3.4105
R9033 GNDA_2.n1471 GNDA_2.n1440 3.4105
R9034 GNDA_2.n1471 GNDA_2.n1453 3.4105
R9035 GNDA_2.n1471 GNDA_2.n1439 3.4105
R9036 GNDA_2.n1471 GNDA_2.n1454 3.4105
R9037 GNDA_2.n1471 GNDA_2.n1438 3.4105
R9038 GNDA_2.n1471 GNDA_2.n1455 3.4105
R9039 GNDA_2.n1471 GNDA_2.n1437 3.4105
R9040 GNDA_2.n1471 GNDA_2.n1456 3.4105
R9041 GNDA_2.n1471 GNDA_2.n1436 3.4105
R9042 GNDA_2.n1471 GNDA_2.n1457 3.4105
R9043 GNDA_2.n1471 GNDA_2.n1435 3.4105
R9044 GNDA_2.n1471 GNDA_2.n1458 3.4105
R9045 GNDA_2.n1471 GNDA_2.n1434 3.4105
R9046 GNDA_2.n1471 GNDA_2.n1459 3.4105
R9047 GNDA_2.n1471 GNDA_2.n1433 3.4105
R9048 GNDA_2.n1471 GNDA_2.n1460 3.4105
R9049 GNDA_2.n1471 GNDA_2.n1432 3.4105
R9050 GNDA_2.n1471 GNDA_2.n1461 3.4105
R9051 GNDA_2.n1471 GNDA_2.n1431 3.4105
R9052 GNDA_2.n1471 GNDA_2.n1462 3.4105
R9053 GNDA_2.n3441 GNDA_2.n1471 3.4105
R9054 GNDA_2.n1545 GNDA_2.n1530 3.4105
R9055 GNDA_2.n1530 GNDA_2.n1447 3.4105
R9056 GNDA_2.n1530 GNDA_2.n1445 3.4105
R9057 GNDA_2.n1530 GNDA_2.n1448 3.4105
R9058 GNDA_2.n1530 GNDA_2.n1444 3.4105
R9059 GNDA_2.n1530 GNDA_2.n1449 3.4105
R9060 GNDA_2.n1530 GNDA_2.n1443 3.4105
R9061 GNDA_2.n1530 GNDA_2.n1450 3.4105
R9062 GNDA_2.n1530 GNDA_2.n1442 3.4105
R9063 GNDA_2.n1530 GNDA_2.n1451 3.4105
R9064 GNDA_2.n1530 GNDA_2.n1441 3.4105
R9065 GNDA_2.n1530 GNDA_2.n1452 3.4105
R9066 GNDA_2.n1530 GNDA_2.n1440 3.4105
R9067 GNDA_2.n1530 GNDA_2.n1453 3.4105
R9068 GNDA_2.n1530 GNDA_2.n1439 3.4105
R9069 GNDA_2.n1530 GNDA_2.n1454 3.4105
R9070 GNDA_2.n1530 GNDA_2.n1438 3.4105
R9071 GNDA_2.n1530 GNDA_2.n1455 3.4105
R9072 GNDA_2.n1530 GNDA_2.n1437 3.4105
R9073 GNDA_2.n1530 GNDA_2.n1456 3.4105
R9074 GNDA_2.n1530 GNDA_2.n1436 3.4105
R9075 GNDA_2.n1530 GNDA_2.n1457 3.4105
R9076 GNDA_2.n1530 GNDA_2.n1435 3.4105
R9077 GNDA_2.n1530 GNDA_2.n1458 3.4105
R9078 GNDA_2.n1530 GNDA_2.n1434 3.4105
R9079 GNDA_2.n1530 GNDA_2.n1459 3.4105
R9080 GNDA_2.n1530 GNDA_2.n1433 3.4105
R9081 GNDA_2.n1530 GNDA_2.n1460 3.4105
R9082 GNDA_2.n1530 GNDA_2.n1432 3.4105
R9083 GNDA_2.n1530 GNDA_2.n1461 3.4105
R9084 GNDA_2.n1530 GNDA_2.n1431 3.4105
R9085 GNDA_2.n1530 GNDA_2.n1462 3.4105
R9086 GNDA_2.n3441 GNDA_2.n1530 3.4105
R9087 GNDA_2.n1545 GNDA_2.n1470 3.4105
R9088 GNDA_2.n1470 GNDA_2.n1447 3.4105
R9089 GNDA_2.n1470 GNDA_2.n1445 3.4105
R9090 GNDA_2.n1470 GNDA_2.n1448 3.4105
R9091 GNDA_2.n1470 GNDA_2.n1444 3.4105
R9092 GNDA_2.n1470 GNDA_2.n1449 3.4105
R9093 GNDA_2.n1470 GNDA_2.n1443 3.4105
R9094 GNDA_2.n1470 GNDA_2.n1450 3.4105
R9095 GNDA_2.n1470 GNDA_2.n1442 3.4105
R9096 GNDA_2.n1470 GNDA_2.n1451 3.4105
R9097 GNDA_2.n1470 GNDA_2.n1441 3.4105
R9098 GNDA_2.n1470 GNDA_2.n1452 3.4105
R9099 GNDA_2.n1470 GNDA_2.n1440 3.4105
R9100 GNDA_2.n1470 GNDA_2.n1453 3.4105
R9101 GNDA_2.n1470 GNDA_2.n1439 3.4105
R9102 GNDA_2.n1470 GNDA_2.n1454 3.4105
R9103 GNDA_2.n1470 GNDA_2.n1438 3.4105
R9104 GNDA_2.n1470 GNDA_2.n1455 3.4105
R9105 GNDA_2.n1470 GNDA_2.n1437 3.4105
R9106 GNDA_2.n1470 GNDA_2.n1456 3.4105
R9107 GNDA_2.n1470 GNDA_2.n1436 3.4105
R9108 GNDA_2.n1470 GNDA_2.n1457 3.4105
R9109 GNDA_2.n1470 GNDA_2.n1435 3.4105
R9110 GNDA_2.n1470 GNDA_2.n1458 3.4105
R9111 GNDA_2.n1470 GNDA_2.n1434 3.4105
R9112 GNDA_2.n1470 GNDA_2.n1459 3.4105
R9113 GNDA_2.n1470 GNDA_2.n1433 3.4105
R9114 GNDA_2.n1470 GNDA_2.n1460 3.4105
R9115 GNDA_2.n1470 GNDA_2.n1432 3.4105
R9116 GNDA_2.n1470 GNDA_2.n1461 3.4105
R9117 GNDA_2.n1470 GNDA_2.n1431 3.4105
R9118 GNDA_2.n1470 GNDA_2.n1462 3.4105
R9119 GNDA_2.n3441 GNDA_2.n1470 3.4105
R9120 GNDA_2.n1545 GNDA_2.n1532 3.4105
R9121 GNDA_2.n1532 GNDA_2.n1447 3.4105
R9122 GNDA_2.n1532 GNDA_2.n1445 3.4105
R9123 GNDA_2.n1532 GNDA_2.n1448 3.4105
R9124 GNDA_2.n1532 GNDA_2.n1444 3.4105
R9125 GNDA_2.n1532 GNDA_2.n1449 3.4105
R9126 GNDA_2.n1532 GNDA_2.n1443 3.4105
R9127 GNDA_2.n1532 GNDA_2.n1450 3.4105
R9128 GNDA_2.n1532 GNDA_2.n1442 3.4105
R9129 GNDA_2.n1532 GNDA_2.n1451 3.4105
R9130 GNDA_2.n1532 GNDA_2.n1441 3.4105
R9131 GNDA_2.n1532 GNDA_2.n1452 3.4105
R9132 GNDA_2.n1532 GNDA_2.n1440 3.4105
R9133 GNDA_2.n1532 GNDA_2.n1453 3.4105
R9134 GNDA_2.n1532 GNDA_2.n1439 3.4105
R9135 GNDA_2.n1532 GNDA_2.n1454 3.4105
R9136 GNDA_2.n1532 GNDA_2.n1438 3.4105
R9137 GNDA_2.n1532 GNDA_2.n1455 3.4105
R9138 GNDA_2.n1532 GNDA_2.n1437 3.4105
R9139 GNDA_2.n1532 GNDA_2.n1456 3.4105
R9140 GNDA_2.n1532 GNDA_2.n1436 3.4105
R9141 GNDA_2.n1532 GNDA_2.n1457 3.4105
R9142 GNDA_2.n1532 GNDA_2.n1435 3.4105
R9143 GNDA_2.n1532 GNDA_2.n1458 3.4105
R9144 GNDA_2.n1532 GNDA_2.n1434 3.4105
R9145 GNDA_2.n1532 GNDA_2.n1459 3.4105
R9146 GNDA_2.n1532 GNDA_2.n1433 3.4105
R9147 GNDA_2.n1532 GNDA_2.n1460 3.4105
R9148 GNDA_2.n1532 GNDA_2.n1432 3.4105
R9149 GNDA_2.n1532 GNDA_2.n1461 3.4105
R9150 GNDA_2.n1532 GNDA_2.n1431 3.4105
R9151 GNDA_2.n1532 GNDA_2.n1462 3.4105
R9152 GNDA_2.n3441 GNDA_2.n1532 3.4105
R9153 GNDA_2.n1545 GNDA_2.n1469 3.4105
R9154 GNDA_2.n1469 GNDA_2.n1447 3.4105
R9155 GNDA_2.n1469 GNDA_2.n1445 3.4105
R9156 GNDA_2.n1469 GNDA_2.n1448 3.4105
R9157 GNDA_2.n1469 GNDA_2.n1444 3.4105
R9158 GNDA_2.n1469 GNDA_2.n1449 3.4105
R9159 GNDA_2.n1469 GNDA_2.n1443 3.4105
R9160 GNDA_2.n1469 GNDA_2.n1450 3.4105
R9161 GNDA_2.n1469 GNDA_2.n1442 3.4105
R9162 GNDA_2.n1469 GNDA_2.n1451 3.4105
R9163 GNDA_2.n1469 GNDA_2.n1441 3.4105
R9164 GNDA_2.n1469 GNDA_2.n1452 3.4105
R9165 GNDA_2.n1469 GNDA_2.n1440 3.4105
R9166 GNDA_2.n1469 GNDA_2.n1453 3.4105
R9167 GNDA_2.n1469 GNDA_2.n1439 3.4105
R9168 GNDA_2.n1469 GNDA_2.n1454 3.4105
R9169 GNDA_2.n1469 GNDA_2.n1438 3.4105
R9170 GNDA_2.n1469 GNDA_2.n1455 3.4105
R9171 GNDA_2.n1469 GNDA_2.n1437 3.4105
R9172 GNDA_2.n1469 GNDA_2.n1456 3.4105
R9173 GNDA_2.n1469 GNDA_2.n1436 3.4105
R9174 GNDA_2.n1469 GNDA_2.n1457 3.4105
R9175 GNDA_2.n1469 GNDA_2.n1435 3.4105
R9176 GNDA_2.n1469 GNDA_2.n1458 3.4105
R9177 GNDA_2.n1469 GNDA_2.n1434 3.4105
R9178 GNDA_2.n1469 GNDA_2.n1459 3.4105
R9179 GNDA_2.n1469 GNDA_2.n1433 3.4105
R9180 GNDA_2.n1469 GNDA_2.n1460 3.4105
R9181 GNDA_2.n1469 GNDA_2.n1432 3.4105
R9182 GNDA_2.n1469 GNDA_2.n1461 3.4105
R9183 GNDA_2.n1469 GNDA_2.n1431 3.4105
R9184 GNDA_2.n1469 GNDA_2.n1462 3.4105
R9185 GNDA_2.n3441 GNDA_2.n1469 3.4105
R9186 GNDA_2.n1545 GNDA_2.n1534 3.4105
R9187 GNDA_2.n1534 GNDA_2.n1447 3.4105
R9188 GNDA_2.n1534 GNDA_2.n1445 3.4105
R9189 GNDA_2.n1534 GNDA_2.n1448 3.4105
R9190 GNDA_2.n1534 GNDA_2.n1444 3.4105
R9191 GNDA_2.n1534 GNDA_2.n1449 3.4105
R9192 GNDA_2.n1534 GNDA_2.n1443 3.4105
R9193 GNDA_2.n1534 GNDA_2.n1450 3.4105
R9194 GNDA_2.n1534 GNDA_2.n1442 3.4105
R9195 GNDA_2.n1534 GNDA_2.n1451 3.4105
R9196 GNDA_2.n1534 GNDA_2.n1441 3.4105
R9197 GNDA_2.n1534 GNDA_2.n1452 3.4105
R9198 GNDA_2.n1534 GNDA_2.n1440 3.4105
R9199 GNDA_2.n1534 GNDA_2.n1453 3.4105
R9200 GNDA_2.n1534 GNDA_2.n1439 3.4105
R9201 GNDA_2.n1534 GNDA_2.n1454 3.4105
R9202 GNDA_2.n1534 GNDA_2.n1438 3.4105
R9203 GNDA_2.n1534 GNDA_2.n1455 3.4105
R9204 GNDA_2.n1534 GNDA_2.n1437 3.4105
R9205 GNDA_2.n1534 GNDA_2.n1456 3.4105
R9206 GNDA_2.n1534 GNDA_2.n1436 3.4105
R9207 GNDA_2.n1534 GNDA_2.n1457 3.4105
R9208 GNDA_2.n1534 GNDA_2.n1435 3.4105
R9209 GNDA_2.n1534 GNDA_2.n1458 3.4105
R9210 GNDA_2.n1534 GNDA_2.n1434 3.4105
R9211 GNDA_2.n1534 GNDA_2.n1459 3.4105
R9212 GNDA_2.n1534 GNDA_2.n1433 3.4105
R9213 GNDA_2.n1534 GNDA_2.n1460 3.4105
R9214 GNDA_2.n1534 GNDA_2.n1432 3.4105
R9215 GNDA_2.n1534 GNDA_2.n1461 3.4105
R9216 GNDA_2.n1534 GNDA_2.n1431 3.4105
R9217 GNDA_2.n1534 GNDA_2.n1462 3.4105
R9218 GNDA_2.n3441 GNDA_2.n1534 3.4105
R9219 GNDA_2.n1545 GNDA_2.n1468 3.4105
R9220 GNDA_2.n1468 GNDA_2.n1447 3.4105
R9221 GNDA_2.n1468 GNDA_2.n1445 3.4105
R9222 GNDA_2.n1468 GNDA_2.n1448 3.4105
R9223 GNDA_2.n1468 GNDA_2.n1444 3.4105
R9224 GNDA_2.n1468 GNDA_2.n1449 3.4105
R9225 GNDA_2.n1468 GNDA_2.n1443 3.4105
R9226 GNDA_2.n1468 GNDA_2.n1450 3.4105
R9227 GNDA_2.n1468 GNDA_2.n1442 3.4105
R9228 GNDA_2.n1468 GNDA_2.n1451 3.4105
R9229 GNDA_2.n1468 GNDA_2.n1441 3.4105
R9230 GNDA_2.n1468 GNDA_2.n1452 3.4105
R9231 GNDA_2.n1468 GNDA_2.n1440 3.4105
R9232 GNDA_2.n1468 GNDA_2.n1453 3.4105
R9233 GNDA_2.n1468 GNDA_2.n1439 3.4105
R9234 GNDA_2.n1468 GNDA_2.n1454 3.4105
R9235 GNDA_2.n1468 GNDA_2.n1438 3.4105
R9236 GNDA_2.n1468 GNDA_2.n1455 3.4105
R9237 GNDA_2.n1468 GNDA_2.n1437 3.4105
R9238 GNDA_2.n1468 GNDA_2.n1456 3.4105
R9239 GNDA_2.n1468 GNDA_2.n1436 3.4105
R9240 GNDA_2.n1468 GNDA_2.n1457 3.4105
R9241 GNDA_2.n1468 GNDA_2.n1435 3.4105
R9242 GNDA_2.n1468 GNDA_2.n1458 3.4105
R9243 GNDA_2.n1468 GNDA_2.n1434 3.4105
R9244 GNDA_2.n1468 GNDA_2.n1459 3.4105
R9245 GNDA_2.n1468 GNDA_2.n1433 3.4105
R9246 GNDA_2.n1468 GNDA_2.n1460 3.4105
R9247 GNDA_2.n1468 GNDA_2.n1432 3.4105
R9248 GNDA_2.n1468 GNDA_2.n1461 3.4105
R9249 GNDA_2.n1468 GNDA_2.n1431 3.4105
R9250 GNDA_2.n1468 GNDA_2.n1462 3.4105
R9251 GNDA_2.n3441 GNDA_2.n1468 3.4105
R9252 GNDA_2.n1545 GNDA_2.n1536 3.4105
R9253 GNDA_2.n1536 GNDA_2.n1447 3.4105
R9254 GNDA_2.n1536 GNDA_2.n1445 3.4105
R9255 GNDA_2.n1536 GNDA_2.n1448 3.4105
R9256 GNDA_2.n1536 GNDA_2.n1444 3.4105
R9257 GNDA_2.n1536 GNDA_2.n1449 3.4105
R9258 GNDA_2.n1536 GNDA_2.n1443 3.4105
R9259 GNDA_2.n1536 GNDA_2.n1450 3.4105
R9260 GNDA_2.n1536 GNDA_2.n1442 3.4105
R9261 GNDA_2.n1536 GNDA_2.n1451 3.4105
R9262 GNDA_2.n1536 GNDA_2.n1441 3.4105
R9263 GNDA_2.n1536 GNDA_2.n1452 3.4105
R9264 GNDA_2.n1536 GNDA_2.n1440 3.4105
R9265 GNDA_2.n1536 GNDA_2.n1453 3.4105
R9266 GNDA_2.n1536 GNDA_2.n1439 3.4105
R9267 GNDA_2.n1536 GNDA_2.n1454 3.4105
R9268 GNDA_2.n1536 GNDA_2.n1438 3.4105
R9269 GNDA_2.n1536 GNDA_2.n1455 3.4105
R9270 GNDA_2.n1536 GNDA_2.n1437 3.4105
R9271 GNDA_2.n1536 GNDA_2.n1456 3.4105
R9272 GNDA_2.n1536 GNDA_2.n1436 3.4105
R9273 GNDA_2.n1536 GNDA_2.n1457 3.4105
R9274 GNDA_2.n1536 GNDA_2.n1435 3.4105
R9275 GNDA_2.n1536 GNDA_2.n1458 3.4105
R9276 GNDA_2.n1536 GNDA_2.n1434 3.4105
R9277 GNDA_2.n1536 GNDA_2.n1459 3.4105
R9278 GNDA_2.n1536 GNDA_2.n1433 3.4105
R9279 GNDA_2.n1536 GNDA_2.n1460 3.4105
R9280 GNDA_2.n1536 GNDA_2.n1432 3.4105
R9281 GNDA_2.n1536 GNDA_2.n1461 3.4105
R9282 GNDA_2.n1536 GNDA_2.n1431 3.4105
R9283 GNDA_2.n1536 GNDA_2.n1462 3.4105
R9284 GNDA_2.n3441 GNDA_2.n1536 3.4105
R9285 GNDA_2.n1545 GNDA_2.n1467 3.4105
R9286 GNDA_2.n1467 GNDA_2.n1447 3.4105
R9287 GNDA_2.n1467 GNDA_2.n1445 3.4105
R9288 GNDA_2.n1467 GNDA_2.n1448 3.4105
R9289 GNDA_2.n1467 GNDA_2.n1444 3.4105
R9290 GNDA_2.n1467 GNDA_2.n1449 3.4105
R9291 GNDA_2.n1467 GNDA_2.n1443 3.4105
R9292 GNDA_2.n1467 GNDA_2.n1450 3.4105
R9293 GNDA_2.n1467 GNDA_2.n1442 3.4105
R9294 GNDA_2.n1467 GNDA_2.n1451 3.4105
R9295 GNDA_2.n1467 GNDA_2.n1441 3.4105
R9296 GNDA_2.n1467 GNDA_2.n1452 3.4105
R9297 GNDA_2.n1467 GNDA_2.n1440 3.4105
R9298 GNDA_2.n1467 GNDA_2.n1453 3.4105
R9299 GNDA_2.n1467 GNDA_2.n1439 3.4105
R9300 GNDA_2.n1467 GNDA_2.n1454 3.4105
R9301 GNDA_2.n1467 GNDA_2.n1438 3.4105
R9302 GNDA_2.n1467 GNDA_2.n1455 3.4105
R9303 GNDA_2.n1467 GNDA_2.n1437 3.4105
R9304 GNDA_2.n1467 GNDA_2.n1456 3.4105
R9305 GNDA_2.n1467 GNDA_2.n1436 3.4105
R9306 GNDA_2.n1467 GNDA_2.n1457 3.4105
R9307 GNDA_2.n1467 GNDA_2.n1435 3.4105
R9308 GNDA_2.n1467 GNDA_2.n1458 3.4105
R9309 GNDA_2.n1467 GNDA_2.n1434 3.4105
R9310 GNDA_2.n1467 GNDA_2.n1459 3.4105
R9311 GNDA_2.n1467 GNDA_2.n1433 3.4105
R9312 GNDA_2.n1467 GNDA_2.n1460 3.4105
R9313 GNDA_2.n1467 GNDA_2.n1432 3.4105
R9314 GNDA_2.n1467 GNDA_2.n1461 3.4105
R9315 GNDA_2.n1467 GNDA_2.n1431 3.4105
R9316 GNDA_2.n1467 GNDA_2.n1462 3.4105
R9317 GNDA_2.n3441 GNDA_2.n1467 3.4105
R9318 GNDA_2.n1545 GNDA_2.n1538 3.4105
R9319 GNDA_2.n1538 GNDA_2.n1447 3.4105
R9320 GNDA_2.n1538 GNDA_2.n1445 3.4105
R9321 GNDA_2.n1538 GNDA_2.n1448 3.4105
R9322 GNDA_2.n1538 GNDA_2.n1444 3.4105
R9323 GNDA_2.n1538 GNDA_2.n1449 3.4105
R9324 GNDA_2.n1538 GNDA_2.n1443 3.4105
R9325 GNDA_2.n1538 GNDA_2.n1450 3.4105
R9326 GNDA_2.n1538 GNDA_2.n1442 3.4105
R9327 GNDA_2.n1538 GNDA_2.n1451 3.4105
R9328 GNDA_2.n1538 GNDA_2.n1441 3.4105
R9329 GNDA_2.n1538 GNDA_2.n1452 3.4105
R9330 GNDA_2.n1538 GNDA_2.n1440 3.4105
R9331 GNDA_2.n1538 GNDA_2.n1453 3.4105
R9332 GNDA_2.n1538 GNDA_2.n1439 3.4105
R9333 GNDA_2.n1538 GNDA_2.n1454 3.4105
R9334 GNDA_2.n1538 GNDA_2.n1438 3.4105
R9335 GNDA_2.n1538 GNDA_2.n1455 3.4105
R9336 GNDA_2.n1538 GNDA_2.n1437 3.4105
R9337 GNDA_2.n1538 GNDA_2.n1456 3.4105
R9338 GNDA_2.n1538 GNDA_2.n1436 3.4105
R9339 GNDA_2.n1538 GNDA_2.n1457 3.4105
R9340 GNDA_2.n1538 GNDA_2.n1435 3.4105
R9341 GNDA_2.n1538 GNDA_2.n1458 3.4105
R9342 GNDA_2.n1538 GNDA_2.n1434 3.4105
R9343 GNDA_2.n1538 GNDA_2.n1459 3.4105
R9344 GNDA_2.n1538 GNDA_2.n1433 3.4105
R9345 GNDA_2.n1538 GNDA_2.n1460 3.4105
R9346 GNDA_2.n1538 GNDA_2.n1432 3.4105
R9347 GNDA_2.n1538 GNDA_2.n1461 3.4105
R9348 GNDA_2.n1538 GNDA_2.n1431 3.4105
R9349 GNDA_2.n1538 GNDA_2.n1462 3.4105
R9350 GNDA_2.n3441 GNDA_2.n1538 3.4105
R9351 GNDA_2.n1545 GNDA_2.n1466 3.4105
R9352 GNDA_2.n1466 GNDA_2.n1447 3.4105
R9353 GNDA_2.n1466 GNDA_2.n1445 3.4105
R9354 GNDA_2.n1466 GNDA_2.n1448 3.4105
R9355 GNDA_2.n1466 GNDA_2.n1444 3.4105
R9356 GNDA_2.n1466 GNDA_2.n1449 3.4105
R9357 GNDA_2.n1466 GNDA_2.n1443 3.4105
R9358 GNDA_2.n1466 GNDA_2.n1450 3.4105
R9359 GNDA_2.n1466 GNDA_2.n1442 3.4105
R9360 GNDA_2.n1466 GNDA_2.n1451 3.4105
R9361 GNDA_2.n1466 GNDA_2.n1441 3.4105
R9362 GNDA_2.n1466 GNDA_2.n1452 3.4105
R9363 GNDA_2.n1466 GNDA_2.n1440 3.4105
R9364 GNDA_2.n1466 GNDA_2.n1453 3.4105
R9365 GNDA_2.n1466 GNDA_2.n1439 3.4105
R9366 GNDA_2.n1466 GNDA_2.n1454 3.4105
R9367 GNDA_2.n1466 GNDA_2.n1438 3.4105
R9368 GNDA_2.n1466 GNDA_2.n1455 3.4105
R9369 GNDA_2.n1466 GNDA_2.n1437 3.4105
R9370 GNDA_2.n1466 GNDA_2.n1456 3.4105
R9371 GNDA_2.n1466 GNDA_2.n1436 3.4105
R9372 GNDA_2.n1466 GNDA_2.n1457 3.4105
R9373 GNDA_2.n1466 GNDA_2.n1435 3.4105
R9374 GNDA_2.n1466 GNDA_2.n1458 3.4105
R9375 GNDA_2.n1466 GNDA_2.n1434 3.4105
R9376 GNDA_2.n1466 GNDA_2.n1459 3.4105
R9377 GNDA_2.n1466 GNDA_2.n1433 3.4105
R9378 GNDA_2.n1466 GNDA_2.n1460 3.4105
R9379 GNDA_2.n1466 GNDA_2.n1432 3.4105
R9380 GNDA_2.n1466 GNDA_2.n1461 3.4105
R9381 GNDA_2.n1466 GNDA_2.n1431 3.4105
R9382 GNDA_2.n1466 GNDA_2.n1462 3.4105
R9383 GNDA_2.n3441 GNDA_2.n1466 3.4105
R9384 GNDA_2.n1545 GNDA_2.n1540 3.4105
R9385 GNDA_2.n1540 GNDA_2.n1447 3.4105
R9386 GNDA_2.n1540 GNDA_2.n1445 3.4105
R9387 GNDA_2.n1540 GNDA_2.n1448 3.4105
R9388 GNDA_2.n1540 GNDA_2.n1444 3.4105
R9389 GNDA_2.n1540 GNDA_2.n1449 3.4105
R9390 GNDA_2.n1540 GNDA_2.n1443 3.4105
R9391 GNDA_2.n1540 GNDA_2.n1450 3.4105
R9392 GNDA_2.n1540 GNDA_2.n1442 3.4105
R9393 GNDA_2.n1540 GNDA_2.n1451 3.4105
R9394 GNDA_2.n1540 GNDA_2.n1441 3.4105
R9395 GNDA_2.n1540 GNDA_2.n1452 3.4105
R9396 GNDA_2.n1540 GNDA_2.n1440 3.4105
R9397 GNDA_2.n1540 GNDA_2.n1453 3.4105
R9398 GNDA_2.n1540 GNDA_2.n1439 3.4105
R9399 GNDA_2.n1540 GNDA_2.n1454 3.4105
R9400 GNDA_2.n1540 GNDA_2.n1438 3.4105
R9401 GNDA_2.n1540 GNDA_2.n1455 3.4105
R9402 GNDA_2.n1540 GNDA_2.n1437 3.4105
R9403 GNDA_2.n1540 GNDA_2.n1456 3.4105
R9404 GNDA_2.n1540 GNDA_2.n1436 3.4105
R9405 GNDA_2.n1540 GNDA_2.n1457 3.4105
R9406 GNDA_2.n1540 GNDA_2.n1435 3.4105
R9407 GNDA_2.n1540 GNDA_2.n1458 3.4105
R9408 GNDA_2.n1540 GNDA_2.n1434 3.4105
R9409 GNDA_2.n1540 GNDA_2.n1459 3.4105
R9410 GNDA_2.n1540 GNDA_2.n1433 3.4105
R9411 GNDA_2.n1540 GNDA_2.n1460 3.4105
R9412 GNDA_2.n1540 GNDA_2.n1432 3.4105
R9413 GNDA_2.n1540 GNDA_2.n1461 3.4105
R9414 GNDA_2.n1540 GNDA_2.n1431 3.4105
R9415 GNDA_2.n1540 GNDA_2.n1462 3.4105
R9416 GNDA_2.n3441 GNDA_2.n1540 3.4105
R9417 GNDA_2.n1545 GNDA_2.n1465 3.4105
R9418 GNDA_2.n1465 GNDA_2.n1447 3.4105
R9419 GNDA_2.n1465 GNDA_2.n1445 3.4105
R9420 GNDA_2.n1465 GNDA_2.n1448 3.4105
R9421 GNDA_2.n1465 GNDA_2.n1444 3.4105
R9422 GNDA_2.n1465 GNDA_2.n1449 3.4105
R9423 GNDA_2.n1465 GNDA_2.n1443 3.4105
R9424 GNDA_2.n1465 GNDA_2.n1450 3.4105
R9425 GNDA_2.n1465 GNDA_2.n1442 3.4105
R9426 GNDA_2.n1465 GNDA_2.n1451 3.4105
R9427 GNDA_2.n1465 GNDA_2.n1441 3.4105
R9428 GNDA_2.n1465 GNDA_2.n1452 3.4105
R9429 GNDA_2.n1465 GNDA_2.n1440 3.4105
R9430 GNDA_2.n1465 GNDA_2.n1453 3.4105
R9431 GNDA_2.n1465 GNDA_2.n1439 3.4105
R9432 GNDA_2.n1465 GNDA_2.n1454 3.4105
R9433 GNDA_2.n1465 GNDA_2.n1438 3.4105
R9434 GNDA_2.n1465 GNDA_2.n1455 3.4105
R9435 GNDA_2.n1465 GNDA_2.n1437 3.4105
R9436 GNDA_2.n1465 GNDA_2.n1456 3.4105
R9437 GNDA_2.n1465 GNDA_2.n1436 3.4105
R9438 GNDA_2.n1465 GNDA_2.n1457 3.4105
R9439 GNDA_2.n1465 GNDA_2.n1435 3.4105
R9440 GNDA_2.n1465 GNDA_2.n1458 3.4105
R9441 GNDA_2.n1465 GNDA_2.n1434 3.4105
R9442 GNDA_2.n1465 GNDA_2.n1459 3.4105
R9443 GNDA_2.n1465 GNDA_2.n1433 3.4105
R9444 GNDA_2.n1465 GNDA_2.n1460 3.4105
R9445 GNDA_2.n1465 GNDA_2.n1432 3.4105
R9446 GNDA_2.n1465 GNDA_2.n1461 3.4105
R9447 GNDA_2.n1465 GNDA_2.n1431 3.4105
R9448 GNDA_2.n1465 GNDA_2.n1462 3.4105
R9449 GNDA_2.n3441 GNDA_2.n1465 3.4105
R9450 GNDA_2.n1545 GNDA_2.n1542 3.4105
R9451 GNDA_2.n1542 GNDA_2.n1447 3.4105
R9452 GNDA_2.n1542 GNDA_2.n1445 3.4105
R9453 GNDA_2.n1542 GNDA_2.n1448 3.4105
R9454 GNDA_2.n1542 GNDA_2.n1444 3.4105
R9455 GNDA_2.n1542 GNDA_2.n1449 3.4105
R9456 GNDA_2.n1542 GNDA_2.n1443 3.4105
R9457 GNDA_2.n1542 GNDA_2.n1450 3.4105
R9458 GNDA_2.n1542 GNDA_2.n1442 3.4105
R9459 GNDA_2.n1542 GNDA_2.n1451 3.4105
R9460 GNDA_2.n1542 GNDA_2.n1441 3.4105
R9461 GNDA_2.n1542 GNDA_2.n1452 3.4105
R9462 GNDA_2.n1542 GNDA_2.n1440 3.4105
R9463 GNDA_2.n1542 GNDA_2.n1453 3.4105
R9464 GNDA_2.n1542 GNDA_2.n1439 3.4105
R9465 GNDA_2.n1542 GNDA_2.n1454 3.4105
R9466 GNDA_2.n1542 GNDA_2.n1438 3.4105
R9467 GNDA_2.n1542 GNDA_2.n1455 3.4105
R9468 GNDA_2.n1542 GNDA_2.n1437 3.4105
R9469 GNDA_2.n1542 GNDA_2.n1456 3.4105
R9470 GNDA_2.n1542 GNDA_2.n1436 3.4105
R9471 GNDA_2.n1542 GNDA_2.n1457 3.4105
R9472 GNDA_2.n1542 GNDA_2.n1435 3.4105
R9473 GNDA_2.n1542 GNDA_2.n1458 3.4105
R9474 GNDA_2.n1542 GNDA_2.n1434 3.4105
R9475 GNDA_2.n1542 GNDA_2.n1459 3.4105
R9476 GNDA_2.n1542 GNDA_2.n1433 3.4105
R9477 GNDA_2.n1542 GNDA_2.n1460 3.4105
R9478 GNDA_2.n1542 GNDA_2.n1432 3.4105
R9479 GNDA_2.n1542 GNDA_2.n1461 3.4105
R9480 GNDA_2.n1542 GNDA_2.n1431 3.4105
R9481 GNDA_2.n1542 GNDA_2.n1462 3.4105
R9482 GNDA_2.n3441 GNDA_2.n1542 3.4105
R9483 GNDA_2.n1545 GNDA_2.n1464 3.4105
R9484 GNDA_2.n1464 GNDA_2.n1447 3.4105
R9485 GNDA_2.n1464 GNDA_2.n1445 3.4105
R9486 GNDA_2.n1464 GNDA_2.n1448 3.4105
R9487 GNDA_2.n1464 GNDA_2.n1444 3.4105
R9488 GNDA_2.n1464 GNDA_2.n1449 3.4105
R9489 GNDA_2.n1464 GNDA_2.n1443 3.4105
R9490 GNDA_2.n1464 GNDA_2.n1450 3.4105
R9491 GNDA_2.n1464 GNDA_2.n1442 3.4105
R9492 GNDA_2.n1464 GNDA_2.n1451 3.4105
R9493 GNDA_2.n1464 GNDA_2.n1441 3.4105
R9494 GNDA_2.n1464 GNDA_2.n1452 3.4105
R9495 GNDA_2.n1464 GNDA_2.n1440 3.4105
R9496 GNDA_2.n1464 GNDA_2.n1453 3.4105
R9497 GNDA_2.n1464 GNDA_2.n1439 3.4105
R9498 GNDA_2.n1464 GNDA_2.n1454 3.4105
R9499 GNDA_2.n1464 GNDA_2.n1438 3.4105
R9500 GNDA_2.n1464 GNDA_2.n1455 3.4105
R9501 GNDA_2.n1464 GNDA_2.n1437 3.4105
R9502 GNDA_2.n1464 GNDA_2.n1456 3.4105
R9503 GNDA_2.n1464 GNDA_2.n1436 3.4105
R9504 GNDA_2.n1464 GNDA_2.n1457 3.4105
R9505 GNDA_2.n1464 GNDA_2.n1435 3.4105
R9506 GNDA_2.n1464 GNDA_2.n1458 3.4105
R9507 GNDA_2.n1464 GNDA_2.n1434 3.4105
R9508 GNDA_2.n1464 GNDA_2.n1459 3.4105
R9509 GNDA_2.n1464 GNDA_2.n1433 3.4105
R9510 GNDA_2.n1464 GNDA_2.n1460 3.4105
R9511 GNDA_2.n1464 GNDA_2.n1432 3.4105
R9512 GNDA_2.n1464 GNDA_2.n1461 3.4105
R9513 GNDA_2.n1464 GNDA_2.n1431 3.4105
R9514 GNDA_2.n1464 GNDA_2.n1462 3.4105
R9515 GNDA_2.n3441 GNDA_2.n1464 3.4105
R9516 GNDA_2.n3440 GNDA_2.n1545 3.4105
R9517 GNDA_2.n3440 GNDA_2.n1447 3.4105
R9518 GNDA_2.n3440 GNDA_2.n1445 3.4105
R9519 GNDA_2.n3440 GNDA_2.n1448 3.4105
R9520 GNDA_2.n3440 GNDA_2.n1444 3.4105
R9521 GNDA_2.n3440 GNDA_2.n1449 3.4105
R9522 GNDA_2.n3440 GNDA_2.n1443 3.4105
R9523 GNDA_2.n3440 GNDA_2.n1450 3.4105
R9524 GNDA_2.n3440 GNDA_2.n1442 3.4105
R9525 GNDA_2.n3440 GNDA_2.n1451 3.4105
R9526 GNDA_2.n3440 GNDA_2.n1441 3.4105
R9527 GNDA_2.n3440 GNDA_2.n1452 3.4105
R9528 GNDA_2.n3440 GNDA_2.n1440 3.4105
R9529 GNDA_2.n3440 GNDA_2.n1453 3.4105
R9530 GNDA_2.n3440 GNDA_2.n1439 3.4105
R9531 GNDA_2.n3440 GNDA_2.n1454 3.4105
R9532 GNDA_2.n3440 GNDA_2.n1438 3.4105
R9533 GNDA_2.n3440 GNDA_2.n1455 3.4105
R9534 GNDA_2.n3440 GNDA_2.n1437 3.4105
R9535 GNDA_2.n3440 GNDA_2.n1456 3.4105
R9536 GNDA_2.n3440 GNDA_2.n1436 3.4105
R9537 GNDA_2.n3440 GNDA_2.n1457 3.4105
R9538 GNDA_2.n3440 GNDA_2.n1435 3.4105
R9539 GNDA_2.n3440 GNDA_2.n1458 3.4105
R9540 GNDA_2.n3440 GNDA_2.n1434 3.4105
R9541 GNDA_2.n3440 GNDA_2.n1459 3.4105
R9542 GNDA_2.n3440 GNDA_2.n1433 3.4105
R9543 GNDA_2.n3440 GNDA_2.n1460 3.4105
R9544 GNDA_2.n3440 GNDA_2.n1432 3.4105
R9545 GNDA_2.n3440 GNDA_2.n1461 3.4105
R9546 GNDA_2.n3440 GNDA_2.n1431 3.4105
R9547 GNDA_2.n3440 GNDA_2.n1462 3.4105
R9548 GNDA_2.n3441 GNDA_2.n3440 3.4105
R9549 GNDA_2.n1545 GNDA_2.n1463 3.4105
R9550 GNDA_2.n1463 GNDA_2.n1447 3.4105
R9551 GNDA_2.n1463 GNDA_2.n1445 3.4105
R9552 GNDA_2.n1463 GNDA_2.n1448 3.4105
R9553 GNDA_2.n1463 GNDA_2.n1444 3.4105
R9554 GNDA_2.n1463 GNDA_2.n1449 3.4105
R9555 GNDA_2.n1463 GNDA_2.n1443 3.4105
R9556 GNDA_2.n1463 GNDA_2.n1450 3.4105
R9557 GNDA_2.n1463 GNDA_2.n1442 3.4105
R9558 GNDA_2.n1463 GNDA_2.n1451 3.4105
R9559 GNDA_2.n1463 GNDA_2.n1441 3.4105
R9560 GNDA_2.n1463 GNDA_2.n1452 3.4105
R9561 GNDA_2.n1463 GNDA_2.n1440 3.4105
R9562 GNDA_2.n1463 GNDA_2.n1453 3.4105
R9563 GNDA_2.n1463 GNDA_2.n1439 3.4105
R9564 GNDA_2.n1463 GNDA_2.n1454 3.4105
R9565 GNDA_2.n1463 GNDA_2.n1438 3.4105
R9566 GNDA_2.n1463 GNDA_2.n1455 3.4105
R9567 GNDA_2.n1463 GNDA_2.n1437 3.4105
R9568 GNDA_2.n1463 GNDA_2.n1456 3.4105
R9569 GNDA_2.n1463 GNDA_2.n1436 3.4105
R9570 GNDA_2.n1463 GNDA_2.n1457 3.4105
R9571 GNDA_2.n1463 GNDA_2.n1435 3.4105
R9572 GNDA_2.n1463 GNDA_2.n1458 3.4105
R9573 GNDA_2.n1463 GNDA_2.n1434 3.4105
R9574 GNDA_2.n1463 GNDA_2.n1459 3.4105
R9575 GNDA_2.n1463 GNDA_2.n1433 3.4105
R9576 GNDA_2.n1463 GNDA_2.n1460 3.4105
R9577 GNDA_2.n1463 GNDA_2.n1432 3.4105
R9578 GNDA_2.n1463 GNDA_2.n1461 3.4105
R9579 GNDA_2.n1463 GNDA_2.n1431 3.4105
R9580 GNDA_2.n1463 GNDA_2.n1462 3.4105
R9581 GNDA_2.n3441 GNDA_2.n1463 3.4105
R9582 GNDA_2.n3442 GNDA_2.n1447 3.4105
R9583 GNDA_2.n3442 GNDA_2.n1445 3.4105
R9584 GNDA_2.n3442 GNDA_2.n1448 3.4105
R9585 GNDA_2.n3442 GNDA_2.n1444 3.4105
R9586 GNDA_2.n3442 GNDA_2.n1449 3.4105
R9587 GNDA_2.n3442 GNDA_2.n1443 3.4105
R9588 GNDA_2.n3442 GNDA_2.n1450 3.4105
R9589 GNDA_2.n3442 GNDA_2.n1442 3.4105
R9590 GNDA_2.n3442 GNDA_2.n1451 3.4105
R9591 GNDA_2.n3442 GNDA_2.n1441 3.4105
R9592 GNDA_2.n3442 GNDA_2.n1452 3.4105
R9593 GNDA_2.n3442 GNDA_2.n1440 3.4105
R9594 GNDA_2.n3442 GNDA_2.n1453 3.4105
R9595 GNDA_2.n3442 GNDA_2.n1439 3.4105
R9596 GNDA_2.n3442 GNDA_2.n1454 3.4105
R9597 GNDA_2.n3442 GNDA_2.n1438 3.4105
R9598 GNDA_2.n3442 GNDA_2.n1455 3.4105
R9599 GNDA_2.n3442 GNDA_2.n1437 3.4105
R9600 GNDA_2.n3442 GNDA_2.n1456 3.4105
R9601 GNDA_2.n3442 GNDA_2.n1436 3.4105
R9602 GNDA_2.n3442 GNDA_2.n1457 3.4105
R9603 GNDA_2.n3442 GNDA_2.n1435 3.4105
R9604 GNDA_2.n3442 GNDA_2.n1458 3.4105
R9605 GNDA_2.n3442 GNDA_2.n1434 3.4105
R9606 GNDA_2.n3442 GNDA_2.n1459 3.4105
R9607 GNDA_2.n3442 GNDA_2.n1433 3.4105
R9608 GNDA_2.n3442 GNDA_2.n1460 3.4105
R9609 GNDA_2.n3442 GNDA_2.n1432 3.4105
R9610 GNDA_2.n3442 GNDA_2.n1461 3.4105
R9611 GNDA_2.n3442 GNDA_2.n1431 3.4105
R9612 GNDA_2.n3442 GNDA_2.n1462 3.4105
R9613 GNDA_2.n3442 GNDA_2.n3441 3.4105
R9614 GNDA_2.n3492 GNDA_2.n3459 3.4105
R9615 GNDA_2.n3512 GNDA_2.n3459 3.4105
R9616 GNDA_2.n3512 GNDA_2.n1428 3.4105
R9617 GNDA_2.n3492 GNDA_2.n3461 3.4105
R9618 GNDA_2.n3461 GNDA_2.n1381 3.4105
R9619 GNDA_2.n3461 GNDA_2.n1379 3.4105
R9620 GNDA_2.n3461 GNDA_2.n1382 3.4105
R9621 GNDA_2.n3461 GNDA_2.n1378 3.4105
R9622 GNDA_2.n3461 GNDA_2.n1383 3.4105
R9623 GNDA_2.n3461 GNDA_2.n1377 3.4105
R9624 GNDA_2.n3461 GNDA_2.n1384 3.4105
R9625 GNDA_2.n3461 GNDA_2.n1376 3.4105
R9626 GNDA_2.n3461 GNDA_2.n1385 3.4105
R9627 GNDA_2.n3461 GNDA_2.n1375 3.4105
R9628 GNDA_2.n3461 GNDA_2.n1386 3.4105
R9629 GNDA_2.n3461 GNDA_2.n1374 3.4105
R9630 GNDA_2.n3461 GNDA_2.n1387 3.4105
R9631 GNDA_2.n3461 GNDA_2.n1373 3.4105
R9632 GNDA_2.n3461 GNDA_2.n1388 3.4105
R9633 GNDA_2.n3461 GNDA_2.n1372 3.4105
R9634 GNDA_2.n3461 GNDA_2.n1389 3.4105
R9635 GNDA_2.n3461 GNDA_2.n1371 3.4105
R9636 GNDA_2.n3461 GNDA_2.n1390 3.4105
R9637 GNDA_2.n3461 GNDA_2.n1370 3.4105
R9638 GNDA_2.n3461 GNDA_2.n1391 3.4105
R9639 GNDA_2.n3461 GNDA_2.n1369 3.4105
R9640 GNDA_2.n3461 GNDA_2.n1392 3.4105
R9641 GNDA_2.n3461 GNDA_2.n1368 3.4105
R9642 GNDA_2.n3461 GNDA_2.n1393 3.4105
R9643 GNDA_2.n3461 GNDA_2.n1367 3.4105
R9644 GNDA_2.n3461 GNDA_2.n1394 3.4105
R9645 GNDA_2.n3461 GNDA_2.n1366 3.4105
R9646 GNDA_2.n3461 GNDA_2.n1395 3.4105
R9647 GNDA_2.n3461 GNDA_2.n1365 3.4105
R9648 GNDA_2.n3461 GNDA_2.n1396 3.4105
R9649 GNDA_2.n3512 GNDA_2.n3461 3.4105
R9650 GNDA_2.n3492 GNDA_2.n1412 3.4105
R9651 GNDA_2.n1412 GNDA_2.n1381 3.4105
R9652 GNDA_2.n1412 GNDA_2.n1379 3.4105
R9653 GNDA_2.n1412 GNDA_2.n1382 3.4105
R9654 GNDA_2.n1412 GNDA_2.n1378 3.4105
R9655 GNDA_2.n1412 GNDA_2.n1383 3.4105
R9656 GNDA_2.n1412 GNDA_2.n1377 3.4105
R9657 GNDA_2.n1412 GNDA_2.n1384 3.4105
R9658 GNDA_2.n1412 GNDA_2.n1376 3.4105
R9659 GNDA_2.n1412 GNDA_2.n1385 3.4105
R9660 GNDA_2.n1412 GNDA_2.n1375 3.4105
R9661 GNDA_2.n1412 GNDA_2.n1386 3.4105
R9662 GNDA_2.n1412 GNDA_2.n1374 3.4105
R9663 GNDA_2.n1412 GNDA_2.n1387 3.4105
R9664 GNDA_2.n1412 GNDA_2.n1373 3.4105
R9665 GNDA_2.n1412 GNDA_2.n1388 3.4105
R9666 GNDA_2.n1412 GNDA_2.n1372 3.4105
R9667 GNDA_2.n1412 GNDA_2.n1389 3.4105
R9668 GNDA_2.n1412 GNDA_2.n1371 3.4105
R9669 GNDA_2.n1412 GNDA_2.n1390 3.4105
R9670 GNDA_2.n1412 GNDA_2.n1370 3.4105
R9671 GNDA_2.n1412 GNDA_2.n1391 3.4105
R9672 GNDA_2.n1412 GNDA_2.n1369 3.4105
R9673 GNDA_2.n1412 GNDA_2.n1392 3.4105
R9674 GNDA_2.n1412 GNDA_2.n1368 3.4105
R9675 GNDA_2.n1412 GNDA_2.n1393 3.4105
R9676 GNDA_2.n1412 GNDA_2.n1367 3.4105
R9677 GNDA_2.n1412 GNDA_2.n1394 3.4105
R9678 GNDA_2.n1412 GNDA_2.n1366 3.4105
R9679 GNDA_2.n1412 GNDA_2.n1395 3.4105
R9680 GNDA_2.n1412 GNDA_2.n1365 3.4105
R9681 GNDA_2.n1412 GNDA_2.n1396 3.4105
R9682 GNDA_2.n3512 GNDA_2.n1412 3.4105
R9683 GNDA_2.n3492 GNDA_2.n3463 3.4105
R9684 GNDA_2.n3463 GNDA_2.n1381 3.4105
R9685 GNDA_2.n3463 GNDA_2.n1379 3.4105
R9686 GNDA_2.n3463 GNDA_2.n1382 3.4105
R9687 GNDA_2.n3463 GNDA_2.n1378 3.4105
R9688 GNDA_2.n3463 GNDA_2.n1383 3.4105
R9689 GNDA_2.n3463 GNDA_2.n1377 3.4105
R9690 GNDA_2.n3463 GNDA_2.n1384 3.4105
R9691 GNDA_2.n3463 GNDA_2.n1376 3.4105
R9692 GNDA_2.n3463 GNDA_2.n1385 3.4105
R9693 GNDA_2.n3463 GNDA_2.n1375 3.4105
R9694 GNDA_2.n3463 GNDA_2.n1386 3.4105
R9695 GNDA_2.n3463 GNDA_2.n1374 3.4105
R9696 GNDA_2.n3463 GNDA_2.n1387 3.4105
R9697 GNDA_2.n3463 GNDA_2.n1373 3.4105
R9698 GNDA_2.n3463 GNDA_2.n1388 3.4105
R9699 GNDA_2.n3463 GNDA_2.n1372 3.4105
R9700 GNDA_2.n3463 GNDA_2.n1389 3.4105
R9701 GNDA_2.n3463 GNDA_2.n1371 3.4105
R9702 GNDA_2.n3463 GNDA_2.n1390 3.4105
R9703 GNDA_2.n3463 GNDA_2.n1370 3.4105
R9704 GNDA_2.n3463 GNDA_2.n1391 3.4105
R9705 GNDA_2.n3463 GNDA_2.n1369 3.4105
R9706 GNDA_2.n3463 GNDA_2.n1392 3.4105
R9707 GNDA_2.n3463 GNDA_2.n1368 3.4105
R9708 GNDA_2.n3463 GNDA_2.n1393 3.4105
R9709 GNDA_2.n3463 GNDA_2.n1367 3.4105
R9710 GNDA_2.n3463 GNDA_2.n1394 3.4105
R9711 GNDA_2.n3463 GNDA_2.n1366 3.4105
R9712 GNDA_2.n3463 GNDA_2.n1395 3.4105
R9713 GNDA_2.n3463 GNDA_2.n1365 3.4105
R9714 GNDA_2.n3463 GNDA_2.n1396 3.4105
R9715 GNDA_2.n3512 GNDA_2.n3463 3.4105
R9716 GNDA_2.n3492 GNDA_2.n1411 3.4105
R9717 GNDA_2.n1411 GNDA_2.n1381 3.4105
R9718 GNDA_2.n1411 GNDA_2.n1379 3.4105
R9719 GNDA_2.n1411 GNDA_2.n1382 3.4105
R9720 GNDA_2.n1411 GNDA_2.n1378 3.4105
R9721 GNDA_2.n1411 GNDA_2.n1383 3.4105
R9722 GNDA_2.n1411 GNDA_2.n1377 3.4105
R9723 GNDA_2.n1411 GNDA_2.n1384 3.4105
R9724 GNDA_2.n1411 GNDA_2.n1376 3.4105
R9725 GNDA_2.n1411 GNDA_2.n1385 3.4105
R9726 GNDA_2.n1411 GNDA_2.n1375 3.4105
R9727 GNDA_2.n1411 GNDA_2.n1386 3.4105
R9728 GNDA_2.n1411 GNDA_2.n1374 3.4105
R9729 GNDA_2.n1411 GNDA_2.n1387 3.4105
R9730 GNDA_2.n1411 GNDA_2.n1373 3.4105
R9731 GNDA_2.n1411 GNDA_2.n1388 3.4105
R9732 GNDA_2.n1411 GNDA_2.n1372 3.4105
R9733 GNDA_2.n1411 GNDA_2.n1389 3.4105
R9734 GNDA_2.n1411 GNDA_2.n1371 3.4105
R9735 GNDA_2.n1411 GNDA_2.n1390 3.4105
R9736 GNDA_2.n1411 GNDA_2.n1370 3.4105
R9737 GNDA_2.n1411 GNDA_2.n1391 3.4105
R9738 GNDA_2.n1411 GNDA_2.n1369 3.4105
R9739 GNDA_2.n1411 GNDA_2.n1392 3.4105
R9740 GNDA_2.n1411 GNDA_2.n1368 3.4105
R9741 GNDA_2.n1411 GNDA_2.n1393 3.4105
R9742 GNDA_2.n1411 GNDA_2.n1367 3.4105
R9743 GNDA_2.n1411 GNDA_2.n1394 3.4105
R9744 GNDA_2.n1411 GNDA_2.n1366 3.4105
R9745 GNDA_2.n1411 GNDA_2.n1395 3.4105
R9746 GNDA_2.n1411 GNDA_2.n1365 3.4105
R9747 GNDA_2.n1411 GNDA_2.n1396 3.4105
R9748 GNDA_2.n3512 GNDA_2.n1411 3.4105
R9749 GNDA_2.n3492 GNDA_2.n3465 3.4105
R9750 GNDA_2.n3465 GNDA_2.n1381 3.4105
R9751 GNDA_2.n3465 GNDA_2.n1379 3.4105
R9752 GNDA_2.n3465 GNDA_2.n1382 3.4105
R9753 GNDA_2.n3465 GNDA_2.n1378 3.4105
R9754 GNDA_2.n3465 GNDA_2.n1383 3.4105
R9755 GNDA_2.n3465 GNDA_2.n1377 3.4105
R9756 GNDA_2.n3465 GNDA_2.n1384 3.4105
R9757 GNDA_2.n3465 GNDA_2.n1376 3.4105
R9758 GNDA_2.n3465 GNDA_2.n1385 3.4105
R9759 GNDA_2.n3465 GNDA_2.n1375 3.4105
R9760 GNDA_2.n3465 GNDA_2.n1386 3.4105
R9761 GNDA_2.n3465 GNDA_2.n1374 3.4105
R9762 GNDA_2.n3465 GNDA_2.n1387 3.4105
R9763 GNDA_2.n3465 GNDA_2.n1373 3.4105
R9764 GNDA_2.n3465 GNDA_2.n1388 3.4105
R9765 GNDA_2.n3465 GNDA_2.n1372 3.4105
R9766 GNDA_2.n3465 GNDA_2.n1389 3.4105
R9767 GNDA_2.n3465 GNDA_2.n1371 3.4105
R9768 GNDA_2.n3465 GNDA_2.n1390 3.4105
R9769 GNDA_2.n3465 GNDA_2.n1370 3.4105
R9770 GNDA_2.n3465 GNDA_2.n1391 3.4105
R9771 GNDA_2.n3465 GNDA_2.n1369 3.4105
R9772 GNDA_2.n3465 GNDA_2.n1392 3.4105
R9773 GNDA_2.n3465 GNDA_2.n1368 3.4105
R9774 GNDA_2.n3465 GNDA_2.n1393 3.4105
R9775 GNDA_2.n3465 GNDA_2.n1367 3.4105
R9776 GNDA_2.n3465 GNDA_2.n1394 3.4105
R9777 GNDA_2.n3465 GNDA_2.n1366 3.4105
R9778 GNDA_2.n3465 GNDA_2.n1395 3.4105
R9779 GNDA_2.n3465 GNDA_2.n1365 3.4105
R9780 GNDA_2.n3465 GNDA_2.n1396 3.4105
R9781 GNDA_2.n3512 GNDA_2.n3465 3.4105
R9782 GNDA_2.n3492 GNDA_2.n1410 3.4105
R9783 GNDA_2.n1410 GNDA_2.n1381 3.4105
R9784 GNDA_2.n1410 GNDA_2.n1379 3.4105
R9785 GNDA_2.n1410 GNDA_2.n1382 3.4105
R9786 GNDA_2.n1410 GNDA_2.n1378 3.4105
R9787 GNDA_2.n1410 GNDA_2.n1383 3.4105
R9788 GNDA_2.n1410 GNDA_2.n1377 3.4105
R9789 GNDA_2.n1410 GNDA_2.n1384 3.4105
R9790 GNDA_2.n1410 GNDA_2.n1376 3.4105
R9791 GNDA_2.n1410 GNDA_2.n1385 3.4105
R9792 GNDA_2.n1410 GNDA_2.n1375 3.4105
R9793 GNDA_2.n1410 GNDA_2.n1386 3.4105
R9794 GNDA_2.n1410 GNDA_2.n1374 3.4105
R9795 GNDA_2.n1410 GNDA_2.n1387 3.4105
R9796 GNDA_2.n1410 GNDA_2.n1373 3.4105
R9797 GNDA_2.n1410 GNDA_2.n1388 3.4105
R9798 GNDA_2.n1410 GNDA_2.n1372 3.4105
R9799 GNDA_2.n1410 GNDA_2.n1389 3.4105
R9800 GNDA_2.n1410 GNDA_2.n1371 3.4105
R9801 GNDA_2.n1410 GNDA_2.n1390 3.4105
R9802 GNDA_2.n1410 GNDA_2.n1370 3.4105
R9803 GNDA_2.n1410 GNDA_2.n1391 3.4105
R9804 GNDA_2.n1410 GNDA_2.n1369 3.4105
R9805 GNDA_2.n1410 GNDA_2.n1392 3.4105
R9806 GNDA_2.n1410 GNDA_2.n1368 3.4105
R9807 GNDA_2.n1410 GNDA_2.n1393 3.4105
R9808 GNDA_2.n1410 GNDA_2.n1367 3.4105
R9809 GNDA_2.n1410 GNDA_2.n1394 3.4105
R9810 GNDA_2.n1410 GNDA_2.n1366 3.4105
R9811 GNDA_2.n1410 GNDA_2.n1395 3.4105
R9812 GNDA_2.n1410 GNDA_2.n1365 3.4105
R9813 GNDA_2.n1410 GNDA_2.n1396 3.4105
R9814 GNDA_2.n3512 GNDA_2.n1410 3.4105
R9815 GNDA_2.n3492 GNDA_2.n3467 3.4105
R9816 GNDA_2.n3467 GNDA_2.n1381 3.4105
R9817 GNDA_2.n3467 GNDA_2.n1379 3.4105
R9818 GNDA_2.n3467 GNDA_2.n1382 3.4105
R9819 GNDA_2.n3467 GNDA_2.n1378 3.4105
R9820 GNDA_2.n3467 GNDA_2.n1383 3.4105
R9821 GNDA_2.n3467 GNDA_2.n1377 3.4105
R9822 GNDA_2.n3467 GNDA_2.n1384 3.4105
R9823 GNDA_2.n3467 GNDA_2.n1376 3.4105
R9824 GNDA_2.n3467 GNDA_2.n1385 3.4105
R9825 GNDA_2.n3467 GNDA_2.n1375 3.4105
R9826 GNDA_2.n3467 GNDA_2.n1386 3.4105
R9827 GNDA_2.n3467 GNDA_2.n1374 3.4105
R9828 GNDA_2.n3467 GNDA_2.n1387 3.4105
R9829 GNDA_2.n3467 GNDA_2.n1373 3.4105
R9830 GNDA_2.n3467 GNDA_2.n1388 3.4105
R9831 GNDA_2.n3467 GNDA_2.n1372 3.4105
R9832 GNDA_2.n3467 GNDA_2.n1389 3.4105
R9833 GNDA_2.n3467 GNDA_2.n1371 3.4105
R9834 GNDA_2.n3467 GNDA_2.n1390 3.4105
R9835 GNDA_2.n3467 GNDA_2.n1370 3.4105
R9836 GNDA_2.n3467 GNDA_2.n1391 3.4105
R9837 GNDA_2.n3467 GNDA_2.n1369 3.4105
R9838 GNDA_2.n3467 GNDA_2.n1392 3.4105
R9839 GNDA_2.n3467 GNDA_2.n1368 3.4105
R9840 GNDA_2.n3467 GNDA_2.n1393 3.4105
R9841 GNDA_2.n3467 GNDA_2.n1367 3.4105
R9842 GNDA_2.n3467 GNDA_2.n1394 3.4105
R9843 GNDA_2.n3467 GNDA_2.n1366 3.4105
R9844 GNDA_2.n3467 GNDA_2.n1395 3.4105
R9845 GNDA_2.n3467 GNDA_2.n1365 3.4105
R9846 GNDA_2.n3467 GNDA_2.n1396 3.4105
R9847 GNDA_2.n3512 GNDA_2.n3467 3.4105
R9848 GNDA_2.n3492 GNDA_2.n1409 3.4105
R9849 GNDA_2.n1409 GNDA_2.n1381 3.4105
R9850 GNDA_2.n1409 GNDA_2.n1379 3.4105
R9851 GNDA_2.n1409 GNDA_2.n1382 3.4105
R9852 GNDA_2.n1409 GNDA_2.n1378 3.4105
R9853 GNDA_2.n1409 GNDA_2.n1383 3.4105
R9854 GNDA_2.n1409 GNDA_2.n1377 3.4105
R9855 GNDA_2.n1409 GNDA_2.n1384 3.4105
R9856 GNDA_2.n1409 GNDA_2.n1376 3.4105
R9857 GNDA_2.n1409 GNDA_2.n1385 3.4105
R9858 GNDA_2.n1409 GNDA_2.n1375 3.4105
R9859 GNDA_2.n1409 GNDA_2.n1386 3.4105
R9860 GNDA_2.n1409 GNDA_2.n1374 3.4105
R9861 GNDA_2.n1409 GNDA_2.n1387 3.4105
R9862 GNDA_2.n1409 GNDA_2.n1373 3.4105
R9863 GNDA_2.n1409 GNDA_2.n1388 3.4105
R9864 GNDA_2.n1409 GNDA_2.n1372 3.4105
R9865 GNDA_2.n1409 GNDA_2.n1389 3.4105
R9866 GNDA_2.n1409 GNDA_2.n1371 3.4105
R9867 GNDA_2.n1409 GNDA_2.n1390 3.4105
R9868 GNDA_2.n1409 GNDA_2.n1370 3.4105
R9869 GNDA_2.n1409 GNDA_2.n1391 3.4105
R9870 GNDA_2.n1409 GNDA_2.n1369 3.4105
R9871 GNDA_2.n1409 GNDA_2.n1392 3.4105
R9872 GNDA_2.n1409 GNDA_2.n1368 3.4105
R9873 GNDA_2.n1409 GNDA_2.n1393 3.4105
R9874 GNDA_2.n1409 GNDA_2.n1367 3.4105
R9875 GNDA_2.n1409 GNDA_2.n1394 3.4105
R9876 GNDA_2.n1409 GNDA_2.n1366 3.4105
R9877 GNDA_2.n1409 GNDA_2.n1395 3.4105
R9878 GNDA_2.n1409 GNDA_2.n1365 3.4105
R9879 GNDA_2.n1409 GNDA_2.n1396 3.4105
R9880 GNDA_2.n3512 GNDA_2.n1409 3.4105
R9881 GNDA_2.n3492 GNDA_2.n3469 3.4105
R9882 GNDA_2.n3469 GNDA_2.n1381 3.4105
R9883 GNDA_2.n3469 GNDA_2.n1379 3.4105
R9884 GNDA_2.n3469 GNDA_2.n1382 3.4105
R9885 GNDA_2.n3469 GNDA_2.n1378 3.4105
R9886 GNDA_2.n3469 GNDA_2.n1383 3.4105
R9887 GNDA_2.n3469 GNDA_2.n1377 3.4105
R9888 GNDA_2.n3469 GNDA_2.n1384 3.4105
R9889 GNDA_2.n3469 GNDA_2.n1376 3.4105
R9890 GNDA_2.n3469 GNDA_2.n1385 3.4105
R9891 GNDA_2.n3469 GNDA_2.n1375 3.4105
R9892 GNDA_2.n3469 GNDA_2.n1386 3.4105
R9893 GNDA_2.n3469 GNDA_2.n1374 3.4105
R9894 GNDA_2.n3469 GNDA_2.n1387 3.4105
R9895 GNDA_2.n3469 GNDA_2.n1373 3.4105
R9896 GNDA_2.n3469 GNDA_2.n1388 3.4105
R9897 GNDA_2.n3469 GNDA_2.n1372 3.4105
R9898 GNDA_2.n3469 GNDA_2.n1389 3.4105
R9899 GNDA_2.n3469 GNDA_2.n1371 3.4105
R9900 GNDA_2.n3469 GNDA_2.n1390 3.4105
R9901 GNDA_2.n3469 GNDA_2.n1370 3.4105
R9902 GNDA_2.n3469 GNDA_2.n1391 3.4105
R9903 GNDA_2.n3469 GNDA_2.n1369 3.4105
R9904 GNDA_2.n3469 GNDA_2.n1392 3.4105
R9905 GNDA_2.n3469 GNDA_2.n1368 3.4105
R9906 GNDA_2.n3469 GNDA_2.n1393 3.4105
R9907 GNDA_2.n3469 GNDA_2.n1367 3.4105
R9908 GNDA_2.n3469 GNDA_2.n1394 3.4105
R9909 GNDA_2.n3469 GNDA_2.n1366 3.4105
R9910 GNDA_2.n3469 GNDA_2.n1395 3.4105
R9911 GNDA_2.n3469 GNDA_2.n1365 3.4105
R9912 GNDA_2.n3469 GNDA_2.n1396 3.4105
R9913 GNDA_2.n3512 GNDA_2.n3469 3.4105
R9914 GNDA_2.n3492 GNDA_2.n1408 3.4105
R9915 GNDA_2.n1408 GNDA_2.n1381 3.4105
R9916 GNDA_2.n1408 GNDA_2.n1379 3.4105
R9917 GNDA_2.n1408 GNDA_2.n1382 3.4105
R9918 GNDA_2.n1408 GNDA_2.n1378 3.4105
R9919 GNDA_2.n1408 GNDA_2.n1383 3.4105
R9920 GNDA_2.n1408 GNDA_2.n1377 3.4105
R9921 GNDA_2.n1408 GNDA_2.n1384 3.4105
R9922 GNDA_2.n1408 GNDA_2.n1376 3.4105
R9923 GNDA_2.n1408 GNDA_2.n1385 3.4105
R9924 GNDA_2.n1408 GNDA_2.n1375 3.4105
R9925 GNDA_2.n1408 GNDA_2.n1386 3.4105
R9926 GNDA_2.n1408 GNDA_2.n1374 3.4105
R9927 GNDA_2.n1408 GNDA_2.n1387 3.4105
R9928 GNDA_2.n1408 GNDA_2.n1373 3.4105
R9929 GNDA_2.n1408 GNDA_2.n1388 3.4105
R9930 GNDA_2.n1408 GNDA_2.n1372 3.4105
R9931 GNDA_2.n1408 GNDA_2.n1389 3.4105
R9932 GNDA_2.n1408 GNDA_2.n1371 3.4105
R9933 GNDA_2.n1408 GNDA_2.n1390 3.4105
R9934 GNDA_2.n1408 GNDA_2.n1370 3.4105
R9935 GNDA_2.n1408 GNDA_2.n1391 3.4105
R9936 GNDA_2.n1408 GNDA_2.n1369 3.4105
R9937 GNDA_2.n1408 GNDA_2.n1392 3.4105
R9938 GNDA_2.n1408 GNDA_2.n1368 3.4105
R9939 GNDA_2.n1408 GNDA_2.n1393 3.4105
R9940 GNDA_2.n1408 GNDA_2.n1367 3.4105
R9941 GNDA_2.n1408 GNDA_2.n1394 3.4105
R9942 GNDA_2.n1408 GNDA_2.n1366 3.4105
R9943 GNDA_2.n1408 GNDA_2.n1395 3.4105
R9944 GNDA_2.n1408 GNDA_2.n1365 3.4105
R9945 GNDA_2.n1408 GNDA_2.n1396 3.4105
R9946 GNDA_2.n3512 GNDA_2.n1408 3.4105
R9947 GNDA_2.n3492 GNDA_2.n3471 3.4105
R9948 GNDA_2.n3471 GNDA_2.n1381 3.4105
R9949 GNDA_2.n3471 GNDA_2.n1379 3.4105
R9950 GNDA_2.n3471 GNDA_2.n1382 3.4105
R9951 GNDA_2.n3471 GNDA_2.n1378 3.4105
R9952 GNDA_2.n3471 GNDA_2.n1383 3.4105
R9953 GNDA_2.n3471 GNDA_2.n1377 3.4105
R9954 GNDA_2.n3471 GNDA_2.n1384 3.4105
R9955 GNDA_2.n3471 GNDA_2.n1376 3.4105
R9956 GNDA_2.n3471 GNDA_2.n1385 3.4105
R9957 GNDA_2.n3471 GNDA_2.n1375 3.4105
R9958 GNDA_2.n3471 GNDA_2.n1386 3.4105
R9959 GNDA_2.n3471 GNDA_2.n1374 3.4105
R9960 GNDA_2.n3471 GNDA_2.n1387 3.4105
R9961 GNDA_2.n3471 GNDA_2.n1373 3.4105
R9962 GNDA_2.n3471 GNDA_2.n1388 3.4105
R9963 GNDA_2.n3471 GNDA_2.n1372 3.4105
R9964 GNDA_2.n3471 GNDA_2.n1389 3.4105
R9965 GNDA_2.n3471 GNDA_2.n1371 3.4105
R9966 GNDA_2.n3471 GNDA_2.n1390 3.4105
R9967 GNDA_2.n3471 GNDA_2.n1370 3.4105
R9968 GNDA_2.n3471 GNDA_2.n1391 3.4105
R9969 GNDA_2.n3471 GNDA_2.n1369 3.4105
R9970 GNDA_2.n3471 GNDA_2.n1392 3.4105
R9971 GNDA_2.n3471 GNDA_2.n1368 3.4105
R9972 GNDA_2.n3471 GNDA_2.n1393 3.4105
R9973 GNDA_2.n3471 GNDA_2.n1367 3.4105
R9974 GNDA_2.n3471 GNDA_2.n1394 3.4105
R9975 GNDA_2.n3471 GNDA_2.n1366 3.4105
R9976 GNDA_2.n3471 GNDA_2.n1395 3.4105
R9977 GNDA_2.n3471 GNDA_2.n1365 3.4105
R9978 GNDA_2.n3471 GNDA_2.n1396 3.4105
R9979 GNDA_2.n3512 GNDA_2.n3471 3.4105
R9980 GNDA_2.n3492 GNDA_2.n1407 3.4105
R9981 GNDA_2.n1407 GNDA_2.n1381 3.4105
R9982 GNDA_2.n1407 GNDA_2.n1379 3.4105
R9983 GNDA_2.n1407 GNDA_2.n1382 3.4105
R9984 GNDA_2.n1407 GNDA_2.n1378 3.4105
R9985 GNDA_2.n1407 GNDA_2.n1383 3.4105
R9986 GNDA_2.n1407 GNDA_2.n1377 3.4105
R9987 GNDA_2.n1407 GNDA_2.n1384 3.4105
R9988 GNDA_2.n1407 GNDA_2.n1376 3.4105
R9989 GNDA_2.n1407 GNDA_2.n1385 3.4105
R9990 GNDA_2.n1407 GNDA_2.n1375 3.4105
R9991 GNDA_2.n1407 GNDA_2.n1386 3.4105
R9992 GNDA_2.n1407 GNDA_2.n1374 3.4105
R9993 GNDA_2.n1407 GNDA_2.n1387 3.4105
R9994 GNDA_2.n1407 GNDA_2.n1373 3.4105
R9995 GNDA_2.n1407 GNDA_2.n1388 3.4105
R9996 GNDA_2.n1407 GNDA_2.n1372 3.4105
R9997 GNDA_2.n1407 GNDA_2.n1389 3.4105
R9998 GNDA_2.n1407 GNDA_2.n1371 3.4105
R9999 GNDA_2.n1407 GNDA_2.n1390 3.4105
R10000 GNDA_2.n1407 GNDA_2.n1370 3.4105
R10001 GNDA_2.n1407 GNDA_2.n1391 3.4105
R10002 GNDA_2.n1407 GNDA_2.n1369 3.4105
R10003 GNDA_2.n1407 GNDA_2.n1392 3.4105
R10004 GNDA_2.n1407 GNDA_2.n1368 3.4105
R10005 GNDA_2.n1407 GNDA_2.n1393 3.4105
R10006 GNDA_2.n1407 GNDA_2.n1367 3.4105
R10007 GNDA_2.n1407 GNDA_2.n1394 3.4105
R10008 GNDA_2.n1407 GNDA_2.n1366 3.4105
R10009 GNDA_2.n1407 GNDA_2.n1395 3.4105
R10010 GNDA_2.n1407 GNDA_2.n1365 3.4105
R10011 GNDA_2.n1407 GNDA_2.n1396 3.4105
R10012 GNDA_2.n3512 GNDA_2.n1407 3.4105
R10013 GNDA_2.n3492 GNDA_2.n3473 3.4105
R10014 GNDA_2.n3473 GNDA_2.n1381 3.4105
R10015 GNDA_2.n3473 GNDA_2.n1379 3.4105
R10016 GNDA_2.n3473 GNDA_2.n1382 3.4105
R10017 GNDA_2.n3473 GNDA_2.n1378 3.4105
R10018 GNDA_2.n3473 GNDA_2.n1383 3.4105
R10019 GNDA_2.n3473 GNDA_2.n1377 3.4105
R10020 GNDA_2.n3473 GNDA_2.n1384 3.4105
R10021 GNDA_2.n3473 GNDA_2.n1376 3.4105
R10022 GNDA_2.n3473 GNDA_2.n1385 3.4105
R10023 GNDA_2.n3473 GNDA_2.n1375 3.4105
R10024 GNDA_2.n3473 GNDA_2.n1386 3.4105
R10025 GNDA_2.n3473 GNDA_2.n1374 3.4105
R10026 GNDA_2.n3473 GNDA_2.n1387 3.4105
R10027 GNDA_2.n3473 GNDA_2.n1373 3.4105
R10028 GNDA_2.n3473 GNDA_2.n1388 3.4105
R10029 GNDA_2.n3473 GNDA_2.n1372 3.4105
R10030 GNDA_2.n3473 GNDA_2.n1389 3.4105
R10031 GNDA_2.n3473 GNDA_2.n1371 3.4105
R10032 GNDA_2.n3473 GNDA_2.n1390 3.4105
R10033 GNDA_2.n3473 GNDA_2.n1370 3.4105
R10034 GNDA_2.n3473 GNDA_2.n1391 3.4105
R10035 GNDA_2.n3473 GNDA_2.n1369 3.4105
R10036 GNDA_2.n3473 GNDA_2.n1392 3.4105
R10037 GNDA_2.n3473 GNDA_2.n1368 3.4105
R10038 GNDA_2.n3473 GNDA_2.n1393 3.4105
R10039 GNDA_2.n3473 GNDA_2.n1367 3.4105
R10040 GNDA_2.n3473 GNDA_2.n1394 3.4105
R10041 GNDA_2.n3473 GNDA_2.n1366 3.4105
R10042 GNDA_2.n3473 GNDA_2.n1395 3.4105
R10043 GNDA_2.n3473 GNDA_2.n1365 3.4105
R10044 GNDA_2.n3473 GNDA_2.n1396 3.4105
R10045 GNDA_2.n3512 GNDA_2.n3473 3.4105
R10046 GNDA_2.n3492 GNDA_2.n1406 3.4105
R10047 GNDA_2.n1406 GNDA_2.n1381 3.4105
R10048 GNDA_2.n1406 GNDA_2.n1379 3.4105
R10049 GNDA_2.n1406 GNDA_2.n1382 3.4105
R10050 GNDA_2.n1406 GNDA_2.n1378 3.4105
R10051 GNDA_2.n1406 GNDA_2.n1383 3.4105
R10052 GNDA_2.n1406 GNDA_2.n1377 3.4105
R10053 GNDA_2.n1406 GNDA_2.n1384 3.4105
R10054 GNDA_2.n1406 GNDA_2.n1376 3.4105
R10055 GNDA_2.n1406 GNDA_2.n1385 3.4105
R10056 GNDA_2.n1406 GNDA_2.n1375 3.4105
R10057 GNDA_2.n1406 GNDA_2.n1386 3.4105
R10058 GNDA_2.n1406 GNDA_2.n1374 3.4105
R10059 GNDA_2.n1406 GNDA_2.n1387 3.4105
R10060 GNDA_2.n1406 GNDA_2.n1373 3.4105
R10061 GNDA_2.n1406 GNDA_2.n1388 3.4105
R10062 GNDA_2.n1406 GNDA_2.n1372 3.4105
R10063 GNDA_2.n1406 GNDA_2.n1389 3.4105
R10064 GNDA_2.n1406 GNDA_2.n1371 3.4105
R10065 GNDA_2.n1406 GNDA_2.n1390 3.4105
R10066 GNDA_2.n1406 GNDA_2.n1370 3.4105
R10067 GNDA_2.n1406 GNDA_2.n1391 3.4105
R10068 GNDA_2.n1406 GNDA_2.n1369 3.4105
R10069 GNDA_2.n1406 GNDA_2.n1392 3.4105
R10070 GNDA_2.n1406 GNDA_2.n1368 3.4105
R10071 GNDA_2.n1406 GNDA_2.n1393 3.4105
R10072 GNDA_2.n1406 GNDA_2.n1367 3.4105
R10073 GNDA_2.n1406 GNDA_2.n1394 3.4105
R10074 GNDA_2.n1406 GNDA_2.n1366 3.4105
R10075 GNDA_2.n1406 GNDA_2.n1395 3.4105
R10076 GNDA_2.n1406 GNDA_2.n1365 3.4105
R10077 GNDA_2.n1406 GNDA_2.n1396 3.4105
R10078 GNDA_2.n3512 GNDA_2.n1406 3.4105
R10079 GNDA_2.n3492 GNDA_2.n3475 3.4105
R10080 GNDA_2.n3475 GNDA_2.n1381 3.4105
R10081 GNDA_2.n3475 GNDA_2.n1379 3.4105
R10082 GNDA_2.n3475 GNDA_2.n1382 3.4105
R10083 GNDA_2.n3475 GNDA_2.n1378 3.4105
R10084 GNDA_2.n3475 GNDA_2.n1383 3.4105
R10085 GNDA_2.n3475 GNDA_2.n1377 3.4105
R10086 GNDA_2.n3475 GNDA_2.n1384 3.4105
R10087 GNDA_2.n3475 GNDA_2.n1376 3.4105
R10088 GNDA_2.n3475 GNDA_2.n1385 3.4105
R10089 GNDA_2.n3475 GNDA_2.n1375 3.4105
R10090 GNDA_2.n3475 GNDA_2.n1386 3.4105
R10091 GNDA_2.n3475 GNDA_2.n1374 3.4105
R10092 GNDA_2.n3475 GNDA_2.n1387 3.4105
R10093 GNDA_2.n3475 GNDA_2.n1373 3.4105
R10094 GNDA_2.n3475 GNDA_2.n1388 3.4105
R10095 GNDA_2.n3475 GNDA_2.n1372 3.4105
R10096 GNDA_2.n3475 GNDA_2.n1389 3.4105
R10097 GNDA_2.n3475 GNDA_2.n1371 3.4105
R10098 GNDA_2.n3475 GNDA_2.n1390 3.4105
R10099 GNDA_2.n3475 GNDA_2.n1370 3.4105
R10100 GNDA_2.n3475 GNDA_2.n1391 3.4105
R10101 GNDA_2.n3475 GNDA_2.n1369 3.4105
R10102 GNDA_2.n3475 GNDA_2.n1392 3.4105
R10103 GNDA_2.n3475 GNDA_2.n1368 3.4105
R10104 GNDA_2.n3475 GNDA_2.n1393 3.4105
R10105 GNDA_2.n3475 GNDA_2.n1367 3.4105
R10106 GNDA_2.n3475 GNDA_2.n1394 3.4105
R10107 GNDA_2.n3475 GNDA_2.n1366 3.4105
R10108 GNDA_2.n3475 GNDA_2.n1395 3.4105
R10109 GNDA_2.n3475 GNDA_2.n1365 3.4105
R10110 GNDA_2.n3475 GNDA_2.n1396 3.4105
R10111 GNDA_2.n3512 GNDA_2.n3475 3.4105
R10112 GNDA_2.n3492 GNDA_2.n1405 3.4105
R10113 GNDA_2.n1405 GNDA_2.n1381 3.4105
R10114 GNDA_2.n1405 GNDA_2.n1379 3.4105
R10115 GNDA_2.n1405 GNDA_2.n1382 3.4105
R10116 GNDA_2.n1405 GNDA_2.n1378 3.4105
R10117 GNDA_2.n1405 GNDA_2.n1383 3.4105
R10118 GNDA_2.n1405 GNDA_2.n1377 3.4105
R10119 GNDA_2.n1405 GNDA_2.n1384 3.4105
R10120 GNDA_2.n1405 GNDA_2.n1376 3.4105
R10121 GNDA_2.n1405 GNDA_2.n1385 3.4105
R10122 GNDA_2.n1405 GNDA_2.n1375 3.4105
R10123 GNDA_2.n1405 GNDA_2.n1386 3.4105
R10124 GNDA_2.n1405 GNDA_2.n1374 3.4105
R10125 GNDA_2.n1405 GNDA_2.n1387 3.4105
R10126 GNDA_2.n1405 GNDA_2.n1373 3.4105
R10127 GNDA_2.n1405 GNDA_2.n1388 3.4105
R10128 GNDA_2.n1405 GNDA_2.n1372 3.4105
R10129 GNDA_2.n1405 GNDA_2.n1389 3.4105
R10130 GNDA_2.n1405 GNDA_2.n1371 3.4105
R10131 GNDA_2.n1405 GNDA_2.n1390 3.4105
R10132 GNDA_2.n1405 GNDA_2.n1370 3.4105
R10133 GNDA_2.n1405 GNDA_2.n1391 3.4105
R10134 GNDA_2.n1405 GNDA_2.n1369 3.4105
R10135 GNDA_2.n1405 GNDA_2.n1392 3.4105
R10136 GNDA_2.n1405 GNDA_2.n1368 3.4105
R10137 GNDA_2.n1405 GNDA_2.n1393 3.4105
R10138 GNDA_2.n1405 GNDA_2.n1367 3.4105
R10139 GNDA_2.n1405 GNDA_2.n1394 3.4105
R10140 GNDA_2.n1405 GNDA_2.n1366 3.4105
R10141 GNDA_2.n1405 GNDA_2.n1395 3.4105
R10142 GNDA_2.n1405 GNDA_2.n1365 3.4105
R10143 GNDA_2.n1405 GNDA_2.n1396 3.4105
R10144 GNDA_2.n3512 GNDA_2.n1405 3.4105
R10145 GNDA_2.n3492 GNDA_2.n3477 3.4105
R10146 GNDA_2.n3477 GNDA_2.n1381 3.4105
R10147 GNDA_2.n3477 GNDA_2.n1379 3.4105
R10148 GNDA_2.n3477 GNDA_2.n1382 3.4105
R10149 GNDA_2.n3477 GNDA_2.n1378 3.4105
R10150 GNDA_2.n3477 GNDA_2.n1383 3.4105
R10151 GNDA_2.n3477 GNDA_2.n1377 3.4105
R10152 GNDA_2.n3477 GNDA_2.n1384 3.4105
R10153 GNDA_2.n3477 GNDA_2.n1376 3.4105
R10154 GNDA_2.n3477 GNDA_2.n1385 3.4105
R10155 GNDA_2.n3477 GNDA_2.n1375 3.4105
R10156 GNDA_2.n3477 GNDA_2.n1386 3.4105
R10157 GNDA_2.n3477 GNDA_2.n1374 3.4105
R10158 GNDA_2.n3477 GNDA_2.n1387 3.4105
R10159 GNDA_2.n3477 GNDA_2.n1373 3.4105
R10160 GNDA_2.n3477 GNDA_2.n1388 3.4105
R10161 GNDA_2.n3477 GNDA_2.n1372 3.4105
R10162 GNDA_2.n3477 GNDA_2.n1389 3.4105
R10163 GNDA_2.n3477 GNDA_2.n1371 3.4105
R10164 GNDA_2.n3477 GNDA_2.n1390 3.4105
R10165 GNDA_2.n3477 GNDA_2.n1370 3.4105
R10166 GNDA_2.n3477 GNDA_2.n1391 3.4105
R10167 GNDA_2.n3477 GNDA_2.n1369 3.4105
R10168 GNDA_2.n3477 GNDA_2.n1392 3.4105
R10169 GNDA_2.n3477 GNDA_2.n1368 3.4105
R10170 GNDA_2.n3477 GNDA_2.n1393 3.4105
R10171 GNDA_2.n3477 GNDA_2.n1367 3.4105
R10172 GNDA_2.n3477 GNDA_2.n1394 3.4105
R10173 GNDA_2.n3477 GNDA_2.n1366 3.4105
R10174 GNDA_2.n3477 GNDA_2.n1395 3.4105
R10175 GNDA_2.n3477 GNDA_2.n1365 3.4105
R10176 GNDA_2.n3477 GNDA_2.n1396 3.4105
R10177 GNDA_2.n3512 GNDA_2.n3477 3.4105
R10178 GNDA_2.n3492 GNDA_2.n1404 3.4105
R10179 GNDA_2.n1404 GNDA_2.n1381 3.4105
R10180 GNDA_2.n1404 GNDA_2.n1379 3.4105
R10181 GNDA_2.n1404 GNDA_2.n1382 3.4105
R10182 GNDA_2.n1404 GNDA_2.n1378 3.4105
R10183 GNDA_2.n1404 GNDA_2.n1383 3.4105
R10184 GNDA_2.n1404 GNDA_2.n1377 3.4105
R10185 GNDA_2.n1404 GNDA_2.n1384 3.4105
R10186 GNDA_2.n1404 GNDA_2.n1376 3.4105
R10187 GNDA_2.n1404 GNDA_2.n1385 3.4105
R10188 GNDA_2.n1404 GNDA_2.n1375 3.4105
R10189 GNDA_2.n1404 GNDA_2.n1386 3.4105
R10190 GNDA_2.n1404 GNDA_2.n1374 3.4105
R10191 GNDA_2.n1404 GNDA_2.n1387 3.4105
R10192 GNDA_2.n1404 GNDA_2.n1373 3.4105
R10193 GNDA_2.n1404 GNDA_2.n1388 3.4105
R10194 GNDA_2.n1404 GNDA_2.n1372 3.4105
R10195 GNDA_2.n1404 GNDA_2.n1389 3.4105
R10196 GNDA_2.n1404 GNDA_2.n1371 3.4105
R10197 GNDA_2.n1404 GNDA_2.n1390 3.4105
R10198 GNDA_2.n1404 GNDA_2.n1370 3.4105
R10199 GNDA_2.n1404 GNDA_2.n1391 3.4105
R10200 GNDA_2.n1404 GNDA_2.n1369 3.4105
R10201 GNDA_2.n1404 GNDA_2.n1392 3.4105
R10202 GNDA_2.n1404 GNDA_2.n1368 3.4105
R10203 GNDA_2.n1404 GNDA_2.n1393 3.4105
R10204 GNDA_2.n1404 GNDA_2.n1367 3.4105
R10205 GNDA_2.n1404 GNDA_2.n1394 3.4105
R10206 GNDA_2.n1404 GNDA_2.n1366 3.4105
R10207 GNDA_2.n1404 GNDA_2.n1395 3.4105
R10208 GNDA_2.n1404 GNDA_2.n1365 3.4105
R10209 GNDA_2.n1404 GNDA_2.n1396 3.4105
R10210 GNDA_2.n3512 GNDA_2.n1404 3.4105
R10211 GNDA_2.n3492 GNDA_2.n3479 3.4105
R10212 GNDA_2.n3479 GNDA_2.n1381 3.4105
R10213 GNDA_2.n3479 GNDA_2.n1379 3.4105
R10214 GNDA_2.n3479 GNDA_2.n1382 3.4105
R10215 GNDA_2.n3479 GNDA_2.n1378 3.4105
R10216 GNDA_2.n3479 GNDA_2.n1383 3.4105
R10217 GNDA_2.n3479 GNDA_2.n1377 3.4105
R10218 GNDA_2.n3479 GNDA_2.n1384 3.4105
R10219 GNDA_2.n3479 GNDA_2.n1376 3.4105
R10220 GNDA_2.n3479 GNDA_2.n1385 3.4105
R10221 GNDA_2.n3479 GNDA_2.n1375 3.4105
R10222 GNDA_2.n3479 GNDA_2.n1386 3.4105
R10223 GNDA_2.n3479 GNDA_2.n1374 3.4105
R10224 GNDA_2.n3479 GNDA_2.n1387 3.4105
R10225 GNDA_2.n3479 GNDA_2.n1373 3.4105
R10226 GNDA_2.n3479 GNDA_2.n1388 3.4105
R10227 GNDA_2.n3479 GNDA_2.n1372 3.4105
R10228 GNDA_2.n3479 GNDA_2.n1389 3.4105
R10229 GNDA_2.n3479 GNDA_2.n1371 3.4105
R10230 GNDA_2.n3479 GNDA_2.n1390 3.4105
R10231 GNDA_2.n3479 GNDA_2.n1370 3.4105
R10232 GNDA_2.n3479 GNDA_2.n1391 3.4105
R10233 GNDA_2.n3479 GNDA_2.n1369 3.4105
R10234 GNDA_2.n3479 GNDA_2.n1392 3.4105
R10235 GNDA_2.n3479 GNDA_2.n1368 3.4105
R10236 GNDA_2.n3479 GNDA_2.n1393 3.4105
R10237 GNDA_2.n3479 GNDA_2.n1367 3.4105
R10238 GNDA_2.n3479 GNDA_2.n1394 3.4105
R10239 GNDA_2.n3479 GNDA_2.n1366 3.4105
R10240 GNDA_2.n3479 GNDA_2.n1395 3.4105
R10241 GNDA_2.n3479 GNDA_2.n1365 3.4105
R10242 GNDA_2.n3479 GNDA_2.n1396 3.4105
R10243 GNDA_2.n3512 GNDA_2.n3479 3.4105
R10244 GNDA_2.n3492 GNDA_2.n1403 3.4105
R10245 GNDA_2.n1403 GNDA_2.n1381 3.4105
R10246 GNDA_2.n1403 GNDA_2.n1379 3.4105
R10247 GNDA_2.n1403 GNDA_2.n1382 3.4105
R10248 GNDA_2.n1403 GNDA_2.n1378 3.4105
R10249 GNDA_2.n1403 GNDA_2.n1383 3.4105
R10250 GNDA_2.n1403 GNDA_2.n1377 3.4105
R10251 GNDA_2.n1403 GNDA_2.n1384 3.4105
R10252 GNDA_2.n1403 GNDA_2.n1376 3.4105
R10253 GNDA_2.n1403 GNDA_2.n1385 3.4105
R10254 GNDA_2.n1403 GNDA_2.n1375 3.4105
R10255 GNDA_2.n1403 GNDA_2.n1386 3.4105
R10256 GNDA_2.n1403 GNDA_2.n1374 3.4105
R10257 GNDA_2.n1403 GNDA_2.n1387 3.4105
R10258 GNDA_2.n1403 GNDA_2.n1373 3.4105
R10259 GNDA_2.n1403 GNDA_2.n1388 3.4105
R10260 GNDA_2.n1403 GNDA_2.n1372 3.4105
R10261 GNDA_2.n1403 GNDA_2.n1389 3.4105
R10262 GNDA_2.n1403 GNDA_2.n1371 3.4105
R10263 GNDA_2.n1403 GNDA_2.n1390 3.4105
R10264 GNDA_2.n1403 GNDA_2.n1370 3.4105
R10265 GNDA_2.n1403 GNDA_2.n1391 3.4105
R10266 GNDA_2.n1403 GNDA_2.n1369 3.4105
R10267 GNDA_2.n1403 GNDA_2.n1392 3.4105
R10268 GNDA_2.n1403 GNDA_2.n1368 3.4105
R10269 GNDA_2.n1403 GNDA_2.n1393 3.4105
R10270 GNDA_2.n1403 GNDA_2.n1367 3.4105
R10271 GNDA_2.n1403 GNDA_2.n1394 3.4105
R10272 GNDA_2.n1403 GNDA_2.n1366 3.4105
R10273 GNDA_2.n1403 GNDA_2.n1395 3.4105
R10274 GNDA_2.n1403 GNDA_2.n1365 3.4105
R10275 GNDA_2.n1403 GNDA_2.n1396 3.4105
R10276 GNDA_2.n3512 GNDA_2.n1403 3.4105
R10277 GNDA_2.n3492 GNDA_2.n3481 3.4105
R10278 GNDA_2.n3481 GNDA_2.n1381 3.4105
R10279 GNDA_2.n3481 GNDA_2.n1379 3.4105
R10280 GNDA_2.n3481 GNDA_2.n1382 3.4105
R10281 GNDA_2.n3481 GNDA_2.n1378 3.4105
R10282 GNDA_2.n3481 GNDA_2.n1383 3.4105
R10283 GNDA_2.n3481 GNDA_2.n1377 3.4105
R10284 GNDA_2.n3481 GNDA_2.n1384 3.4105
R10285 GNDA_2.n3481 GNDA_2.n1376 3.4105
R10286 GNDA_2.n3481 GNDA_2.n1385 3.4105
R10287 GNDA_2.n3481 GNDA_2.n1375 3.4105
R10288 GNDA_2.n3481 GNDA_2.n1386 3.4105
R10289 GNDA_2.n3481 GNDA_2.n1374 3.4105
R10290 GNDA_2.n3481 GNDA_2.n1387 3.4105
R10291 GNDA_2.n3481 GNDA_2.n1373 3.4105
R10292 GNDA_2.n3481 GNDA_2.n1388 3.4105
R10293 GNDA_2.n3481 GNDA_2.n1372 3.4105
R10294 GNDA_2.n3481 GNDA_2.n1389 3.4105
R10295 GNDA_2.n3481 GNDA_2.n1371 3.4105
R10296 GNDA_2.n3481 GNDA_2.n1390 3.4105
R10297 GNDA_2.n3481 GNDA_2.n1370 3.4105
R10298 GNDA_2.n3481 GNDA_2.n1391 3.4105
R10299 GNDA_2.n3481 GNDA_2.n1369 3.4105
R10300 GNDA_2.n3481 GNDA_2.n1392 3.4105
R10301 GNDA_2.n3481 GNDA_2.n1368 3.4105
R10302 GNDA_2.n3481 GNDA_2.n1393 3.4105
R10303 GNDA_2.n3481 GNDA_2.n1367 3.4105
R10304 GNDA_2.n3481 GNDA_2.n1394 3.4105
R10305 GNDA_2.n3481 GNDA_2.n1366 3.4105
R10306 GNDA_2.n3481 GNDA_2.n1395 3.4105
R10307 GNDA_2.n3481 GNDA_2.n1365 3.4105
R10308 GNDA_2.n3481 GNDA_2.n1396 3.4105
R10309 GNDA_2.n3512 GNDA_2.n3481 3.4105
R10310 GNDA_2.n3492 GNDA_2.n1402 3.4105
R10311 GNDA_2.n1402 GNDA_2.n1381 3.4105
R10312 GNDA_2.n1402 GNDA_2.n1379 3.4105
R10313 GNDA_2.n1402 GNDA_2.n1382 3.4105
R10314 GNDA_2.n1402 GNDA_2.n1378 3.4105
R10315 GNDA_2.n1402 GNDA_2.n1383 3.4105
R10316 GNDA_2.n1402 GNDA_2.n1377 3.4105
R10317 GNDA_2.n1402 GNDA_2.n1384 3.4105
R10318 GNDA_2.n1402 GNDA_2.n1376 3.4105
R10319 GNDA_2.n1402 GNDA_2.n1385 3.4105
R10320 GNDA_2.n1402 GNDA_2.n1375 3.4105
R10321 GNDA_2.n1402 GNDA_2.n1386 3.4105
R10322 GNDA_2.n1402 GNDA_2.n1374 3.4105
R10323 GNDA_2.n1402 GNDA_2.n1387 3.4105
R10324 GNDA_2.n1402 GNDA_2.n1373 3.4105
R10325 GNDA_2.n1402 GNDA_2.n1388 3.4105
R10326 GNDA_2.n1402 GNDA_2.n1372 3.4105
R10327 GNDA_2.n1402 GNDA_2.n1389 3.4105
R10328 GNDA_2.n1402 GNDA_2.n1371 3.4105
R10329 GNDA_2.n1402 GNDA_2.n1390 3.4105
R10330 GNDA_2.n1402 GNDA_2.n1370 3.4105
R10331 GNDA_2.n1402 GNDA_2.n1391 3.4105
R10332 GNDA_2.n1402 GNDA_2.n1369 3.4105
R10333 GNDA_2.n1402 GNDA_2.n1392 3.4105
R10334 GNDA_2.n1402 GNDA_2.n1368 3.4105
R10335 GNDA_2.n1402 GNDA_2.n1393 3.4105
R10336 GNDA_2.n1402 GNDA_2.n1367 3.4105
R10337 GNDA_2.n1402 GNDA_2.n1394 3.4105
R10338 GNDA_2.n1402 GNDA_2.n1366 3.4105
R10339 GNDA_2.n1402 GNDA_2.n1395 3.4105
R10340 GNDA_2.n1402 GNDA_2.n1365 3.4105
R10341 GNDA_2.n1402 GNDA_2.n1396 3.4105
R10342 GNDA_2.n3512 GNDA_2.n1402 3.4105
R10343 GNDA_2.n3492 GNDA_2.n3483 3.4105
R10344 GNDA_2.n3483 GNDA_2.n1381 3.4105
R10345 GNDA_2.n3483 GNDA_2.n1379 3.4105
R10346 GNDA_2.n3483 GNDA_2.n1382 3.4105
R10347 GNDA_2.n3483 GNDA_2.n1378 3.4105
R10348 GNDA_2.n3483 GNDA_2.n1383 3.4105
R10349 GNDA_2.n3483 GNDA_2.n1377 3.4105
R10350 GNDA_2.n3483 GNDA_2.n1384 3.4105
R10351 GNDA_2.n3483 GNDA_2.n1376 3.4105
R10352 GNDA_2.n3483 GNDA_2.n1385 3.4105
R10353 GNDA_2.n3483 GNDA_2.n1375 3.4105
R10354 GNDA_2.n3483 GNDA_2.n1386 3.4105
R10355 GNDA_2.n3483 GNDA_2.n1374 3.4105
R10356 GNDA_2.n3483 GNDA_2.n1387 3.4105
R10357 GNDA_2.n3483 GNDA_2.n1373 3.4105
R10358 GNDA_2.n3483 GNDA_2.n1388 3.4105
R10359 GNDA_2.n3483 GNDA_2.n1372 3.4105
R10360 GNDA_2.n3483 GNDA_2.n1389 3.4105
R10361 GNDA_2.n3483 GNDA_2.n1371 3.4105
R10362 GNDA_2.n3483 GNDA_2.n1390 3.4105
R10363 GNDA_2.n3483 GNDA_2.n1370 3.4105
R10364 GNDA_2.n3483 GNDA_2.n1391 3.4105
R10365 GNDA_2.n3483 GNDA_2.n1369 3.4105
R10366 GNDA_2.n3483 GNDA_2.n1392 3.4105
R10367 GNDA_2.n3483 GNDA_2.n1368 3.4105
R10368 GNDA_2.n3483 GNDA_2.n1393 3.4105
R10369 GNDA_2.n3483 GNDA_2.n1367 3.4105
R10370 GNDA_2.n3483 GNDA_2.n1394 3.4105
R10371 GNDA_2.n3483 GNDA_2.n1366 3.4105
R10372 GNDA_2.n3483 GNDA_2.n1395 3.4105
R10373 GNDA_2.n3483 GNDA_2.n1365 3.4105
R10374 GNDA_2.n3483 GNDA_2.n1396 3.4105
R10375 GNDA_2.n3512 GNDA_2.n3483 3.4105
R10376 GNDA_2.n3492 GNDA_2.n1401 3.4105
R10377 GNDA_2.n1401 GNDA_2.n1381 3.4105
R10378 GNDA_2.n1401 GNDA_2.n1379 3.4105
R10379 GNDA_2.n1401 GNDA_2.n1382 3.4105
R10380 GNDA_2.n1401 GNDA_2.n1378 3.4105
R10381 GNDA_2.n1401 GNDA_2.n1383 3.4105
R10382 GNDA_2.n1401 GNDA_2.n1377 3.4105
R10383 GNDA_2.n1401 GNDA_2.n1384 3.4105
R10384 GNDA_2.n1401 GNDA_2.n1376 3.4105
R10385 GNDA_2.n1401 GNDA_2.n1385 3.4105
R10386 GNDA_2.n1401 GNDA_2.n1375 3.4105
R10387 GNDA_2.n1401 GNDA_2.n1386 3.4105
R10388 GNDA_2.n1401 GNDA_2.n1374 3.4105
R10389 GNDA_2.n1401 GNDA_2.n1387 3.4105
R10390 GNDA_2.n1401 GNDA_2.n1373 3.4105
R10391 GNDA_2.n1401 GNDA_2.n1388 3.4105
R10392 GNDA_2.n1401 GNDA_2.n1372 3.4105
R10393 GNDA_2.n1401 GNDA_2.n1389 3.4105
R10394 GNDA_2.n1401 GNDA_2.n1371 3.4105
R10395 GNDA_2.n1401 GNDA_2.n1390 3.4105
R10396 GNDA_2.n1401 GNDA_2.n1370 3.4105
R10397 GNDA_2.n1401 GNDA_2.n1391 3.4105
R10398 GNDA_2.n1401 GNDA_2.n1369 3.4105
R10399 GNDA_2.n1401 GNDA_2.n1392 3.4105
R10400 GNDA_2.n1401 GNDA_2.n1368 3.4105
R10401 GNDA_2.n1401 GNDA_2.n1393 3.4105
R10402 GNDA_2.n1401 GNDA_2.n1367 3.4105
R10403 GNDA_2.n1401 GNDA_2.n1394 3.4105
R10404 GNDA_2.n1401 GNDA_2.n1366 3.4105
R10405 GNDA_2.n1401 GNDA_2.n1395 3.4105
R10406 GNDA_2.n1401 GNDA_2.n1365 3.4105
R10407 GNDA_2.n1401 GNDA_2.n1396 3.4105
R10408 GNDA_2.n3512 GNDA_2.n1401 3.4105
R10409 GNDA_2.n3492 GNDA_2.n3485 3.4105
R10410 GNDA_2.n3485 GNDA_2.n1381 3.4105
R10411 GNDA_2.n3485 GNDA_2.n1379 3.4105
R10412 GNDA_2.n3485 GNDA_2.n1382 3.4105
R10413 GNDA_2.n3485 GNDA_2.n1378 3.4105
R10414 GNDA_2.n3485 GNDA_2.n1383 3.4105
R10415 GNDA_2.n3485 GNDA_2.n1377 3.4105
R10416 GNDA_2.n3485 GNDA_2.n1384 3.4105
R10417 GNDA_2.n3485 GNDA_2.n1376 3.4105
R10418 GNDA_2.n3485 GNDA_2.n1385 3.4105
R10419 GNDA_2.n3485 GNDA_2.n1375 3.4105
R10420 GNDA_2.n3485 GNDA_2.n1386 3.4105
R10421 GNDA_2.n3485 GNDA_2.n1374 3.4105
R10422 GNDA_2.n3485 GNDA_2.n1387 3.4105
R10423 GNDA_2.n3485 GNDA_2.n1373 3.4105
R10424 GNDA_2.n3485 GNDA_2.n1388 3.4105
R10425 GNDA_2.n3485 GNDA_2.n1372 3.4105
R10426 GNDA_2.n3485 GNDA_2.n1389 3.4105
R10427 GNDA_2.n3485 GNDA_2.n1371 3.4105
R10428 GNDA_2.n3485 GNDA_2.n1390 3.4105
R10429 GNDA_2.n3485 GNDA_2.n1370 3.4105
R10430 GNDA_2.n3485 GNDA_2.n1391 3.4105
R10431 GNDA_2.n3485 GNDA_2.n1369 3.4105
R10432 GNDA_2.n3485 GNDA_2.n1392 3.4105
R10433 GNDA_2.n3485 GNDA_2.n1368 3.4105
R10434 GNDA_2.n3485 GNDA_2.n1393 3.4105
R10435 GNDA_2.n3485 GNDA_2.n1367 3.4105
R10436 GNDA_2.n3485 GNDA_2.n1394 3.4105
R10437 GNDA_2.n3485 GNDA_2.n1366 3.4105
R10438 GNDA_2.n3485 GNDA_2.n1395 3.4105
R10439 GNDA_2.n3485 GNDA_2.n1365 3.4105
R10440 GNDA_2.n3485 GNDA_2.n1396 3.4105
R10441 GNDA_2.n3512 GNDA_2.n3485 3.4105
R10442 GNDA_2.n3492 GNDA_2.n1400 3.4105
R10443 GNDA_2.n1400 GNDA_2.n1381 3.4105
R10444 GNDA_2.n1400 GNDA_2.n1379 3.4105
R10445 GNDA_2.n1400 GNDA_2.n1382 3.4105
R10446 GNDA_2.n1400 GNDA_2.n1378 3.4105
R10447 GNDA_2.n1400 GNDA_2.n1383 3.4105
R10448 GNDA_2.n1400 GNDA_2.n1377 3.4105
R10449 GNDA_2.n1400 GNDA_2.n1384 3.4105
R10450 GNDA_2.n1400 GNDA_2.n1376 3.4105
R10451 GNDA_2.n1400 GNDA_2.n1385 3.4105
R10452 GNDA_2.n1400 GNDA_2.n1375 3.4105
R10453 GNDA_2.n1400 GNDA_2.n1386 3.4105
R10454 GNDA_2.n1400 GNDA_2.n1374 3.4105
R10455 GNDA_2.n1400 GNDA_2.n1387 3.4105
R10456 GNDA_2.n1400 GNDA_2.n1373 3.4105
R10457 GNDA_2.n1400 GNDA_2.n1388 3.4105
R10458 GNDA_2.n1400 GNDA_2.n1372 3.4105
R10459 GNDA_2.n1400 GNDA_2.n1389 3.4105
R10460 GNDA_2.n1400 GNDA_2.n1371 3.4105
R10461 GNDA_2.n1400 GNDA_2.n1390 3.4105
R10462 GNDA_2.n1400 GNDA_2.n1370 3.4105
R10463 GNDA_2.n1400 GNDA_2.n1391 3.4105
R10464 GNDA_2.n1400 GNDA_2.n1369 3.4105
R10465 GNDA_2.n1400 GNDA_2.n1392 3.4105
R10466 GNDA_2.n1400 GNDA_2.n1368 3.4105
R10467 GNDA_2.n1400 GNDA_2.n1393 3.4105
R10468 GNDA_2.n1400 GNDA_2.n1367 3.4105
R10469 GNDA_2.n1400 GNDA_2.n1394 3.4105
R10470 GNDA_2.n1400 GNDA_2.n1366 3.4105
R10471 GNDA_2.n1400 GNDA_2.n1395 3.4105
R10472 GNDA_2.n1400 GNDA_2.n1365 3.4105
R10473 GNDA_2.n1400 GNDA_2.n1396 3.4105
R10474 GNDA_2.n3512 GNDA_2.n1400 3.4105
R10475 GNDA_2.n3492 GNDA_2.n3487 3.4105
R10476 GNDA_2.n3487 GNDA_2.n1381 3.4105
R10477 GNDA_2.n3487 GNDA_2.n1379 3.4105
R10478 GNDA_2.n3487 GNDA_2.n1382 3.4105
R10479 GNDA_2.n3487 GNDA_2.n1378 3.4105
R10480 GNDA_2.n3487 GNDA_2.n1383 3.4105
R10481 GNDA_2.n3487 GNDA_2.n1377 3.4105
R10482 GNDA_2.n3487 GNDA_2.n1384 3.4105
R10483 GNDA_2.n3487 GNDA_2.n1376 3.4105
R10484 GNDA_2.n3487 GNDA_2.n1385 3.4105
R10485 GNDA_2.n3487 GNDA_2.n1375 3.4105
R10486 GNDA_2.n3487 GNDA_2.n1386 3.4105
R10487 GNDA_2.n3487 GNDA_2.n1374 3.4105
R10488 GNDA_2.n3487 GNDA_2.n1387 3.4105
R10489 GNDA_2.n3487 GNDA_2.n1373 3.4105
R10490 GNDA_2.n3487 GNDA_2.n1388 3.4105
R10491 GNDA_2.n3487 GNDA_2.n1372 3.4105
R10492 GNDA_2.n3487 GNDA_2.n1389 3.4105
R10493 GNDA_2.n3487 GNDA_2.n1371 3.4105
R10494 GNDA_2.n3487 GNDA_2.n1390 3.4105
R10495 GNDA_2.n3487 GNDA_2.n1370 3.4105
R10496 GNDA_2.n3487 GNDA_2.n1391 3.4105
R10497 GNDA_2.n3487 GNDA_2.n1369 3.4105
R10498 GNDA_2.n3487 GNDA_2.n1392 3.4105
R10499 GNDA_2.n3487 GNDA_2.n1368 3.4105
R10500 GNDA_2.n3487 GNDA_2.n1393 3.4105
R10501 GNDA_2.n3487 GNDA_2.n1367 3.4105
R10502 GNDA_2.n3487 GNDA_2.n1394 3.4105
R10503 GNDA_2.n3487 GNDA_2.n1366 3.4105
R10504 GNDA_2.n3487 GNDA_2.n1395 3.4105
R10505 GNDA_2.n3487 GNDA_2.n1365 3.4105
R10506 GNDA_2.n3487 GNDA_2.n1396 3.4105
R10507 GNDA_2.n3512 GNDA_2.n3487 3.4105
R10508 GNDA_2.n3492 GNDA_2.n1399 3.4105
R10509 GNDA_2.n1399 GNDA_2.n1381 3.4105
R10510 GNDA_2.n1399 GNDA_2.n1379 3.4105
R10511 GNDA_2.n1399 GNDA_2.n1382 3.4105
R10512 GNDA_2.n1399 GNDA_2.n1378 3.4105
R10513 GNDA_2.n1399 GNDA_2.n1383 3.4105
R10514 GNDA_2.n1399 GNDA_2.n1377 3.4105
R10515 GNDA_2.n1399 GNDA_2.n1384 3.4105
R10516 GNDA_2.n1399 GNDA_2.n1376 3.4105
R10517 GNDA_2.n1399 GNDA_2.n1385 3.4105
R10518 GNDA_2.n1399 GNDA_2.n1375 3.4105
R10519 GNDA_2.n1399 GNDA_2.n1386 3.4105
R10520 GNDA_2.n1399 GNDA_2.n1374 3.4105
R10521 GNDA_2.n1399 GNDA_2.n1387 3.4105
R10522 GNDA_2.n1399 GNDA_2.n1373 3.4105
R10523 GNDA_2.n1399 GNDA_2.n1388 3.4105
R10524 GNDA_2.n1399 GNDA_2.n1372 3.4105
R10525 GNDA_2.n1399 GNDA_2.n1389 3.4105
R10526 GNDA_2.n1399 GNDA_2.n1371 3.4105
R10527 GNDA_2.n1399 GNDA_2.n1390 3.4105
R10528 GNDA_2.n1399 GNDA_2.n1370 3.4105
R10529 GNDA_2.n1399 GNDA_2.n1391 3.4105
R10530 GNDA_2.n1399 GNDA_2.n1369 3.4105
R10531 GNDA_2.n1399 GNDA_2.n1392 3.4105
R10532 GNDA_2.n1399 GNDA_2.n1368 3.4105
R10533 GNDA_2.n1399 GNDA_2.n1393 3.4105
R10534 GNDA_2.n1399 GNDA_2.n1367 3.4105
R10535 GNDA_2.n1399 GNDA_2.n1394 3.4105
R10536 GNDA_2.n1399 GNDA_2.n1366 3.4105
R10537 GNDA_2.n1399 GNDA_2.n1395 3.4105
R10538 GNDA_2.n1399 GNDA_2.n1365 3.4105
R10539 GNDA_2.n1399 GNDA_2.n1396 3.4105
R10540 GNDA_2.n3512 GNDA_2.n1399 3.4105
R10541 GNDA_2.n3492 GNDA_2.n3489 3.4105
R10542 GNDA_2.n3489 GNDA_2.n1381 3.4105
R10543 GNDA_2.n3489 GNDA_2.n1379 3.4105
R10544 GNDA_2.n3489 GNDA_2.n1382 3.4105
R10545 GNDA_2.n3489 GNDA_2.n1378 3.4105
R10546 GNDA_2.n3489 GNDA_2.n1383 3.4105
R10547 GNDA_2.n3489 GNDA_2.n1377 3.4105
R10548 GNDA_2.n3489 GNDA_2.n1384 3.4105
R10549 GNDA_2.n3489 GNDA_2.n1376 3.4105
R10550 GNDA_2.n3489 GNDA_2.n1385 3.4105
R10551 GNDA_2.n3489 GNDA_2.n1375 3.4105
R10552 GNDA_2.n3489 GNDA_2.n1386 3.4105
R10553 GNDA_2.n3489 GNDA_2.n1374 3.4105
R10554 GNDA_2.n3489 GNDA_2.n1387 3.4105
R10555 GNDA_2.n3489 GNDA_2.n1373 3.4105
R10556 GNDA_2.n3489 GNDA_2.n1388 3.4105
R10557 GNDA_2.n3489 GNDA_2.n1372 3.4105
R10558 GNDA_2.n3489 GNDA_2.n1389 3.4105
R10559 GNDA_2.n3489 GNDA_2.n1371 3.4105
R10560 GNDA_2.n3489 GNDA_2.n1390 3.4105
R10561 GNDA_2.n3489 GNDA_2.n1370 3.4105
R10562 GNDA_2.n3489 GNDA_2.n1391 3.4105
R10563 GNDA_2.n3489 GNDA_2.n1369 3.4105
R10564 GNDA_2.n3489 GNDA_2.n1392 3.4105
R10565 GNDA_2.n3489 GNDA_2.n1368 3.4105
R10566 GNDA_2.n3489 GNDA_2.n1393 3.4105
R10567 GNDA_2.n3489 GNDA_2.n1367 3.4105
R10568 GNDA_2.n3489 GNDA_2.n1394 3.4105
R10569 GNDA_2.n3489 GNDA_2.n1366 3.4105
R10570 GNDA_2.n3489 GNDA_2.n1395 3.4105
R10571 GNDA_2.n3489 GNDA_2.n1365 3.4105
R10572 GNDA_2.n3489 GNDA_2.n1396 3.4105
R10573 GNDA_2.n3512 GNDA_2.n3489 3.4105
R10574 GNDA_2.n3492 GNDA_2.n1398 3.4105
R10575 GNDA_2.n1398 GNDA_2.n1381 3.4105
R10576 GNDA_2.n1398 GNDA_2.n1379 3.4105
R10577 GNDA_2.n1398 GNDA_2.n1382 3.4105
R10578 GNDA_2.n1398 GNDA_2.n1378 3.4105
R10579 GNDA_2.n1398 GNDA_2.n1383 3.4105
R10580 GNDA_2.n1398 GNDA_2.n1377 3.4105
R10581 GNDA_2.n1398 GNDA_2.n1384 3.4105
R10582 GNDA_2.n1398 GNDA_2.n1376 3.4105
R10583 GNDA_2.n1398 GNDA_2.n1385 3.4105
R10584 GNDA_2.n1398 GNDA_2.n1375 3.4105
R10585 GNDA_2.n1398 GNDA_2.n1386 3.4105
R10586 GNDA_2.n1398 GNDA_2.n1374 3.4105
R10587 GNDA_2.n1398 GNDA_2.n1387 3.4105
R10588 GNDA_2.n1398 GNDA_2.n1373 3.4105
R10589 GNDA_2.n1398 GNDA_2.n1388 3.4105
R10590 GNDA_2.n1398 GNDA_2.n1372 3.4105
R10591 GNDA_2.n1398 GNDA_2.n1389 3.4105
R10592 GNDA_2.n1398 GNDA_2.n1371 3.4105
R10593 GNDA_2.n1398 GNDA_2.n1390 3.4105
R10594 GNDA_2.n1398 GNDA_2.n1370 3.4105
R10595 GNDA_2.n1398 GNDA_2.n1391 3.4105
R10596 GNDA_2.n1398 GNDA_2.n1369 3.4105
R10597 GNDA_2.n1398 GNDA_2.n1392 3.4105
R10598 GNDA_2.n1398 GNDA_2.n1368 3.4105
R10599 GNDA_2.n1398 GNDA_2.n1393 3.4105
R10600 GNDA_2.n1398 GNDA_2.n1367 3.4105
R10601 GNDA_2.n1398 GNDA_2.n1394 3.4105
R10602 GNDA_2.n1398 GNDA_2.n1366 3.4105
R10603 GNDA_2.n1398 GNDA_2.n1395 3.4105
R10604 GNDA_2.n1398 GNDA_2.n1365 3.4105
R10605 GNDA_2.n1398 GNDA_2.n1396 3.4105
R10606 GNDA_2.n3512 GNDA_2.n1398 3.4105
R10607 GNDA_2.n3511 GNDA_2.n3492 3.4105
R10608 GNDA_2.n3511 GNDA_2.n1381 3.4105
R10609 GNDA_2.n3511 GNDA_2.n1379 3.4105
R10610 GNDA_2.n3511 GNDA_2.n1382 3.4105
R10611 GNDA_2.n3511 GNDA_2.n1378 3.4105
R10612 GNDA_2.n3511 GNDA_2.n1383 3.4105
R10613 GNDA_2.n3511 GNDA_2.n1377 3.4105
R10614 GNDA_2.n3511 GNDA_2.n1384 3.4105
R10615 GNDA_2.n3511 GNDA_2.n1376 3.4105
R10616 GNDA_2.n3511 GNDA_2.n1385 3.4105
R10617 GNDA_2.n3511 GNDA_2.n1375 3.4105
R10618 GNDA_2.n3511 GNDA_2.n1386 3.4105
R10619 GNDA_2.n3511 GNDA_2.n1374 3.4105
R10620 GNDA_2.n3511 GNDA_2.n1387 3.4105
R10621 GNDA_2.n3511 GNDA_2.n1373 3.4105
R10622 GNDA_2.n3511 GNDA_2.n1388 3.4105
R10623 GNDA_2.n3511 GNDA_2.n1372 3.4105
R10624 GNDA_2.n3511 GNDA_2.n1389 3.4105
R10625 GNDA_2.n3511 GNDA_2.n1371 3.4105
R10626 GNDA_2.n3511 GNDA_2.n1390 3.4105
R10627 GNDA_2.n3511 GNDA_2.n1370 3.4105
R10628 GNDA_2.n3511 GNDA_2.n1391 3.4105
R10629 GNDA_2.n3511 GNDA_2.n1369 3.4105
R10630 GNDA_2.n3511 GNDA_2.n1392 3.4105
R10631 GNDA_2.n3511 GNDA_2.n1368 3.4105
R10632 GNDA_2.n3511 GNDA_2.n1393 3.4105
R10633 GNDA_2.n3511 GNDA_2.n1367 3.4105
R10634 GNDA_2.n3511 GNDA_2.n1394 3.4105
R10635 GNDA_2.n3511 GNDA_2.n1366 3.4105
R10636 GNDA_2.n3511 GNDA_2.n1395 3.4105
R10637 GNDA_2.n3511 GNDA_2.n1365 3.4105
R10638 GNDA_2.n3511 GNDA_2.n1396 3.4105
R10639 GNDA_2.n3512 GNDA_2.n3511 3.4105
R10640 GNDA_2.n3492 GNDA_2.n1397 3.4105
R10641 GNDA_2.n1397 GNDA_2.n1381 3.4105
R10642 GNDA_2.n1397 GNDA_2.n1379 3.4105
R10643 GNDA_2.n1397 GNDA_2.n1382 3.4105
R10644 GNDA_2.n1397 GNDA_2.n1378 3.4105
R10645 GNDA_2.n1397 GNDA_2.n1383 3.4105
R10646 GNDA_2.n1397 GNDA_2.n1377 3.4105
R10647 GNDA_2.n1397 GNDA_2.n1384 3.4105
R10648 GNDA_2.n1397 GNDA_2.n1376 3.4105
R10649 GNDA_2.n1397 GNDA_2.n1385 3.4105
R10650 GNDA_2.n1397 GNDA_2.n1375 3.4105
R10651 GNDA_2.n1397 GNDA_2.n1386 3.4105
R10652 GNDA_2.n1397 GNDA_2.n1374 3.4105
R10653 GNDA_2.n1397 GNDA_2.n1387 3.4105
R10654 GNDA_2.n1397 GNDA_2.n1373 3.4105
R10655 GNDA_2.n1397 GNDA_2.n1388 3.4105
R10656 GNDA_2.n1397 GNDA_2.n1372 3.4105
R10657 GNDA_2.n1397 GNDA_2.n1389 3.4105
R10658 GNDA_2.n1397 GNDA_2.n1371 3.4105
R10659 GNDA_2.n1397 GNDA_2.n1390 3.4105
R10660 GNDA_2.n1397 GNDA_2.n1370 3.4105
R10661 GNDA_2.n1397 GNDA_2.n1391 3.4105
R10662 GNDA_2.n1397 GNDA_2.n1369 3.4105
R10663 GNDA_2.n1397 GNDA_2.n1392 3.4105
R10664 GNDA_2.n1397 GNDA_2.n1368 3.4105
R10665 GNDA_2.n1397 GNDA_2.n1393 3.4105
R10666 GNDA_2.n1397 GNDA_2.n1367 3.4105
R10667 GNDA_2.n1397 GNDA_2.n1394 3.4105
R10668 GNDA_2.n1397 GNDA_2.n1366 3.4105
R10669 GNDA_2.n1397 GNDA_2.n1395 3.4105
R10670 GNDA_2.n1397 GNDA_2.n1365 3.4105
R10671 GNDA_2.n1397 GNDA_2.n1396 3.4105
R10672 GNDA_2.n3512 GNDA_2.n1397 3.4105
R10673 GNDA_2.n3513 GNDA_2.n1381 3.4105
R10674 GNDA_2.n3513 GNDA_2.n1379 3.4105
R10675 GNDA_2.n3513 GNDA_2.n1382 3.4105
R10676 GNDA_2.n3513 GNDA_2.n1378 3.4105
R10677 GNDA_2.n3513 GNDA_2.n1383 3.4105
R10678 GNDA_2.n3513 GNDA_2.n1377 3.4105
R10679 GNDA_2.n3513 GNDA_2.n1384 3.4105
R10680 GNDA_2.n3513 GNDA_2.n1376 3.4105
R10681 GNDA_2.n3513 GNDA_2.n1385 3.4105
R10682 GNDA_2.n3513 GNDA_2.n1375 3.4105
R10683 GNDA_2.n3513 GNDA_2.n1386 3.4105
R10684 GNDA_2.n3513 GNDA_2.n1374 3.4105
R10685 GNDA_2.n3513 GNDA_2.n1387 3.4105
R10686 GNDA_2.n3513 GNDA_2.n1373 3.4105
R10687 GNDA_2.n3513 GNDA_2.n1388 3.4105
R10688 GNDA_2.n3513 GNDA_2.n1372 3.4105
R10689 GNDA_2.n3513 GNDA_2.n1389 3.4105
R10690 GNDA_2.n3513 GNDA_2.n1371 3.4105
R10691 GNDA_2.n3513 GNDA_2.n1390 3.4105
R10692 GNDA_2.n3513 GNDA_2.n1370 3.4105
R10693 GNDA_2.n3513 GNDA_2.n1391 3.4105
R10694 GNDA_2.n3513 GNDA_2.n1369 3.4105
R10695 GNDA_2.n3513 GNDA_2.n1392 3.4105
R10696 GNDA_2.n3513 GNDA_2.n1368 3.4105
R10697 GNDA_2.n3513 GNDA_2.n1393 3.4105
R10698 GNDA_2.n3513 GNDA_2.n1367 3.4105
R10699 GNDA_2.n3513 GNDA_2.n1394 3.4105
R10700 GNDA_2.n3513 GNDA_2.n1366 3.4105
R10701 GNDA_2.n3513 GNDA_2.n1395 3.4105
R10702 GNDA_2.n3513 GNDA_2.n1365 3.4105
R10703 GNDA_2.n3513 GNDA_2.n1396 3.4105
R10704 GNDA_2.n3513 GNDA_2.n3512 3.4105
R10705 GNDA_2.n1363 GNDA_2.n1331 3.4105
R10706 GNDA_2.n1363 GNDA_2.n1347 3.4105
R10707 GNDA_2.n3551 GNDA_2.n1363 3.4105
R10708 GNDA_2.n3550 GNDA_2.n1332 3.4105
R10709 GNDA_2.n3550 GNDA_2.n1330 3.4105
R10710 GNDA_2.n3550 GNDA_2.n1333 3.4105
R10711 GNDA_2.n3550 GNDA_2.n1329 3.4105
R10712 GNDA_2.n3550 GNDA_2.n1334 3.4105
R10713 GNDA_2.n3550 GNDA_2.n1328 3.4105
R10714 GNDA_2.n3550 GNDA_2.n1335 3.4105
R10715 GNDA_2.n3550 GNDA_2.n1327 3.4105
R10716 GNDA_2.n3550 GNDA_2.n1336 3.4105
R10717 GNDA_2.n3550 GNDA_2.n1326 3.4105
R10718 GNDA_2.n3550 GNDA_2.n1337 3.4105
R10719 GNDA_2.n3550 GNDA_2.n1325 3.4105
R10720 GNDA_2.n3550 GNDA_2.n1338 3.4105
R10721 GNDA_2.n3550 GNDA_2.n1324 3.4105
R10722 GNDA_2.n3550 GNDA_2.n1339 3.4105
R10723 GNDA_2.n3550 GNDA_2.n1323 3.4105
R10724 GNDA_2.n3550 GNDA_2.n1340 3.4105
R10725 GNDA_2.n3550 GNDA_2.n1322 3.4105
R10726 GNDA_2.n3550 GNDA_2.n1341 3.4105
R10727 GNDA_2.n3550 GNDA_2.n1321 3.4105
R10728 GNDA_2.n3550 GNDA_2.n1342 3.4105
R10729 GNDA_2.n3550 GNDA_2.n1320 3.4105
R10730 GNDA_2.n3550 GNDA_2.n1343 3.4105
R10731 GNDA_2.n3550 GNDA_2.n1319 3.4105
R10732 GNDA_2.n3550 GNDA_2.n1344 3.4105
R10733 GNDA_2.n3550 GNDA_2.n1318 3.4105
R10734 GNDA_2.n3550 GNDA_2.n1345 3.4105
R10735 GNDA_2.n3550 GNDA_2.n1317 3.4105
R10736 GNDA_2.n3550 GNDA_2.n1346 3.4105
R10737 GNDA_2.n3550 GNDA_2.n1347 3.4105
R10738 GNDA_2.n3551 GNDA_2.n3550 3.4105
R10739 GNDA_2.n3553 GNDA_2.n1282 3.4105
R10740 GNDA_2.n1331 GNDA_2.n1282 3.4105
R10741 GNDA_2.n1332 GNDA_2.n1282 3.4105
R10742 GNDA_2.n1330 GNDA_2.n1282 3.4105
R10743 GNDA_2.n1333 GNDA_2.n1282 3.4105
R10744 GNDA_2.n1329 GNDA_2.n1282 3.4105
R10745 GNDA_2.n1334 GNDA_2.n1282 3.4105
R10746 GNDA_2.n1328 GNDA_2.n1282 3.4105
R10747 GNDA_2.n1335 GNDA_2.n1282 3.4105
R10748 GNDA_2.n1327 GNDA_2.n1282 3.4105
R10749 GNDA_2.n1336 GNDA_2.n1282 3.4105
R10750 GNDA_2.n1326 GNDA_2.n1282 3.4105
R10751 GNDA_2.n1337 GNDA_2.n1282 3.4105
R10752 GNDA_2.n1325 GNDA_2.n1282 3.4105
R10753 GNDA_2.n1338 GNDA_2.n1282 3.4105
R10754 GNDA_2.n1324 GNDA_2.n1282 3.4105
R10755 GNDA_2.n1339 GNDA_2.n1282 3.4105
R10756 GNDA_2.n1323 GNDA_2.n1282 3.4105
R10757 GNDA_2.n1340 GNDA_2.n1282 3.4105
R10758 GNDA_2.n1322 GNDA_2.n1282 3.4105
R10759 GNDA_2.n1341 GNDA_2.n1282 3.4105
R10760 GNDA_2.n1321 GNDA_2.n1282 3.4105
R10761 GNDA_2.n1342 GNDA_2.n1282 3.4105
R10762 GNDA_2.n1320 GNDA_2.n1282 3.4105
R10763 GNDA_2.n1343 GNDA_2.n1282 3.4105
R10764 GNDA_2.n1319 GNDA_2.n1282 3.4105
R10765 GNDA_2.n1344 GNDA_2.n1282 3.4105
R10766 GNDA_2.n1318 GNDA_2.n1282 3.4105
R10767 GNDA_2.n1345 GNDA_2.n1282 3.4105
R10768 GNDA_2.n1317 GNDA_2.n1282 3.4105
R10769 GNDA_2.n1346 GNDA_2.n1282 3.4105
R10770 GNDA_2.n1347 GNDA_2.n1282 3.4105
R10771 GNDA_2.n3551 GNDA_2.n1282 3.4105
R10772 GNDA_2.n3553 GNDA_2.n1285 3.4105
R10773 GNDA_2.n1331 GNDA_2.n1285 3.4105
R10774 GNDA_2.n1332 GNDA_2.n1285 3.4105
R10775 GNDA_2.n1330 GNDA_2.n1285 3.4105
R10776 GNDA_2.n1333 GNDA_2.n1285 3.4105
R10777 GNDA_2.n1329 GNDA_2.n1285 3.4105
R10778 GNDA_2.n1334 GNDA_2.n1285 3.4105
R10779 GNDA_2.n1328 GNDA_2.n1285 3.4105
R10780 GNDA_2.n1335 GNDA_2.n1285 3.4105
R10781 GNDA_2.n1327 GNDA_2.n1285 3.4105
R10782 GNDA_2.n1336 GNDA_2.n1285 3.4105
R10783 GNDA_2.n1326 GNDA_2.n1285 3.4105
R10784 GNDA_2.n1337 GNDA_2.n1285 3.4105
R10785 GNDA_2.n1325 GNDA_2.n1285 3.4105
R10786 GNDA_2.n1338 GNDA_2.n1285 3.4105
R10787 GNDA_2.n1324 GNDA_2.n1285 3.4105
R10788 GNDA_2.n1339 GNDA_2.n1285 3.4105
R10789 GNDA_2.n1323 GNDA_2.n1285 3.4105
R10790 GNDA_2.n1340 GNDA_2.n1285 3.4105
R10791 GNDA_2.n1322 GNDA_2.n1285 3.4105
R10792 GNDA_2.n1341 GNDA_2.n1285 3.4105
R10793 GNDA_2.n1321 GNDA_2.n1285 3.4105
R10794 GNDA_2.n1342 GNDA_2.n1285 3.4105
R10795 GNDA_2.n1320 GNDA_2.n1285 3.4105
R10796 GNDA_2.n1343 GNDA_2.n1285 3.4105
R10797 GNDA_2.n1319 GNDA_2.n1285 3.4105
R10798 GNDA_2.n1344 GNDA_2.n1285 3.4105
R10799 GNDA_2.n1318 GNDA_2.n1285 3.4105
R10800 GNDA_2.n1345 GNDA_2.n1285 3.4105
R10801 GNDA_2.n1317 GNDA_2.n1285 3.4105
R10802 GNDA_2.n1346 GNDA_2.n1285 3.4105
R10803 GNDA_2.n1347 GNDA_2.n1285 3.4105
R10804 GNDA_2.n3551 GNDA_2.n1285 3.4105
R10805 GNDA_2.n3553 GNDA_2.n1281 3.4105
R10806 GNDA_2.n1331 GNDA_2.n1281 3.4105
R10807 GNDA_2.n1332 GNDA_2.n1281 3.4105
R10808 GNDA_2.n1330 GNDA_2.n1281 3.4105
R10809 GNDA_2.n1333 GNDA_2.n1281 3.4105
R10810 GNDA_2.n1329 GNDA_2.n1281 3.4105
R10811 GNDA_2.n1334 GNDA_2.n1281 3.4105
R10812 GNDA_2.n1328 GNDA_2.n1281 3.4105
R10813 GNDA_2.n1335 GNDA_2.n1281 3.4105
R10814 GNDA_2.n1327 GNDA_2.n1281 3.4105
R10815 GNDA_2.n1336 GNDA_2.n1281 3.4105
R10816 GNDA_2.n1326 GNDA_2.n1281 3.4105
R10817 GNDA_2.n1337 GNDA_2.n1281 3.4105
R10818 GNDA_2.n1325 GNDA_2.n1281 3.4105
R10819 GNDA_2.n1338 GNDA_2.n1281 3.4105
R10820 GNDA_2.n1324 GNDA_2.n1281 3.4105
R10821 GNDA_2.n1339 GNDA_2.n1281 3.4105
R10822 GNDA_2.n1323 GNDA_2.n1281 3.4105
R10823 GNDA_2.n1340 GNDA_2.n1281 3.4105
R10824 GNDA_2.n1322 GNDA_2.n1281 3.4105
R10825 GNDA_2.n1341 GNDA_2.n1281 3.4105
R10826 GNDA_2.n1321 GNDA_2.n1281 3.4105
R10827 GNDA_2.n1342 GNDA_2.n1281 3.4105
R10828 GNDA_2.n1320 GNDA_2.n1281 3.4105
R10829 GNDA_2.n1343 GNDA_2.n1281 3.4105
R10830 GNDA_2.n1319 GNDA_2.n1281 3.4105
R10831 GNDA_2.n1344 GNDA_2.n1281 3.4105
R10832 GNDA_2.n1318 GNDA_2.n1281 3.4105
R10833 GNDA_2.n1345 GNDA_2.n1281 3.4105
R10834 GNDA_2.n1317 GNDA_2.n1281 3.4105
R10835 GNDA_2.n1346 GNDA_2.n1281 3.4105
R10836 GNDA_2.n1347 GNDA_2.n1281 3.4105
R10837 GNDA_2.n3551 GNDA_2.n1281 3.4105
R10838 GNDA_2.n3553 GNDA_2.n1286 3.4105
R10839 GNDA_2.n1331 GNDA_2.n1286 3.4105
R10840 GNDA_2.n1332 GNDA_2.n1286 3.4105
R10841 GNDA_2.n1330 GNDA_2.n1286 3.4105
R10842 GNDA_2.n1333 GNDA_2.n1286 3.4105
R10843 GNDA_2.n1329 GNDA_2.n1286 3.4105
R10844 GNDA_2.n1334 GNDA_2.n1286 3.4105
R10845 GNDA_2.n1328 GNDA_2.n1286 3.4105
R10846 GNDA_2.n1335 GNDA_2.n1286 3.4105
R10847 GNDA_2.n1327 GNDA_2.n1286 3.4105
R10848 GNDA_2.n1336 GNDA_2.n1286 3.4105
R10849 GNDA_2.n1326 GNDA_2.n1286 3.4105
R10850 GNDA_2.n1337 GNDA_2.n1286 3.4105
R10851 GNDA_2.n1325 GNDA_2.n1286 3.4105
R10852 GNDA_2.n1338 GNDA_2.n1286 3.4105
R10853 GNDA_2.n1324 GNDA_2.n1286 3.4105
R10854 GNDA_2.n1339 GNDA_2.n1286 3.4105
R10855 GNDA_2.n1323 GNDA_2.n1286 3.4105
R10856 GNDA_2.n1340 GNDA_2.n1286 3.4105
R10857 GNDA_2.n1322 GNDA_2.n1286 3.4105
R10858 GNDA_2.n1341 GNDA_2.n1286 3.4105
R10859 GNDA_2.n1321 GNDA_2.n1286 3.4105
R10860 GNDA_2.n1342 GNDA_2.n1286 3.4105
R10861 GNDA_2.n1320 GNDA_2.n1286 3.4105
R10862 GNDA_2.n1343 GNDA_2.n1286 3.4105
R10863 GNDA_2.n1319 GNDA_2.n1286 3.4105
R10864 GNDA_2.n1344 GNDA_2.n1286 3.4105
R10865 GNDA_2.n1318 GNDA_2.n1286 3.4105
R10866 GNDA_2.n1345 GNDA_2.n1286 3.4105
R10867 GNDA_2.n1317 GNDA_2.n1286 3.4105
R10868 GNDA_2.n1346 GNDA_2.n1286 3.4105
R10869 GNDA_2.n1347 GNDA_2.n1286 3.4105
R10870 GNDA_2.n3551 GNDA_2.n1286 3.4105
R10871 GNDA_2.n3553 GNDA_2.n1280 3.4105
R10872 GNDA_2.n1331 GNDA_2.n1280 3.4105
R10873 GNDA_2.n1332 GNDA_2.n1280 3.4105
R10874 GNDA_2.n1330 GNDA_2.n1280 3.4105
R10875 GNDA_2.n1333 GNDA_2.n1280 3.4105
R10876 GNDA_2.n1329 GNDA_2.n1280 3.4105
R10877 GNDA_2.n1334 GNDA_2.n1280 3.4105
R10878 GNDA_2.n1328 GNDA_2.n1280 3.4105
R10879 GNDA_2.n1335 GNDA_2.n1280 3.4105
R10880 GNDA_2.n1327 GNDA_2.n1280 3.4105
R10881 GNDA_2.n1336 GNDA_2.n1280 3.4105
R10882 GNDA_2.n1326 GNDA_2.n1280 3.4105
R10883 GNDA_2.n1337 GNDA_2.n1280 3.4105
R10884 GNDA_2.n1325 GNDA_2.n1280 3.4105
R10885 GNDA_2.n1338 GNDA_2.n1280 3.4105
R10886 GNDA_2.n1324 GNDA_2.n1280 3.4105
R10887 GNDA_2.n1339 GNDA_2.n1280 3.4105
R10888 GNDA_2.n1323 GNDA_2.n1280 3.4105
R10889 GNDA_2.n1340 GNDA_2.n1280 3.4105
R10890 GNDA_2.n1322 GNDA_2.n1280 3.4105
R10891 GNDA_2.n1341 GNDA_2.n1280 3.4105
R10892 GNDA_2.n1321 GNDA_2.n1280 3.4105
R10893 GNDA_2.n1342 GNDA_2.n1280 3.4105
R10894 GNDA_2.n1320 GNDA_2.n1280 3.4105
R10895 GNDA_2.n1343 GNDA_2.n1280 3.4105
R10896 GNDA_2.n1319 GNDA_2.n1280 3.4105
R10897 GNDA_2.n1344 GNDA_2.n1280 3.4105
R10898 GNDA_2.n1318 GNDA_2.n1280 3.4105
R10899 GNDA_2.n1345 GNDA_2.n1280 3.4105
R10900 GNDA_2.n1317 GNDA_2.n1280 3.4105
R10901 GNDA_2.n1346 GNDA_2.n1280 3.4105
R10902 GNDA_2.n1347 GNDA_2.n1280 3.4105
R10903 GNDA_2.n3551 GNDA_2.n1280 3.4105
R10904 GNDA_2.n3553 GNDA_2.n1287 3.4105
R10905 GNDA_2.n1331 GNDA_2.n1287 3.4105
R10906 GNDA_2.n1332 GNDA_2.n1287 3.4105
R10907 GNDA_2.n1330 GNDA_2.n1287 3.4105
R10908 GNDA_2.n1333 GNDA_2.n1287 3.4105
R10909 GNDA_2.n1329 GNDA_2.n1287 3.4105
R10910 GNDA_2.n1334 GNDA_2.n1287 3.4105
R10911 GNDA_2.n1328 GNDA_2.n1287 3.4105
R10912 GNDA_2.n1335 GNDA_2.n1287 3.4105
R10913 GNDA_2.n1327 GNDA_2.n1287 3.4105
R10914 GNDA_2.n1336 GNDA_2.n1287 3.4105
R10915 GNDA_2.n1326 GNDA_2.n1287 3.4105
R10916 GNDA_2.n1337 GNDA_2.n1287 3.4105
R10917 GNDA_2.n1325 GNDA_2.n1287 3.4105
R10918 GNDA_2.n1338 GNDA_2.n1287 3.4105
R10919 GNDA_2.n1324 GNDA_2.n1287 3.4105
R10920 GNDA_2.n1339 GNDA_2.n1287 3.4105
R10921 GNDA_2.n1323 GNDA_2.n1287 3.4105
R10922 GNDA_2.n1340 GNDA_2.n1287 3.4105
R10923 GNDA_2.n1322 GNDA_2.n1287 3.4105
R10924 GNDA_2.n1341 GNDA_2.n1287 3.4105
R10925 GNDA_2.n1321 GNDA_2.n1287 3.4105
R10926 GNDA_2.n1342 GNDA_2.n1287 3.4105
R10927 GNDA_2.n1320 GNDA_2.n1287 3.4105
R10928 GNDA_2.n1343 GNDA_2.n1287 3.4105
R10929 GNDA_2.n1319 GNDA_2.n1287 3.4105
R10930 GNDA_2.n1344 GNDA_2.n1287 3.4105
R10931 GNDA_2.n1318 GNDA_2.n1287 3.4105
R10932 GNDA_2.n1345 GNDA_2.n1287 3.4105
R10933 GNDA_2.n1317 GNDA_2.n1287 3.4105
R10934 GNDA_2.n1346 GNDA_2.n1287 3.4105
R10935 GNDA_2.n1347 GNDA_2.n1287 3.4105
R10936 GNDA_2.n3551 GNDA_2.n1287 3.4105
R10937 GNDA_2.n3553 GNDA_2.n1279 3.4105
R10938 GNDA_2.n1331 GNDA_2.n1279 3.4105
R10939 GNDA_2.n1332 GNDA_2.n1279 3.4105
R10940 GNDA_2.n1330 GNDA_2.n1279 3.4105
R10941 GNDA_2.n1333 GNDA_2.n1279 3.4105
R10942 GNDA_2.n1329 GNDA_2.n1279 3.4105
R10943 GNDA_2.n1334 GNDA_2.n1279 3.4105
R10944 GNDA_2.n1328 GNDA_2.n1279 3.4105
R10945 GNDA_2.n1335 GNDA_2.n1279 3.4105
R10946 GNDA_2.n1327 GNDA_2.n1279 3.4105
R10947 GNDA_2.n1336 GNDA_2.n1279 3.4105
R10948 GNDA_2.n1326 GNDA_2.n1279 3.4105
R10949 GNDA_2.n1337 GNDA_2.n1279 3.4105
R10950 GNDA_2.n1325 GNDA_2.n1279 3.4105
R10951 GNDA_2.n1338 GNDA_2.n1279 3.4105
R10952 GNDA_2.n1324 GNDA_2.n1279 3.4105
R10953 GNDA_2.n1339 GNDA_2.n1279 3.4105
R10954 GNDA_2.n1323 GNDA_2.n1279 3.4105
R10955 GNDA_2.n1340 GNDA_2.n1279 3.4105
R10956 GNDA_2.n1322 GNDA_2.n1279 3.4105
R10957 GNDA_2.n1341 GNDA_2.n1279 3.4105
R10958 GNDA_2.n1321 GNDA_2.n1279 3.4105
R10959 GNDA_2.n1342 GNDA_2.n1279 3.4105
R10960 GNDA_2.n1320 GNDA_2.n1279 3.4105
R10961 GNDA_2.n1343 GNDA_2.n1279 3.4105
R10962 GNDA_2.n1319 GNDA_2.n1279 3.4105
R10963 GNDA_2.n1344 GNDA_2.n1279 3.4105
R10964 GNDA_2.n1318 GNDA_2.n1279 3.4105
R10965 GNDA_2.n1345 GNDA_2.n1279 3.4105
R10966 GNDA_2.n1317 GNDA_2.n1279 3.4105
R10967 GNDA_2.n1346 GNDA_2.n1279 3.4105
R10968 GNDA_2.n1347 GNDA_2.n1279 3.4105
R10969 GNDA_2.n3551 GNDA_2.n1279 3.4105
R10970 GNDA_2.n3553 GNDA_2.n1288 3.4105
R10971 GNDA_2.n1331 GNDA_2.n1288 3.4105
R10972 GNDA_2.n1332 GNDA_2.n1288 3.4105
R10973 GNDA_2.n1330 GNDA_2.n1288 3.4105
R10974 GNDA_2.n1333 GNDA_2.n1288 3.4105
R10975 GNDA_2.n1329 GNDA_2.n1288 3.4105
R10976 GNDA_2.n1334 GNDA_2.n1288 3.4105
R10977 GNDA_2.n1328 GNDA_2.n1288 3.4105
R10978 GNDA_2.n1335 GNDA_2.n1288 3.4105
R10979 GNDA_2.n1327 GNDA_2.n1288 3.4105
R10980 GNDA_2.n1336 GNDA_2.n1288 3.4105
R10981 GNDA_2.n1326 GNDA_2.n1288 3.4105
R10982 GNDA_2.n1337 GNDA_2.n1288 3.4105
R10983 GNDA_2.n1325 GNDA_2.n1288 3.4105
R10984 GNDA_2.n1338 GNDA_2.n1288 3.4105
R10985 GNDA_2.n1324 GNDA_2.n1288 3.4105
R10986 GNDA_2.n1339 GNDA_2.n1288 3.4105
R10987 GNDA_2.n1323 GNDA_2.n1288 3.4105
R10988 GNDA_2.n1340 GNDA_2.n1288 3.4105
R10989 GNDA_2.n1322 GNDA_2.n1288 3.4105
R10990 GNDA_2.n1341 GNDA_2.n1288 3.4105
R10991 GNDA_2.n1321 GNDA_2.n1288 3.4105
R10992 GNDA_2.n1342 GNDA_2.n1288 3.4105
R10993 GNDA_2.n1320 GNDA_2.n1288 3.4105
R10994 GNDA_2.n1343 GNDA_2.n1288 3.4105
R10995 GNDA_2.n1319 GNDA_2.n1288 3.4105
R10996 GNDA_2.n1344 GNDA_2.n1288 3.4105
R10997 GNDA_2.n1318 GNDA_2.n1288 3.4105
R10998 GNDA_2.n1345 GNDA_2.n1288 3.4105
R10999 GNDA_2.n1317 GNDA_2.n1288 3.4105
R11000 GNDA_2.n1346 GNDA_2.n1288 3.4105
R11001 GNDA_2.n1347 GNDA_2.n1288 3.4105
R11002 GNDA_2.n3551 GNDA_2.n1288 3.4105
R11003 GNDA_2.n3553 GNDA_2.n1278 3.4105
R11004 GNDA_2.n1331 GNDA_2.n1278 3.4105
R11005 GNDA_2.n1332 GNDA_2.n1278 3.4105
R11006 GNDA_2.n1330 GNDA_2.n1278 3.4105
R11007 GNDA_2.n1333 GNDA_2.n1278 3.4105
R11008 GNDA_2.n1329 GNDA_2.n1278 3.4105
R11009 GNDA_2.n1334 GNDA_2.n1278 3.4105
R11010 GNDA_2.n1328 GNDA_2.n1278 3.4105
R11011 GNDA_2.n1335 GNDA_2.n1278 3.4105
R11012 GNDA_2.n1327 GNDA_2.n1278 3.4105
R11013 GNDA_2.n1336 GNDA_2.n1278 3.4105
R11014 GNDA_2.n1326 GNDA_2.n1278 3.4105
R11015 GNDA_2.n1337 GNDA_2.n1278 3.4105
R11016 GNDA_2.n1325 GNDA_2.n1278 3.4105
R11017 GNDA_2.n1338 GNDA_2.n1278 3.4105
R11018 GNDA_2.n1324 GNDA_2.n1278 3.4105
R11019 GNDA_2.n1339 GNDA_2.n1278 3.4105
R11020 GNDA_2.n1323 GNDA_2.n1278 3.4105
R11021 GNDA_2.n1340 GNDA_2.n1278 3.4105
R11022 GNDA_2.n1322 GNDA_2.n1278 3.4105
R11023 GNDA_2.n1341 GNDA_2.n1278 3.4105
R11024 GNDA_2.n1321 GNDA_2.n1278 3.4105
R11025 GNDA_2.n1342 GNDA_2.n1278 3.4105
R11026 GNDA_2.n1320 GNDA_2.n1278 3.4105
R11027 GNDA_2.n1343 GNDA_2.n1278 3.4105
R11028 GNDA_2.n1319 GNDA_2.n1278 3.4105
R11029 GNDA_2.n1344 GNDA_2.n1278 3.4105
R11030 GNDA_2.n1318 GNDA_2.n1278 3.4105
R11031 GNDA_2.n1345 GNDA_2.n1278 3.4105
R11032 GNDA_2.n1317 GNDA_2.n1278 3.4105
R11033 GNDA_2.n1346 GNDA_2.n1278 3.4105
R11034 GNDA_2.n1347 GNDA_2.n1278 3.4105
R11035 GNDA_2.n3551 GNDA_2.n1278 3.4105
R11036 GNDA_2.n3553 GNDA_2.n1289 3.4105
R11037 GNDA_2.n1331 GNDA_2.n1289 3.4105
R11038 GNDA_2.n1332 GNDA_2.n1289 3.4105
R11039 GNDA_2.n1330 GNDA_2.n1289 3.4105
R11040 GNDA_2.n1333 GNDA_2.n1289 3.4105
R11041 GNDA_2.n1329 GNDA_2.n1289 3.4105
R11042 GNDA_2.n1334 GNDA_2.n1289 3.4105
R11043 GNDA_2.n1328 GNDA_2.n1289 3.4105
R11044 GNDA_2.n1335 GNDA_2.n1289 3.4105
R11045 GNDA_2.n1327 GNDA_2.n1289 3.4105
R11046 GNDA_2.n1336 GNDA_2.n1289 3.4105
R11047 GNDA_2.n1326 GNDA_2.n1289 3.4105
R11048 GNDA_2.n1337 GNDA_2.n1289 3.4105
R11049 GNDA_2.n1325 GNDA_2.n1289 3.4105
R11050 GNDA_2.n1338 GNDA_2.n1289 3.4105
R11051 GNDA_2.n1324 GNDA_2.n1289 3.4105
R11052 GNDA_2.n1339 GNDA_2.n1289 3.4105
R11053 GNDA_2.n1323 GNDA_2.n1289 3.4105
R11054 GNDA_2.n1340 GNDA_2.n1289 3.4105
R11055 GNDA_2.n1322 GNDA_2.n1289 3.4105
R11056 GNDA_2.n1341 GNDA_2.n1289 3.4105
R11057 GNDA_2.n1321 GNDA_2.n1289 3.4105
R11058 GNDA_2.n1342 GNDA_2.n1289 3.4105
R11059 GNDA_2.n1320 GNDA_2.n1289 3.4105
R11060 GNDA_2.n1343 GNDA_2.n1289 3.4105
R11061 GNDA_2.n1319 GNDA_2.n1289 3.4105
R11062 GNDA_2.n1344 GNDA_2.n1289 3.4105
R11063 GNDA_2.n1318 GNDA_2.n1289 3.4105
R11064 GNDA_2.n1345 GNDA_2.n1289 3.4105
R11065 GNDA_2.n1317 GNDA_2.n1289 3.4105
R11066 GNDA_2.n1346 GNDA_2.n1289 3.4105
R11067 GNDA_2.n1347 GNDA_2.n1289 3.4105
R11068 GNDA_2.n3551 GNDA_2.n1289 3.4105
R11069 GNDA_2.n3553 GNDA_2.n1277 3.4105
R11070 GNDA_2.n1331 GNDA_2.n1277 3.4105
R11071 GNDA_2.n1332 GNDA_2.n1277 3.4105
R11072 GNDA_2.n1330 GNDA_2.n1277 3.4105
R11073 GNDA_2.n1333 GNDA_2.n1277 3.4105
R11074 GNDA_2.n1329 GNDA_2.n1277 3.4105
R11075 GNDA_2.n1334 GNDA_2.n1277 3.4105
R11076 GNDA_2.n1328 GNDA_2.n1277 3.4105
R11077 GNDA_2.n1335 GNDA_2.n1277 3.4105
R11078 GNDA_2.n1327 GNDA_2.n1277 3.4105
R11079 GNDA_2.n1336 GNDA_2.n1277 3.4105
R11080 GNDA_2.n1326 GNDA_2.n1277 3.4105
R11081 GNDA_2.n1337 GNDA_2.n1277 3.4105
R11082 GNDA_2.n1325 GNDA_2.n1277 3.4105
R11083 GNDA_2.n1338 GNDA_2.n1277 3.4105
R11084 GNDA_2.n1324 GNDA_2.n1277 3.4105
R11085 GNDA_2.n1339 GNDA_2.n1277 3.4105
R11086 GNDA_2.n1323 GNDA_2.n1277 3.4105
R11087 GNDA_2.n1340 GNDA_2.n1277 3.4105
R11088 GNDA_2.n1322 GNDA_2.n1277 3.4105
R11089 GNDA_2.n1341 GNDA_2.n1277 3.4105
R11090 GNDA_2.n1321 GNDA_2.n1277 3.4105
R11091 GNDA_2.n1342 GNDA_2.n1277 3.4105
R11092 GNDA_2.n1320 GNDA_2.n1277 3.4105
R11093 GNDA_2.n1343 GNDA_2.n1277 3.4105
R11094 GNDA_2.n1319 GNDA_2.n1277 3.4105
R11095 GNDA_2.n1344 GNDA_2.n1277 3.4105
R11096 GNDA_2.n1318 GNDA_2.n1277 3.4105
R11097 GNDA_2.n1345 GNDA_2.n1277 3.4105
R11098 GNDA_2.n1317 GNDA_2.n1277 3.4105
R11099 GNDA_2.n1346 GNDA_2.n1277 3.4105
R11100 GNDA_2.n1347 GNDA_2.n1277 3.4105
R11101 GNDA_2.n3551 GNDA_2.n1277 3.4105
R11102 GNDA_2.n3553 GNDA_2.n1290 3.4105
R11103 GNDA_2.n1331 GNDA_2.n1290 3.4105
R11104 GNDA_2.n1332 GNDA_2.n1290 3.4105
R11105 GNDA_2.n1330 GNDA_2.n1290 3.4105
R11106 GNDA_2.n1333 GNDA_2.n1290 3.4105
R11107 GNDA_2.n1329 GNDA_2.n1290 3.4105
R11108 GNDA_2.n1334 GNDA_2.n1290 3.4105
R11109 GNDA_2.n1328 GNDA_2.n1290 3.4105
R11110 GNDA_2.n1335 GNDA_2.n1290 3.4105
R11111 GNDA_2.n1327 GNDA_2.n1290 3.4105
R11112 GNDA_2.n1336 GNDA_2.n1290 3.4105
R11113 GNDA_2.n1326 GNDA_2.n1290 3.4105
R11114 GNDA_2.n1337 GNDA_2.n1290 3.4105
R11115 GNDA_2.n1325 GNDA_2.n1290 3.4105
R11116 GNDA_2.n1338 GNDA_2.n1290 3.4105
R11117 GNDA_2.n1324 GNDA_2.n1290 3.4105
R11118 GNDA_2.n1339 GNDA_2.n1290 3.4105
R11119 GNDA_2.n1323 GNDA_2.n1290 3.4105
R11120 GNDA_2.n1340 GNDA_2.n1290 3.4105
R11121 GNDA_2.n1322 GNDA_2.n1290 3.4105
R11122 GNDA_2.n1341 GNDA_2.n1290 3.4105
R11123 GNDA_2.n1321 GNDA_2.n1290 3.4105
R11124 GNDA_2.n1342 GNDA_2.n1290 3.4105
R11125 GNDA_2.n1320 GNDA_2.n1290 3.4105
R11126 GNDA_2.n1343 GNDA_2.n1290 3.4105
R11127 GNDA_2.n1319 GNDA_2.n1290 3.4105
R11128 GNDA_2.n1344 GNDA_2.n1290 3.4105
R11129 GNDA_2.n1318 GNDA_2.n1290 3.4105
R11130 GNDA_2.n1345 GNDA_2.n1290 3.4105
R11131 GNDA_2.n1317 GNDA_2.n1290 3.4105
R11132 GNDA_2.n1346 GNDA_2.n1290 3.4105
R11133 GNDA_2.n1347 GNDA_2.n1290 3.4105
R11134 GNDA_2.n3551 GNDA_2.n1290 3.4105
R11135 GNDA_2.n3553 GNDA_2.n1276 3.4105
R11136 GNDA_2.n1331 GNDA_2.n1276 3.4105
R11137 GNDA_2.n1332 GNDA_2.n1276 3.4105
R11138 GNDA_2.n1330 GNDA_2.n1276 3.4105
R11139 GNDA_2.n1333 GNDA_2.n1276 3.4105
R11140 GNDA_2.n1329 GNDA_2.n1276 3.4105
R11141 GNDA_2.n1334 GNDA_2.n1276 3.4105
R11142 GNDA_2.n1328 GNDA_2.n1276 3.4105
R11143 GNDA_2.n1335 GNDA_2.n1276 3.4105
R11144 GNDA_2.n1327 GNDA_2.n1276 3.4105
R11145 GNDA_2.n1336 GNDA_2.n1276 3.4105
R11146 GNDA_2.n1326 GNDA_2.n1276 3.4105
R11147 GNDA_2.n1337 GNDA_2.n1276 3.4105
R11148 GNDA_2.n1325 GNDA_2.n1276 3.4105
R11149 GNDA_2.n1338 GNDA_2.n1276 3.4105
R11150 GNDA_2.n1324 GNDA_2.n1276 3.4105
R11151 GNDA_2.n1339 GNDA_2.n1276 3.4105
R11152 GNDA_2.n1323 GNDA_2.n1276 3.4105
R11153 GNDA_2.n1340 GNDA_2.n1276 3.4105
R11154 GNDA_2.n1322 GNDA_2.n1276 3.4105
R11155 GNDA_2.n1341 GNDA_2.n1276 3.4105
R11156 GNDA_2.n1321 GNDA_2.n1276 3.4105
R11157 GNDA_2.n1342 GNDA_2.n1276 3.4105
R11158 GNDA_2.n1320 GNDA_2.n1276 3.4105
R11159 GNDA_2.n1343 GNDA_2.n1276 3.4105
R11160 GNDA_2.n1319 GNDA_2.n1276 3.4105
R11161 GNDA_2.n1344 GNDA_2.n1276 3.4105
R11162 GNDA_2.n1318 GNDA_2.n1276 3.4105
R11163 GNDA_2.n1345 GNDA_2.n1276 3.4105
R11164 GNDA_2.n1317 GNDA_2.n1276 3.4105
R11165 GNDA_2.n1346 GNDA_2.n1276 3.4105
R11166 GNDA_2.n1347 GNDA_2.n1276 3.4105
R11167 GNDA_2.n3551 GNDA_2.n1276 3.4105
R11168 GNDA_2.n3553 GNDA_2.n1291 3.4105
R11169 GNDA_2.n1331 GNDA_2.n1291 3.4105
R11170 GNDA_2.n1332 GNDA_2.n1291 3.4105
R11171 GNDA_2.n1330 GNDA_2.n1291 3.4105
R11172 GNDA_2.n1333 GNDA_2.n1291 3.4105
R11173 GNDA_2.n1329 GNDA_2.n1291 3.4105
R11174 GNDA_2.n1334 GNDA_2.n1291 3.4105
R11175 GNDA_2.n1328 GNDA_2.n1291 3.4105
R11176 GNDA_2.n1335 GNDA_2.n1291 3.4105
R11177 GNDA_2.n1327 GNDA_2.n1291 3.4105
R11178 GNDA_2.n1336 GNDA_2.n1291 3.4105
R11179 GNDA_2.n1326 GNDA_2.n1291 3.4105
R11180 GNDA_2.n1337 GNDA_2.n1291 3.4105
R11181 GNDA_2.n1325 GNDA_2.n1291 3.4105
R11182 GNDA_2.n1338 GNDA_2.n1291 3.4105
R11183 GNDA_2.n1324 GNDA_2.n1291 3.4105
R11184 GNDA_2.n1339 GNDA_2.n1291 3.4105
R11185 GNDA_2.n1323 GNDA_2.n1291 3.4105
R11186 GNDA_2.n1340 GNDA_2.n1291 3.4105
R11187 GNDA_2.n1322 GNDA_2.n1291 3.4105
R11188 GNDA_2.n1341 GNDA_2.n1291 3.4105
R11189 GNDA_2.n1321 GNDA_2.n1291 3.4105
R11190 GNDA_2.n1342 GNDA_2.n1291 3.4105
R11191 GNDA_2.n1320 GNDA_2.n1291 3.4105
R11192 GNDA_2.n1343 GNDA_2.n1291 3.4105
R11193 GNDA_2.n1319 GNDA_2.n1291 3.4105
R11194 GNDA_2.n1344 GNDA_2.n1291 3.4105
R11195 GNDA_2.n1318 GNDA_2.n1291 3.4105
R11196 GNDA_2.n1345 GNDA_2.n1291 3.4105
R11197 GNDA_2.n1317 GNDA_2.n1291 3.4105
R11198 GNDA_2.n1346 GNDA_2.n1291 3.4105
R11199 GNDA_2.n1347 GNDA_2.n1291 3.4105
R11200 GNDA_2.n3551 GNDA_2.n1291 3.4105
R11201 GNDA_2.n3553 GNDA_2.n1275 3.4105
R11202 GNDA_2.n1331 GNDA_2.n1275 3.4105
R11203 GNDA_2.n1332 GNDA_2.n1275 3.4105
R11204 GNDA_2.n1330 GNDA_2.n1275 3.4105
R11205 GNDA_2.n1333 GNDA_2.n1275 3.4105
R11206 GNDA_2.n1329 GNDA_2.n1275 3.4105
R11207 GNDA_2.n1334 GNDA_2.n1275 3.4105
R11208 GNDA_2.n1328 GNDA_2.n1275 3.4105
R11209 GNDA_2.n1335 GNDA_2.n1275 3.4105
R11210 GNDA_2.n1327 GNDA_2.n1275 3.4105
R11211 GNDA_2.n1336 GNDA_2.n1275 3.4105
R11212 GNDA_2.n1326 GNDA_2.n1275 3.4105
R11213 GNDA_2.n1337 GNDA_2.n1275 3.4105
R11214 GNDA_2.n1325 GNDA_2.n1275 3.4105
R11215 GNDA_2.n1338 GNDA_2.n1275 3.4105
R11216 GNDA_2.n1324 GNDA_2.n1275 3.4105
R11217 GNDA_2.n1339 GNDA_2.n1275 3.4105
R11218 GNDA_2.n1323 GNDA_2.n1275 3.4105
R11219 GNDA_2.n1340 GNDA_2.n1275 3.4105
R11220 GNDA_2.n1322 GNDA_2.n1275 3.4105
R11221 GNDA_2.n1341 GNDA_2.n1275 3.4105
R11222 GNDA_2.n1321 GNDA_2.n1275 3.4105
R11223 GNDA_2.n1342 GNDA_2.n1275 3.4105
R11224 GNDA_2.n1320 GNDA_2.n1275 3.4105
R11225 GNDA_2.n1343 GNDA_2.n1275 3.4105
R11226 GNDA_2.n1319 GNDA_2.n1275 3.4105
R11227 GNDA_2.n1344 GNDA_2.n1275 3.4105
R11228 GNDA_2.n1318 GNDA_2.n1275 3.4105
R11229 GNDA_2.n1345 GNDA_2.n1275 3.4105
R11230 GNDA_2.n1317 GNDA_2.n1275 3.4105
R11231 GNDA_2.n1346 GNDA_2.n1275 3.4105
R11232 GNDA_2.n1347 GNDA_2.n1275 3.4105
R11233 GNDA_2.n3551 GNDA_2.n1275 3.4105
R11234 GNDA_2.n3553 GNDA_2.n1292 3.4105
R11235 GNDA_2.n1331 GNDA_2.n1292 3.4105
R11236 GNDA_2.n1332 GNDA_2.n1292 3.4105
R11237 GNDA_2.n1330 GNDA_2.n1292 3.4105
R11238 GNDA_2.n1333 GNDA_2.n1292 3.4105
R11239 GNDA_2.n1329 GNDA_2.n1292 3.4105
R11240 GNDA_2.n1334 GNDA_2.n1292 3.4105
R11241 GNDA_2.n1328 GNDA_2.n1292 3.4105
R11242 GNDA_2.n1335 GNDA_2.n1292 3.4105
R11243 GNDA_2.n1327 GNDA_2.n1292 3.4105
R11244 GNDA_2.n1336 GNDA_2.n1292 3.4105
R11245 GNDA_2.n1326 GNDA_2.n1292 3.4105
R11246 GNDA_2.n1337 GNDA_2.n1292 3.4105
R11247 GNDA_2.n1325 GNDA_2.n1292 3.4105
R11248 GNDA_2.n1338 GNDA_2.n1292 3.4105
R11249 GNDA_2.n1324 GNDA_2.n1292 3.4105
R11250 GNDA_2.n1339 GNDA_2.n1292 3.4105
R11251 GNDA_2.n1323 GNDA_2.n1292 3.4105
R11252 GNDA_2.n1340 GNDA_2.n1292 3.4105
R11253 GNDA_2.n1322 GNDA_2.n1292 3.4105
R11254 GNDA_2.n1341 GNDA_2.n1292 3.4105
R11255 GNDA_2.n1321 GNDA_2.n1292 3.4105
R11256 GNDA_2.n1342 GNDA_2.n1292 3.4105
R11257 GNDA_2.n1320 GNDA_2.n1292 3.4105
R11258 GNDA_2.n1343 GNDA_2.n1292 3.4105
R11259 GNDA_2.n1319 GNDA_2.n1292 3.4105
R11260 GNDA_2.n1344 GNDA_2.n1292 3.4105
R11261 GNDA_2.n1318 GNDA_2.n1292 3.4105
R11262 GNDA_2.n1345 GNDA_2.n1292 3.4105
R11263 GNDA_2.n1317 GNDA_2.n1292 3.4105
R11264 GNDA_2.n1346 GNDA_2.n1292 3.4105
R11265 GNDA_2.n1347 GNDA_2.n1292 3.4105
R11266 GNDA_2.n3551 GNDA_2.n1292 3.4105
R11267 GNDA_2.n3553 GNDA_2.n1274 3.4105
R11268 GNDA_2.n1331 GNDA_2.n1274 3.4105
R11269 GNDA_2.n1332 GNDA_2.n1274 3.4105
R11270 GNDA_2.n1330 GNDA_2.n1274 3.4105
R11271 GNDA_2.n1333 GNDA_2.n1274 3.4105
R11272 GNDA_2.n1329 GNDA_2.n1274 3.4105
R11273 GNDA_2.n1334 GNDA_2.n1274 3.4105
R11274 GNDA_2.n1328 GNDA_2.n1274 3.4105
R11275 GNDA_2.n1335 GNDA_2.n1274 3.4105
R11276 GNDA_2.n1327 GNDA_2.n1274 3.4105
R11277 GNDA_2.n1336 GNDA_2.n1274 3.4105
R11278 GNDA_2.n1326 GNDA_2.n1274 3.4105
R11279 GNDA_2.n1337 GNDA_2.n1274 3.4105
R11280 GNDA_2.n1325 GNDA_2.n1274 3.4105
R11281 GNDA_2.n1338 GNDA_2.n1274 3.4105
R11282 GNDA_2.n1324 GNDA_2.n1274 3.4105
R11283 GNDA_2.n1339 GNDA_2.n1274 3.4105
R11284 GNDA_2.n1323 GNDA_2.n1274 3.4105
R11285 GNDA_2.n1340 GNDA_2.n1274 3.4105
R11286 GNDA_2.n1322 GNDA_2.n1274 3.4105
R11287 GNDA_2.n1341 GNDA_2.n1274 3.4105
R11288 GNDA_2.n1321 GNDA_2.n1274 3.4105
R11289 GNDA_2.n1342 GNDA_2.n1274 3.4105
R11290 GNDA_2.n1320 GNDA_2.n1274 3.4105
R11291 GNDA_2.n1343 GNDA_2.n1274 3.4105
R11292 GNDA_2.n1319 GNDA_2.n1274 3.4105
R11293 GNDA_2.n1344 GNDA_2.n1274 3.4105
R11294 GNDA_2.n1318 GNDA_2.n1274 3.4105
R11295 GNDA_2.n1345 GNDA_2.n1274 3.4105
R11296 GNDA_2.n1317 GNDA_2.n1274 3.4105
R11297 GNDA_2.n1346 GNDA_2.n1274 3.4105
R11298 GNDA_2.n1347 GNDA_2.n1274 3.4105
R11299 GNDA_2.n3551 GNDA_2.n1274 3.4105
R11300 GNDA_2.n3553 GNDA_2.n1293 3.4105
R11301 GNDA_2.n1331 GNDA_2.n1293 3.4105
R11302 GNDA_2.n1332 GNDA_2.n1293 3.4105
R11303 GNDA_2.n1330 GNDA_2.n1293 3.4105
R11304 GNDA_2.n1333 GNDA_2.n1293 3.4105
R11305 GNDA_2.n1329 GNDA_2.n1293 3.4105
R11306 GNDA_2.n1334 GNDA_2.n1293 3.4105
R11307 GNDA_2.n1328 GNDA_2.n1293 3.4105
R11308 GNDA_2.n1335 GNDA_2.n1293 3.4105
R11309 GNDA_2.n1327 GNDA_2.n1293 3.4105
R11310 GNDA_2.n1336 GNDA_2.n1293 3.4105
R11311 GNDA_2.n1326 GNDA_2.n1293 3.4105
R11312 GNDA_2.n1337 GNDA_2.n1293 3.4105
R11313 GNDA_2.n1325 GNDA_2.n1293 3.4105
R11314 GNDA_2.n1338 GNDA_2.n1293 3.4105
R11315 GNDA_2.n1324 GNDA_2.n1293 3.4105
R11316 GNDA_2.n1339 GNDA_2.n1293 3.4105
R11317 GNDA_2.n1323 GNDA_2.n1293 3.4105
R11318 GNDA_2.n1340 GNDA_2.n1293 3.4105
R11319 GNDA_2.n1322 GNDA_2.n1293 3.4105
R11320 GNDA_2.n1341 GNDA_2.n1293 3.4105
R11321 GNDA_2.n1321 GNDA_2.n1293 3.4105
R11322 GNDA_2.n1342 GNDA_2.n1293 3.4105
R11323 GNDA_2.n1320 GNDA_2.n1293 3.4105
R11324 GNDA_2.n1343 GNDA_2.n1293 3.4105
R11325 GNDA_2.n1319 GNDA_2.n1293 3.4105
R11326 GNDA_2.n1344 GNDA_2.n1293 3.4105
R11327 GNDA_2.n1318 GNDA_2.n1293 3.4105
R11328 GNDA_2.n1345 GNDA_2.n1293 3.4105
R11329 GNDA_2.n1317 GNDA_2.n1293 3.4105
R11330 GNDA_2.n1346 GNDA_2.n1293 3.4105
R11331 GNDA_2.n1347 GNDA_2.n1293 3.4105
R11332 GNDA_2.n3551 GNDA_2.n1293 3.4105
R11333 GNDA_2.n3553 GNDA_2.n1273 3.4105
R11334 GNDA_2.n1331 GNDA_2.n1273 3.4105
R11335 GNDA_2.n1332 GNDA_2.n1273 3.4105
R11336 GNDA_2.n1330 GNDA_2.n1273 3.4105
R11337 GNDA_2.n1333 GNDA_2.n1273 3.4105
R11338 GNDA_2.n1329 GNDA_2.n1273 3.4105
R11339 GNDA_2.n1334 GNDA_2.n1273 3.4105
R11340 GNDA_2.n1328 GNDA_2.n1273 3.4105
R11341 GNDA_2.n1335 GNDA_2.n1273 3.4105
R11342 GNDA_2.n1327 GNDA_2.n1273 3.4105
R11343 GNDA_2.n1336 GNDA_2.n1273 3.4105
R11344 GNDA_2.n1326 GNDA_2.n1273 3.4105
R11345 GNDA_2.n1337 GNDA_2.n1273 3.4105
R11346 GNDA_2.n1325 GNDA_2.n1273 3.4105
R11347 GNDA_2.n1338 GNDA_2.n1273 3.4105
R11348 GNDA_2.n1324 GNDA_2.n1273 3.4105
R11349 GNDA_2.n1339 GNDA_2.n1273 3.4105
R11350 GNDA_2.n1323 GNDA_2.n1273 3.4105
R11351 GNDA_2.n1340 GNDA_2.n1273 3.4105
R11352 GNDA_2.n1322 GNDA_2.n1273 3.4105
R11353 GNDA_2.n1341 GNDA_2.n1273 3.4105
R11354 GNDA_2.n1321 GNDA_2.n1273 3.4105
R11355 GNDA_2.n1342 GNDA_2.n1273 3.4105
R11356 GNDA_2.n1320 GNDA_2.n1273 3.4105
R11357 GNDA_2.n1343 GNDA_2.n1273 3.4105
R11358 GNDA_2.n1319 GNDA_2.n1273 3.4105
R11359 GNDA_2.n1344 GNDA_2.n1273 3.4105
R11360 GNDA_2.n1318 GNDA_2.n1273 3.4105
R11361 GNDA_2.n1345 GNDA_2.n1273 3.4105
R11362 GNDA_2.n1317 GNDA_2.n1273 3.4105
R11363 GNDA_2.n1346 GNDA_2.n1273 3.4105
R11364 GNDA_2.n1347 GNDA_2.n1273 3.4105
R11365 GNDA_2.n3551 GNDA_2.n1273 3.4105
R11366 GNDA_2.n3553 GNDA_2.n1294 3.4105
R11367 GNDA_2.n1331 GNDA_2.n1294 3.4105
R11368 GNDA_2.n1332 GNDA_2.n1294 3.4105
R11369 GNDA_2.n1330 GNDA_2.n1294 3.4105
R11370 GNDA_2.n1333 GNDA_2.n1294 3.4105
R11371 GNDA_2.n1329 GNDA_2.n1294 3.4105
R11372 GNDA_2.n1334 GNDA_2.n1294 3.4105
R11373 GNDA_2.n1328 GNDA_2.n1294 3.4105
R11374 GNDA_2.n1335 GNDA_2.n1294 3.4105
R11375 GNDA_2.n1327 GNDA_2.n1294 3.4105
R11376 GNDA_2.n1336 GNDA_2.n1294 3.4105
R11377 GNDA_2.n1326 GNDA_2.n1294 3.4105
R11378 GNDA_2.n1337 GNDA_2.n1294 3.4105
R11379 GNDA_2.n1325 GNDA_2.n1294 3.4105
R11380 GNDA_2.n1338 GNDA_2.n1294 3.4105
R11381 GNDA_2.n1324 GNDA_2.n1294 3.4105
R11382 GNDA_2.n1339 GNDA_2.n1294 3.4105
R11383 GNDA_2.n1323 GNDA_2.n1294 3.4105
R11384 GNDA_2.n1340 GNDA_2.n1294 3.4105
R11385 GNDA_2.n1322 GNDA_2.n1294 3.4105
R11386 GNDA_2.n1341 GNDA_2.n1294 3.4105
R11387 GNDA_2.n1321 GNDA_2.n1294 3.4105
R11388 GNDA_2.n1342 GNDA_2.n1294 3.4105
R11389 GNDA_2.n1320 GNDA_2.n1294 3.4105
R11390 GNDA_2.n1343 GNDA_2.n1294 3.4105
R11391 GNDA_2.n1319 GNDA_2.n1294 3.4105
R11392 GNDA_2.n1344 GNDA_2.n1294 3.4105
R11393 GNDA_2.n1318 GNDA_2.n1294 3.4105
R11394 GNDA_2.n1345 GNDA_2.n1294 3.4105
R11395 GNDA_2.n1317 GNDA_2.n1294 3.4105
R11396 GNDA_2.n1346 GNDA_2.n1294 3.4105
R11397 GNDA_2.n1347 GNDA_2.n1294 3.4105
R11398 GNDA_2.n3551 GNDA_2.n1294 3.4105
R11399 GNDA_2.n3553 GNDA_2.n1272 3.4105
R11400 GNDA_2.n1331 GNDA_2.n1272 3.4105
R11401 GNDA_2.n1332 GNDA_2.n1272 3.4105
R11402 GNDA_2.n1330 GNDA_2.n1272 3.4105
R11403 GNDA_2.n1333 GNDA_2.n1272 3.4105
R11404 GNDA_2.n1329 GNDA_2.n1272 3.4105
R11405 GNDA_2.n1334 GNDA_2.n1272 3.4105
R11406 GNDA_2.n1328 GNDA_2.n1272 3.4105
R11407 GNDA_2.n1335 GNDA_2.n1272 3.4105
R11408 GNDA_2.n1327 GNDA_2.n1272 3.4105
R11409 GNDA_2.n1336 GNDA_2.n1272 3.4105
R11410 GNDA_2.n1326 GNDA_2.n1272 3.4105
R11411 GNDA_2.n1337 GNDA_2.n1272 3.4105
R11412 GNDA_2.n1325 GNDA_2.n1272 3.4105
R11413 GNDA_2.n1338 GNDA_2.n1272 3.4105
R11414 GNDA_2.n1324 GNDA_2.n1272 3.4105
R11415 GNDA_2.n1339 GNDA_2.n1272 3.4105
R11416 GNDA_2.n1323 GNDA_2.n1272 3.4105
R11417 GNDA_2.n1340 GNDA_2.n1272 3.4105
R11418 GNDA_2.n1322 GNDA_2.n1272 3.4105
R11419 GNDA_2.n1341 GNDA_2.n1272 3.4105
R11420 GNDA_2.n1321 GNDA_2.n1272 3.4105
R11421 GNDA_2.n1342 GNDA_2.n1272 3.4105
R11422 GNDA_2.n1320 GNDA_2.n1272 3.4105
R11423 GNDA_2.n1343 GNDA_2.n1272 3.4105
R11424 GNDA_2.n1319 GNDA_2.n1272 3.4105
R11425 GNDA_2.n1344 GNDA_2.n1272 3.4105
R11426 GNDA_2.n1318 GNDA_2.n1272 3.4105
R11427 GNDA_2.n1345 GNDA_2.n1272 3.4105
R11428 GNDA_2.n1317 GNDA_2.n1272 3.4105
R11429 GNDA_2.n1346 GNDA_2.n1272 3.4105
R11430 GNDA_2.n1347 GNDA_2.n1272 3.4105
R11431 GNDA_2.n3551 GNDA_2.n1272 3.4105
R11432 GNDA_2.n3553 GNDA_2.n1295 3.4105
R11433 GNDA_2.n1331 GNDA_2.n1295 3.4105
R11434 GNDA_2.n1332 GNDA_2.n1295 3.4105
R11435 GNDA_2.n1330 GNDA_2.n1295 3.4105
R11436 GNDA_2.n1333 GNDA_2.n1295 3.4105
R11437 GNDA_2.n1329 GNDA_2.n1295 3.4105
R11438 GNDA_2.n1334 GNDA_2.n1295 3.4105
R11439 GNDA_2.n1328 GNDA_2.n1295 3.4105
R11440 GNDA_2.n1335 GNDA_2.n1295 3.4105
R11441 GNDA_2.n1327 GNDA_2.n1295 3.4105
R11442 GNDA_2.n1336 GNDA_2.n1295 3.4105
R11443 GNDA_2.n1326 GNDA_2.n1295 3.4105
R11444 GNDA_2.n1337 GNDA_2.n1295 3.4105
R11445 GNDA_2.n1325 GNDA_2.n1295 3.4105
R11446 GNDA_2.n1338 GNDA_2.n1295 3.4105
R11447 GNDA_2.n1324 GNDA_2.n1295 3.4105
R11448 GNDA_2.n1339 GNDA_2.n1295 3.4105
R11449 GNDA_2.n1323 GNDA_2.n1295 3.4105
R11450 GNDA_2.n1340 GNDA_2.n1295 3.4105
R11451 GNDA_2.n1322 GNDA_2.n1295 3.4105
R11452 GNDA_2.n1341 GNDA_2.n1295 3.4105
R11453 GNDA_2.n1321 GNDA_2.n1295 3.4105
R11454 GNDA_2.n1342 GNDA_2.n1295 3.4105
R11455 GNDA_2.n1320 GNDA_2.n1295 3.4105
R11456 GNDA_2.n1343 GNDA_2.n1295 3.4105
R11457 GNDA_2.n1319 GNDA_2.n1295 3.4105
R11458 GNDA_2.n1344 GNDA_2.n1295 3.4105
R11459 GNDA_2.n1318 GNDA_2.n1295 3.4105
R11460 GNDA_2.n1345 GNDA_2.n1295 3.4105
R11461 GNDA_2.n1317 GNDA_2.n1295 3.4105
R11462 GNDA_2.n1346 GNDA_2.n1295 3.4105
R11463 GNDA_2.n1347 GNDA_2.n1295 3.4105
R11464 GNDA_2.n3551 GNDA_2.n1295 3.4105
R11465 GNDA_2.n3553 GNDA_2.n1271 3.4105
R11466 GNDA_2.n1331 GNDA_2.n1271 3.4105
R11467 GNDA_2.n1332 GNDA_2.n1271 3.4105
R11468 GNDA_2.n1330 GNDA_2.n1271 3.4105
R11469 GNDA_2.n1333 GNDA_2.n1271 3.4105
R11470 GNDA_2.n1329 GNDA_2.n1271 3.4105
R11471 GNDA_2.n1334 GNDA_2.n1271 3.4105
R11472 GNDA_2.n1328 GNDA_2.n1271 3.4105
R11473 GNDA_2.n1335 GNDA_2.n1271 3.4105
R11474 GNDA_2.n1327 GNDA_2.n1271 3.4105
R11475 GNDA_2.n1336 GNDA_2.n1271 3.4105
R11476 GNDA_2.n1326 GNDA_2.n1271 3.4105
R11477 GNDA_2.n1337 GNDA_2.n1271 3.4105
R11478 GNDA_2.n1325 GNDA_2.n1271 3.4105
R11479 GNDA_2.n1338 GNDA_2.n1271 3.4105
R11480 GNDA_2.n1324 GNDA_2.n1271 3.4105
R11481 GNDA_2.n1339 GNDA_2.n1271 3.4105
R11482 GNDA_2.n1323 GNDA_2.n1271 3.4105
R11483 GNDA_2.n1340 GNDA_2.n1271 3.4105
R11484 GNDA_2.n1322 GNDA_2.n1271 3.4105
R11485 GNDA_2.n1341 GNDA_2.n1271 3.4105
R11486 GNDA_2.n1321 GNDA_2.n1271 3.4105
R11487 GNDA_2.n1342 GNDA_2.n1271 3.4105
R11488 GNDA_2.n1320 GNDA_2.n1271 3.4105
R11489 GNDA_2.n1343 GNDA_2.n1271 3.4105
R11490 GNDA_2.n1319 GNDA_2.n1271 3.4105
R11491 GNDA_2.n1344 GNDA_2.n1271 3.4105
R11492 GNDA_2.n1318 GNDA_2.n1271 3.4105
R11493 GNDA_2.n1345 GNDA_2.n1271 3.4105
R11494 GNDA_2.n1317 GNDA_2.n1271 3.4105
R11495 GNDA_2.n1346 GNDA_2.n1271 3.4105
R11496 GNDA_2.n1347 GNDA_2.n1271 3.4105
R11497 GNDA_2.n3551 GNDA_2.n1271 3.4105
R11498 GNDA_2.n3553 GNDA_2.n1296 3.4105
R11499 GNDA_2.n1331 GNDA_2.n1296 3.4105
R11500 GNDA_2.n1332 GNDA_2.n1296 3.4105
R11501 GNDA_2.n1330 GNDA_2.n1296 3.4105
R11502 GNDA_2.n1333 GNDA_2.n1296 3.4105
R11503 GNDA_2.n1329 GNDA_2.n1296 3.4105
R11504 GNDA_2.n1334 GNDA_2.n1296 3.4105
R11505 GNDA_2.n1328 GNDA_2.n1296 3.4105
R11506 GNDA_2.n1335 GNDA_2.n1296 3.4105
R11507 GNDA_2.n1327 GNDA_2.n1296 3.4105
R11508 GNDA_2.n1336 GNDA_2.n1296 3.4105
R11509 GNDA_2.n1326 GNDA_2.n1296 3.4105
R11510 GNDA_2.n1337 GNDA_2.n1296 3.4105
R11511 GNDA_2.n1325 GNDA_2.n1296 3.4105
R11512 GNDA_2.n1338 GNDA_2.n1296 3.4105
R11513 GNDA_2.n1324 GNDA_2.n1296 3.4105
R11514 GNDA_2.n1339 GNDA_2.n1296 3.4105
R11515 GNDA_2.n1323 GNDA_2.n1296 3.4105
R11516 GNDA_2.n1340 GNDA_2.n1296 3.4105
R11517 GNDA_2.n1322 GNDA_2.n1296 3.4105
R11518 GNDA_2.n1341 GNDA_2.n1296 3.4105
R11519 GNDA_2.n1321 GNDA_2.n1296 3.4105
R11520 GNDA_2.n1342 GNDA_2.n1296 3.4105
R11521 GNDA_2.n1320 GNDA_2.n1296 3.4105
R11522 GNDA_2.n1343 GNDA_2.n1296 3.4105
R11523 GNDA_2.n1319 GNDA_2.n1296 3.4105
R11524 GNDA_2.n1344 GNDA_2.n1296 3.4105
R11525 GNDA_2.n1318 GNDA_2.n1296 3.4105
R11526 GNDA_2.n1345 GNDA_2.n1296 3.4105
R11527 GNDA_2.n1317 GNDA_2.n1296 3.4105
R11528 GNDA_2.n1346 GNDA_2.n1296 3.4105
R11529 GNDA_2.n1347 GNDA_2.n1296 3.4105
R11530 GNDA_2.n3551 GNDA_2.n1296 3.4105
R11531 GNDA_2.n3553 GNDA_2.n1270 3.4105
R11532 GNDA_2.n1331 GNDA_2.n1270 3.4105
R11533 GNDA_2.n1332 GNDA_2.n1270 3.4105
R11534 GNDA_2.n1330 GNDA_2.n1270 3.4105
R11535 GNDA_2.n1333 GNDA_2.n1270 3.4105
R11536 GNDA_2.n1329 GNDA_2.n1270 3.4105
R11537 GNDA_2.n1334 GNDA_2.n1270 3.4105
R11538 GNDA_2.n1328 GNDA_2.n1270 3.4105
R11539 GNDA_2.n1335 GNDA_2.n1270 3.4105
R11540 GNDA_2.n1327 GNDA_2.n1270 3.4105
R11541 GNDA_2.n1336 GNDA_2.n1270 3.4105
R11542 GNDA_2.n1326 GNDA_2.n1270 3.4105
R11543 GNDA_2.n1337 GNDA_2.n1270 3.4105
R11544 GNDA_2.n1325 GNDA_2.n1270 3.4105
R11545 GNDA_2.n1338 GNDA_2.n1270 3.4105
R11546 GNDA_2.n1324 GNDA_2.n1270 3.4105
R11547 GNDA_2.n1339 GNDA_2.n1270 3.4105
R11548 GNDA_2.n1323 GNDA_2.n1270 3.4105
R11549 GNDA_2.n1340 GNDA_2.n1270 3.4105
R11550 GNDA_2.n1322 GNDA_2.n1270 3.4105
R11551 GNDA_2.n1341 GNDA_2.n1270 3.4105
R11552 GNDA_2.n1321 GNDA_2.n1270 3.4105
R11553 GNDA_2.n1342 GNDA_2.n1270 3.4105
R11554 GNDA_2.n1320 GNDA_2.n1270 3.4105
R11555 GNDA_2.n1343 GNDA_2.n1270 3.4105
R11556 GNDA_2.n1319 GNDA_2.n1270 3.4105
R11557 GNDA_2.n1344 GNDA_2.n1270 3.4105
R11558 GNDA_2.n1318 GNDA_2.n1270 3.4105
R11559 GNDA_2.n1345 GNDA_2.n1270 3.4105
R11560 GNDA_2.n1317 GNDA_2.n1270 3.4105
R11561 GNDA_2.n1346 GNDA_2.n1270 3.4105
R11562 GNDA_2.n1347 GNDA_2.n1270 3.4105
R11563 GNDA_2.n3551 GNDA_2.n1270 3.4105
R11564 GNDA_2.n3553 GNDA_2.n1297 3.4105
R11565 GNDA_2.n1331 GNDA_2.n1297 3.4105
R11566 GNDA_2.n1332 GNDA_2.n1297 3.4105
R11567 GNDA_2.n1330 GNDA_2.n1297 3.4105
R11568 GNDA_2.n1333 GNDA_2.n1297 3.4105
R11569 GNDA_2.n1329 GNDA_2.n1297 3.4105
R11570 GNDA_2.n1334 GNDA_2.n1297 3.4105
R11571 GNDA_2.n1328 GNDA_2.n1297 3.4105
R11572 GNDA_2.n1335 GNDA_2.n1297 3.4105
R11573 GNDA_2.n1327 GNDA_2.n1297 3.4105
R11574 GNDA_2.n1336 GNDA_2.n1297 3.4105
R11575 GNDA_2.n1326 GNDA_2.n1297 3.4105
R11576 GNDA_2.n1337 GNDA_2.n1297 3.4105
R11577 GNDA_2.n1325 GNDA_2.n1297 3.4105
R11578 GNDA_2.n1338 GNDA_2.n1297 3.4105
R11579 GNDA_2.n1324 GNDA_2.n1297 3.4105
R11580 GNDA_2.n1339 GNDA_2.n1297 3.4105
R11581 GNDA_2.n1323 GNDA_2.n1297 3.4105
R11582 GNDA_2.n1340 GNDA_2.n1297 3.4105
R11583 GNDA_2.n1322 GNDA_2.n1297 3.4105
R11584 GNDA_2.n1341 GNDA_2.n1297 3.4105
R11585 GNDA_2.n1321 GNDA_2.n1297 3.4105
R11586 GNDA_2.n1342 GNDA_2.n1297 3.4105
R11587 GNDA_2.n1320 GNDA_2.n1297 3.4105
R11588 GNDA_2.n1343 GNDA_2.n1297 3.4105
R11589 GNDA_2.n1319 GNDA_2.n1297 3.4105
R11590 GNDA_2.n1344 GNDA_2.n1297 3.4105
R11591 GNDA_2.n1318 GNDA_2.n1297 3.4105
R11592 GNDA_2.n1345 GNDA_2.n1297 3.4105
R11593 GNDA_2.n1317 GNDA_2.n1297 3.4105
R11594 GNDA_2.n1346 GNDA_2.n1297 3.4105
R11595 GNDA_2.n1347 GNDA_2.n1297 3.4105
R11596 GNDA_2.n3551 GNDA_2.n1297 3.4105
R11597 GNDA_2.n3553 GNDA_2.n1269 3.4105
R11598 GNDA_2.n1331 GNDA_2.n1269 3.4105
R11599 GNDA_2.n1332 GNDA_2.n1269 3.4105
R11600 GNDA_2.n1330 GNDA_2.n1269 3.4105
R11601 GNDA_2.n1333 GNDA_2.n1269 3.4105
R11602 GNDA_2.n1329 GNDA_2.n1269 3.4105
R11603 GNDA_2.n1334 GNDA_2.n1269 3.4105
R11604 GNDA_2.n1328 GNDA_2.n1269 3.4105
R11605 GNDA_2.n1335 GNDA_2.n1269 3.4105
R11606 GNDA_2.n1327 GNDA_2.n1269 3.4105
R11607 GNDA_2.n1336 GNDA_2.n1269 3.4105
R11608 GNDA_2.n1326 GNDA_2.n1269 3.4105
R11609 GNDA_2.n1337 GNDA_2.n1269 3.4105
R11610 GNDA_2.n1325 GNDA_2.n1269 3.4105
R11611 GNDA_2.n1338 GNDA_2.n1269 3.4105
R11612 GNDA_2.n1324 GNDA_2.n1269 3.4105
R11613 GNDA_2.n1339 GNDA_2.n1269 3.4105
R11614 GNDA_2.n1323 GNDA_2.n1269 3.4105
R11615 GNDA_2.n1340 GNDA_2.n1269 3.4105
R11616 GNDA_2.n1322 GNDA_2.n1269 3.4105
R11617 GNDA_2.n1341 GNDA_2.n1269 3.4105
R11618 GNDA_2.n1321 GNDA_2.n1269 3.4105
R11619 GNDA_2.n1342 GNDA_2.n1269 3.4105
R11620 GNDA_2.n1320 GNDA_2.n1269 3.4105
R11621 GNDA_2.n1343 GNDA_2.n1269 3.4105
R11622 GNDA_2.n1319 GNDA_2.n1269 3.4105
R11623 GNDA_2.n1344 GNDA_2.n1269 3.4105
R11624 GNDA_2.n1318 GNDA_2.n1269 3.4105
R11625 GNDA_2.n1345 GNDA_2.n1269 3.4105
R11626 GNDA_2.n1317 GNDA_2.n1269 3.4105
R11627 GNDA_2.n1346 GNDA_2.n1269 3.4105
R11628 GNDA_2.n1347 GNDA_2.n1269 3.4105
R11629 GNDA_2.n3551 GNDA_2.n1269 3.4105
R11630 GNDA_2.n3553 GNDA_2.n1298 3.4105
R11631 GNDA_2.n1331 GNDA_2.n1298 3.4105
R11632 GNDA_2.n1332 GNDA_2.n1298 3.4105
R11633 GNDA_2.n1330 GNDA_2.n1298 3.4105
R11634 GNDA_2.n1333 GNDA_2.n1298 3.4105
R11635 GNDA_2.n1329 GNDA_2.n1298 3.4105
R11636 GNDA_2.n1334 GNDA_2.n1298 3.4105
R11637 GNDA_2.n1328 GNDA_2.n1298 3.4105
R11638 GNDA_2.n1335 GNDA_2.n1298 3.4105
R11639 GNDA_2.n1327 GNDA_2.n1298 3.4105
R11640 GNDA_2.n1336 GNDA_2.n1298 3.4105
R11641 GNDA_2.n1326 GNDA_2.n1298 3.4105
R11642 GNDA_2.n1337 GNDA_2.n1298 3.4105
R11643 GNDA_2.n1325 GNDA_2.n1298 3.4105
R11644 GNDA_2.n1338 GNDA_2.n1298 3.4105
R11645 GNDA_2.n1324 GNDA_2.n1298 3.4105
R11646 GNDA_2.n1339 GNDA_2.n1298 3.4105
R11647 GNDA_2.n1323 GNDA_2.n1298 3.4105
R11648 GNDA_2.n1340 GNDA_2.n1298 3.4105
R11649 GNDA_2.n1322 GNDA_2.n1298 3.4105
R11650 GNDA_2.n1341 GNDA_2.n1298 3.4105
R11651 GNDA_2.n1321 GNDA_2.n1298 3.4105
R11652 GNDA_2.n1342 GNDA_2.n1298 3.4105
R11653 GNDA_2.n1320 GNDA_2.n1298 3.4105
R11654 GNDA_2.n1343 GNDA_2.n1298 3.4105
R11655 GNDA_2.n1319 GNDA_2.n1298 3.4105
R11656 GNDA_2.n1344 GNDA_2.n1298 3.4105
R11657 GNDA_2.n1318 GNDA_2.n1298 3.4105
R11658 GNDA_2.n1345 GNDA_2.n1298 3.4105
R11659 GNDA_2.n1317 GNDA_2.n1298 3.4105
R11660 GNDA_2.n1346 GNDA_2.n1298 3.4105
R11661 GNDA_2.n1347 GNDA_2.n1298 3.4105
R11662 GNDA_2.n3551 GNDA_2.n1298 3.4105
R11663 GNDA_2.n3553 GNDA_2.n1268 3.4105
R11664 GNDA_2.n1331 GNDA_2.n1268 3.4105
R11665 GNDA_2.n1332 GNDA_2.n1268 3.4105
R11666 GNDA_2.n1330 GNDA_2.n1268 3.4105
R11667 GNDA_2.n1333 GNDA_2.n1268 3.4105
R11668 GNDA_2.n1329 GNDA_2.n1268 3.4105
R11669 GNDA_2.n1334 GNDA_2.n1268 3.4105
R11670 GNDA_2.n1328 GNDA_2.n1268 3.4105
R11671 GNDA_2.n1335 GNDA_2.n1268 3.4105
R11672 GNDA_2.n1327 GNDA_2.n1268 3.4105
R11673 GNDA_2.n1336 GNDA_2.n1268 3.4105
R11674 GNDA_2.n1326 GNDA_2.n1268 3.4105
R11675 GNDA_2.n1337 GNDA_2.n1268 3.4105
R11676 GNDA_2.n1325 GNDA_2.n1268 3.4105
R11677 GNDA_2.n1338 GNDA_2.n1268 3.4105
R11678 GNDA_2.n1324 GNDA_2.n1268 3.4105
R11679 GNDA_2.n1339 GNDA_2.n1268 3.4105
R11680 GNDA_2.n1323 GNDA_2.n1268 3.4105
R11681 GNDA_2.n1340 GNDA_2.n1268 3.4105
R11682 GNDA_2.n1322 GNDA_2.n1268 3.4105
R11683 GNDA_2.n1341 GNDA_2.n1268 3.4105
R11684 GNDA_2.n1321 GNDA_2.n1268 3.4105
R11685 GNDA_2.n1342 GNDA_2.n1268 3.4105
R11686 GNDA_2.n1320 GNDA_2.n1268 3.4105
R11687 GNDA_2.n1343 GNDA_2.n1268 3.4105
R11688 GNDA_2.n1319 GNDA_2.n1268 3.4105
R11689 GNDA_2.n1344 GNDA_2.n1268 3.4105
R11690 GNDA_2.n1318 GNDA_2.n1268 3.4105
R11691 GNDA_2.n1345 GNDA_2.n1268 3.4105
R11692 GNDA_2.n1317 GNDA_2.n1268 3.4105
R11693 GNDA_2.n1346 GNDA_2.n1268 3.4105
R11694 GNDA_2.n1347 GNDA_2.n1268 3.4105
R11695 GNDA_2.n3551 GNDA_2.n1268 3.4105
R11696 GNDA_2.n3553 GNDA_2.n1299 3.4105
R11697 GNDA_2.n1331 GNDA_2.n1299 3.4105
R11698 GNDA_2.n1332 GNDA_2.n1299 3.4105
R11699 GNDA_2.n1330 GNDA_2.n1299 3.4105
R11700 GNDA_2.n1333 GNDA_2.n1299 3.4105
R11701 GNDA_2.n1329 GNDA_2.n1299 3.4105
R11702 GNDA_2.n1334 GNDA_2.n1299 3.4105
R11703 GNDA_2.n1328 GNDA_2.n1299 3.4105
R11704 GNDA_2.n1335 GNDA_2.n1299 3.4105
R11705 GNDA_2.n1327 GNDA_2.n1299 3.4105
R11706 GNDA_2.n1336 GNDA_2.n1299 3.4105
R11707 GNDA_2.n1326 GNDA_2.n1299 3.4105
R11708 GNDA_2.n1337 GNDA_2.n1299 3.4105
R11709 GNDA_2.n1325 GNDA_2.n1299 3.4105
R11710 GNDA_2.n1338 GNDA_2.n1299 3.4105
R11711 GNDA_2.n1324 GNDA_2.n1299 3.4105
R11712 GNDA_2.n1339 GNDA_2.n1299 3.4105
R11713 GNDA_2.n1323 GNDA_2.n1299 3.4105
R11714 GNDA_2.n1340 GNDA_2.n1299 3.4105
R11715 GNDA_2.n1322 GNDA_2.n1299 3.4105
R11716 GNDA_2.n1341 GNDA_2.n1299 3.4105
R11717 GNDA_2.n1321 GNDA_2.n1299 3.4105
R11718 GNDA_2.n1342 GNDA_2.n1299 3.4105
R11719 GNDA_2.n1320 GNDA_2.n1299 3.4105
R11720 GNDA_2.n1343 GNDA_2.n1299 3.4105
R11721 GNDA_2.n1319 GNDA_2.n1299 3.4105
R11722 GNDA_2.n1344 GNDA_2.n1299 3.4105
R11723 GNDA_2.n1318 GNDA_2.n1299 3.4105
R11724 GNDA_2.n1345 GNDA_2.n1299 3.4105
R11725 GNDA_2.n1317 GNDA_2.n1299 3.4105
R11726 GNDA_2.n1346 GNDA_2.n1299 3.4105
R11727 GNDA_2.n1347 GNDA_2.n1299 3.4105
R11728 GNDA_2.n3551 GNDA_2.n1299 3.4105
R11729 GNDA_2.n3553 GNDA_2.n1267 3.4105
R11730 GNDA_2.n1331 GNDA_2.n1267 3.4105
R11731 GNDA_2.n1332 GNDA_2.n1267 3.4105
R11732 GNDA_2.n1330 GNDA_2.n1267 3.4105
R11733 GNDA_2.n1333 GNDA_2.n1267 3.4105
R11734 GNDA_2.n1329 GNDA_2.n1267 3.4105
R11735 GNDA_2.n1334 GNDA_2.n1267 3.4105
R11736 GNDA_2.n1328 GNDA_2.n1267 3.4105
R11737 GNDA_2.n1335 GNDA_2.n1267 3.4105
R11738 GNDA_2.n1327 GNDA_2.n1267 3.4105
R11739 GNDA_2.n1336 GNDA_2.n1267 3.4105
R11740 GNDA_2.n1326 GNDA_2.n1267 3.4105
R11741 GNDA_2.n1337 GNDA_2.n1267 3.4105
R11742 GNDA_2.n1325 GNDA_2.n1267 3.4105
R11743 GNDA_2.n1338 GNDA_2.n1267 3.4105
R11744 GNDA_2.n1324 GNDA_2.n1267 3.4105
R11745 GNDA_2.n1339 GNDA_2.n1267 3.4105
R11746 GNDA_2.n1323 GNDA_2.n1267 3.4105
R11747 GNDA_2.n1340 GNDA_2.n1267 3.4105
R11748 GNDA_2.n1322 GNDA_2.n1267 3.4105
R11749 GNDA_2.n1341 GNDA_2.n1267 3.4105
R11750 GNDA_2.n1321 GNDA_2.n1267 3.4105
R11751 GNDA_2.n1342 GNDA_2.n1267 3.4105
R11752 GNDA_2.n1320 GNDA_2.n1267 3.4105
R11753 GNDA_2.n1343 GNDA_2.n1267 3.4105
R11754 GNDA_2.n1319 GNDA_2.n1267 3.4105
R11755 GNDA_2.n1344 GNDA_2.n1267 3.4105
R11756 GNDA_2.n1318 GNDA_2.n1267 3.4105
R11757 GNDA_2.n1345 GNDA_2.n1267 3.4105
R11758 GNDA_2.n1317 GNDA_2.n1267 3.4105
R11759 GNDA_2.n1346 GNDA_2.n1267 3.4105
R11760 GNDA_2.n1347 GNDA_2.n1267 3.4105
R11761 GNDA_2.n3551 GNDA_2.n1267 3.4105
R11762 GNDA_2.n3553 GNDA_2.n3552 3.4105
R11763 GNDA_2.n3552 GNDA_2.n1331 3.4105
R11764 GNDA_2.n3552 GNDA_2.n1332 3.4105
R11765 GNDA_2.n3552 GNDA_2.n1330 3.4105
R11766 GNDA_2.n3552 GNDA_2.n1333 3.4105
R11767 GNDA_2.n3552 GNDA_2.n1329 3.4105
R11768 GNDA_2.n3552 GNDA_2.n1334 3.4105
R11769 GNDA_2.n3552 GNDA_2.n1328 3.4105
R11770 GNDA_2.n3552 GNDA_2.n1335 3.4105
R11771 GNDA_2.n3552 GNDA_2.n1327 3.4105
R11772 GNDA_2.n3552 GNDA_2.n1336 3.4105
R11773 GNDA_2.n3552 GNDA_2.n1326 3.4105
R11774 GNDA_2.n3552 GNDA_2.n1337 3.4105
R11775 GNDA_2.n3552 GNDA_2.n1325 3.4105
R11776 GNDA_2.n3552 GNDA_2.n1338 3.4105
R11777 GNDA_2.n3552 GNDA_2.n1324 3.4105
R11778 GNDA_2.n3552 GNDA_2.n1339 3.4105
R11779 GNDA_2.n3552 GNDA_2.n1323 3.4105
R11780 GNDA_2.n3552 GNDA_2.n1340 3.4105
R11781 GNDA_2.n3552 GNDA_2.n1322 3.4105
R11782 GNDA_2.n3552 GNDA_2.n1341 3.4105
R11783 GNDA_2.n3552 GNDA_2.n1321 3.4105
R11784 GNDA_2.n3552 GNDA_2.n1342 3.4105
R11785 GNDA_2.n3552 GNDA_2.n1320 3.4105
R11786 GNDA_2.n3552 GNDA_2.n1343 3.4105
R11787 GNDA_2.n3552 GNDA_2.n1319 3.4105
R11788 GNDA_2.n3552 GNDA_2.n1344 3.4105
R11789 GNDA_2.n3552 GNDA_2.n1318 3.4105
R11790 GNDA_2.n3552 GNDA_2.n1345 3.4105
R11791 GNDA_2.n3552 GNDA_2.n1317 3.4105
R11792 GNDA_2.n3552 GNDA_2.n1346 3.4105
R11793 GNDA_2.n3552 GNDA_2.n1316 3.4105
R11794 GNDA_2.n3552 GNDA_2.n1347 3.4105
R11795 GNDA_2.n3552 GNDA_2.n3551 3.4105
R11796 GNDA_2.n3954 GNDA_2.n3953 3.4105
R11797 GNDA_2.n3953 GNDA_2.n3952 3.4105
R11798 GNDA_2.n3888 GNDA_2.n3565 3.4105
R11799 GNDA_2.n3888 GNDA_2.n3887 3.4105
R11800 GNDA_2.n3819 GNDA_2.n3577 3.4105
R11801 GNDA_2.n3819 GNDA_2.n3818 3.4105
R11802 GNDA_2.n3750 GNDA_2.n3589 3.4105
R11803 GNDA_2.n3750 GNDA_2.n3749 3.4105
R11804 GNDA_2.n3681 GNDA_2.n3601 3.4105
R11805 GNDA_2.n3681 GNDA_2.n3680 3.4105
R11806 GNDA_2.n1162 GNDA_2.n1122 3.4105
R11807 GNDA_2.n1206 GNDA_2.n1122 3.4105
R11808 GNDA_2.n4074 GNDA_2.n1123 3.4105
R11809 GNDA_2.n4074 GNDA_2.n4073 3.4105
R11810 GNDA_2.n4155 GNDA_2.n4075 3.4105
R11811 GNDA_2.n4155 GNDA_2.n4154 3.4105
R11812 GNDA_2.n4264 GNDA_2.n4172 3.4105
R11813 GNDA_2.n4264 GNDA_2.n4263 3.4105
R11814 GNDA_2.n4265 GNDA_2.n1094 3.4105
R11815 GNDA_2.n4266 GNDA_2.n4265 3.4105
R11816 GNDA_2.n4535 GNDA_2.n188 3.4105
R11817 GNDA_2.n4535 GNDA_2.n4534 3.4105
R11818 GNDA_2.n4702 GNDA_2.n147 3.4105
R11819 GNDA_2.n4668 GNDA_2.n147 3.4105
R11820 GNDA_2.n4772 GNDA_2.n148 3.4105
R11821 GNDA_2.n4772 GNDA_2.n4771 3.4105
R11822 GNDA_2.n5213 GNDA_2.n5212 3.4105
R11823 GNDA_2.n5212 GNDA_2.n5211 3.4105
R11824 GNDA_2.n4612 GNDA_2.n4611 3.4105
R11825 GNDA_2.n4611 GNDA_2.n4610 3.4105
R11826 GNDA_2.n5147 GNDA_2.n4784 3.4105
R11827 GNDA_2.n5147 GNDA_2.n5146 3.4105
R11828 GNDA_2.n4890 GNDA_2.n4796 3.4105
R11829 GNDA_2.n4856 GNDA_2.n4796 3.4105
R11830 GNDA_2.n4987 GNDA_2.n4906 3.4105
R11831 GNDA_2.n4987 GNDA_2.n4986 3.4105
R11832 GNDA_2.n5064 GNDA_2.n5063 3.4105
R11833 GNDA_2.n5063 GNDA_2.n5062 3.4105
R11834 GNDA_2.n261 GNDA_2.n258 3.4105
R11835 GNDA_2.n262 GNDA_2.n257 3.4105
R11836 GNDA_2.n263 GNDA_2.n255 3.4105
R11837 GNDA_2.n254 GNDA_2.n251 3.4105
R11838 GNDA_2.n267 GNDA_2.n250 3.4105
R11839 GNDA_2.n268 GNDA_2.n249 3.4105
R11840 GNDA_2.n269 GNDA_2.n247 3.4105
R11841 GNDA_2.n246 GNDA_2.n243 3.4105
R11842 GNDA_2.n273 GNDA_2.n242 3.4105
R11843 GNDA_2.n274 GNDA_2.n241 3.4105
R11844 GNDA_2.n275 GNDA_2.n239 3.4105
R11845 GNDA_2.n238 GNDA_2.n235 3.4105
R11846 GNDA_2.n279 GNDA_2.n234 3.4105
R11847 GNDA_2.n280 GNDA_2.n233 3.4105
R11848 GNDA_2.n281 GNDA_2.n231 3.4105
R11849 GNDA_2.n230 GNDA_2.n227 3.4105
R11850 GNDA_2.n285 GNDA_2.n226 3.4105
R11851 GNDA_2.n286 GNDA_2.n225 3.4105
R11852 GNDA_2.n287 GNDA_2.n223 3.4105
R11853 GNDA_2.n222 GNDA_2.n219 3.4105
R11854 GNDA_2.n291 GNDA_2.n218 3.4105
R11855 GNDA_2.n292 GNDA_2.n217 3.4105
R11856 GNDA_2.n630 GNDA_2.n629 3.4105
R11857 GNDA_2.n694 GNDA_2.n693 3.4105
R11858 GNDA_2.n692 GNDA_2.n691 3.4105
R11859 GNDA_2.n690 GNDA_2.n634 3.4105
R11860 GNDA_2.n633 GNDA_2.n632 3.4105
R11861 GNDA_2.n686 GNDA_2.n685 3.4105
R11862 GNDA_2.n684 GNDA_2.n683 3.4105
R11863 GNDA_2.n682 GNDA_2.n638 3.4105
R11864 GNDA_2.n637 GNDA_2.n636 3.4105
R11865 GNDA_2.n678 GNDA_2.n677 3.4105
R11866 GNDA_2.n676 GNDA_2.n675 3.4105
R11867 GNDA_2.n674 GNDA_2.n642 3.4105
R11868 GNDA_2.n641 GNDA_2.n640 3.4105
R11869 GNDA_2.n670 GNDA_2.n669 3.4105
R11870 GNDA_2.n668 GNDA_2.n667 3.4105
R11871 GNDA_2.n666 GNDA_2.n646 3.4105
R11872 GNDA_2.n645 GNDA_2.n644 3.4105
R11873 GNDA_2.n662 GNDA_2.n661 3.4105
R11874 GNDA_2.n660 GNDA_2.n659 3.4105
R11875 GNDA_2.n658 GNDA_2.n650 3.4105
R11876 GNDA_2.n649 GNDA_2.n648 3.4105
R11877 GNDA_2.n654 GNDA_2.n653 3.4105
R11878 GNDA_2.n652 GNDA_2.n617 3.4105
R11879 GNDA_2.n444 GNDA_2.n443 3.4105
R11880 GNDA_2.n1010 GNDA_2.n1009 3.4105
R11881 GNDA_2.n1008 GNDA_2.n1007 3.4105
R11882 GNDA_2.n1006 GNDA_2.n448 3.4105
R11883 GNDA_2.n447 GNDA_2.n446 3.4105
R11884 GNDA_2.n1002 GNDA_2.n1001 3.4105
R11885 GNDA_2.n1000 GNDA_2.n999 3.4105
R11886 GNDA_2.n998 GNDA_2.n452 3.4105
R11887 GNDA_2.n451 GNDA_2.n450 3.4105
R11888 GNDA_2.n994 GNDA_2.n993 3.4105
R11889 GNDA_2.n992 GNDA_2.n991 3.4105
R11890 GNDA_2.n990 GNDA_2.n456 3.4105
R11891 GNDA_2.n455 GNDA_2.n454 3.4105
R11892 GNDA_2.n986 GNDA_2.n985 3.4105
R11893 GNDA_2.n984 GNDA_2.n983 3.4105
R11894 GNDA_2.n982 GNDA_2.n460 3.4105
R11895 GNDA_2.n459 GNDA_2.n458 3.4105
R11896 GNDA_2.n978 GNDA_2.n977 3.4105
R11897 GNDA_2.n976 GNDA_2.n975 3.4105
R11898 GNDA_2.n974 GNDA_2.n464 3.4105
R11899 GNDA_2.n463 GNDA_2.n462 3.4105
R11900 GNDA_2.n970 GNDA_2.n969 3.4105
R11901 GNDA_2.n968 GNDA_2.n431 3.4105
R11902 GNDA_2.n516 GNDA_2.n513 3.4105
R11903 GNDA_2.n517 GNDA_2.n511 3.4105
R11904 GNDA_2.n518 GNDA_2.n510 3.4105
R11905 GNDA_2.n508 GNDA_2.n506 3.4105
R11906 GNDA_2.n522 GNDA_2.n505 3.4105
R11907 GNDA_2.n523 GNDA_2.n503 3.4105
R11908 GNDA_2.n524 GNDA_2.n502 3.4105
R11909 GNDA_2.n500 GNDA_2.n498 3.4105
R11910 GNDA_2.n528 GNDA_2.n497 3.4105
R11911 GNDA_2.n529 GNDA_2.n495 3.4105
R11912 GNDA_2.n530 GNDA_2.n494 3.4105
R11913 GNDA_2.n492 GNDA_2.n490 3.4105
R11914 GNDA_2.n534 GNDA_2.n489 3.4105
R11915 GNDA_2.n535 GNDA_2.n487 3.4105
R11916 GNDA_2.n536 GNDA_2.n486 3.4105
R11917 GNDA_2.n484 GNDA_2.n482 3.4105
R11918 GNDA_2.n540 GNDA_2.n481 3.4105
R11919 GNDA_2.n541 GNDA_2.n479 3.4105
R11920 GNDA_2.n542 GNDA_2.n478 3.4105
R11921 GNDA_2.n476 GNDA_2.n474 3.4105
R11922 GNDA_2.n546 GNDA_2.n473 3.4105
R11923 GNDA_2.n547 GNDA_2.n471 3.4105
R11924 GNDA_2.n548 GNDA_2.n470 3.4105
R11925 GNDA_2.n735 GNDA_2.n734 3.4105
R11926 GNDA_2.n798 GNDA_2.n797 3.4105
R11927 GNDA_2.n796 GNDA_2.n795 3.4105
R11928 GNDA_2.n794 GNDA_2.n739 3.4105
R11929 GNDA_2.n738 GNDA_2.n737 3.4105
R11930 GNDA_2.n790 GNDA_2.n789 3.4105
R11931 GNDA_2.n788 GNDA_2.n787 3.4105
R11932 GNDA_2.n786 GNDA_2.n743 3.4105
R11933 GNDA_2.n742 GNDA_2.n741 3.4105
R11934 GNDA_2.n782 GNDA_2.n781 3.4105
R11935 GNDA_2.n780 GNDA_2.n779 3.4105
R11936 GNDA_2.n778 GNDA_2.n747 3.4105
R11937 GNDA_2.n746 GNDA_2.n745 3.4105
R11938 GNDA_2.n774 GNDA_2.n773 3.4105
R11939 GNDA_2.n772 GNDA_2.n771 3.4105
R11940 GNDA_2.n770 GNDA_2.n751 3.4105
R11941 GNDA_2.n750 GNDA_2.n749 3.4105
R11942 GNDA_2.n766 GNDA_2.n765 3.4105
R11943 GNDA_2.n764 GNDA_2.n763 3.4105
R11944 GNDA_2.n762 GNDA_2.n755 3.4105
R11945 GNDA_2.n754 GNDA_2.n753 3.4105
R11946 GNDA_2.n758 GNDA_2.n757 3.4105
R11947 GNDA_2.n756 GNDA_2.n722 3.4105
R11948 GNDA_2.n804 GNDA_2.n803 3.4105
R11949 GNDA_2.n867 GNDA_2.n866 3.4105
R11950 GNDA_2.n865 GNDA_2.n864 3.4105
R11951 GNDA_2.n863 GNDA_2.n808 3.4105
R11952 GNDA_2.n807 GNDA_2.n806 3.4105
R11953 GNDA_2.n859 GNDA_2.n858 3.4105
R11954 GNDA_2.n857 GNDA_2.n856 3.4105
R11955 GNDA_2.n855 GNDA_2.n812 3.4105
R11956 GNDA_2.n811 GNDA_2.n810 3.4105
R11957 GNDA_2.n851 GNDA_2.n850 3.4105
R11958 GNDA_2.n849 GNDA_2.n848 3.4105
R11959 GNDA_2.n847 GNDA_2.n816 3.4105
R11960 GNDA_2.n815 GNDA_2.n814 3.4105
R11961 GNDA_2.n843 GNDA_2.n842 3.4105
R11962 GNDA_2.n841 GNDA_2.n840 3.4105
R11963 GNDA_2.n839 GNDA_2.n820 3.4105
R11964 GNDA_2.n819 GNDA_2.n818 3.4105
R11965 GNDA_2.n835 GNDA_2.n834 3.4105
R11966 GNDA_2.n833 GNDA_2.n832 3.4105
R11967 GNDA_2.n831 GNDA_2.n824 3.4105
R11968 GNDA_2.n823 GNDA_2.n822 3.4105
R11969 GNDA_2.n827 GNDA_2.n826 3.4105
R11970 GNDA_2.n825 GNDA_2.n710 3.4105
R11971 GNDA_2.n873 GNDA_2.n872 3.4105
R11972 GNDA_2.n932 GNDA_2.n931 3.4105
R11973 GNDA_2.n930 GNDA_2.n929 3.4105
R11974 GNDA_2.n928 GNDA_2.n927 3.4105
R11975 GNDA_2.n926 GNDA_2.n875 3.4105
R11976 GNDA_2.n922 GNDA_2.n921 3.4105
R11977 GNDA_2.n920 GNDA_2.n919 3.4105
R11978 GNDA_2.n918 GNDA_2.n917 3.4105
R11979 GNDA_2.n916 GNDA_2.n877 3.4105
R11980 GNDA_2.n912 GNDA_2.n911 3.4105
R11981 GNDA_2.n910 GNDA_2.n909 3.4105
R11982 GNDA_2.n908 GNDA_2.n907 3.4105
R11983 GNDA_2.n906 GNDA_2.n879 3.4105
R11984 GNDA_2.n902 GNDA_2.n901 3.4105
R11985 GNDA_2.n900 GNDA_2.n899 3.4105
R11986 GNDA_2.n898 GNDA_2.n897 3.4105
R11987 GNDA_2.n896 GNDA_2.n881 3.4105
R11988 GNDA_2.n892 GNDA_2.n891 3.4105
R11989 GNDA_2.n890 GNDA_2.n889 3.4105
R11990 GNDA_2.n888 GNDA_2.n887 3.4105
R11991 GNDA_2.n886 GNDA_2.n883 3.4105
R11992 GNDA_2.n616 GNDA_2.n615 3.4105
R11993 GNDA_2.n938 GNDA_2.n937 3.4105
R11994 GNDA_2.n937 GNDA_2.n936 3.4105
R11995 GNDA_2.n936 GNDA_2.n935 3.4105
R11996 GNDA_2.n871 GNDA_2.n710 3.4105
R11997 GNDA_2.n871 GNDA_2.n870 3.4105
R11998 GNDA_2.n802 GNDA_2.n722 3.4105
R11999 GNDA_2.n802 GNDA_2.n801 3.4105
R12000 GNDA_2.n470 GNDA_2.n430 3.4105
R12001 GNDA_2.n514 GNDA_2.n430 3.4105
R12002 GNDA_2.n1014 GNDA_2.n431 3.4105
R12003 GNDA_2.n1014 GNDA_2.n1013 3.4105
R12004 GNDA_2.n698 GNDA_2.n617 3.4105
R12005 GNDA_2.n698 GNDA_2.n697 3.4105
R12006 GNDA_2.n1031 GNDA_2.n402 3.4105
R12007 GNDA_2.n1032 GNDA_2.n1031 3.4105
R12008 GNDA_2.n4351 GNDA_2.n4350 3.08383
R12009 GNDA_2.n378 GNDA_2.n377 3.08383
R12010 GNDA_2.n3388 GNDA_2.n1679 3.04346
R12011 GNDA_2.n2653 GNDA_2.n2617 3.00528
R12012 GNDA_2.n2702 GNDA_2.n2701 3.00528
R12013 GNDA_2.n3357 GNDA_2.t48 3.00528
R12014 GNDA_2.n1703 GNDA_2.t165 3.00528
R12015 GNDA_2.n3375 GNDA_2.n1684 2.86505
R12016 GNDA_2.n3376 GNDA_2.n3375 2.86505
R12017 GNDA_2.n3374 GNDA_2.n3370 2.86505
R12018 GNDA_2.n3371 GNDA_2.n3370 2.86505
R12019 GNDA_2.n3377 GNDA_2.n3376 2.86505
R12020 GNDA_2.n3372 GNDA_2.n3371 2.86505
R12021 GNDA_2.n3381 GNDA_2.n1684 2.86505
R12022 GNDA_2.n3377 GNDA_2.n3374 2.86505
R12023 GNDA_2.n2835 GNDA_2.n2834 2.86505
R12024 GNDA_2.n2834 GNDA_2.n2832 2.86505
R12025 GNDA_2.n2832 GNDA_2.n2831 2.86505
R12026 GNDA_2.n2836 GNDA_2.n2835 2.86505
R12027 GNDA_2.n3428 GNDA_2.n3426 2.69842
R12028 GNDA_2.n5548 GNDA_2.n5547 2.6629
R12029 GNDA_2.n5461 GNDA_2.n82 2.6629
R12030 GNDA_2.n2603 GNDA_2.n2602 2.6629
R12031 GNDA_2.n2536 GNDA_2.n1913 2.6629
R12032 GNDA_2.n2928 GNDA_2.n2614 2.6629
R12033 GNDA_2.n2641 GNDA_2.n1806 2.6629
R12034 GNDA_2.n2769 GNDA_2.n2767 2.6629
R12035 GNDA_2.n2808 GNDA_2.n1782 2.6629
R12036 GNDA_2.n2106 GNDA_2.n2105 2.6629
R12037 GNDA_2.n2460 GNDA_2.n2143 2.6629
R12038 GNDA_2.n5453 GNDA_2.n5452 2.6629
R12039 GNDA_2.n5361 GNDA_2.n110 2.6629
R12040 GNDA_2.n2326 GNDA_2.n2325 2.6629
R12041 GNDA_2.n1781 GNDA_2.n1780 2.6629
R12042 GNDA_2.n5353 GNDA_2.n5352 2.6629
R12043 GNDA_2.t130 GNDA_2.t73 2.59854
R12044 GNDA_2.n1068 GNDA_2.n1067 2.57978
R12045 GNDA_2.n651 GNDA_2.n613 2.57937
R12046 GNDA_2.n967 GNDA_2.n966 2.54738
R12047 GNDA_2.n959 GNDA_2.n549 2.54738
R12048 GNDA_2.n954 GNDA_2.n553 2.54738
R12049 GNDA_2.n949 GNDA_2.n557 2.54738
R12050 GNDA_2.n940 GNDA_2.n939 2.54738
R12051 GNDA_2.n563 GNDA_2.n562 2.46404
R12052 GNDA_2.n1075 GNDA_2.n1074 2.46404
R12053 GNDA_2.n5462 GNDA_2.n5461 2.4581
R12054 GNDA_2.n2537 GNDA_2.n2536 2.4581
R12055 GNDA_2.n2642 GNDA_2.n2641 2.4581
R12056 GNDA_2.n2767 GNDA_2.n1806 2.4581
R12057 GNDA_2.n2809 GNDA_2.n2808 2.4581
R12058 GNDA_2.n2105 GNDA_2.n1913 2.4581
R12059 GNDA_2.n2143 GNDA_2.n2142 2.4581
R12060 GNDA_2.n5453 GNDA_2.n82 2.4581
R12061 GNDA_2.n5362 GNDA_2.n5361 2.4581
R12062 GNDA_2.n2460 GNDA_2.n2326 2.4581
R12063 GNDA_2.n2235 GNDA_2.n2234 2.4581
R12064 GNDA_2.n1782 GNDA_2.n1781 2.4581
R12065 GNDA_2.n3399 GNDA_2.n3398 2.4581
R12066 GNDA_2.n5353 GNDA_2.n110 2.4581
R12067 GNDA_2.n5286 GNDA_2.n5285 2.4581
R12068 GNDA_2.n3391 GNDA_2.n3390 2.44675
R12069 GNDA_2.n3390 GNDA_2.n3389 2.44675
R12070 GNDA_2.n1590 GNDA_2.n1589 2.39683
R12071 GNDA_2.n1033 GNDA_2.n426 2.30736
R12072 GNDA_2.n5061 GNDA_2.n5060 2.30736
R12073 GNDA_2.n4985 GNDA_2.n4984 2.30736
R12074 GNDA_2.n4855 GNDA_2.n4854 2.30736
R12075 GNDA_2.n5145 GNDA_2.n5144 2.30736
R12076 GNDA_2.n4609 GNDA_2.n4608 2.30736
R12077 GNDA_2.n5210 GNDA_2.n5209 2.30736
R12078 GNDA_2.n4770 GNDA_2.n4769 2.30736
R12079 GNDA_2.n4667 GNDA_2.n4666 2.30736
R12080 GNDA_2.n4533 GNDA_2.n4532 2.30736
R12081 GNDA_2.n4267 GNDA_2.n1118 2.30736
R12082 GNDA_2.n4262 GNDA_2.n4261 2.30736
R12083 GNDA_2.n4153 GNDA_2.n4152 2.30736
R12084 GNDA_2.n4072 GNDA_2.n4071 2.30736
R12085 GNDA_2.n1207 GNDA_2.n1199 2.30736
R12086 GNDA_2.n3679 GNDA_2.n3678 2.30736
R12087 GNDA_2.n3748 GNDA_2.n3747 2.30736
R12088 GNDA_2.n3817 GNDA_2.n3816 2.30736
R12089 GNDA_2.n3886 GNDA_2.n3885 2.30736
R12090 GNDA_2.n3951 GNDA_2.n3950 2.30736
R12091 GNDA_2.n3000 GNDA_2.n2997 2.30736
R12092 GNDA_2.n260 GNDA_2.n252 2.30736
R12093 GNDA_2.n696 GNDA_2.n695 2.30736
R12094 GNDA_2.n1012 GNDA_2.n1011 2.30736
R12095 GNDA_2.n515 GNDA_2.n507 2.30736
R12096 GNDA_2.n800 GNDA_2.n799 2.30736
R12097 GNDA_2.n869 GNDA_2.n868 2.30736
R12098 GNDA_2.n934 GNDA_2.n933 2.30736
R12099 GNDA_2.n5253 GNDA_2.n5252 2.29914
R12100 GNDA_2.n4467 GNDA_2.n133 2.29914
R12101 GNDA_2.n4410 GNDA_2.n4409 2.29914
R12102 GNDA_2.n4315 GNDA_2.n331 2.29914
R12103 GNDA_2.n3434 GNDA_2.n3433 2.29738
R12104 GNDA_2.n357 GNDA_2.n354 2.26187
R12105 GNDA_2.n358 GNDA_2.n357 2.26187
R12106 GNDA_2.n4390 GNDA_2.n342 2.26187
R12107 GNDA_2.n3997 GNDA_2.n3981 2.26187
R12108 GNDA_2.n4004 GNDA_2.n3979 2.26187
R12109 GNDA_2.n3959 GNDA_2.n3958 2.26187
R12110 GNDA_2.n2691 GNDA_2.n2668 2.26187
R12111 GNDA_2.n3385 GNDA_2.n3384 2.26187
R12112 GNDA_2.n3427 GNDA_2.n1641 2.26187
R12113 GNDA_2.n1647 GNDA_2.n1644 2.26187
R12114 GNDA_2.n1648 GNDA_2.n1647 2.26187
R12115 GNDA_2.n5224 GNDA_2.n5222 2.26187
R12116 GNDA_2.n606 GNDA_2.n567 2.26187
R12117 GNDA_2.n5241 GNDA_2.n5228 2.26187
R12118 GNDA_2.n5242 GNDA_2.n5241 2.26187
R12119 GNDA_2.n364 GNDA_2.n363 2.26187
R12120 GNDA_2.n4434 GNDA_2.n4433 2.26187
R12121 GNDA_2.n4448 GNDA_2.n4447 2.26187
R12122 GNDA_2.n4452 GNDA_2.n4451 2.26187
R12123 GNDA_2.n4380 GNDA_2.n4379 2.26187
R12124 GNDA_2.n4387 GNDA_2.n342 2.26187
R12125 GNDA_2.n3994 GNDA_2.n3981 2.26187
R12126 GNDA_2.n3963 GNDA_2.n1258 2.26187
R12127 GNDA_2.n3968 GNDA_2.n1254 2.26187
R12128 GNDA_2.n3973 GNDA_2.n1250 2.26187
R12129 GNDA_2.n4012 GNDA_2.n1243 2.26187
R12130 GNDA_2.n4017 GNDA_2.n1159 2.26187
R12131 GNDA_2.n4024 GNDA_2.n4023 2.26187
R12132 GNDA_2.n4214 GNDA_2.n4213 2.26187
R12133 GNDA_2.n3960 GNDA_2.n3959 2.26187
R12134 GNDA_2.n3386 GNDA_2.n3385 2.26187
R12135 GNDA_2.n2662 GNDA_2.n2661 2.26187
R12136 GNDA_2.n3060 GNDA_2.n3059 2.26187
R12137 GNDA_2.n296 GNDA_2.n213 2.26187
R12138 GNDA_2.n1071 GNDA_2.n1070 2.26187
R12139 GNDA_2.n396 GNDA_2.n395 2.26187
R12140 GNDA_2.n603 GNDA_2.n567 2.26187
R12141 GNDA_2.n947 GNDA_2.n555 2.26187
R12142 GNDA_2.n952 GNDA_2.n551 2.26187
R12143 GNDA_2.n957 GNDA_2.n467 2.26187
R12144 GNDA_2.n964 GNDA_2.n963 2.26187
R12145 GNDA_2.n944 GNDA_2.n943 2.26187
R12146 GNDA_2.n4308 GNDA_2.n4307 2.24241
R12147 GNDA_2.n1090 GNDA_2.n1088 2.24241
R12148 GNDA_2.n4619 GNDA_2.n179 2.24241
R12149 GNDA_2.n181 GNDA_2.n178 2.24241
R12150 GNDA_2.n5245 GNDA_2.n5240 2.24063
R12151 GNDA_2.n5246 GNDA_2.n5228 2.24063
R12152 GNDA_2.n5249 GNDA_2.n5248 2.24063
R12153 GNDA_2.n5227 GNDA_2.n136 2.24063
R12154 GNDA_2.n4437 GNDA_2.n4430 2.24063
R12155 GNDA_2.n4438 GNDA_2.n4428 2.24063
R12156 GNDA_2.n4443 GNDA_2.n317 2.24063
R12157 GNDA_2.n318 GNDA_2.n316 2.24063
R12158 GNDA_2.n4455 GNDA_2.n308 2.24063
R12159 GNDA_2.n4451 GNDA_2.n4450 2.24063
R12160 GNDA_2.n4445 GNDA_2.n4444 2.24063
R12161 GNDA_2.n4447 GNDA_2.n4446 2.24063
R12162 GNDA_2.n367 GNDA_2.n352 2.24063
R12163 GNDA_2.n364 GNDA_2.n362 2.24063
R12164 GNDA_2.n4379 GNDA_2.n4378 2.24063
R12165 GNDA_2.n4377 GNDA_2.n4376 2.24063
R12166 GNDA_2.n4391 GNDA_2.n341 2.24063
R12167 GNDA_2.n4397 GNDA_2.n340 2.24063
R12168 GNDA_2.n4392 GNDA_2.n339 2.24063
R12169 GNDA_2.n4394 GNDA_2.n321 2.24063
R12170 GNDA_2.n4426 GNDA_2.n320 2.24063
R12171 GNDA_2.n322 GNDA_2.n319 2.24063
R12172 GNDA_2.n4423 GNDA_2.n4422 2.24063
R12173 GNDA_2.n4416 GNDA_2.n325 2.24063
R12174 GNDA_2.n4418 GNDA_2.n324 2.24063
R12175 GNDA_2.n4419 GNDA_2.n4417 2.24063
R12176 GNDA_2.n4414 GNDA_2.n4413 2.24063
R12177 GNDA_2.n330 GNDA_2.n329 2.24063
R12178 GNDA_2.n3998 GNDA_2.n3980 2.24063
R12179 GNDA_2.n4005 GNDA_2.n3978 2.24063
R12180 GNDA_2.n3966 GNDA_2.n1258 2.24063
R12181 GNDA_2.n1259 GNDA_2.n1257 2.24063
R12182 GNDA_2.n3971 GNDA_2.n1254 2.24063
R12183 GNDA_2.n1255 GNDA_2.n1253 2.24063
R12184 GNDA_2.n3976 GNDA_2.n1250 2.24063
R12185 GNDA_2.n1251 GNDA_2.n1249 2.24063
R12186 GNDA_2.n4015 GNDA_2.n1243 2.24063
R12187 GNDA_2.n1244 GNDA_2.n1242 2.24063
R12188 GNDA_2.n4020 GNDA_2.n1159 2.24063
R12189 GNDA_2.n1160 GNDA_2.n1158 2.24063
R12190 GNDA_2.n4023 GNDA_2.n1085 2.24063
R12191 GNDA_2.n4022 GNDA_2.n1157 2.24063
R12192 GNDA_2.n4213 GNDA_2.n4207 2.24063
R12193 GNDA_2.n4212 GNDA_2.n4206 2.24063
R12194 GNDA_2.n4010 GNDA_2.n1247 2.24063
R12195 GNDA_2.n1248 GNDA_2.n1246 2.24063
R12196 GNDA_2.n3957 GNDA_2.n1261 2.24063
R12197 GNDA_2.n2692 GNDA_2.n2691 2.24063
R12198 GNDA_2.n2661 GNDA_2.n1683 2.24063
R12199 GNDA_2.n2664 GNDA_2.n2663 2.24063
R12200 GNDA_2.n3063 GNDA_2.n2975 2.24063
R12201 GNDA_2.n3059 GNDA_2.n1679 2.24063
R12202 GNDA_2.n3384 GNDA_2.n3383 2.24063
R12203 GNDA_2.n3429 GNDA_2.n3428 2.24063
R12204 GNDA_2.n299 GNDA_2.n213 2.24063
R12205 GNDA_2.n214 GNDA_2.n212 2.24063
R12206 GNDA_2.n4709 GNDA_2.n176 2.24063
R12207 GNDA_2.n177 GNDA_2.n175 2.24063
R12208 GNDA_2.n4706 GNDA_2.n4705 2.24063
R12209 GNDA_2.n4713 GNDA_2.n142 2.24063
R12210 GNDA_2.n174 GNDA_2.n173 2.24063
R12211 GNDA_2.n4714 GNDA_2.n172 2.24063
R12212 GNDA_2.n5220 GNDA_2.n140 2.24063
R12213 GNDA_2.n141 GNDA_2.n139 2.24063
R12214 GNDA_2.n5217 GNDA_2.n5216 2.24063
R12215 GNDA_2.n4616 GNDA_2.n4615 2.24063
R12216 GNDA_2.n5088 GNDA_2.n5082 2.24063
R12217 GNDA_2.n5084 GNDA_2.n5083 2.24063
R12218 GNDA_2.n5089 GNDA_2.n4809 2.24063
R12219 GNDA_2.n5078 GNDA_2.n4895 2.24063
R12220 GNDA_2.n5079 GNDA_2.n4894 2.24063
R12221 GNDA_2.n5080 GNDA_2.n4893 2.24063
R12222 GNDA_2.n5074 GNDA_2.n4900 2.24063
R12223 GNDA_2.n5075 GNDA_2.n4899 2.24063
R12224 GNDA_2.n5076 GNDA_2.n4898 2.24063
R12225 GNDA_2.n5070 GNDA_2.n5069 2.24063
R12226 GNDA_2.n5071 GNDA_2.n5068 2.24063
R12227 GNDA_2.n5072 GNDA_2.n5067 2.24063
R12228 GNDA_2.n5222 GNDA_2.n138 2.24063
R12229 GNDA_2.n5223 GNDA_2.n137 2.24063
R12230 GNDA_2.n1074 GNDA_2.n389 2.24063
R12231 GNDA_2.n1070 GNDA_2.n1069 2.24063
R12232 GNDA_2.n395 GNDA_2.n392 2.24063
R12233 GNDA_2.n394 GNDA_2.n391 2.24063
R12234 GNDA_2.n607 GNDA_2.n566 2.24063
R12235 GNDA_2.n611 GNDA_2.n563 2.24063
R12236 GNDA_2.n565 GNDA_2.n564 2.24063
R12237 GNDA_2.n612 GNDA_2.n561 2.24063
R12238 GNDA_2.n950 GNDA_2.n555 2.24063
R12239 GNDA_2.n556 GNDA_2.n554 2.24063
R12240 GNDA_2.n955 GNDA_2.n551 2.24063
R12241 GNDA_2.n552 GNDA_2.n550 2.24063
R12242 GNDA_2.n960 GNDA_2.n467 2.24063
R12243 GNDA_2.n468 GNDA_2.n466 2.24063
R12244 GNDA_2.n963 GNDA_2.n400 2.24063
R12245 GNDA_2.n962 GNDA_2.n465 2.24063
R12246 GNDA_2.n942 GNDA_2.n941 2.24063
R12247 GNDA_2.n940 GNDA_2.n558 2.24063
R12248 GNDA_2.n5247 GNDA_2.n135 2.24063
R12249 GNDA_2.n4433 GNDA_2.n4432 2.24063
R12250 GNDA_2.n4440 GNDA_2.n4439 2.24063
R12251 GNDA_2.n4454 GNDA_2.n4453 2.24063
R12252 GNDA_2.n4449 GNDA_2.n312 2.24063
R12253 GNDA_2.n366 GNDA_2.n315 2.24063
R12254 GNDA_2.n361 GNDA_2.n354 2.24063
R12255 GNDA_2.n360 GNDA_2.n359 2.24063
R12256 GNDA_2.n4387 GNDA_2.n4386 2.24063
R12257 GNDA_2.n4415 GNDA_2.n327 2.24063
R12258 GNDA_2.n3994 GNDA_2.n3993 2.24063
R12259 GNDA_2.n3999 GNDA_2.n3979 2.24063
R12260 GNDA_2.n4001 GNDA_2.n4000 2.24063
R12261 GNDA_2.n4306 GNDA_2.n1087 2.24063
R12262 GNDA_2.n4007 GNDA_2.n4006 2.24063
R12263 GNDA_2.n3961 GNDA_2.n3960 2.24063
R12264 GNDA_2.n2825 GNDA_2.n2665 2.24063
R12265 GNDA_2.n2824 GNDA_2.n2823 2.24063
R12266 GNDA_2.n3062 GNDA_2.n3061 2.24063
R12267 GNDA_2.n3387 GNDA_2.n1680 2.24063
R12268 GNDA_2.n3433 GNDA_2.n1641 2.24063
R12269 GNDA_2.n3432 GNDA_2.n3431 2.24063
R12270 GNDA_2.n3426 GNDA_2.n1644 2.24063
R12271 GNDA_2.n3425 GNDA_2.n3424 2.24063
R12272 GNDA_2.n1073 GNDA_2.n1072 2.24063
R12273 GNDA_2.n603 GNDA_2.n602 2.24063
R12274 GNDA_2.n945 GNDA_2.n944 2.24063
R12275 GNDA_2.n374 GNDA_2.n373 2.22018
R12276 GNDA_2.n4358 GNDA_2.n368 2.22018
R12277 GNDA_2.n4401 GNDA_2.n4400 2.22018
R12278 GNDA_2.n4456 GNDA_2.n306 2.22018
R12279 GNDA_2.n2693 GNDA_2.n2689 2.22018
R12280 GNDA_2.n2822 GNDA_2.n2669 2.22018
R12281 GNDA_2.n3068 GNDA_2.n3067 2.22018
R12282 GNDA_2.n601 GNDA_2.n596 2.22018
R12283 GNDA_2.n4340 GNDA_2.n386 2.22018
R12284 GNDA_2.n113 GNDA_2.n110 2.18124
R12285 GNDA_2.n2461 GNDA_2.n2460 2.18124
R12286 GNDA_2.n1785 GNDA_2.n1782 2.18124
R12287 GNDA_2.n1809 GNDA_2.n1806 2.18124
R12288 GNDA_2.n1916 GNDA_2.n1913 2.18124
R12289 GNDA_2.n86 GNDA_2.n82 2.18124
R12290 GNDA_2.n3061 GNDA_2.n3057 2.16717
R12291 GNDA_2.n5480 GNDA_2.n5462 2.1509
R12292 GNDA_2.n2537 GNDA_2.n1912 2.1509
R12293 GNDA_2.n2860 GNDA_2.n2642 2.1509
R12294 GNDA_2.n2810 GNDA_2.n2809 2.1509
R12295 GNDA_2.n2142 GNDA_2.n2141 2.1509
R12296 GNDA_2.n5388 GNDA_2.n5362 2.1509
R12297 GNDA_2.n2261 GNDA_2.n2235 2.1509
R12298 GNDA_2.n3400 GNDA_2.n3399 2.1509
R12299 GNDA_2.n5296 GNDA_2.n5286 2.1509
R12300 GNDA_2.n5547 GNDA_2.n57 2.13383
R12301 GNDA_2.n2602 GNDA_2.n1847 2.13383
R12302 GNDA_2.n2914 GNDA_2.n2614 2.13383
R12303 GNDA_2.n2770 GNDA_2.n2769 2.13383
R12304 GNDA_2.n2106 GNDA_2.n2100 2.13383
R12305 GNDA_2.n5452 GNDA_2.n89 2.13383
R12306 GNDA_2.n2325 GNDA_2.n2144 2.13383
R12307 GNDA_2.n1780 GNDA_2.n1779 2.13383
R12308 GNDA_2.n5352 GNDA_2.n5351 2.13383
R12309 GNDA_2.n4621 GNDA_2.n4620 2.09414
R12310 GNDA_2.n4209 GNDA_2.n4208 2.09414
R12311 GNDA_2.n4313 GNDA_2.n4312 2.09414
R12312 GNDA_2.n4472 GNDA_2.n4471 2.09414
R12313 GNDA_2.n111 GNDA_2.n110 2.08643
R12314 GNDA_2.n2460 GNDA_2.n2459 2.08643
R12315 GNDA_2.n3339 GNDA_2.n1782 2.08643
R12316 GNDA_2.n3332 GNDA_2.n1806 2.08643
R12317 GNDA_2.n1915 GNDA_2.n1913 2.08643
R12318 GNDA_2.n84 GNDA_2.n82 2.08643
R12319 GNDA_2.n5547 GNDA_2.n5546 1.9461
R12320 GNDA_2.n2602 GNDA_2.n2601 1.9461
R12321 GNDA_2.n2619 GNDA_2.n2614 1.9461
R12322 GNDA_2.n2769 GNDA_2.n2768 1.9461
R12323 GNDA_2.n2107 GNDA_2.n2106 1.9461
R12324 GNDA_2.n5452 GNDA_2.n5451 1.9461
R12325 GNDA_2.n2325 GNDA_2.n2324 1.9461
R12326 GNDA_2.n1780 GNDA_2.n1725 1.9461
R12327 GNDA_2.n5352 GNDA_2.n22 1.9461
R12328 GNDA_2.n5254 GNDA_2.n5253 1.93383
R12329 GNDA_2.n4468 GNDA_2.n4467 1.93383
R12330 GNDA_2.n4409 GNDA_2.n4408 1.93383
R12331 GNDA_2.n4316 GNDA_2.n4315 1.93383
R12332 GNDA_2.n5250 GNDA_2.n5226 1.82342
R12333 GNDA_2.n4006 GNDA_2.n4005 1.82342
R12334 GNDA_2.n3383 GNDA_2.n3382 1.71925
R12335 GNDA_2.n1512 GNDA_2.n1511 1.70567
R12336 GNDA_2.n1512 GNDA_2.n1510 1.70567
R12337 GNDA_2.n1512 GNDA_2.n1509 1.70567
R12338 GNDA_2.n1512 GNDA_2.n1508 1.70567
R12339 GNDA_2.n1512 GNDA_2.n1507 1.70567
R12340 GNDA_2.n1512 GNDA_2.n1506 1.70567
R12341 GNDA_2.n1512 GNDA_2.n1505 1.70567
R12342 GNDA_2.n1512 GNDA_2.n1504 1.70567
R12343 GNDA_2.n1512 GNDA_2.n1503 1.70567
R12344 GNDA_2.n1512 GNDA_2.n1502 1.70567
R12345 GNDA_2.n1512 GNDA_2.n1501 1.70567
R12346 GNDA_2.n1512 GNDA_2.n1500 1.70567
R12347 GNDA_2.n1512 GNDA_2.n1499 1.70567
R12348 GNDA_2.n1512 GNDA_2.n1498 1.70567
R12349 GNDA_2.n1512 GNDA_2.n1497 1.70567
R12350 GNDA_2.n1512 GNDA_2.n1496 1.70567
R12351 GNDA_2.n3438 GNDA_2.n1561 1.70567
R12352 GNDA_2.n1544 GNDA_2.n1494 1.70567
R12353 GNDA_2.n1494 GNDA_2.n1493 1.70567
R12354 GNDA_2.n1494 GNDA_2.n1492 1.70567
R12355 GNDA_2.n1494 GNDA_2.n1491 1.70567
R12356 GNDA_2.n1494 GNDA_2.n1490 1.70567
R12357 GNDA_2.n1494 GNDA_2.n1489 1.70567
R12358 GNDA_2.n1494 GNDA_2.n1488 1.70567
R12359 GNDA_2.n1494 GNDA_2.n1487 1.70567
R12360 GNDA_2.n1494 GNDA_2.n1486 1.70567
R12361 GNDA_2.n1494 GNDA_2.n1485 1.70567
R12362 GNDA_2.n1494 GNDA_2.n1484 1.70567
R12363 GNDA_2.n1494 GNDA_2.n1483 1.70567
R12364 GNDA_2.n1494 GNDA_2.n1482 1.70567
R12365 GNDA_2.n1494 GNDA_2.n1481 1.70567
R12366 GNDA_2.n1494 GNDA_2.n1480 1.70567
R12367 GNDA_2.n1494 GNDA_2.n1479 1.70567
R12368 GNDA_2.n1513 GNDA_2.n1495 1.70567
R12369 GNDA_2.n3438 GNDA_2.n1560 1.70567
R12370 GNDA_2.n1515 GNDA_2.n1495 1.70567
R12371 GNDA_2.n3438 GNDA_2.n1559 1.70567
R12372 GNDA_2.n1517 GNDA_2.n1495 1.70567
R12373 GNDA_2.n3438 GNDA_2.n1558 1.70567
R12374 GNDA_2.n1519 GNDA_2.n1495 1.70567
R12375 GNDA_2.n3438 GNDA_2.n1557 1.70567
R12376 GNDA_2.n1521 GNDA_2.n1495 1.70567
R12377 GNDA_2.n3438 GNDA_2.n1556 1.70567
R12378 GNDA_2.n1523 GNDA_2.n1495 1.70567
R12379 GNDA_2.n3438 GNDA_2.n1555 1.70567
R12380 GNDA_2.n1525 GNDA_2.n1495 1.70567
R12381 GNDA_2.n3438 GNDA_2.n1554 1.70567
R12382 GNDA_2.n1527 GNDA_2.n1495 1.70567
R12383 GNDA_2.n3438 GNDA_2.n1553 1.70567
R12384 GNDA_2.n1529 GNDA_2.n1495 1.70567
R12385 GNDA_2.n3438 GNDA_2.n1552 1.70567
R12386 GNDA_2.n1531 GNDA_2.n1495 1.70567
R12387 GNDA_2.n3438 GNDA_2.n1551 1.70567
R12388 GNDA_2.n1533 GNDA_2.n1495 1.70567
R12389 GNDA_2.n3438 GNDA_2.n1550 1.70567
R12390 GNDA_2.n1535 GNDA_2.n1495 1.70567
R12391 GNDA_2.n3438 GNDA_2.n1549 1.70567
R12392 GNDA_2.n1537 GNDA_2.n1495 1.70567
R12393 GNDA_2.n3438 GNDA_2.n1548 1.70567
R12394 GNDA_2.n1539 GNDA_2.n1495 1.70567
R12395 GNDA_2.n3438 GNDA_2.n1547 1.70567
R12396 GNDA_2.n1541 GNDA_2.n1495 1.70567
R12397 GNDA_2.n3438 GNDA_2.n1546 1.70567
R12398 GNDA_2.n1543 GNDA_2.n1495 1.70567
R12399 GNDA_2.n3439 GNDA_2.n3438 1.70567
R12400 GNDA_2.n3442 GNDA_2.n1446 1.70567
R12401 GNDA_2.n1495 GNDA_2.n1430 1.70567
R12402 GNDA_2.n3459 GNDA_2.n3458 1.70567
R12403 GNDA_2.n3459 GNDA_2.n3457 1.70567
R12404 GNDA_2.n3459 GNDA_2.n3456 1.70567
R12405 GNDA_2.n3459 GNDA_2.n3455 1.70567
R12406 GNDA_2.n3459 GNDA_2.n3454 1.70567
R12407 GNDA_2.n3459 GNDA_2.n3453 1.70567
R12408 GNDA_2.n3459 GNDA_2.n3452 1.70567
R12409 GNDA_2.n3459 GNDA_2.n3451 1.70567
R12410 GNDA_2.n3459 GNDA_2.n3450 1.70567
R12411 GNDA_2.n3459 GNDA_2.n3449 1.70567
R12412 GNDA_2.n3459 GNDA_2.n3448 1.70567
R12413 GNDA_2.n3459 GNDA_2.n3447 1.70567
R12414 GNDA_2.n3459 GNDA_2.n3446 1.70567
R12415 GNDA_2.n3459 GNDA_2.n3445 1.70567
R12416 GNDA_2.n3459 GNDA_2.n3444 1.70567
R12417 GNDA_2.n3459 GNDA_2.n3443 1.70567
R12418 GNDA_2.n3509 GNDA_2.n3508 1.70567
R12419 GNDA_2.n3491 GNDA_2.n1428 1.70567
R12420 GNDA_2.n1428 GNDA_2.n1427 1.70567
R12421 GNDA_2.n1428 GNDA_2.n1426 1.70567
R12422 GNDA_2.n1428 GNDA_2.n1425 1.70567
R12423 GNDA_2.n1428 GNDA_2.n1424 1.70567
R12424 GNDA_2.n1428 GNDA_2.n1423 1.70567
R12425 GNDA_2.n1428 GNDA_2.n1422 1.70567
R12426 GNDA_2.n1428 GNDA_2.n1421 1.70567
R12427 GNDA_2.n1428 GNDA_2.n1420 1.70567
R12428 GNDA_2.n1428 GNDA_2.n1419 1.70567
R12429 GNDA_2.n1428 GNDA_2.n1418 1.70567
R12430 GNDA_2.n1428 GNDA_2.n1417 1.70567
R12431 GNDA_2.n1428 GNDA_2.n1416 1.70567
R12432 GNDA_2.n1428 GNDA_2.n1415 1.70567
R12433 GNDA_2.n1428 GNDA_2.n1414 1.70567
R12434 GNDA_2.n1428 GNDA_2.n1413 1.70567
R12435 GNDA_2.n3460 GNDA_2.n1429 1.70567
R12436 GNDA_2.n3509 GNDA_2.n3507 1.70567
R12437 GNDA_2.n3462 GNDA_2.n1429 1.70567
R12438 GNDA_2.n3509 GNDA_2.n3506 1.70567
R12439 GNDA_2.n3464 GNDA_2.n1429 1.70567
R12440 GNDA_2.n3509 GNDA_2.n3505 1.70567
R12441 GNDA_2.n3466 GNDA_2.n1429 1.70567
R12442 GNDA_2.n3509 GNDA_2.n3504 1.70567
R12443 GNDA_2.n3468 GNDA_2.n1429 1.70567
R12444 GNDA_2.n3509 GNDA_2.n3503 1.70567
R12445 GNDA_2.n3470 GNDA_2.n1429 1.70567
R12446 GNDA_2.n3509 GNDA_2.n3502 1.70567
R12447 GNDA_2.n3472 GNDA_2.n1429 1.70567
R12448 GNDA_2.n3509 GNDA_2.n3501 1.70567
R12449 GNDA_2.n3474 GNDA_2.n1429 1.70567
R12450 GNDA_2.n3509 GNDA_2.n3500 1.70567
R12451 GNDA_2.n3476 GNDA_2.n1429 1.70567
R12452 GNDA_2.n3509 GNDA_2.n3499 1.70567
R12453 GNDA_2.n3478 GNDA_2.n1429 1.70567
R12454 GNDA_2.n3509 GNDA_2.n3498 1.70567
R12455 GNDA_2.n3480 GNDA_2.n1429 1.70567
R12456 GNDA_2.n3509 GNDA_2.n3497 1.70567
R12457 GNDA_2.n3482 GNDA_2.n1429 1.70567
R12458 GNDA_2.n3509 GNDA_2.n3496 1.70567
R12459 GNDA_2.n3484 GNDA_2.n1429 1.70567
R12460 GNDA_2.n3509 GNDA_2.n3495 1.70567
R12461 GNDA_2.n3486 GNDA_2.n1429 1.70567
R12462 GNDA_2.n3509 GNDA_2.n3494 1.70567
R12463 GNDA_2.n3488 GNDA_2.n1429 1.70567
R12464 GNDA_2.n3509 GNDA_2.n3493 1.70567
R12465 GNDA_2.n3490 GNDA_2.n1429 1.70567
R12466 GNDA_2.n3510 GNDA_2.n3509 1.70567
R12467 GNDA_2.n3513 GNDA_2.n1380 1.70567
R12468 GNDA_2.n1429 GNDA_2.n1364 1.70567
R12469 GNDA_2.n3553 GNDA_2.n1283 1.70567
R12470 GNDA_2.n3530 GNDA_2.n3529 1.70567
R12471 GNDA_2.n3530 GNDA_2.n3528 1.70567
R12472 GNDA_2.n3530 GNDA_2.n3527 1.70567
R12473 GNDA_2.n3530 GNDA_2.n3526 1.70567
R12474 GNDA_2.n3530 GNDA_2.n3525 1.70567
R12475 GNDA_2.n3530 GNDA_2.n3524 1.70567
R12476 GNDA_2.n3530 GNDA_2.n3523 1.70567
R12477 GNDA_2.n3530 GNDA_2.n3522 1.70567
R12478 GNDA_2.n3530 GNDA_2.n3521 1.70567
R12479 GNDA_2.n3530 GNDA_2.n3520 1.70567
R12480 GNDA_2.n3530 GNDA_2.n3519 1.70567
R12481 GNDA_2.n3530 GNDA_2.n3518 1.70567
R12482 GNDA_2.n3530 GNDA_2.n3517 1.70567
R12483 GNDA_2.n3530 GNDA_2.n3516 1.70567
R12484 GNDA_2.n3530 GNDA_2.n3515 1.70567
R12485 GNDA_2.n3530 GNDA_2.n3514 1.70567
R12486 GNDA_2.n3531 GNDA_2.n3530 1.70567
R12487 GNDA_2.n1363 GNDA_2.n1362 1.70567
R12488 GNDA_2.n1363 GNDA_2.n1361 1.70567
R12489 GNDA_2.n1363 GNDA_2.n1360 1.70567
R12490 GNDA_2.n1363 GNDA_2.n1359 1.70567
R12491 GNDA_2.n1363 GNDA_2.n1358 1.70567
R12492 GNDA_2.n1363 GNDA_2.n1357 1.70567
R12493 GNDA_2.n1363 GNDA_2.n1356 1.70567
R12494 GNDA_2.n1363 GNDA_2.n1355 1.70567
R12495 GNDA_2.n1363 GNDA_2.n1354 1.70567
R12496 GNDA_2.n1363 GNDA_2.n1353 1.70567
R12497 GNDA_2.n1363 GNDA_2.n1352 1.70567
R12498 GNDA_2.n1363 GNDA_2.n1351 1.70567
R12499 GNDA_2.n1363 GNDA_2.n1350 1.70567
R12500 GNDA_2.n1363 GNDA_2.n1349 1.70567
R12501 GNDA_2.n1363 GNDA_2.n1348 1.70567
R12502 GNDA_2.n3550 GNDA_2.n1284 1.70567
R12503 GNDA_2.n3548 GNDA_2.n3547 1.70567
R12504 GNDA_2.n3549 GNDA_2.n1316 1.70567
R12505 GNDA_2.n3547 GNDA_2.n3532 1.70567
R12506 GNDA_2.n1316 GNDA_2.n1315 1.70567
R12507 GNDA_2.n3547 GNDA_2.n3533 1.70567
R12508 GNDA_2.n1316 GNDA_2.n1314 1.70567
R12509 GNDA_2.n3547 GNDA_2.n3534 1.70567
R12510 GNDA_2.n1316 GNDA_2.n1313 1.70567
R12511 GNDA_2.n3547 GNDA_2.n3535 1.70567
R12512 GNDA_2.n1316 GNDA_2.n1312 1.70567
R12513 GNDA_2.n3547 GNDA_2.n3536 1.70567
R12514 GNDA_2.n1316 GNDA_2.n1311 1.70567
R12515 GNDA_2.n3547 GNDA_2.n3537 1.70567
R12516 GNDA_2.n1316 GNDA_2.n1310 1.70567
R12517 GNDA_2.n3547 GNDA_2.n3538 1.70567
R12518 GNDA_2.n1316 GNDA_2.n1309 1.70567
R12519 GNDA_2.n3547 GNDA_2.n3539 1.70567
R12520 GNDA_2.n1316 GNDA_2.n1308 1.70567
R12521 GNDA_2.n3547 GNDA_2.n3540 1.70567
R12522 GNDA_2.n1316 GNDA_2.n1307 1.70567
R12523 GNDA_2.n3547 GNDA_2.n3541 1.70567
R12524 GNDA_2.n1316 GNDA_2.n1306 1.70567
R12525 GNDA_2.n3547 GNDA_2.n3542 1.70567
R12526 GNDA_2.n1316 GNDA_2.n1305 1.70567
R12527 GNDA_2.n3547 GNDA_2.n3543 1.70567
R12528 GNDA_2.n1316 GNDA_2.n1304 1.70567
R12529 GNDA_2.n3547 GNDA_2.n3544 1.70567
R12530 GNDA_2.n1316 GNDA_2.n1303 1.70567
R12531 GNDA_2.n3547 GNDA_2.n3545 1.70567
R12532 GNDA_2.n1316 GNDA_2.n1302 1.70567
R12533 GNDA_2.n3547 GNDA_2.n3546 1.70567
R12534 GNDA_2.n1316 GNDA_2.n1301 1.70567
R12535 GNDA_2.n3547 GNDA_2.n1300 1.70567
R12536 GNDA_2.n3437 GNDA_2.n1571 1.69433
R12537 GNDA_2.n3437 GNDA_2.n1568 1.69433
R12538 GNDA_2.n3437 GNDA_2.n1565 1.69433
R12539 GNDA_2.n3043 GNDA_2.n1574 1.69433
R12540 GNDA_2.n3025 GNDA_2.n1574 1.69433
R12541 GNDA_2.n3013 GNDA_2.n1574 1.69433
R12542 GNDA_2.n3953 GNDA_2.n3562 1.69433
R12543 GNDA_2.n3953 GNDA_2.n3559 1.69433
R12544 GNDA_2.n3953 GNDA_2.n3556 1.69433
R12545 GNDA_2.n3888 GNDA_2.n3574 1.69433
R12546 GNDA_2.n3888 GNDA_2.n3571 1.69433
R12547 GNDA_2.n3888 GNDA_2.n3568 1.69433
R12548 GNDA_2.n3819 GNDA_2.n3586 1.69433
R12549 GNDA_2.n3819 GNDA_2.n3583 1.69433
R12550 GNDA_2.n3819 GNDA_2.n3580 1.69433
R12551 GNDA_2.n3750 GNDA_2.n3598 1.69433
R12552 GNDA_2.n3750 GNDA_2.n3595 1.69433
R12553 GNDA_2.n3750 GNDA_2.n3592 1.69433
R12554 GNDA_2.n3681 GNDA_2.n3610 1.69433
R12555 GNDA_2.n3681 GNDA_2.n3607 1.69433
R12556 GNDA_2.n3681 GNDA_2.n3604 1.69433
R12557 GNDA_2.n1196 GNDA_2.n1122 1.69433
R12558 GNDA_2.n1185 GNDA_2.n1122 1.69433
R12559 GNDA_2.n1172 GNDA_2.n1122 1.69433
R12560 GNDA_2.n4074 GNDA_2.n1132 1.69433
R12561 GNDA_2.n4074 GNDA_2.n1129 1.69433
R12562 GNDA_2.n4074 GNDA_2.n1126 1.69433
R12563 GNDA_2.n4155 GNDA_2.n4084 1.69433
R12564 GNDA_2.n4155 GNDA_2.n4081 1.69433
R12565 GNDA_2.n4155 GNDA_2.n4078 1.69433
R12566 GNDA_2.n4264 GNDA_2.n4181 1.69433
R12567 GNDA_2.n4264 GNDA_2.n4178 1.69433
R12568 GNDA_2.n4264 GNDA_2.n4175 1.69433
R12569 GNDA_2.n4265 GNDA_2.n4168 1.69433
R12570 GNDA_2.n4265 GNDA_2.n4164 1.69433
R12571 GNDA_2.n4265 GNDA_2.n4159 1.69433
R12572 GNDA_2.n4535 GNDA_2.n197 1.69433
R12573 GNDA_2.n4535 GNDA_2.n194 1.69433
R12574 GNDA_2.n4535 GNDA_2.n191 1.69433
R12575 GNDA_2.n4676 GNDA_2.n147 1.69433
R12576 GNDA_2.n4685 GNDA_2.n147 1.69433
R12577 GNDA_2.n4694 GNDA_2.n147 1.69433
R12578 GNDA_2.n4772 GNDA_2.n157 1.69433
R12579 GNDA_2.n4772 GNDA_2.n154 1.69433
R12580 GNDA_2.n4772 GNDA_2.n151 1.69433
R12581 GNDA_2.n5212 GNDA_2.n4781 1.69433
R12582 GNDA_2.n5212 GNDA_2.n4778 1.69433
R12583 GNDA_2.n5212 GNDA_2.n4775 1.69433
R12584 GNDA_2.n4611 GNDA_2.n4544 1.69433
R12585 GNDA_2.n4611 GNDA_2.n4541 1.69433
R12586 GNDA_2.n4611 GNDA_2.n4538 1.69433
R12587 GNDA_2.n5147 GNDA_2.n4793 1.69433
R12588 GNDA_2.n5147 GNDA_2.n4790 1.69433
R12589 GNDA_2.n5147 GNDA_2.n4787 1.69433
R12590 GNDA_2.n4864 GNDA_2.n4796 1.69433
R12591 GNDA_2.n4873 GNDA_2.n4796 1.69433
R12592 GNDA_2.n4882 GNDA_2.n4796 1.69433
R12593 GNDA_2.n4987 GNDA_2.n4915 1.69433
R12594 GNDA_2.n4987 GNDA_2.n4912 1.69433
R12595 GNDA_2.n4987 GNDA_2.n4909 1.69433
R12596 GNDA_2.n5063 GNDA_2.n4996 1.69433
R12597 GNDA_2.n5063 GNDA_2.n4993 1.69433
R12598 GNDA_2.n5063 GNDA_2.n4990 1.69433
R12599 GNDA_2.n936 GNDA_2.n707 1.69433
R12600 GNDA_2.n936 GNDA_2.n704 1.69433
R12601 GNDA_2.n936 GNDA_2.n701 1.69433
R12602 GNDA_2.n871 GNDA_2.n719 1.69433
R12603 GNDA_2.n871 GNDA_2.n716 1.69433
R12604 GNDA_2.n871 GNDA_2.n713 1.69433
R12605 GNDA_2.n802 GNDA_2.n731 1.69433
R12606 GNDA_2.n802 GNDA_2.n728 1.69433
R12607 GNDA_2.n802 GNDA_2.n725 1.69433
R12608 GNDA_2.n504 GNDA_2.n430 1.69433
R12609 GNDA_2.n493 GNDA_2.n430 1.69433
R12610 GNDA_2.n480 GNDA_2.n430 1.69433
R12611 GNDA_2.n1014 GNDA_2.n440 1.69433
R12612 GNDA_2.n1014 GNDA_2.n437 1.69433
R12613 GNDA_2.n1014 GNDA_2.n434 1.69433
R12614 GNDA_2.n698 GNDA_2.n626 1.69433
R12615 GNDA_2.n698 GNDA_2.n623 1.69433
R12616 GNDA_2.n698 GNDA_2.n620 1.69433
R12617 GNDA_2.n1031 GNDA_2.n1027 1.69433
R12618 GNDA_2.n1031 GNDA_2.n1023 1.69433
R12619 GNDA_2.n1031 GNDA_2.n1018 1.69433
R12620 GNDA_2.n253 GNDA_2.n187 1.69337
R12621 GNDA_2.n248 GNDA_2.n187 1.69337
R12622 GNDA_2.n240 GNDA_2.n187 1.69337
R12623 GNDA_2.n237 GNDA_2.n187 1.69337
R12624 GNDA_2.n229 GNDA_2.n187 1.69337
R12625 GNDA_2.n224 GNDA_2.n187 1.69337
R12626 GNDA_2.n216 GNDA_2.n187 1.69337
R12627 GNDA_2.n259 GNDA_2.n187 1.69337
R12628 GNDA_2.n3437 GNDA_2.n1573 1.6924
R12629 GNDA_2.n3437 GNDA_2.n1572 1.6924
R12630 GNDA_2.n3437 GNDA_2.n1570 1.6924
R12631 GNDA_2.n3437 GNDA_2.n1569 1.6924
R12632 GNDA_2.n3437 GNDA_2.n1567 1.6924
R12633 GNDA_2.n3437 GNDA_2.n1566 1.6924
R12634 GNDA_2.n3437 GNDA_2.n1564 1.6924
R12635 GNDA_2.n3437 GNDA_2.n1563 1.6924
R12636 GNDA_2.n3053 GNDA_2.n1574 1.6924
R12637 GNDA_2.n3045 GNDA_2.n1574 1.6924
R12638 GNDA_2.n3035 GNDA_2.n1574 1.6924
R12639 GNDA_2.n3033 GNDA_2.n1574 1.6924
R12640 GNDA_2.n3023 GNDA_2.n1574 1.6924
R12641 GNDA_2.n3015 GNDA_2.n1574 1.6924
R12642 GNDA_2.n3005 GNDA_2.n1574 1.6924
R12643 GNDA_2.n3003 GNDA_2.n1574 1.6924
R12644 GNDA_2.n3953 GNDA_2.n3564 1.6924
R12645 GNDA_2.n3953 GNDA_2.n3563 1.6924
R12646 GNDA_2.n3953 GNDA_2.n3561 1.6924
R12647 GNDA_2.n3953 GNDA_2.n3560 1.6924
R12648 GNDA_2.n3953 GNDA_2.n3558 1.6924
R12649 GNDA_2.n3953 GNDA_2.n3557 1.6924
R12650 GNDA_2.n3953 GNDA_2.n3555 1.6924
R12651 GNDA_2.n3953 GNDA_2.n3554 1.6924
R12652 GNDA_2.n3888 GNDA_2.n3576 1.6924
R12653 GNDA_2.n3888 GNDA_2.n3575 1.6924
R12654 GNDA_2.n3888 GNDA_2.n3573 1.6924
R12655 GNDA_2.n3888 GNDA_2.n3572 1.6924
R12656 GNDA_2.n3888 GNDA_2.n3570 1.6924
R12657 GNDA_2.n3888 GNDA_2.n3569 1.6924
R12658 GNDA_2.n3888 GNDA_2.n3567 1.6924
R12659 GNDA_2.n3888 GNDA_2.n3566 1.6924
R12660 GNDA_2.n3819 GNDA_2.n3588 1.6924
R12661 GNDA_2.n3819 GNDA_2.n3587 1.6924
R12662 GNDA_2.n3819 GNDA_2.n3585 1.6924
R12663 GNDA_2.n3819 GNDA_2.n3584 1.6924
R12664 GNDA_2.n3819 GNDA_2.n3582 1.6924
R12665 GNDA_2.n3819 GNDA_2.n3581 1.6924
R12666 GNDA_2.n3819 GNDA_2.n3579 1.6924
R12667 GNDA_2.n3819 GNDA_2.n3578 1.6924
R12668 GNDA_2.n3750 GNDA_2.n3600 1.6924
R12669 GNDA_2.n3750 GNDA_2.n3599 1.6924
R12670 GNDA_2.n3750 GNDA_2.n3597 1.6924
R12671 GNDA_2.n3750 GNDA_2.n3596 1.6924
R12672 GNDA_2.n3750 GNDA_2.n3594 1.6924
R12673 GNDA_2.n3750 GNDA_2.n3593 1.6924
R12674 GNDA_2.n3750 GNDA_2.n3591 1.6924
R12675 GNDA_2.n3750 GNDA_2.n3590 1.6924
R12676 GNDA_2.n3681 GNDA_2.n3612 1.6924
R12677 GNDA_2.n3681 GNDA_2.n3611 1.6924
R12678 GNDA_2.n3681 GNDA_2.n3609 1.6924
R12679 GNDA_2.n3681 GNDA_2.n3608 1.6924
R12680 GNDA_2.n3681 GNDA_2.n3606 1.6924
R12681 GNDA_2.n3681 GNDA_2.n3605 1.6924
R12682 GNDA_2.n3681 GNDA_2.n3603 1.6924
R12683 GNDA_2.n3681 GNDA_2.n3602 1.6924
R12684 GNDA_2.n1204 GNDA_2.n1122 1.6924
R12685 GNDA_2.n1201 GNDA_2.n1122 1.6924
R12686 GNDA_2.n1193 GNDA_2.n1122 1.6924
R12687 GNDA_2.n1188 GNDA_2.n1122 1.6924
R12688 GNDA_2.n1180 GNDA_2.n1122 1.6924
R12689 GNDA_2.n1177 GNDA_2.n1122 1.6924
R12690 GNDA_2.n1169 GNDA_2.n1122 1.6924
R12691 GNDA_2.n1164 GNDA_2.n1122 1.6924
R12692 GNDA_2.n4074 GNDA_2.n1134 1.6924
R12693 GNDA_2.n4074 GNDA_2.n1133 1.6924
R12694 GNDA_2.n4074 GNDA_2.n1131 1.6924
R12695 GNDA_2.n4074 GNDA_2.n1130 1.6924
R12696 GNDA_2.n4074 GNDA_2.n1128 1.6924
R12697 GNDA_2.n4074 GNDA_2.n1127 1.6924
R12698 GNDA_2.n4074 GNDA_2.n1125 1.6924
R12699 GNDA_2.n4074 GNDA_2.n1124 1.6924
R12700 GNDA_2.n4155 GNDA_2.n4086 1.6924
R12701 GNDA_2.n4155 GNDA_2.n4085 1.6924
R12702 GNDA_2.n4155 GNDA_2.n4083 1.6924
R12703 GNDA_2.n4155 GNDA_2.n4082 1.6924
R12704 GNDA_2.n4155 GNDA_2.n4080 1.6924
R12705 GNDA_2.n4155 GNDA_2.n4079 1.6924
R12706 GNDA_2.n4155 GNDA_2.n4077 1.6924
R12707 GNDA_2.n4155 GNDA_2.n4076 1.6924
R12708 GNDA_2.n4264 GNDA_2.n4183 1.6924
R12709 GNDA_2.n4264 GNDA_2.n4182 1.6924
R12710 GNDA_2.n4264 GNDA_2.n4180 1.6924
R12711 GNDA_2.n4264 GNDA_2.n4179 1.6924
R12712 GNDA_2.n4264 GNDA_2.n4177 1.6924
R12713 GNDA_2.n4264 GNDA_2.n4176 1.6924
R12714 GNDA_2.n4264 GNDA_2.n4174 1.6924
R12715 GNDA_2.n4264 GNDA_2.n4173 1.6924
R12716 GNDA_2.n4265 GNDA_2.n4171 1.6924
R12717 GNDA_2.n4265 GNDA_2.n4170 1.6924
R12718 GNDA_2.n4265 GNDA_2.n4167 1.6924
R12719 GNDA_2.n4265 GNDA_2.n4165 1.6924
R12720 GNDA_2.n4265 GNDA_2.n4162 1.6924
R12721 GNDA_2.n4265 GNDA_2.n4161 1.6924
R12722 GNDA_2.n4265 GNDA_2.n4158 1.6924
R12723 GNDA_2.n4265 GNDA_2.n4156 1.6924
R12724 GNDA_2.n4535 GNDA_2.n199 1.6924
R12725 GNDA_2.n4535 GNDA_2.n198 1.6924
R12726 GNDA_2.n4535 GNDA_2.n196 1.6924
R12727 GNDA_2.n4535 GNDA_2.n195 1.6924
R12728 GNDA_2.n4535 GNDA_2.n193 1.6924
R12729 GNDA_2.n4535 GNDA_2.n192 1.6924
R12730 GNDA_2.n4535 GNDA_2.n190 1.6924
R12731 GNDA_2.n4535 GNDA_2.n189 1.6924
R12732 GNDA_2.n4670 GNDA_2.n147 1.6924
R12733 GNDA_2.n4673 GNDA_2.n147 1.6924
R12734 GNDA_2.n4679 GNDA_2.n147 1.6924
R12735 GNDA_2.n4682 GNDA_2.n147 1.6924
R12736 GNDA_2.n4688 GNDA_2.n147 1.6924
R12737 GNDA_2.n4691 GNDA_2.n147 1.6924
R12738 GNDA_2.n4697 GNDA_2.n147 1.6924
R12739 GNDA_2.n4700 GNDA_2.n147 1.6924
R12740 GNDA_2.n4772 GNDA_2.n159 1.6924
R12741 GNDA_2.n4772 GNDA_2.n158 1.6924
R12742 GNDA_2.n4772 GNDA_2.n156 1.6924
R12743 GNDA_2.n4772 GNDA_2.n155 1.6924
R12744 GNDA_2.n4772 GNDA_2.n153 1.6924
R12745 GNDA_2.n4772 GNDA_2.n152 1.6924
R12746 GNDA_2.n4772 GNDA_2.n150 1.6924
R12747 GNDA_2.n4772 GNDA_2.n149 1.6924
R12748 GNDA_2.n5212 GNDA_2.n4783 1.6924
R12749 GNDA_2.n5212 GNDA_2.n4782 1.6924
R12750 GNDA_2.n5212 GNDA_2.n4780 1.6924
R12751 GNDA_2.n5212 GNDA_2.n4779 1.6924
R12752 GNDA_2.n5212 GNDA_2.n4777 1.6924
R12753 GNDA_2.n5212 GNDA_2.n4776 1.6924
R12754 GNDA_2.n5212 GNDA_2.n4774 1.6924
R12755 GNDA_2.n5212 GNDA_2.n4773 1.6924
R12756 GNDA_2.n4611 GNDA_2.n4546 1.6924
R12757 GNDA_2.n4611 GNDA_2.n4545 1.6924
R12758 GNDA_2.n4611 GNDA_2.n4543 1.6924
R12759 GNDA_2.n4611 GNDA_2.n4542 1.6924
R12760 GNDA_2.n4611 GNDA_2.n4540 1.6924
R12761 GNDA_2.n4611 GNDA_2.n4539 1.6924
R12762 GNDA_2.n4611 GNDA_2.n4537 1.6924
R12763 GNDA_2.n4611 GNDA_2.n4536 1.6924
R12764 GNDA_2.n5147 GNDA_2.n4795 1.6924
R12765 GNDA_2.n5147 GNDA_2.n4794 1.6924
R12766 GNDA_2.n5147 GNDA_2.n4792 1.6924
R12767 GNDA_2.n5147 GNDA_2.n4791 1.6924
R12768 GNDA_2.n5147 GNDA_2.n4789 1.6924
R12769 GNDA_2.n5147 GNDA_2.n4788 1.6924
R12770 GNDA_2.n5147 GNDA_2.n4786 1.6924
R12771 GNDA_2.n5147 GNDA_2.n4785 1.6924
R12772 GNDA_2.n4858 GNDA_2.n4796 1.6924
R12773 GNDA_2.n4861 GNDA_2.n4796 1.6924
R12774 GNDA_2.n4867 GNDA_2.n4796 1.6924
R12775 GNDA_2.n4870 GNDA_2.n4796 1.6924
R12776 GNDA_2.n4876 GNDA_2.n4796 1.6924
R12777 GNDA_2.n4879 GNDA_2.n4796 1.6924
R12778 GNDA_2.n4885 GNDA_2.n4796 1.6924
R12779 GNDA_2.n4888 GNDA_2.n4796 1.6924
R12780 GNDA_2.n4987 GNDA_2.n4917 1.6924
R12781 GNDA_2.n4987 GNDA_2.n4916 1.6924
R12782 GNDA_2.n4987 GNDA_2.n4914 1.6924
R12783 GNDA_2.n4987 GNDA_2.n4913 1.6924
R12784 GNDA_2.n4987 GNDA_2.n4911 1.6924
R12785 GNDA_2.n4987 GNDA_2.n4910 1.6924
R12786 GNDA_2.n4987 GNDA_2.n4908 1.6924
R12787 GNDA_2.n4987 GNDA_2.n4907 1.6924
R12788 GNDA_2.n5063 GNDA_2.n4998 1.6924
R12789 GNDA_2.n5063 GNDA_2.n4997 1.6924
R12790 GNDA_2.n5063 GNDA_2.n4995 1.6924
R12791 GNDA_2.n5063 GNDA_2.n4994 1.6924
R12792 GNDA_2.n5063 GNDA_2.n4992 1.6924
R12793 GNDA_2.n5063 GNDA_2.n4991 1.6924
R12794 GNDA_2.n5063 GNDA_2.n4989 1.6924
R12795 GNDA_2.n5063 GNDA_2.n4988 1.6924
R12796 GNDA_2.n936 GNDA_2.n709 1.6924
R12797 GNDA_2.n936 GNDA_2.n708 1.6924
R12798 GNDA_2.n936 GNDA_2.n706 1.6924
R12799 GNDA_2.n936 GNDA_2.n705 1.6924
R12800 GNDA_2.n936 GNDA_2.n703 1.6924
R12801 GNDA_2.n936 GNDA_2.n702 1.6924
R12802 GNDA_2.n936 GNDA_2.n700 1.6924
R12803 GNDA_2.n936 GNDA_2.n699 1.6924
R12804 GNDA_2.n871 GNDA_2.n721 1.6924
R12805 GNDA_2.n871 GNDA_2.n720 1.6924
R12806 GNDA_2.n871 GNDA_2.n718 1.6924
R12807 GNDA_2.n871 GNDA_2.n717 1.6924
R12808 GNDA_2.n871 GNDA_2.n715 1.6924
R12809 GNDA_2.n871 GNDA_2.n714 1.6924
R12810 GNDA_2.n871 GNDA_2.n712 1.6924
R12811 GNDA_2.n871 GNDA_2.n711 1.6924
R12812 GNDA_2.n802 GNDA_2.n733 1.6924
R12813 GNDA_2.n802 GNDA_2.n732 1.6924
R12814 GNDA_2.n802 GNDA_2.n730 1.6924
R12815 GNDA_2.n802 GNDA_2.n729 1.6924
R12816 GNDA_2.n802 GNDA_2.n727 1.6924
R12817 GNDA_2.n802 GNDA_2.n726 1.6924
R12818 GNDA_2.n802 GNDA_2.n724 1.6924
R12819 GNDA_2.n802 GNDA_2.n723 1.6924
R12820 GNDA_2.n512 GNDA_2.n430 1.6924
R12821 GNDA_2.n509 GNDA_2.n430 1.6924
R12822 GNDA_2.n501 GNDA_2.n430 1.6924
R12823 GNDA_2.n496 GNDA_2.n430 1.6924
R12824 GNDA_2.n488 GNDA_2.n430 1.6924
R12825 GNDA_2.n485 GNDA_2.n430 1.6924
R12826 GNDA_2.n477 GNDA_2.n430 1.6924
R12827 GNDA_2.n472 GNDA_2.n430 1.6924
R12828 GNDA_2.n1014 GNDA_2.n442 1.6924
R12829 GNDA_2.n1014 GNDA_2.n441 1.6924
R12830 GNDA_2.n1014 GNDA_2.n439 1.6924
R12831 GNDA_2.n1014 GNDA_2.n438 1.6924
R12832 GNDA_2.n1014 GNDA_2.n436 1.6924
R12833 GNDA_2.n1014 GNDA_2.n435 1.6924
R12834 GNDA_2.n1014 GNDA_2.n433 1.6924
R12835 GNDA_2.n1014 GNDA_2.n432 1.6924
R12836 GNDA_2.n698 GNDA_2.n628 1.6924
R12837 GNDA_2.n698 GNDA_2.n627 1.6924
R12838 GNDA_2.n698 GNDA_2.n625 1.6924
R12839 GNDA_2.n698 GNDA_2.n624 1.6924
R12840 GNDA_2.n698 GNDA_2.n622 1.6924
R12841 GNDA_2.n698 GNDA_2.n621 1.6924
R12842 GNDA_2.n698 GNDA_2.n619 1.6924
R12843 GNDA_2.n698 GNDA_2.n618 1.6924
R12844 GNDA_2.n1031 GNDA_2.n1030 1.6924
R12845 GNDA_2.n1031 GNDA_2.n1029 1.6924
R12846 GNDA_2.n1031 GNDA_2.n1026 1.6924
R12847 GNDA_2.n1031 GNDA_2.n1024 1.6924
R12848 GNDA_2.n1031 GNDA_2.n1021 1.6924
R12849 GNDA_2.n1031 GNDA_2.n1020 1.6924
R12850 GNDA_2.n1031 GNDA_2.n1017 1.6924
R12851 GNDA_2.n1031 GNDA_2.n1015 1.6924
R12852 GNDA_2.n256 GNDA_2.n187 1.6924
R12853 GNDA_2.n245 GNDA_2.n187 1.6924
R12854 GNDA_2.n232 GNDA_2.n187 1.6924
R12855 GNDA_2.n221 GNDA_2.n187 1.6924
R12856 GNDA_2.n4430 GNDA_2.n4429 1.65675
R12857 GNDA_2.n4432 GNDA_2.n4431 1.65675
R12858 GNDA_2.t158 GNDA_2.t288 1.65215
R12859 GNDA_2.t21 GNDA_2.t134 1.65215
R12860 GNDA_2.t112 GNDA_2.t199 1.65215
R12861 GNDA_2.t220 GNDA_2.t90 1.65215
R12862 GNDA_2.n595 GNDA_2.n568 1.56997
R12863 GNDA_2.n570 GNDA_2.n569 1.56997
R12864 GNDA_2.n1833 GNDA_2.t263 1.51652
R12865 GNDA_2.n4304 GNDA_2.n4303 1.5005
R12866 GNDA_2.n4476 GNDA_2.n182 1.5005
R12867 GNDA_2.n3246 GNDA_2.n56 1.47392
R12868 GNDA_2.n2604 GNDA_2.n1846 1.47392
R12869 GNDA_2.n2930 GNDA_2.n2929 1.47392
R12870 GNDA_2.n2224 GNDA_2.n2165 1.47392
R12871 GNDA_2.n3397 GNDA_2.n1673 1.47392
R12872 GNDA_2.n5275 GNDA_2.n116 1.47392
R12873 GNDA_2.n4385 GNDA_2.n344 1.44719
R12874 GNDA_2.n4382 GNDA_2.n4374 1.44719
R12875 GNDA_2.n1031 GNDA_2 1.24042
R12876 GNDA_2.n3068 GNDA_2.n3065 1.22446
R12877 GNDA_2.n5240 GNDA_2.n5239 1.15154
R12878 GNDA_2.n3993 GNDA_2.n3992 1.15154
R12879 GNDA_2.n4441 GNDA_2.n4426 1.13592
R12880 GNDA_2.n4444 GNDA_2.n4443 1.13592
R12881 GNDA_2.n5252 GNDA_2.n5251 1.09425
R12882 GNDA_2.n4000 GNDA_2.n331 1.09425
R12883 GNDA_2.n5247 GNDA_2.n5246 1.07342
R12884 GNDA_2.n3999 GNDA_2.n3998 1.06821
R12885 GNDA_2.n4386 GNDA_2.n4385 1.063
R12886 GNDA_2.n4382 GNDA_2.n4381 1.063
R12887 GNDA_2.n3424 GNDA_2.n3423 1.05258
R12888 GNDA_2.n4446 GNDA_2.n315 0.984875
R12889 GNDA_2.n4422 GNDA_2.n4421 0.984875
R12890 GNDA_2.n562 GNDA_2.n388 0.975928
R12891 GNDA_2.n1076 GNDA_2.n1075 0.975928
R12892 GNDA_2.n3064 GNDA_2.n3063 0.854667
R12893 GNDA_2.n5545 GNDA_2.n59 0.8197
R12894 GNDA_2.n5542 GNDA_2.n5541 0.8197
R12895 GNDA_2.n5538 GNDA_2.n62 0.8197
R12896 GNDA_2.n5537 GNDA_2.n63 0.8197
R12897 GNDA_2.n5472 GNDA_2.n5469 0.8197
R12898 GNDA_2.n5473 GNDA_2.n5463 0.8197
R12899 GNDA_2.n5477 GNDA_2.n5476 0.8197
R12900 GNDA_2.n5481 GNDA_2.n5480 0.8197
R12901 GNDA_2.n1868 GNDA_2.n1848 0.8197
R12902 GNDA_2.n2595 GNDA_2.n1869 0.8197
R12903 GNDA_2.n2594 GNDA_2.n1870 0.8197
R12904 GNDA_2.n1895 GNDA_2.n1893 0.8197
R12905 GNDA_2.n1902 GNDA_2.n1901 0.8197
R12906 GNDA_2.n1890 GNDA_2.n1889 0.8197
R12907 GNDA_2.n1909 GNDA_2.n1908 0.8197
R12908 GNDA_2.n1912 GNDA_2.n1888 0.8197
R12909 GNDA_2.n2920 GNDA_2.n2620 0.8197
R12910 GNDA_2.n2919 GNDA_2.n2621 0.8197
R12911 GNDA_2.n2651 GNDA_2.n2648 0.8197
R12912 GNDA_2.n2650 GNDA_2.n2647 0.8197
R12913 GNDA_2.n2848 GNDA_2.n2847 0.8197
R12914 GNDA_2.n2853 GNDA_2.n2849 0.8197
R12915 GNDA_2.n2852 GNDA_2.n2643 0.8197
R12916 GNDA_2.n2861 GNDA_2.n2860 0.8197
R12917 GNDA_2.n2777 GNDA_2.n2704 0.8197
R12918 GNDA_2.n2776 GNDA_2.n2705 0.8197
R12919 GNDA_2.n2784 GNDA_2.n2684 0.8197
R12920 GNDA_2.n2786 GNDA_2.n2785 0.8197
R12921 GNDA_2.n2792 GNDA_2.n2681 0.8197
R12922 GNDA_2.n2800 GNDA_2.n2678 0.8197
R12923 GNDA_2.n2802 GNDA_2.n2801 0.8197
R12924 GNDA_2.n2810 GNDA_2.n2674 0.8197
R12925 GNDA_2.n2132 GNDA_2.n2131 0.8197
R12926 GNDA_2.n2128 GNDA_2.n2127 0.8197
R12927 GNDA_2.n2124 GNDA_2.n2108 0.8197
R12928 GNDA_2.n2123 GNDA_2.n2120 0.8197
R12929 GNDA_2.n2116 GNDA_2.n2113 0.8197
R12930 GNDA_2.n2110 GNDA_2.n2028 0.8197
R12931 GNDA_2.n2138 GNDA_2.n2137 0.8197
R12932 GNDA_2.n2141 GNDA_2.n2027 0.8197
R12933 GNDA_2.n5448 GNDA_2.n90 0.8197
R12934 GNDA_2.n5447 GNDA_2.n91 0.8197
R12935 GNDA_2.n5367 GNDA_2.n5364 0.8197
R12936 GNDA_2.n5370 GNDA_2.n5369 0.8197
R12937 GNDA_2.n5380 GNDA_2.n5377 0.8197
R12938 GNDA_2.n5381 GNDA_2.n5363 0.8197
R12939 GNDA_2.n5385 GNDA_2.n5384 0.8197
R12940 GNDA_2.n5389 GNDA_2.n5388 0.8197
R12941 GNDA_2.n2321 GNDA_2.n2145 0.8197
R12942 GNDA_2.n2320 GNDA_2.n2146 0.8197
R12943 GNDA_2.n2240 GNDA_2.n2237 0.8197
R12944 GNDA_2.n2243 GNDA_2.n2242 0.8197
R12945 GNDA_2.n2253 GNDA_2.n2250 0.8197
R12946 GNDA_2.n2254 GNDA_2.n2236 0.8197
R12947 GNDA_2.n2258 GNDA_2.n2257 0.8197
R12948 GNDA_2.n2262 GNDA_2.n2261 0.8197
R12949 GNDA_2.n3360 GNDA_2.n3359 0.8197
R12950 GNDA_2.n3346 GNDA_2.n1726 0.8197
R12951 GNDA_2.n3353 GNDA_2.n3347 0.8197
R12952 GNDA_2.n3352 GNDA_2.n3349 0.8197
R12953 GNDA_2.n3365 GNDA_2.n1694 0.8197
R12954 GNDA_2.n1705 GNDA_2.n1701 0.8197
R12955 GNDA_2.n1707 GNDA_2.n1706 0.8197
R12956 GNDA_2.n3400 GNDA_2.n1671 0.8197
R12957 GNDA_2.n5555 GNDA_2.n5554 0.8197
R12958 GNDA_2.n32 GNDA_2.n23 0.8197
R12959 GNDA_2.n39 GNDA_2.n33 0.8197
R12960 GNDA_2.n38 GNDA_2.n35 0.8197
R12961 GNDA_2.n5560 GNDA_2.n1 0.8197
R12962 GNDA_2.n5290 GNDA_2.n5287 0.8197
R12963 GNDA_2.n5293 GNDA_2.n5292 0.8197
R12964 GNDA_2.n5297 GNDA_2.n5296 0.8197
R12965 GNDA_2.n5067 GNDA_2.n5066 0.776542
R12966 GNDA_2.n4930 GNDA_2.n4898 0.776542
R12967 GNDA_2.n4893 GNDA_2.n4892 0.776542
R12968 GNDA_2.n5090 GNDA_2.n5089 0.776542
R12969 GNDA_2.n5216 GNDA_2.n5215 0.776542
R12970 GNDA_2.n4715 GNDA_2.n4714 0.776542
R12971 GNDA_2.n4705 GNDA_2.n4704 0.776542
R12972 GNDA_2.n4217 GNDA_2.n4216 0.776542
R12973 GNDA_2.n4019 GNDA_2.n1241 0.776542
R12974 GNDA_2.n4014 GNDA_2.n1245 0.776542
R12975 GNDA_2.n3975 GNDA_2.n1252 0.776542
R12976 GNDA_2.n3970 GNDA_2.n1256 0.776542
R12977 GNDA_2.n3965 GNDA_2.n1260 0.776542
R12978 GNDA_2.n3957 GNDA_2.n3956 0.776542
R12979 GNDA_2.n2826 GNDA_2.n2825 0.776542
R12980 GNDA_2.n298 GNDA_2.n294 0.776542
R12981 GNDA_2.n4027 GNDA_2.n4026 0.776542
R12982 GNDA_2.n4615 GNDA_2.n4614 0.77295
R12983 GNDA_2.n4309 GNDA_2.n1089 0.77295
R12984 GNDA_2.n4478 GNDA_2.n4477 0.755708
R12985 GNDA_2.n4302 GNDA_2.n4301 0.755708
R12986 GNDA_2.n4302 GNDA_2.n1091 0.751386
R12987 GNDA_2.n4477 GNDA_2.n4474 0.751
R12988 GNDA_2.n3438 GNDA_2.n3437 0.723198
R12989 GNDA_2.n3431 GNDA_2.n3430 0.71925
R12990 GNDA_2.n5252 GNDA_2.n133 0.688
R12991 GNDA_2.n4410 GNDA_2.n331 0.688
R12992 GNDA_2.n3382 GNDA_2.n1683 0.65675
R12993 GNDA_2.n3953 GNDA_2.n3553 0.655048
R12994 GNDA_2.n1069 GNDA_2.n1068 0.577365
R12995 GNDA_2.n613 GNDA_2.n612 0.576819
R12996 GNDA_2.n942 GNDA_2.n613 0.5696
R12997 GNDA_2.n1068 GNDA_2.n400 0.567414
R12998 GNDA_2 GNDA_2.n5464 0.5637
R12999 GNDA_2.n1894 GNDA_2 0.5637
R13000 GNDA_2.n2844 GNDA_2 0.5637
R13001 GNDA_2.n2682 GNDA_2 0.5637
R13002 GNDA_2 GNDA_2.n2109 0.5637
R13003 GNDA_2.n5374 GNDA_2 0.5637
R13004 GNDA_2.n2247 GNDA_2 0.5637
R13005 GNDA_2.n3348 GNDA_2 0.5637
R13006 GNDA_2.n34 GNDA_2 0.5637
R13007 GNDA_2.n4352 GNDA_2.n4351 0.5005
R13008 GNDA_2.n4350 GNDA_2.n4349 0.5005
R13009 GNDA_2.n379 GNDA_2.n378 0.5005
R13010 GNDA_2.n377 GNDA_2.n376 0.5005
R13011 GNDA_2.n602 GNDA_2.n601 0.427583
R13012 GNDA_2.n397 GNDA_2.n386 0.427583
R13013 GNDA_2.n359 GNDA_2.n133 0.40675
R13014 GNDA_2.n4411 GNDA_2.n4410 0.40675
R13015 GNDA_2.n1072 GNDA_2.n398 0.40675
R13016 GNDA_2.n608 GNDA_2.n607 0.40675
R13017 GNDA_2.n3266 GNDA_2.n1833 0.383687
R13018 GNDA_2.n4453 GNDA_2.n310 0.359875
R13019 GNDA_2.n4396 GNDA_2.n4391 0.359875
R13020 GNDA_2.n3065 GNDA_2.n3064 0.339042
R13021 GNDA_2.n3459 GNDA_2.n3442 0.286759
R13022 GNDA_2.n3964 GNDA_2.n3961 0.28175
R13023 GNDA_2.n3969 GNDA_2.n3966 0.28175
R13024 GNDA_2.n3974 GNDA_2.n3971 0.28175
R13025 GNDA_2.n4018 GNDA_2.n4015 0.28175
R13026 GNDA_2.n4308 GNDA_2.n4304 0.28175
R13027 GNDA_2.n4617 GNDA_2.n182 0.28175
R13028 GNDA_2.n4711 GNDA_2.n4709 0.28175
R13029 GNDA_2.n5218 GNDA_2.n142 0.28175
R13030 GNDA_2.n5082 GNDA_2.n5081 0.28175
R13031 GNDA_2.n5078 GNDA_2.n5077 0.28175
R13032 GNDA_2.n5074 GNDA_2.n5073 0.28175
R13033 GNDA_2.n948 GNDA_2.n945 0.28175
R13034 GNDA_2.n953 GNDA_2.n950 0.28175
R13035 GNDA_2.n958 GNDA_2.n955 0.28175
R13036 GNDA_2.n965 GNDA_2.n960 0.28175
R13037 GNDA_2.n4311 GNDA_2.n1085 0.271333
R13038 GNDA_2.n5467 GNDA_2 0.2565
R13039 GNDA_2.n1898 GNDA_2 0.2565
R13040 GNDA_2 GNDA_2.n2843 0.2565
R13041 GNDA_2.n2793 GNDA_2 0.2565
R13042 GNDA_2.n2117 GNDA_2 0.2565
R13043 GNDA_2 GNDA_2.n5373 0.2565
R13044 GNDA_2 GNDA_2.n2246 0.2565
R13045 GNDA_2.n3366 GNDA_2 0.2565
R13046 GNDA_2 GNDA_2.n0 0.2565
R13047 GNDA_2.n3530 GNDA_2.n3513 0.230359
R13048 GNDA_2.n373 GNDA_2.n325 0.229667
R13049 GNDA_2.n368 GNDA_2.n367 0.229667
R13050 GNDA_2.n4400 GNDA_2.n4397 0.229667
R13051 GNDA_2.n4456 GNDA_2.n4455 0.229667
R13052 GNDA_2.n4439 GNDA_2.n4438 0.214042
R13053 GNDA_2.n4450 GNDA_2.n4449 0.214042
R13054 GNDA_2.n4425 GNDA_2.n321 0.214042
R13055 GNDA_2.n4025 GNDA_2.n4020 0.198417
R13056 GNDA_2.n4215 GNDA_2.n4210 0.198417
R13057 GNDA_2.n4473 GNDA_2.n299 0.198417
R13058 GNDA_2.n2693 GNDA_2.n2692 0.188
R13059 GNDA_2.n2823 GNDA_2.n2822 0.188
R13060 GNDA_2.n4707 GNDA_2.n4622 0.188
R13061 GNDA_2.n3415 GNDA_2.n3414 0.15675
R13062 GNDA_2.n3420 GNDA_2.n3419 0.151542
R13063 GNDA_2.n3410 GNDA_2.n3409 0.151542
R13064 GNDA_2.n3388 GNDA_2.n3387 0.147453
R13065 GNDA_2.n1065 GNDA_2.n1064 0.146333
R13066 GNDA_2.n1064 GNDA_2.n405 0.146333
R13067 GNDA_2.n1060 GNDA_2.n405 0.146333
R13068 GNDA_2.n1054 GNDA_2.n410 0.146333
R13069 GNDA_2.n1054 GNDA_2.n1053 0.146333
R13070 GNDA_2.n1053 GNDA_2.n1052 0.146333
R13071 GNDA_2.n1047 GNDA_2.n1046 0.146333
R13072 GNDA_2.n1046 GNDA_2.n420 0.146333
R13073 GNDA_2.n1042 GNDA_2.n420 0.146333
R13074 GNDA_2.n1036 GNDA_2.n425 0.146333
R13075 GNDA_2.n1036 GNDA_2.n1035 0.146333
R13076 GNDA_2.n1035 GNDA_2.n1034 0.146333
R13077 GNDA_2.n5010 GNDA_2.n4904 0.146333
R13078 GNDA_2.n5015 GNDA_2.n5010 0.146333
R13079 GNDA_2.n5016 GNDA_2.n5015 0.146333
R13080 GNDA_2.n5026 GNDA_2.n5025 0.146333
R13081 GNDA_2.n5029 GNDA_2.n5026 0.146333
R13082 GNDA_2.n5029 GNDA_2.n5006 0.146333
R13083 GNDA_2.n5039 GNDA_2.n5004 0.146333
R13084 GNDA_2.n5045 GNDA_2.n5004 0.146333
R13085 GNDA_2.n5046 GNDA_2.n5045 0.146333
R13086 GNDA_2.n5056 GNDA_2.n5055 0.146333
R13087 GNDA_2.n5059 GNDA_2.n5056 0.146333
R13088 GNDA_2.n5059 GNDA_2.n5000 0.146333
R13089 GNDA_2.n4933 GNDA_2.n4929 0.146333
R13090 GNDA_2.n4939 GNDA_2.n4929 0.146333
R13091 GNDA_2.n4940 GNDA_2.n4939 0.146333
R13092 GNDA_2.n4950 GNDA_2.n4949 0.146333
R13093 GNDA_2.n4953 GNDA_2.n4950 0.146333
R13094 GNDA_2.n4953 GNDA_2.n4925 0.146333
R13095 GNDA_2.n4963 GNDA_2.n4923 0.146333
R13096 GNDA_2.n4969 GNDA_2.n4923 0.146333
R13097 GNDA_2.n4970 GNDA_2.n4969 0.146333
R13098 GNDA_2.n4980 GNDA_2.n4979 0.146333
R13099 GNDA_2.n4983 GNDA_2.n4980 0.146333
R13100 GNDA_2.n4983 GNDA_2.n4919 0.146333
R13101 GNDA_2.n4814 GNDA_2.n4813 0.146333
R13102 GNDA_2.n4815 GNDA_2.n4814 0.146333
R13103 GNDA_2.n4816 GNDA_2.n4815 0.146333
R13104 GNDA_2.n4820 GNDA_2.n4819 0.146333
R13105 GNDA_2.n4821 GNDA_2.n4820 0.146333
R13106 GNDA_2.n4822 GNDA_2.n4821 0.146333
R13107 GNDA_2.n4826 GNDA_2.n4825 0.146333
R13108 GNDA_2.n4827 GNDA_2.n4826 0.146333
R13109 GNDA_2.n4828 GNDA_2.n4827 0.146333
R13110 GNDA_2.n4832 GNDA_2.n4831 0.146333
R13111 GNDA_2.n4833 GNDA_2.n4832 0.146333
R13112 GNDA_2.n4834 GNDA_2.n4833 0.146333
R13113 GNDA_2.n5093 GNDA_2.n4808 0.146333
R13114 GNDA_2.n5099 GNDA_2.n4808 0.146333
R13115 GNDA_2.n5100 GNDA_2.n5099 0.146333
R13116 GNDA_2.n5110 GNDA_2.n5109 0.146333
R13117 GNDA_2.n5113 GNDA_2.n5110 0.146333
R13118 GNDA_2.n5113 GNDA_2.n4804 0.146333
R13119 GNDA_2.n5123 GNDA_2.n4802 0.146333
R13120 GNDA_2.n5129 GNDA_2.n4802 0.146333
R13121 GNDA_2.n5130 GNDA_2.n5129 0.146333
R13122 GNDA_2.n5140 GNDA_2.n5139 0.146333
R13123 GNDA_2.n5143 GNDA_2.n5140 0.146333
R13124 GNDA_2.n5143 GNDA_2.n4798 0.146333
R13125 GNDA_2.n4558 GNDA_2.n185 0.146333
R13126 GNDA_2.n4563 GNDA_2.n4558 0.146333
R13127 GNDA_2.n4564 GNDA_2.n4563 0.146333
R13128 GNDA_2.n4574 GNDA_2.n4573 0.146333
R13129 GNDA_2.n4577 GNDA_2.n4574 0.146333
R13130 GNDA_2.n4577 GNDA_2.n4554 0.146333
R13131 GNDA_2.n4587 GNDA_2.n4552 0.146333
R13132 GNDA_2.n4593 GNDA_2.n4552 0.146333
R13133 GNDA_2.n4594 GNDA_2.n4593 0.146333
R13134 GNDA_2.n4604 GNDA_2.n4603 0.146333
R13135 GNDA_2.n4607 GNDA_2.n4604 0.146333
R13136 GNDA_2.n4607 GNDA_2.n4548 0.146333
R13137 GNDA_2.n5159 GNDA_2.n145 0.146333
R13138 GNDA_2.n5164 GNDA_2.n5159 0.146333
R13139 GNDA_2.n5165 GNDA_2.n5164 0.146333
R13140 GNDA_2.n5175 GNDA_2.n5174 0.146333
R13141 GNDA_2.n5178 GNDA_2.n5175 0.146333
R13142 GNDA_2.n5178 GNDA_2.n5155 0.146333
R13143 GNDA_2.n5188 GNDA_2.n5153 0.146333
R13144 GNDA_2.n5194 GNDA_2.n5153 0.146333
R13145 GNDA_2.n5195 GNDA_2.n5194 0.146333
R13146 GNDA_2.n5205 GNDA_2.n5204 0.146333
R13147 GNDA_2.n5208 GNDA_2.n5205 0.146333
R13148 GNDA_2.n5208 GNDA_2.n5149 0.146333
R13149 GNDA_2.n4718 GNDA_2.n171 0.146333
R13150 GNDA_2.n4724 GNDA_2.n171 0.146333
R13151 GNDA_2.n4725 GNDA_2.n4724 0.146333
R13152 GNDA_2.n4735 GNDA_2.n4734 0.146333
R13153 GNDA_2.n4738 GNDA_2.n4735 0.146333
R13154 GNDA_2.n4738 GNDA_2.n167 0.146333
R13155 GNDA_2.n4748 GNDA_2.n165 0.146333
R13156 GNDA_2.n4754 GNDA_2.n165 0.146333
R13157 GNDA_2.n4755 GNDA_2.n4754 0.146333
R13158 GNDA_2.n4765 GNDA_2.n4764 0.146333
R13159 GNDA_2.n4768 GNDA_2.n4765 0.146333
R13160 GNDA_2.n4768 GNDA_2.n161 0.146333
R13161 GNDA_2.n4626 GNDA_2.n4625 0.146333
R13162 GNDA_2.n4627 GNDA_2.n4626 0.146333
R13163 GNDA_2.n4628 GNDA_2.n4627 0.146333
R13164 GNDA_2.n4632 GNDA_2.n4631 0.146333
R13165 GNDA_2.n4633 GNDA_2.n4632 0.146333
R13166 GNDA_2.n4634 GNDA_2.n4633 0.146333
R13167 GNDA_2.n4638 GNDA_2.n4637 0.146333
R13168 GNDA_2.n4639 GNDA_2.n4638 0.146333
R13169 GNDA_2.n4640 GNDA_2.n4639 0.146333
R13170 GNDA_2.n4644 GNDA_2.n4643 0.146333
R13171 GNDA_2.n4645 GNDA_2.n4644 0.146333
R13172 GNDA_2.n4646 GNDA_2.n4645 0.146333
R13173 GNDA_2.n4481 GNDA_2.n211 0.146333
R13174 GNDA_2.n4487 GNDA_2.n211 0.146333
R13175 GNDA_2.n4488 GNDA_2.n4487 0.146333
R13176 GNDA_2.n4498 GNDA_2.n4497 0.146333
R13177 GNDA_2.n4501 GNDA_2.n4498 0.146333
R13178 GNDA_2.n4501 GNDA_2.n207 0.146333
R13179 GNDA_2.n4511 GNDA_2.n205 0.146333
R13180 GNDA_2.n4517 GNDA_2.n205 0.146333
R13181 GNDA_2.n4518 GNDA_2.n4517 0.146333
R13182 GNDA_2.n4528 GNDA_2.n4527 0.146333
R13183 GNDA_2.n4531 GNDA_2.n4528 0.146333
R13184 GNDA_2.n4531 GNDA_2.n201 0.146333
R13185 GNDA_2.n4299 GNDA_2.n4298 0.146333
R13186 GNDA_2.n4298 GNDA_2.n1097 0.146333
R13187 GNDA_2.n4294 GNDA_2.n1097 0.146333
R13188 GNDA_2.n4288 GNDA_2.n1102 0.146333
R13189 GNDA_2.n4288 GNDA_2.n4287 0.146333
R13190 GNDA_2.n4287 GNDA_2.n4286 0.146333
R13191 GNDA_2.n4281 GNDA_2.n4280 0.146333
R13192 GNDA_2.n4280 GNDA_2.n1112 0.146333
R13193 GNDA_2.n4276 GNDA_2.n1112 0.146333
R13194 GNDA_2.n4270 GNDA_2.n1117 0.146333
R13195 GNDA_2.n4270 GNDA_2.n4269 0.146333
R13196 GNDA_2.n4269 GNDA_2.n4268 0.146333
R13197 GNDA_2.n4220 GNDA_2.n4203 0.146333
R13198 GNDA_2.n4224 GNDA_2.n4203 0.146333
R13199 GNDA_2.n4225 GNDA_2.n4224 0.146333
R13200 GNDA_2.n4233 GNDA_2.n4232 0.146333
R13201 GNDA_2.n4236 GNDA_2.n4233 0.146333
R13202 GNDA_2.n4236 GNDA_2.n4195 0.146333
R13203 GNDA_2.n4244 GNDA_2.n4191 0.146333
R13204 GNDA_2.n4248 GNDA_2.n4191 0.146333
R13205 GNDA_2.n4249 GNDA_2.n4248 0.146333
R13206 GNDA_2.n4257 GNDA_2.n4256 0.146333
R13207 GNDA_2.n4260 GNDA_2.n4257 0.146333
R13208 GNDA_2.n4260 GNDA_2.n4185 0.146333
R13209 GNDA_2.n4111 GNDA_2.n4106 0.146333
R13210 GNDA_2.n4115 GNDA_2.n4106 0.146333
R13211 GNDA_2.n4116 GNDA_2.n4115 0.146333
R13212 GNDA_2.n4124 GNDA_2.n4123 0.146333
R13213 GNDA_2.n4127 GNDA_2.n4124 0.146333
R13214 GNDA_2.n4127 GNDA_2.n4098 0.146333
R13215 GNDA_2.n4135 GNDA_2.n4094 0.146333
R13216 GNDA_2.n4139 GNDA_2.n4094 0.146333
R13217 GNDA_2.n4140 GNDA_2.n4139 0.146333
R13218 GNDA_2.n4148 GNDA_2.n4147 0.146333
R13219 GNDA_2.n4151 GNDA_2.n4148 0.146333
R13220 GNDA_2.n4151 GNDA_2.n4088 0.146333
R13221 GNDA_2.n4030 GNDA_2.n1154 0.146333
R13222 GNDA_2.n4034 GNDA_2.n1154 0.146333
R13223 GNDA_2.n4035 GNDA_2.n4034 0.146333
R13224 GNDA_2.n4043 GNDA_2.n4042 0.146333
R13225 GNDA_2.n4046 GNDA_2.n4043 0.146333
R13226 GNDA_2.n4046 GNDA_2.n1146 0.146333
R13227 GNDA_2.n4054 GNDA_2.n1142 0.146333
R13228 GNDA_2.n4058 GNDA_2.n1142 0.146333
R13229 GNDA_2.n4059 GNDA_2.n4058 0.146333
R13230 GNDA_2.n4067 GNDA_2.n4066 0.146333
R13231 GNDA_2.n4070 GNDA_2.n4067 0.146333
R13232 GNDA_2.n4070 GNDA_2.n1136 0.146333
R13233 GNDA_2.n1239 GNDA_2.n1238 0.146333
R13234 GNDA_2.n1238 GNDA_2.n1166 0.146333
R13235 GNDA_2.n1234 GNDA_2.n1166 0.146333
R13236 GNDA_2.n1228 GNDA_2.n1174 0.146333
R13237 GNDA_2.n1228 GNDA_2.n1227 0.146333
R13238 GNDA_2.n1227 GNDA_2.n1226 0.146333
R13239 GNDA_2.n1221 GNDA_2.n1220 0.146333
R13240 GNDA_2.n1220 GNDA_2.n1190 0.146333
R13241 GNDA_2.n1216 GNDA_2.n1190 0.146333
R13242 GNDA_2.n1210 GNDA_2.n1198 0.146333
R13243 GNDA_2.n1210 GNDA_2.n1209 0.146333
R13244 GNDA_2.n1209 GNDA_2.n1208 0.146333
R13245 GNDA_2.n3637 GNDA_2.n3632 0.146333
R13246 GNDA_2.n3641 GNDA_2.n3632 0.146333
R13247 GNDA_2.n3642 GNDA_2.n3641 0.146333
R13248 GNDA_2.n3650 GNDA_2.n3649 0.146333
R13249 GNDA_2.n3653 GNDA_2.n3650 0.146333
R13250 GNDA_2.n3653 GNDA_2.n3624 0.146333
R13251 GNDA_2.n3661 GNDA_2.n3620 0.146333
R13252 GNDA_2.n3665 GNDA_2.n3620 0.146333
R13253 GNDA_2.n3666 GNDA_2.n3665 0.146333
R13254 GNDA_2.n3674 GNDA_2.n3673 0.146333
R13255 GNDA_2.n3677 GNDA_2.n3674 0.146333
R13256 GNDA_2.n3677 GNDA_2.n3614 0.146333
R13257 GNDA_2.n3706 GNDA_2.n3701 0.146333
R13258 GNDA_2.n3710 GNDA_2.n3701 0.146333
R13259 GNDA_2.n3711 GNDA_2.n3710 0.146333
R13260 GNDA_2.n3719 GNDA_2.n3718 0.146333
R13261 GNDA_2.n3722 GNDA_2.n3719 0.146333
R13262 GNDA_2.n3722 GNDA_2.n3693 0.146333
R13263 GNDA_2.n3730 GNDA_2.n3689 0.146333
R13264 GNDA_2.n3734 GNDA_2.n3689 0.146333
R13265 GNDA_2.n3735 GNDA_2.n3734 0.146333
R13266 GNDA_2.n3743 GNDA_2.n3742 0.146333
R13267 GNDA_2.n3746 GNDA_2.n3743 0.146333
R13268 GNDA_2.n3746 GNDA_2.n3683 0.146333
R13269 GNDA_2.n3775 GNDA_2.n3770 0.146333
R13270 GNDA_2.n3779 GNDA_2.n3770 0.146333
R13271 GNDA_2.n3780 GNDA_2.n3779 0.146333
R13272 GNDA_2.n3788 GNDA_2.n3787 0.146333
R13273 GNDA_2.n3791 GNDA_2.n3788 0.146333
R13274 GNDA_2.n3791 GNDA_2.n3762 0.146333
R13275 GNDA_2.n3799 GNDA_2.n3758 0.146333
R13276 GNDA_2.n3803 GNDA_2.n3758 0.146333
R13277 GNDA_2.n3804 GNDA_2.n3803 0.146333
R13278 GNDA_2.n3812 GNDA_2.n3811 0.146333
R13279 GNDA_2.n3815 GNDA_2.n3812 0.146333
R13280 GNDA_2.n3815 GNDA_2.n3752 0.146333
R13281 GNDA_2.n3844 GNDA_2.n3839 0.146333
R13282 GNDA_2.n3848 GNDA_2.n3839 0.146333
R13283 GNDA_2.n3849 GNDA_2.n3848 0.146333
R13284 GNDA_2.n3857 GNDA_2.n3856 0.146333
R13285 GNDA_2.n3860 GNDA_2.n3857 0.146333
R13286 GNDA_2.n3860 GNDA_2.n3831 0.146333
R13287 GNDA_2.n3868 GNDA_2.n3827 0.146333
R13288 GNDA_2.n3872 GNDA_2.n3827 0.146333
R13289 GNDA_2.n3873 GNDA_2.n3872 0.146333
R13290 GNDA_2.n3881 GNDA_2.n3880 0.146333
R13291 GNDA_2.n3884 GNDA_2.n3881 0.146333
R13292 GNDA_2.n3884 GNDA_2.n3821 0.146333
R13293 GNDA_2.n3900 GNDA_2.n1265 0.146333
R13294 GNDA_2.n3905 GNDA_2.n3900 0.146333
R13295 GNDA_2.n3906 GNDA_2.n3905 0.146333
R13296 GNDA_2.n3916 GNDA_2.n3915 0.146333
R13297 GNDA_2.n3919 GNDA_2.n3916 0.146333
R13298 GNDA_2.n3919 GNDA_2.n3896 0.146333
R13299 GNDA_2.n3929 GNDA_2.n3894 0.146333
R13300 GNDA_2.n3935 GNDA_2.n3894 0.146333
R13301 GNDA_2.n3936 GNDA_2.n3935 0.146333
R13302 GNDA_2.n3946 GNDA_2.n3945 0.146333
R13303 GNDA_2.n3949 GNDA_2.n3946 0.146333
R13304 GNDA_2.n3949 GNDA_2.n3890 0.146333
R13305 GNDA_2.n3001 GNDA_2.n2998 0.146333
R13306 GNDA_2.n3007 GNDA_2.n2998 0.146333
R13307 GNDA_2.n3007 GNDA_2.n2996 0.146333
R13308 GNDA_2.n3017 GNDA_2.n2992 0.146333
R13309 GNDA_2.n3021 GNDA_2.n2992 0.146333
R13310 GNDA_2.n3021 GNDA_2.n2990 0.146333
R13311 GNDA_2.n3031 GNDA_2.n2986 0.146333
R13312 GNDA_2.n3037 GNDA_2.n2986 0.146333
R13313 GNDA_2.n3037 GNDA_2.n2984 0.146333
R13314 GNDA_2.n3047 GNDA_2.n2980 0.146333
R13315 GNDA_2.n3051 GNDA_2.n2980 0.146333
R13316 GNDA_2.n3051 GNDA_2.n2978 0.146333
R13317 GNDA_2.n1591 GNDA_2.n1590 0.146333
R13318 GNDA_2.n1591 GNDA_2.n1585 0.146333
R13319 GNDA_2.n1601 GNDA_2.n1583 0.146333
R13320 GNDA_2.n1609 GNDA_2.n1583 0.146333
R13321 GNDA_2.n1610 GNDA_2.n1609 0.146333
R13322 GNDA_2.n1620 GNDA_2.n1619 0.146333
R13323 GNDA_2.n1621 GNDA_2.n1620 0.146333
R13324 GNDA_2.n1621 GNDA_2.n1579 0.146333
R13325 GNDA_2.n1631 GNDA_2.n1577 0.146333
R13326 GNDA_2.n1639 GNDA_2.n1577 0.146333
R13327 GNDA_2.n1640 GNDA_2.n1639 0.146333
R13328 GNDA_2.n1588 GNDA_2.n1586 0.146333
R13329 GNDA_2.n1594 GNDA_2.n1586 0.146333
R13330 GNDA_2.n1595 GNDA_2.n1594 0.146333
R13331 GNDA_2.n1605 GNDA_2.n1604 0.146333
R13332 GNDA_2.n1608 GNDA_2.n1605 0.146333
R13333 GNDA_2.n1608 GNDA_2.n1582 0.146333
R13334 GNDA_2.n1618 GNDA_2.n1580 0.146333
R13335 GNDA_2.n1624 GNDA_2.n1580 0.146333
R13336 GNDA_2.n1625 GNDA_2.n1624 0.146333
R13337 GNDA_2.n1635 GNDA_2.n1634 0.146333
R13338 GNDA_2.n1638 GNDA_2.n1635 0.146333
R13339 GNDA_2.n1638 GNDA_2.n1576 0.146333
R13340 GNDA_2.n292 GNDA_2.n291 0.146333
R13341 GNDA_2.n291 GNDA_2.n219 0.146333
R13342 GNDA_2.n287 GNDA_2.n219 0.146333
R13343 GNDA_2.n281 GNDA_2.n227 0.146333
R13344 GNDA_2.n281 GNDA_2.n280 0.146333
R13345 GNDA_2.n280 GNDA_2.n279 0.146333
R13346 GNDA_2.n274 GNDA_2.n273 0.146333
R13347 GNDA_2.n273 GNDA_2.n243 0.146333
R13348 GNDA_2.n269 GNDA_2.n243 0.146333
R13349 GNDA_2.n263 GNDA_2.n251 0.146333
R13350 GNDA_2.n263 GNDA_2.n262 0.146333
R13351 GNDA_2.n262 GNDA_2.n261 0.146333
R13352 GNDA_2.n654 GNDA_2.n648 0.146333
R13353 GNDA_2.n658 GNDA_2.n648 0.146333
R13354 GNDA_2.n659 GNDA_2.n658 0.146333
R13355 GNDA_2.n667 GNDA_2.n666 0.146333
R13356 GNDA_2.n670 GNDA_2.n667 0.146333
R13357 GNDA_2.n670 GNDA_2.n640 0.146333
R13358 GNDA_2.n678 GNDA_2.n636 0.146333
R13359 GNDA_2.n682 GNDA_2.n636 0.146333
R13360 GNDA_2.n683 GNDA_2.n682 0.146333
R13361 GNDA_2.n691 GNDA_2.n690 0.146333
R13362 GNDA_2.n694 GNDA_2.n691 0.146333
R13363 GNDA_2.n694 GNDA_2.n630 0.146333
R13364 GNDA_2.n970 GNDA_2.n462 0.146333
R13365 GNDA_2.n974 GNDA_2.n462 0.146333
R13366 GNDA_2.n975 GNDA_2.n974 0.146333
R13367 GNDA_2.n983 GNDA_2.n982 0.146333
R13368 GNDA_2.n986 GNDA_2.n983 0.146333
R13369 GNDA_2.n986 GNDA_2.n454 0.146333
R13370 GNDA_2.n994 GNDA_2.n450 0.146333
R13371 GNDA_2.n998 GNDA_2.n450 0.146333
R13372 GNDA_2.n999 GNDA_2.n998 0.146333
R13373 GNDA_2.n1007 GNDA_2.n1006 0.146333
R13374 GNDA_2.n1010 GNDA_2.n1007 0.146333
R13375 GNDA_2.n1010 GNDA_2.n444 0.146333
R13376 GNDA_2.n547 GNDA_2.n546 0.146333
R13377 GNDA_2.n546 GNDA_2.n474 0.146333
R13378 GNDA_2.n542 GNDA_2.n474 0.146333
R13379 GNDA_2.n536 GNDA_2.n482 0.146333
R13380 GNDA_2.n536 GNDA_2.n535 0.146333
R13381 GNDA_2.n535 GNDA_2.n534 0.146333
R13382 GNDA_2.n529 GNDA_2.n528 0.146333
R13383 GNDA_2.n528 GNDA_2.n498 0.146333
R13384 GNDA_2.n524 GNDA_2.n498 0.146333
R13385 GNDA_2.n518 GNDA_2.n506 0.146333
R13386 GNDA_2.n518 GNDA_2.n517 0.146333
R13387 GNDA_2.n517 GNDA_2.n516 0.146333
R13388 GNDA_2.n758 GNDA_2.n753 0.146333
R13389 GNDA_2.n762 GNDA_2.n753 0.146333
R13390 GNDA_2.n763 GNDA_2.n762 0.146333
R13391 GNDA_2.n771 GNDA_2.n770 0.146333
R13392 GNDA_2.n774 GNDA_2.n771 0.146333
R13393 GNDA_2.n774 GNDA_2.n745 0.146333
R13394 GNDA_2.n782 GNDA_2.n741 0.146333
R13395 GNDA_2.n786 GNDA_2.n741 0.146333
R13396 GNDA_2.n787 GNDA_2.n786 0.146333
R13397 GNDA_2.n795 GNDA_2.n794 0.146333
R13398 GNDA_2.n798 GNDA_2.n795 0.146333
R13399 GNDA_2.n798 GNDA_2.n735 0.146333
R13400 GNDA_2.n827 GNDA_2.n822 0.146333
R13401 GNDA_2.n831 GNDA_2.n822 0.146333
R13402 GNDA_2.n832 GNDA_2.n831 0.146333
R13403 GNDA_2.n840 GNDA_2.n839 0.146333
R13404 GNDA_2.n843 GNDA_2.n840 0.146333
R13405 GNDA_2.n843 GNDA_2.n814 0.146333
R13406 GNDA_2.n851 GNDA_2.n810 0.146333
R13407 GNDA_2.n855 GNDA_2.n810 0.146333
R13408 GNDA_2.n856 GNDA_2.n855 0.146333
R13409 GNDA_2.n864 GNDA_2.n863 0.146333
R13410 GNDA_2.n867 GNDA_2.n864 0.146333
R13411 GNDA_2.n867 GNDA_2.n804 0.146333
R13412 GNDA_2.n883 GNDA_2.n615 0.146333
R13413 GNDA_2.n888 GNDA_2.n883 0.146333
R13414 GNDA_2.n889 GNDA_2.n888 0.146333
R13415 GNDA_2.n899 GNDA_2.n898 0.146333
R13416 GNDA_2.n902 GNDA_2.n899 0.146333
R13417 GNDA_2.n902 GNDA_2.n879 0.146333
R13418 GNDA_2.n912 GNDA_2.n877 0.146333
R13419 GNDA_2.n918 GNDA_2.n877 0.146333
R13420 GNDA_2.n919 GNDA_2.n918 0.146333
R13421 GNDA_2.n929 GNDA_2.n928 0.146333
R13422 GNDA_2.n932 GNDA_2.n929 0.146333
R13423 GNDA_2.n932 GNDA_2.n873 0.146333
R13424 GNDA_2.n1066 GNDA_2.n1065 0.135917
R13425 GNDA_2.n1060 GNDA_2.n1059 0.135917
R13426 GNDA_2.n1058 GNDA_2.n410 0.135917
R13427 GNDA_2.n1052 GNDA_2.n415 0.135917
R13428 GNDA_2.n1048 GNDA_2.n1047 0.135917
R13429 GNDA_2.n1042 GNDA_2.n1041 0.135917
R13430 GNDA_2.n1040 GNDA_2.n425 0.135917
R13431 GNDA_2.n5065 GNDA_2.n4904 0.135917
R13432 GNDA_2.n5019 GNDA_2.n5016 0.135917
R13433 GNDA_2.n5025 GNDA_2.n5008 0.135917
R13434 GNDA_2.n5035 GNDA_2.n5006 0.135917
R13435 GNDA_2.n5039 GNDA_2.n5036 0.135917
R13436 GNDA_2.n5049 GNDA_2.n5046 0.135917
R13437 GNDA_2.n5055 GNDA_2.n5002 0.135917
R13438 GNDA_2.n4933 GNDA_2.n4931 0.135917
R13439 GNDA_2.n4943 GNDA_2.n4940 0.135917
R13440 GNDA_2.n4949 GNDA_2.n4927 0.135917
R13441 GNDA_2.n4959 GNDA_2.n4925 0.135917
R13442 GNDA_2.n4963 GNDA_2.n4960 0.135917
R13443 GNDA_2.n4973 GNDA_2.n4970 0.135917
R13444 GNDA_2.n4979 GNDA_2.n4921 0.135917
R13445 GNDA_2.n4891 GNDA_2.n4813 0.135917
R13446 GNDA_2.n4817 GNDA_2.n4816 0.135917
R13447 GNDA_2.n4819 GNDA_2.n4818 0.135917
R13448 GNDA_2.n4823 GNDA_2.n4822 0.135917
R13449 GNDA_2.n4825 GNDA_2.n4824 0.135917
R13450 GNDA_2.n4829 GNDA_2.n4828 0.135917
R13451 GNDA_2.n4831 GNDA_2.n4830 0.135917
R13452 GNDA_2.n5093 GNDA_2.n5091 0.135917
R13453 GNDA_2.n5103 GNDA_2.n5100 0.135917
R13454 GNDA_2.n5109 GNDA_2.n4806 0.135917
R13455 GNDA_2.n5119 GNDA_2.n4804 0.135917
R13456 GNDA_2.n5123 GNDA_2.n5120 0.135917
R13457 GNDA_2.n5133 GNDA_2.n5130 0.135917
R13458 GNDA_2.n5139 GNDA_2.n4800 0.135917
R13459 GNDA_2.n4613 GNDA_2.n185 0.135917
R13460 GNDA_2.n4567 GNDA_2.n4564 0.135917
R13461 GNDA_2.n4573 GNDA_2.n4556 0.135917
R13462 GNDA_2.n4583 GNDA_2.n4554 0.135917
R13463 GNDA_2.n4587 GNDA_2.n4584 0.135917
R13464 GNDA_2.n4597 GNDA_2.n4594 0.135917
R13465 GNDA_2.n4603 GNDA_2.n4550 0.135917
R13466 GNDA_2.n5214 GNDA_2.n145 0.135917
R13467 GNDA_2.n5168 GNDA_2.n5165 0.135917
R13468 GNDA_2.n5174 GNDA_2.n5157 0.135917
R13469 GNDA_2.n5184 GNDA_2.n5155 0.135917
R13470 GNDA_2.n5188 GNDA_2.n5185 0.135917
R13471 GNDA_2.n5198 GNDA_2.n5195 0.135917
R13472 GNDA_2.n5204 GNDA_2.n5151 0.135917
R13473 GNDA_2.n4718 GNDA_2.n4716 0.135917
R13474 GNDA_2.n4728 GNDA_2.n4725 0.135917
R13475 GNDA_2.n4734 GNDA_2.n169 0.135917
R13476 GNDA_2.n4744 GNDA_2.n167 0.135917
R13477 GNDA_2.n4748 GNDA_2.n4745 0.135917
R13478 GNDA_2.n4758 GNDA_2.n4755 0.135917
R13479 GNDA_2.n4764 GNDA_2.n163 0.135917
R13480 GNDA_2.n4703 GNDA_2.n4625 0.135917
R13481 GNDA_2.n4629 GNDA_2.n4628 0.135917
R13482 GNDA_2.n4631 GNDA_2.n4630 0.135917
R13483 GNDA_2.n4635 GNDA_2.n4634 0.135917
R13484 GNDA_2.n4637 GNDA_2.n4636 0.135917
R13485 GNDA_2.n4641 GNDA_2.n4640 0.135917
R13486 GNDA_2.n4643 GNDA_2.n4642 0.135917
R13487 GNDA_2.n4481 GNDA_2.n4479 0.135917
R13488 GNDA_2.n4491 GNDA_2.n4488 0.135917
R13489 GNDA_2.n4497 GNDA_2.n209 0.135917
R13490 GNDA_2.n4507 GNDA_2.n207 0.135917
R13491 GNDA_2.n4511 GNDA_2.n4508 0.135917
R13492 GNDA_2.n4521 GNDA_2.n4518 0.135917
R13493 GNDA_2.n4527 GNDA_2.n203 0.135917
R13494 GNDA_2.n4300 GNDA_2.n4299 0.135917
R13495 GNDA_2.n4294 GNDA_2.n4293 0.135917
R13496 GNDA_2.n4292 GNDA_2.n1102 0.135917
R13497 GNDA_2.n4286 GNDA_2.n1107 0.135917
R13498 GNDA_2.n4282 GNDA_2.n4281 0.135917
R13499 GNDA_2.n4276 GNDA_2.n4275 0.135917
R13500 GNDA_2.n4274 GNDA_2.n1117 0.135917
R13501 GNDA_2.n4220 GNDA_2.n4218 0.135917
R13502 GNDA_2.n4228 GNDA_2.n4225 0.135917
R13503 GNDA_2.n4232 GNDA_2.n4199 0.135917
R13504 GNDA_2.n4240 GNDA_2.n4195 0.135917
R13505 GNDA_2.n4244 GNDA_2.n4241 0.135917
R13506 GNDA_2.n4252 GNDA_2.n4249 0.135917
R13507 GNDA_2.n4256 GNDA_2.n4187 0.135917
R13508 GNDA_2.n4111 GNDA_2.n4109 0.135917
R13509 GNDA_2.n4119 GNDA_2.n4116 0.135917
R13510 GNDA_2.n4123 GNDA_2.n4102 0.135917
R13511 GNDA_2.n4131 GNDA_2.n4098 0.135917
R13512 GNDA_2.n4135 GNDA_2.n4132 0.135917
R13513 GNDA_2.n4143 GNDA_2.n4140 0.135917
R13514 GNDA_2.n4147 GNDA_2.n4090 0.135917
R13515 GNDA_2.n4030 GNDA_2.n4028 0.135917
R13516 GNDA_2.n4038 GNDA_2.n4035 0.135917
R13517 GNDA_2.n4042 GNDA_2.n1150 0.135917
R13518 GNDA_2.n4050 GNDA_2.n1146 0.135917
R13519 GNDA_2.n4054 GNDA_2.n4051 0.135917
R13520 GNDA_2.n4062 GNDA_2.n4059 0.135917
R13521 GNDA_2.n4066 GNDA_2.n1138 0.135917
R13522 GNDA_2.n1240 GNDA_2.n1239 0.135917
R13523 GNDA_2.n1234 GNDA_2.n1233 0.135917
R13524 GNDA_2.n1232 GNDA_2.n1174 0.135917
R13525 GNDA_2.n1226 GNDA_2.n1182 0.135917
R13526 GNDA_2.n1222 GNDA_2.n1221 0.135917
R13527 GNDA_2.n1216 GNDA_2.n1215 0.135917
R13528 GNDA_2.n1214 GNDA_2.n1198 0.135917
R13529 GNDA_2.n3637 GNDA_2.n3635 0.135917
R13530 GNDA_2.n3645 GNDA_2.n3642 0.135917
R13531 GNDA_2.n3649 GNDA_2.n3628 0.135917
R13532 GNDA_2.n3657 GNDA_2.n3624 0.135917
R13533 GNDA_2.n3661 GNDA_2.n3658 0.135917
R13534 GNDA_2.n3669 GNDA_2.n3666 0.135917
R13535 GNDA_2.n3673 GNDA_2.n3616 0.135917
R13536 GNDA_2.n3706 GNDA_2.n3704 0.135917
R13537 GNDA_2.n3714 GNDA_2.n3711 0.135917
R13538 GNDA_2.n3718 GNDA_2.n3697 0.135917
R13539 GNDA_2.n3726 GNDA_2.n3693 0.135917
R13540 GNDA_2.n3730 GNDA_2.n3727 0.135917
R13541 GNDA_2.n3738 GNDA_2.n3735 0.135917
R13542 GNDA_2.n3742 GNDA_2.n3685 0.135917
R13543 GNDA_2.n3775 GNDA_2.n3773 0.135917
R13544 GNDA_2.n3783 GNDA_2.n3780 0.135917
R13545 GNDA_2.n3787 GNDA_2.n3766 0.135917
R13546 GNDA_2.n3795 GNDA_2.n3762 0.135917
R13547 GNDA_2.n3799 GNDA_2.n3796 0.135917
R13548 GNDA_2.n3807 GNDA_2.n3804 0.135917
R13549 GNDA_2.n3811 GNDA_2.n3754 0.135917
R13550 GNDA_2.n3844 GNDA_2.n3842 0.135917
R13551 GNDA_2.n3852 GNDA_2.n3849 0.135917
R13552 GNDA_2.n3856 GNDA_2.n3835 0.135917
R13553 GNDA_2.n3864 GNDA_2.n3831 0.135917
R13554 GNDA_2.n3868 GNDA_2.n3865 0.135917
R13555 GNDA_2.n3876 GNDA_2.n3873 0.135917
R13556 GNDA_2.n3880 GNDA_2.n3823 0.135917
R13557 GNDA_2.n3955 GNDA_2.n1265 0.135917
R13558 GNDA_2.n3909 GNDA_2.n3906 0.135917
R13559 GNDA_2.n3915 GNDA_2.n3898 0.135917
R13560 GNDA_2.n3925 GNDA_2.n3896 0.135917
R13561 GNDA_2.n3929 GNDA_2.n3926 0.135917
R13562 GNDA_2.n3939 GNDA_2.n3936 0.135917
R13563 GNDA_2.n3945 GNDA_2.n3892 0.135917
R13564 GNDA_2.n3011 GNDA_2.n2996 0.135917
R13565 GNDA_2.n3017 GNDA_2.n2994 0.135917
R13566 GNDA_2.n3027 GNDA_2.n2990 0.135917
R13567 GNDA_2.n3031 GNDA_2.n2988 0.135917
R13568 GNDA_2.n3041 GNDA_2.n2984 0.135917
R13569 GNDA_2.n3047 GNDA_2.n2982 0.135917
R13570 GNDA_2.n3056 GNDA_2.n2978 0.135917
R13571 GNDA_2.n1599 GNDA_2.n1585 0.135917
R13572 GNDA_2.n1601 GNDA_2.n1600 0.135917
R13573 GNDA_2.n1611 GNDA_2.n1610 0.135917
R13574 GNDA_2.n1619 GNDA_2.n1581 0.135917
R13575 GNDA_2.n1629 GNDA_2.n1579 0.135917
R13576 GNDA_2.n1631 GNDA_2.n1630 0.135917
R13577 GNDA_2.n3434 GNDA_2.n1640 0.135917
R13578 GNDA_2.n1598 GNDA_2.n1595 0.135917
R13579 GNDA_2.n1604 GNDA_2.n1584 0.135917
R13580 GNDA_2.n1614 GNDA_2.n1582 0.135917
R13581 GNDA_2.n1618 GNDA_2.n1615 0.135917
R13582 GNDA_2.n1628 GNDA_2.n1625 0.135917
R13583 GNDA_2.n1634 GNDA_2.n1578 0.135917
R13584 GNDA_2.n3435 GNDA_2.n1576 0.135917
R13585 GNDA_2.n293 GNDA_2.n292 0.135917
R13586 GNDA_2.n287 GNDA_2.n286 0.135917
R13587 GNDA_2.n285 GNDA_2.n227 0.135917
R13588 GNDA_2.n279 GNDA_2.n235 0.135917
R13589 GNDA_2.n275 GNDA_2.n274 0.135917
R13590 GNDA_2.n269 GNDA_2.n268 0.135917
R13591 GNDA_2.n267 GNDA_2.n251 0.135917
R13592 GNDA_2.n654 GNDA_2.n652 0.135917
R13593 GNDA_2.n662 GNDA_2.n659 0.135917
R13594 GNDA_2.n666 GNDA_2.n644 0.135917
R13595 GNDA_2.n674 GNDA_2.n640 0.135917
R13596 GNDA_2.n678 GNDA_2.n675 0.135917
R13597 GNDA_2.n686 GNDA_2.n683 0.135917
R13598 GNDA_2.n690 GNDA_2.n632 0.135917
R13599 GNDA_2.n970 GNDA_2.n968 0.135917
R13600 GNDA_2.n978 GNDA_2.n975 0.135917
R13601 GNDA_2.n982 GNDA_2.n458 0.135917
R13602 GNDA_2.n990 GNDA_2.n454 0.135917
R13603 GNDA_2.n994 GNDA_2.n991 0.135917
R13604 GNDA_2.n1002 GNDA_2.n999 0.135917
R13605 GNDA_2.n1006 GNDA_2.n446 0.135917
R13606 GNDA_2.n548 GNDA_2.n547 0.135917
R13607 GNDA_2.n542 GNDA_2.n541 0.135917
R13608 GNDA_2.n540 GNDA_2.n482 0.135917
R13609 GNDA_2.n534 GNDA_2.n490 0.135917
R13610 GNDA_2.n530 GNDA_2.n529 0.135917
R13611 GNDA_2.n524 GNDA_2.n523 0.135917
R13612 GNDA_2.n522 GNDA_2.n506 0.135917
R13613 GNDA_2.n758 GNDA_2.n756 0.135917
R13614 GNDA_2.n766 GNDA_2.n763 0.135917
R13615 GNDA_2.n770 GNDA_2.n749 0.135917
R13616 GNDA_2.n778 GNDA_2.n745 0.135917
R13617 GNDA_2.n782 GNDA_2.n779 0.135917
R13618 GNDA_2.n790 GNDA_2.n787 0.135917
R13619 GNDA_2.n794 GNDA_2.n737 0.135917
R13620 GNDA_2.n827 GNDA_2.n825 0.135917
R13621 GNDA_2.n835 GNDA_2.n832 0.135917
R13622 GNDA_2.n839 GNDA_2.n818 0.135917
R13623 GNDA_2.n847 GNDA_2.n814 0.135917
R13624 GNDA_2.n851 GNDA_2.n848 0.135917
R13625 GNDA_2.n859 GNDA_2.n856 0.135917
R13626 GNDA_2.n863 GNDA_2.n806 0.135917
R13627 GNDA_2.n938 GNDA_2.n615 0.135917
R13628 GNDA_2.n892 GNDA_2.n889 0.135917
R13629 GNDA_2.n898 GNDA_2.n881 0.135917
R13630 GNDA_2.n908 GNDA_2.n879 0.135917
R13631 GNDA_2.n912 GNDA_2.n909 0.135917
R13632 GNDA_2.n922 GNDA_2.n919 0.135917
R13633 GNDA_2.n928 GNDA_2.n875 0.135917
R13634 GNDA_2.n3437 GNDA_2.n1574 0.135331
R13635 GNDA_2.n1059 GNDA_2.n1058 0.1255
R13636 GNDA_2.n1048 GNDA_2.n415 0.1255
R13637 GNDA_2.n1041 GNDA_2.n1040 0.1255
R13638 GNDA_2.n600 GNDA_2.n599 0.1255
R13639 GNDA_2.n4339 GNDA_2.n4338 0.1255
R13640 GNDA_2.n5019 GNDA_2.n5008 0.1255
R13641 GNDA_2.n5036 GNDA_2.n5035 0.1255
R13642 GNDA_2.n5049 GNDA_2.n5002 0.1255
R13643 GNDA_2.n4943 GNDA_2.n4927 0.1255
R13644 GNDA_2.n4960 GNDA_2.n4959 0.1255
R13645 GNDA_2.n4973 GNDA_2.n4921 0.1255
R13646 GNDA_2.n4818 GNDA_2.n4817 0.1255
R13647 GNDA_2.n4824 GNDA_2.n4823 0.1255
R13648 GNDA_2.n4830 GNDA_2.n4829 0.1255
R13649 GNDA_2.n5103 GNDA_2.n4806 0.1255
R13650 GNDA_2.n5120 GNDA_2.n5119 0.1255
R13651 GNDA_2.n5133 GNDA_2.n4800 0.1255
R13652 GNDA_2.n4567 GNDA_2.n4556 0.1255
R13653 GNDA_2.n4584 GNDA_2.n4583 0.1255
R13654 GNDA_2.n4597 GNDA_2.n4550 0.1255
R13655 GNDA_2.n5168 GNDA_2.n5157 0.1255
R13656 GNDA_2.n5185 GNDA_2.n5184 0.1255
R13657 GNDA_2.n5198 GNDA_2.n5151 0.1255
R13658 GNDA_2.n4728 GNDA_2.n169 0.1255
R13659 GNDA_2.n4745 GNDA_2.n4744 0.1255
R13660 GNDA_2.n4758 GNDA_2.n163 0.1255
R13661 GNDA_2.n4630 GNDA_2.n4629 0.1255
R13662 GNDA_2.n4636 GNDA_2.n4635 0.1255
R13663 GNDA_2.n4642 GNDA_2.n4641 0.1255
R13664 GNDA_2.n4491 GNDA_2.n209 0.1255
R13665 GNDA_2.n4508 GNDA_2.n4507 0.1255
R13666 GNDA_2.n4521 GNDA_2.n203 0.1255
R13667 GNDA_2.n371 GNDA_2.n370 0.1255
R13668 GNDA_2.n4357 GNDA_2.n4356 0.1255
R13669 GNDA_2.n4398 GNDA_2.n337 0.1255
R13670 GNDA_2.n4458 GNDA_2.n4457 0.1255
R13671 GNDA_2.n4293 GNDA_2.n4292 0.1255
R13672 GNDA_2.n4282 GNDA_2.n1107 0.1255
R13673 GNDA_2.n4275 GNDA_2.n4274 0.1255
R13674 GNDA_2.n4228 GNDA_2.n4199 0.1255
R13675 GNDA_2.n4241 GNDA_2.n4240 0.1255
R13676 GNDA_2.n4252 GNDA_2.n4187 0.1255
R13677 GNDA_2.n4119 GNDA_2.n4102 0.1255
R13678 GNDA_2.n4132 GNDA_2.n4131 0.1255
R13679 GNDA_2.n4143 GNDA_2.n4090 0.1255
R13680 GNDA_2.n4038 GNDA_2.n1150 0.1255
R13681 GNDA_2.n4051 GNDA_2.n4050 0.1255
R13682 GNDA_2.n4062 GNDA_2.n1138 0.1255
R13683 GNDA_2.n1233 GNDA_2.n1232 0.1255
R13684 GNDA_2.n1222 GNDA_2.n1182 0.1255
R13685 GNDA_2.n1215 GNDA_2.n1214 0.1255
R13686 GNDA_2.n3645 GNDA_2.n3628 0.1255
R13687 GNDA_2.n3658 GNDA_2.n3657 0.1255
R13688 GNDA_2.n3669 GNDA_2.n3616 0.1255
R13689 GNDA_2.n3714 GNDA_2.n3697 0.1255
R13690 GNDA_2.n3727 GNDA_2.n3726 0.1255
R13691 GNDA_2.n3738 GNDA_2.n3685 0.1255
R13692 GNDA_2.n3783 GNDA_2.n3766 0.1255
R13693 GNDA_2.n3796 GNDA_2.n3795 0.1255
R13694 GNDA_2.n3807 GNDA_2.n3754 0.1255
R13695 GNDA_2.n3852 GNDA_2.n3835 0.1255
R13696 GNDA_2.n3865 GNDA_2.n3864 0.1255
R13697 GNDA_2.n3876 GNDA_2.n3823 0.1255
R13698 GNDA_2.n4013 GNDA_2.n4010 0.1255
R13699 GNDA_2.n3909 GNDA_2.n3898 0.1255
R13700 GNDA_2.n3926 GNDA_2.n3925 0.1255
R13701 GNDA_2.n3939 GNDA_2.n3892 0.1255
R13702 GNDA_2.n2821 GNDA_2.n2670 0.1255
R13703 GNDA_2.n2695 GNDA_2.n2694 0.1255
R13704 GNDA_2.n3069 GNDA_2.n2974 0.1255
R13705 GNDA_2.n3011 GNDA_2.n2994 0.1255
R13706 GNDA_2.n3027 GNDA_2.n2988 0.1255
R13707 GNDA_2.n3041 GNDA_2.n2982 0.1255
R13708 GNDA_2.n1600 GNDA_2.n1599 0.1255
R13709 GNDA_2.n1611 GNDA_2.n1581 0.1255
R13710 GNDA_2.n1630 GNDA_2.n1629 0.1255
R13711 GNDA_2.n1598 GNDA_2.n1584 0.1255
R13712 GNDA_2.n1615 GNDA_2.n1614 0.1255
R13713 GNDA_2.n1628 GNDA_2.n1578 0.1255
R13714 GNDA_2.n286 GNDA_2.n285 0.1255
R13715 GNDA_2.n275 GNDA_2.n235 0.1255
R13716 GNDA_2.n268 GNDA_2.n267 0.1255
R13717 GNDA_2.n5225 GNDA_2.n5220 0.1255
R13718 GNDA_2.n662 GNDA_2.n644 0.1255
R13719 GNDA_2.n675 GNDA_2.n674 0.1255
R13720 GNDA_2.n686 GNDA_2.n632 0.1255
R13721 GNDA_2.n978 GNDA_2.n458 0.1255
R13722 GNDA_2.n991 GNDA_2.n990 0.1255
R13723 GNDA_2.n1002 GNDA_2.n446 0.1255
R13724 GNDA_2.n541 GNDA_2.n540 0.1255
R13725 GNDA_2.n530 GNDA_2.n490 0.1255
R13726 GNDA_2.n523 GNDA_2.n522 0.1255
R13727 GNDA_2.n766 GNDA_2.n749 0.1255
R13728 GNDA_2.n779 GNDA_2.n778 0.1255
R13729 GNDA_2.n790 GNDA_2.n737 0.1255
R13730 GNDA_2.n835 GNDA_2.n818 0.1255
R13731 GNDA_2.n848 GNDA_2.n847 0.1255
R13732 GNDA_2.n859 GNDA_2.n806 0.1255
R13733 GNDA_2.n892 GNDA_2.n881 0.1255
R13734 GNDA_2.n909 GNDA_2.n908 0.1255
R13735 GNDA_2.n922 GNDA_2.n875 0.1255
R13736 GNDA_2.n344 GNDA_2.n343 0.123287
R13737 GNDA_2.n4374 GNDA_2.n4373 0.12293
R13738 GNDA_2.n5233 GNDA_2.n5231 0.115083
R13739 GNDA_2.n5235 GNDA_2.n5233 0.115083
R13740 GNDA_2.n5237 GNDA_2.n5235 0.115083
R13741 GNDA_2.n5239 GNDA_2.n5237 0.115083
R13742 GNDA_2.n4385 GNDA_2.n4384 0.115083
R13743 GNDA_2.n4384 GNDA_2.n4382 0.115083
R13744 GNDA_2.n3992 GNDA_2.n3990 0.115083
R13745 GNDA_2.n3990 GNDA_2.n3988 0.115083
R13746 GNDA_2.n3988 GNDA_2.n3986 0.115083
R13747 GNDA_2.n3986 GNDA_2.n3984 0.115083
R13748 GNDA_2.n3423 GNDA_2.n3422 0.115083
R13749 GNDA_2.n3422 GNDA_2.n3421 0.115083
R13750 GNDA_2.n3419 GNDA_2.n3418 0.115083
R13751 GNDA_2.n3418 GNDA_2.n3417 0.115083
R13752 GNDA_2.n3417 GNDA_2.n3416 0.115083
R13753 GNDA_2.n3416 GNDA_2.n3415 0.115083
R13754 GNDA_2.n3414 GNDA_2.n3413 0.115083
R13755 GNDA_2.n3413 GNDA_2.n3412 0.115083
R13756 GNDA_2.n3412 GNDA_2.n3411 0.115083
R13757 GNDA_2.n3409 GNDA_2.n3408 0.115083
R13758 GNDA_2.n3408 GNDA_2.n3407 0.115083
R13759 GNDA_2.n3407 GNDA_2.n3406 0.115083
R13760 GNDA_2.n594 GNDA_2.n592 0.115083
R13761 GNDA_2.n592 GNDA_2.n590 0.115083
R13762 GNDA_2.n590 GNDA_2.n588 0.115083
R13763 GNDA_2.n588 GNDA_2.n586 0.115083
R13764 GNDA_2.n586 GNDA_2.n584 0.115083
R13765 GNDA_2.n584 GNDA_2.n582 0.115083
R13766 GNDA_2.n582 GNDA_2.n580 0.115083
R13767 GNDA_2.n580 GNDA_2.n578 0.115083
R13768 GNDA_2.n578 GNDA_2.n576 0.115083
R13769 GNDA_2.n576 GNDA_2.n574 0.115083
R13770 GNDA_2.n574 GNDA_2.n572 0.115083
R13771 GNDA_2.n4210 GNDA_2.n1091 0.10642
R13772 GNDA_2.n4474 GNDA_2.n4473 0.105167
R13773 GNDA_2.n362 GNDA_2.n361 0.0994583
R13774 GNDA_2.n4417 GNDA_2.n4415 0.0994583
R13775 GNDA_2.n4311 GNDA_2.n4310 0.09425
R13776 GNDA_2.n4622 GNDA_2.n4619 0.09425
R13777 GNDA_2.n4264 GNDA_2.n187 0.08275
R13778 GNDA_2.n3512 GNDA 0.0817953
R13779 GNDA_2.n1063 GNDA_2.n401 0.0734167
R13780 GNDA_2.n1063 GNDA_2.n1062 0.0734167
R13781 GNDA_2.n1062 GNDA_2.n1061 0.0734167
R13782 GNDA_2.n1056 GNDA_2.n1055 0.0734167
R13783 GNDA_2.n1055 GNDA_2.n411 0.0734167
R13784 GNDA_2.n1051 GNDA_2.n411 0.0734167
R13785 GNDA_2.n1045 GNDA_2.n416 0.0734167
R13786 GNDA_2.n1045 GNDA_2.n1044 0.0734167
R13787 GNDA_2.n1044 GNDA_2.n1043 0.0734167
R13788 GNDA_2.n1038 GNDA_2.n1037 0.0734167
R13789 GNDA_2.n1037 GNDA_2.n426 0.0734167
R13790 GNDA_2.n5011 GNDA_2.n4903 0.0734167
R13791 GNDA_2.n5012 GNDA_2.n5011 0.0734167
R13792 GNDA_2.n5012 GNDA_2.n5009 0.0734167
R13793 GNDA_2.n5022 GNDA_2.n5007 0.0734167
R13794 GNDA_2.n5030 GNDA_2.n5007 0.0734167
R13795 GNDA_2.n5031 GNDA_2.n5030 0.0734167
R13796 GNDA_2.n5041 GNDA_2.n5040 0.0734167
R13797 GNDA_2.n5042 GNDA_2.n5041 0.0734167
R13798 GNDA_2.n5042 GNDA_2.n5003 0.0734167
R13799 GNDA_2.n5052 GNDA_2.n5001 0.0734167
R13800 GNDA_2.n5060 GNDA_2.n5001 0.0734167
R13801 GNDA_2.n4935 GNDA_2.n4934 0.0734167
R13802 GNDA_2.n4936 GNDA_2.n4935 0.0734167
R13803 GNDA_2.n4936 GNDA_2.n4928 0.0734167
R13804 GNDA_2.n4946 GNDA_2.n4926 0.0734167
R13805 GNDA_2.n4954 GNDA_2.n4926 0.0734167
R13806 GNDA_2.n4955 GNDA_2.n4954 0.0734167
R13807 GNDA_2.n4965 GNDA_2.n4964 0.0734167
R13808 GNDA_2.n4966 GNDA_2.n4965 0.0734167
R13809 GNDA_2.n4966 GNDA_2.n4922 0.0734167
R13810 GNDA_2.n4976 GNDA_2.n4920 0.0734167
R13811 GNDA_2.n4984 GNDA_2.n4920 0.0734167
R13812 GNDA_2.n4835 GNDA_2.n4812 0.0734167
R13813 GNDA_2.n4836 GNDA_2.n4835 0.0734167
R13814 GNDA_2.n4837 GNDA_2.n4836 0.0734167
R13815 GNDA_2.n4841 GNDA_2.n4840 0.0734167
R13816 GNDA_2.n4842 GNDA_2.n4841 0.0734167
R13817 GNDA_2.n4843 GNDA_2.n4842 0.0734167
R13818 GNDA_2.n4847 GNDA_2.n4846 0.0734167
R13819 GNDA_2.n4848 GNDA_2.n4847 0.0734167
R13820 GNDA_2.n4849 GNDA_2.n4848 0.0734167
R13821 GNDA_2.n4853 GNDA_2.n4852 0.0734167
R13822 GNDA_2.n4854 GNDA_2.n4853 0.0734167
R13823 GNDA_2.n5095 GNDA_2.n5094 0.0734167
R13824 GNDA_2.n5096 GNDA_2.n5095 0.0734167
R13825 GNDA_2.n5096 GNDA_2.n4807 0.0734167
R13826 GNDA_2.n5106 GNDA_2.n4805 0.0734167
R13827 GNDA_2.n5114 GNDA_2.n4805 0.0734167
R13828 GNDA_2.n5115 GNDA_2.n5114 0.0734167
R13829 GNDA_2.n5125 GNDA_2.n5124 0.0734167
R13830 GNDA_2.n5126 GNDA_2.n5125 0.0734167
R13831 GNDA_2.n5126 GNDA_2.n4801 0.0734167
R13832 GNDA_2.n5136 GNDA_2.n4799 0.0734167
R13833 GNDA_2.n5144 GNDA_2.n4799 0.0734167
R13834 GNDA_2.n4559 GNDA_2.n184 0.0734167
R13835 GNDA_2.n4560 GNDA_2.n4559 0.0734167
R13836 GNDA_2.n4560 GNDA_2.n4557 0.0734167
R13837 GNDA_2.n4570 GNDA_2.n4555 0.0734167
R13838 GNDA_2.n4578 GNDA_2.n4555 0.0734167
R13839 GNDA_2.n4579 GNDA_2.n4578 0.0734167
R13840 GNDA_2.n4589 GNDA_2.n4588 0.0734167
R13841 GNDA_2.n4590 GNDA_2.n4589 0.0734167
R13842 GNDA_2.n4590 GNDA_2.n4551 0.0734167
R13843 GNDA_2.n4600 GNDA_2.n4549 0.0734167
R13844 GNDA_2.n4608 GNDA_2.n4549 0.0734167
R13845 GNDA_2.n5160 GNDA_2.n144 0.0734167
R13846 GNDA_2.n5161 GNDA_2.n5160 0.0734167
R13847 GNDA_2.n5161 GNDA_2.n5158 0.0734167
R13848 GNDA_2.n5171 GNDA_2.n5156 0.0734167
R13849 GNDA_2.n5179 GNDA_2.n5156 0.0734167
R13850 GNDA_2.n5180 GNDA_2.n5179 0.0734167
R13851 GNDA_2.n5190 GNDA_2.n5189 0.0734167
R13852 GNDA_2.n5191 GNDA_2.n5190 0.0734167
R13853 GNDA_2.n5191 GNDA_2.n5152 0.0734167
R13854 GNDA_2.n5201 GNDA_2.n5150 0.0734167
R13855 GNDA_2.n5209 GNDA_2.n5150 0.0734167
R13856 GNDA_2.n4720 GNDA_2.n4719 0.0734167
R13857 GNDA_2.n4721 GNDA_2.n4720 0.0734167
R13858 GNDA_2.n4721 GNDA_2.n170 0.0734167
R13859 GNDA_2.n4731 GNDA_2.n168 0.0734167
R13860 GNDA_2.n4739 GNDA_2.n168 0.0734167
R13861 GNDA_2.n4740 GNDA_2.n4739 0.0734167
R13862 GNDA_2.n4750 GNDA_2.n4749 0.0734167
R13863 GNDA_2.n4751 GNDA_2.n4750 0.0734167
R13864 GNDA_2.n4751 GNDA_2.n164 0.0734167
R13865 GNDA_2.n4761 GNDA_2.n162 0.0734167
R13866 GNDA_2.n4769 GNDA_2.n162 0.0734167
R13867 GNDA_2.n4647 GNDA_2.n4624 0.0734167
R13868 GNDA_2.n4648 GNDA_2.n4647 0.0734167
R13869 GNDA_2.n4649 GNDA_2.n4648 0.0734167
R13870 GNDA_2.n4653 GNDA_2.n4652 0.0734167
R13871 GNDA_2.n4654 GNDA_2.n4653 0.0734167
R13872 GNDA_2.n4655 GNDA_2.n4654 0.0734167
R13873 GNDA_2.n4659 GNDA_2.n4658 0.0734167
R13874 GNDA_2.n4660 GNDA_2.n4659 0.0734167
R13875 GNDA_2.n4661 GNDA_2.n4660 0.0734167
R13876 GNDA_2.n4665 GNDA_2.n4664 0.0734167
R13877 GNDA_2.n4666 GNDA_2.n4665 0.0734167
R13878 GNDA_2.n4483 GNDA_2.n4482 0.0734167
R13879 GNDA_2.n4484 GNDA_2.n4483 0.0734167
R13880 GNDA_2.n4484 GNDA_2.n210 0.0734167
R13881 GNDA_2.n4494 GNDA_2.n208 0.0734167
R13882 GNDA_2.n4502 GNDA_2.n208 0.0734167
R13883 GNDA_2.n4503 GNDA_2.n4502 0.0734167
R13884 GNDA_2.n4513 GNDA_2.n4512 0.0734167
R13885 GNDA_2.n4514 GNDA_2.n4513 0.0734167
R13886 GNDA_2.n4514 GNDA_2.n204 0.0734167
R13887 GNDA_2.n4524 GNDA_2.n202 0.0734167
R13888 GNDA_2.n4532 GNDA_2.n202 0.0734167
R13889 GNDA_2.n4297 GNDA_2.n1093 0.0734167
R13890 GNDA_2.n4297 GNDA_2.n4296 0.0734167
R13891 GNDA_2.n4296 GNDA_2.n4295 0.0734167
R13892 GNDA_2.n4290 GNDA_2.n4289 0.0734167
R13893 GNDA_2.n4289 GNDA_2.n1103 0.0734167
R13894 GNDA_2.n4285 GNDA_2.n1103 0.0734167
R13895 GNDA_2.n4279 GNDA_2.n1108 0.0734167
R13896 GNDA_2.n4279 GNDA_2.n4278 0.0734167
R13897 GNDA_2.n4278 GNDA_2.n4277 0.0734167
R13898 GNDA_2.n4272 GNDA_2.n4271 0.0734167
R13899 GNDA_2.n4271 GNDA_2.n1118 0.0734167
R13900 GNDA_2.n4222 GNDA_2.n4221 0.0734167
R13901 GNDA_2.n4223 GNDA_2.n4222 0.0734167
R13902 GNDA_2.n4223 GNDA_2.n4202 0.0734167
R13903 GNDA_2.n4231 GNDA_2.n4198 0.0734167
R13904 GNDA_2.n4237 GNDA_2.n4198 0.0734167
R13905 GNDA_2.n4238 GNDA_2.n4237 0.0734167
R13906 GNDA_2.n4246 GNDA_2.n4245 0.0734167
R13907 GNDA_2.n4247 GNDA_2.n4246 0.0734167
R13908 GNDA_2.n4247 GNDA_2.n4190 0.0734167
R13909 GNDA_2.n4255 GNDA_2.n4186 0.0734167
R13910 GNDA_2.n4261 GNDA_2.n4186 0.0734167
R13911 GNDA_2.n4113 GNDA_2.n4112 0.0734167
R13912 GNDA_2.n4114 GNDA_2.n4113 0.0734167
R13913 GNDA_2.n4114 GNDA_2.n4105 0.0734167
R13914 GNDA_2.n4122 GNDA_2.n4101 0.0734167
R13915 GNDA_2.n4128 GNDA_2.n4101 0.0734167
R13916 GNDA_2.n4129 GNDA_2.n4128 0.0734167
R13917 GNDA_2.n4137 GNDA_2.n4136 0.0734167
R13918 GNDA_2.n4138 GNDA_2.n4137 0.0734167
R13919 GNDA_2.n4138 GNDA_2.n4093 0.0734167
R13920 GNDA_2.n4146 GNDA_2.n4089 0.0734167
R13921 GNDA_2.n4152 GNDA_2.n4089 0.0734167
R13922 GNDA_2.n4032 GNDA_2.n4031 0.0734167
R13923 GNDA_2.n4033 GNDA_2.n4032 0.0734167
R13924 GNDA_2.n4033 GNDA_2.n1153 0.0734167
R13925 GNDA_2.n4041 GNDA_2.n1149 0.0734167
R13926 GNDA_2.n4047 GNDA_2.n1149 0.0734167
R13927 GNDA_2.n4048 GNDA_2.n4047 0.0734167
R13928 GNDA_2.n4056 GNDA_2.n4055 0.0734167
R13929 GNDA_2.n4057 GNDA_2.n4056 0.0734167
R13930 GNDA_2.n4057 GNDA_2.n1141 0.0734167
R13931 GNDA_2.n4065 GNDA_2.n1137 0.0734167
R13932 GNDA_2.n4071 GNDA_2.n1137 0.0734167
R13933 GNDA_2.n1237 GNDA_2.n1161 0.0734167
R13934 GNDA_2.n1237 GNDA_2.n1236 0.0734167
R13935 GNDA_2.n1236 GNDA_2.n1235 0.0734167
R13936 GNDA_2.n1230 GNDA_2.n1229 0.0734167
R13937 GNDA_2.n1229 GNDA_2.n1175 0.0734167
R13938 GNDA_2.n1225 GNDA_2.n1175 0.0734167
R13939 GNDA_2.n1219 GNDA_2.n1183 0.0734167
R13940 GNDA_2.n1219 GNDA_2.n1218 0.0734167
R13941 GNDA_2.n1218 GNDA_2.n1217 0.0734167
R13942 GNDA_2.n1212 GNDA_2.n1211 0.0734167
R13943 GNDA_2.n1211 GNDA_2.n1199 0.0734167
R13944 GNDA_2.n3639 GNDA_2.n3638 0.0734167
R13945 GNDA_2.n3640 GNDA_2.n3639 0.0734167
R13946 GNDA_2.n3640 GNDA_2.n3631 0.0734167
R13947 GNDA_2.n3648 GNDA_2.n3627 0.0734167
R13948 GNDA_2.n3654 GNDA_2.n3627 0.0734167
R13949 GNDA_2.n3655 GNDA_2.n3654 0.0734167
R13950 GNDA_2.n3663 GNDA_2.n3662 0.0734167
R13951 GNDA_2.n3664 GNDA_2.n3663 0.0734167
R13952 GNDA_2.n3664 GNDA_2.n3619 0.0734167
R13953 GNDA_2.n3672 GNDA_2.n3615 0.0734167
R13954 GNDA_2.n3678 GNDA_2.n3615 0.0734167
R13955 GNDA_2.n3708 GNDA_2.n3707 0.0734167
R13956 GNDA_2.n3709 GNDA_2.n3708 0.0734167
R13957 GNDA_2.n3709 GNDA_2.n3700 0.0734167
R13958 GNDA_2.n3717 GNDA_2.n3696 0.0734167
R13959 GNDA_2.n3723 GNDA_2.n3696 0.0734167
R13960 GNDA_2.n3724 GNDA_2.n3723 0.0734167
R13961 GNDA_2.n3732 GNDA_2.n3731 0.0734167
R13962 GNDA_2.n3733 GNDA_2.n3732 0.0734167
R13963 GNDA_2.n3733 GNDA_2.n3688 0.0734167
R13964 GNDA_2.n3741 GNDA_2.n3684 0.0734167
R13965 GNDA_2.n3747 GNDA_2.n3684 0.0734167
R13966 GNDA_2.n3777 GNDA_2.n3776 0.0734167
R13967 GNDA_2.n3778 GNDA_2.n3777 0.0734167
R13968 GNDA_2.n3778 GNDA_2.n3769 0.0734167
R13969 GNDA_2.n3786 GNDA_2.n3765 0.0734167
R13970 GNDA_2.n3792 GNDA_2.n3765 0.0734167
R13971 GNDA_2.n3793 GNDA_2.n3792 0.0734167
R13972 GNDA_2.n3801 GNDA_2.n3800 0.0734167
R13973 GNDA_2.n3802 GNDA_2.n3801 0.0734167
R13974 GNDA_2.n3802 GNDA_2.n3757 0.0734167
R13975 GNDA_2.n3810 GNDA_2.n3753 0.0734167
R13976 GNDA_2.n3816 GNDA_2.n3753 0.0734167
R13977 GNDA_2.n3846 GNDA_2.n3845 0.0734167
R13978 GNDA_2.n3847 GNDA_2.n3846 0.0734167
R13979 GNDA_2.n3847 GNDA_2.n3838 0.0734167
R13980 GNDA_2.n3855 GNDA_2.n3834 0.0734167
R13981 GNDA_2.n3861 GNDA_2.n3834 0.0734167
R13982 GNDA_2.n3862 GNDA_2.n3861 0.0734167
R13983 GNDA_2.n3870 GNDA_2.n3869 0.0734167
R13984 GNDA_2.n3871 GNDA_2.n3870 0.0734167
R13985 GNDA_2.n3871 GNDA_2.n3826 0.0734167
R13986 GNDA_2.n3879 GNDA_2.n3822 0.0734167
R13987 GNDA_2.n3885 GNDA_2.n3822 0.0734167
R13988 GNDA_2.n4008 GNDA_2.n3976 0.0734167
R13989 GNDA_2.n3901 GNDA_2.n1264 0.0734167
R13990 GNDA_2.n3902 GNDA_2.n3901 0.0734167
R13991 GNDA_2.n3902 GNDA_2.n3899 0.0734167
R13992 GNDA_2.n3912 GNDA_2.n3897 0.0734167
R13993 GNDA_2.n3920 GNDA_2.n3897 0.0734167
R13994 GNDA_2.n3921 GNDA_2.n3920 0.0734167
R13995 GNDA_2.n3931 GNDA_2.n3930 0.0734167
R13996 GNDA_2.n3932 GNDA_2.n3931 0.0734167
R13997 GNDA_2.n3932 GNDA_2.n3893 0.0734167
R13998 GNDA_2.n3942 GNDA_2.n3891 0.0734167
R13999 GNDA_2.n3950 GNDA_2.n3891 0.0734167
R14000 GNDA_2.n3008 GNDA_2.n2997 0.0734167
R14001 GNDA_2.n3009 GNDA_2.n3008 0.0734167
R14002 GNDA_2.n3019 GNDA_2.n3018 0.0734167
R14003 GNDA_2.n3020 GNDA_2.n3019 0.0734167
R14004 GNDA_2.n3020 GNDA_2.n2989 0.0734167
R14005 GNDA_2.n3030 GNDA_2.n2985 0.0734167
R14006 GNDA_2.n3038 GNDA_2.n2985 0.0734167
R14007 GNDA_2.n3039 GNDA_2.n3038 0.0734167
R14008 GNDA_2.n3049 GNDA_2.n3048 0.0734167
R14009 GNDA_2.n3050 GNDA_2.n3049 0.0734167
R14010 GNDA_2.n3050 GNDA_2.n2977 0.0734167
R14011 GNDA_2.n290 GNDA_2.n215 0.0734167
R14012 GNDA_2.n290 GNDA_2.n289 0.0734167
R14013 GNDA_2.n289 GNDA_2.n288 0.0734167
R14014 GNDA_2.n283 GNDA_2.n282 0.0734167
R14015 GNDA_2.n282 GNDA_2.n228 0.0734167
R14016 GNDA_2.n278 GNDA_2.n228 0.0734167
R14017 GNDA_2.n272 GNDA_2.n236 0.0734167
R14018 GNDA_2.n272 GNDA_2.n271 0.0734167
R14019 GNDA_2.n271 GNDA_2.n270 0.0734167
R14020 GNDA_2.n265 GNDA_2.n264 0.0734167
R14021 GNDA_2.n264 GNDA_2.n252 0.0734167
R14022 GNDA_2.n5086 GNDA_2.n138 0.0734167
R14023 GNDA_2.n656 GNDA_2.n655 0.0734167
R14024 GNDA_2.n657 GNDA_2.n656 0.0734167
R14025 GNDA_2.n657 GNDA_2.n647 0.0734167
R14026 GNDA_2.n665 GNDA_2.n643 0.0734167
R14027 GNDA_2.n671 GNDA_2.n643 0.0734167
R14028 GNDA_2.n672 GNDA_2.n671 0.0734167
R14029 GNDA_2.n680 GNDA_2.n679 0.0734167
R14030 GNDA_2.n681 GNDA_2.n680 0.0734167
R14031 GNDA_2.n681 GNDA_2.n635 0.0734167
R14032 GNDA_2.n689 GNDA_2.n631 0.0734167
R14033 GNDA_2.n695 GNDA_2.n631 0.0734167
R14034 GNDA_2.n972 GNDA_2.n971 0.0734167
R14035 GNDA_2.n973 GNDA_2.n972 0.0734167
R14036 GNDA_2.n973 GNDA_2.n461 0.0734167
R14037 GNDA_2.n981 GNDA_2.n457 0.0734167
R14038 GNDA_2.n987 GNDA_2.n457 0.0734167
R14039 GNDA_2.n988 GNDA_2.n987 0.0734167
R14040 GNDA_2.n996 GNDA_2.n995 0.0734167
R14041 GNDA_2.n997 GNDA_2.n996 0.0734167
R14042 GNDA_2.n997 GNDA_2.n449 0.0734167
R14043 GNDA_2.n1005 GNDA_2.n445 0.0734167
R14044 GNDA_2.n1011 GNDA_2.n445 0.0734167
R14045 GNDA_2.n545 GNDA_2.n469 0.0734167
R14046 GNDA_2.n545 GNDA_2.n544 0.0734167
R14047 GNDA_2.n544 GNDA_2.n543 0.0734167
R14048 GNDA_2.n538 GNDA_2.n537 0.0734167
R14049 GNDA_2.n537 GNDA_2.n483 0.0734167
R14050 GNDA_2.n533 GNDA_2.n483 0.0734167
R14051 GNDA_2.n527 GNDA_2.n491 0.0734167
R14052 GNDA_2.n527 GNDA_2.n526 0.0734167
R14053 GNDA_2.n526 GNDA_2.n525 0.0734167
R14054 GNDA_2.n520 GNDA_2.n519 0.0734167
R14055 GNDA_2.n519 GNDA_2.n507 0.0734167
R14056 GNDA_2.n760 GNDA_2.n759 0.0734167
R14057 GNDA_2.n761 GNDA_2.n760 0.0734167
R14058 GNDA_2.n761 GNDA_2.n752 0.0734167
R14059 GNDA_2.n769 GNDA_2.n748 0.0734167
R14060 GNDA_2.n775 GNDA_2.n748 0.0734167
R14061 GNDA_2.n776 GNDA_2.n775 0.0734167
R14062 GNDA_2.n784 GNDA_2.n783 0.0734167
R14063 GNDA_2.n785 GNDA_2.n784 0.0734167
R14064 GNDA_2.n785 GNDA_2.n740 0.0734167
R14065 GNDA_2.n793 GNDA_2.n736 0.0734167
R14066 GNDA_2.n799 GNDA_2.n736 0.0734167
R14067 GNDA_2.n829 GNDA_2.n828 0.0734167
R14068 GNDA_2.n830 GNDA_2.n829 0.0734167
R14069 GNDA_2.n830 GNDA_2.n821 0.0734167
R14070 GNDA_2.n838 GNDA_2.n817 0.0734167
R14071 GNDA_2.n844 GNDA_2.n817 0.0734167
R14072 GNDA_2.n845 GNDA_2.n844 0.0734167
R14073 GNDA_2.n853 GNDA_2.n852 0.0734167
R14074 GNDA_2.n854 GNDA_2.n853 0.0734167
R14075 GNDA_2.n854 GNDA_2.n809 0.0734167
R14076 GNDA_2.n862 GNDA_2.n805 0.0734167
R14077 GNDA_2.n868 GNDA_2.n805 0.0734167
R14078 GNDA_2.n884 GNDA_2.n614 0.0734167
R14079 GNDA_2.n885 GNDA_2.n884 0.0734167
R14080 GNDA_2.n885 GNDA_2.n882 0.0734167
R14081 GNDA_2.n895 GNDA_2.n880 0.0734167
R14082 GNDA_2.n903 GNDA_2.n880 0.0734167
R14083 GNDA_2.n904 GNDA_2.n903 0.0734167
R14084 GNDA_2.n914 GNDA_2.n913 0.0734167
R14085 GNDA_2.n915 GNDA_2.n914 0.0734167
R14086 GNDA_2.n915 GNDA_2.n876 0.0734167
R14087 GNDA_2.n925 GNDA_2.n874 0.0734167
R14088 GNDA_2.n933 GNDA_2.n874 0.0734167
R14089 GNDA_2.n1067 GNDA_2.n401 0.0682083
R14090 GNDA_2.n1061 GNDA_2.n406 0.0682083
R14091 GNDA_2.n1057 GNDA_2.n1056 0.0682083
R14092 GNDA_2.n1051 GNDA_2.n1050 0.0682083
R14093 GNDA_2.n1049 GNDA_2.n416 0.0682083
R14094 GNDA_2.n1043 GNDA_2.n421 0.0682083
R14095 GNDA_2.n1039 GNDA_2.n1038 0.0682083
R14096 GNDA_2.n5066 GNDA_2.n4903 0.0682083
R14097 GNDA_2.n5020 GNDA_2.n5009 0.0682083
R14098 GNDA_2.n5022 GNDA_2.n5021 0.0682083
R14099 GNDA_2.n5032 GNDA_2.n5031 0.0682083
R14100 GNDA_2.n5040 GNDA_2.n5005 0.0682083
R14101 GNDA_2.n5050 GNDA_2.n5003 0.0682083
R14102 GNDA_2.n5052 GNDA_2.n5051 0.0682083
R14103 GNDA_2.n4934 GNDA_2.n4930 0.0682083
R14104 GNDA_2.n4944 GNDA_2.n4928 0.0682083
R14105 GNDA_2.n4946 GNDA_2.n4945 0.0682083
R14106 GNDA_2.n4956 GNDA_2.n4955 0.0682083
R14107 GNDA_2.n4964 GNDA_2.n4924 0.0682083
R14108 GNDA_2.n4974 GNDA_2.n4922 0.0682083
R14109 GNDA_2.n4976 GNDA_2.n4975 0.0682083
R14110 GNDA_2.n4892 GNDA_2.n4812 0.0682083
R14111 GNDA_2.n4838 GNDA_2.n4837 0.0682083
R14112 GNDA_2.n4840 GNDA_2.n4839 0.0682083
R14113 GNDA_2.n4844 GNDA_2.n4843 0.0682083
R14114 GNDA_2.n4846 GNDA_2.n4845 0.0682083
R14115 GNDA_2.n4850 GNDA_2.n4849 0.0682083
R14116 GNDA_2.n4852 GNDA_2.n4851 0.0682083
R14117 GNDA_2.n5094 GNDA_2.n5090 0.0682083
R14118 GNDA_2.n5104 GNDA_2.n4807 0.0682083
R14119 GNDA_2.n5106 GNDA_2.n5105 0.0682083
R14120 GNDA_2.n5116 GNDA_2.n5115 0.0682083
R14121 GNDA_2.n5124 GNDA_2.n4803 0.0682083
R14122 GNDA_2.n5134 GNDA_2.n4801 0.0682083
R14123 GNDA_2.n5136 GNDA_2.n5135 0.0682083
R14124 GNDA_2.n4614 GNDA_2.n184 0.0682083
R14125 GNDA_2.n4568 GNDA_2.n4557 0.0682083
R14126 GNDA_2.n4570 GNDA_2.n4569 0.0682083
R14127 GNDA_2.n4580 GNDA_2.n4579 0.0682083
R14128 GNDA_2.n4588 GNDA_2.n4553 0.0682083
R14129 GNDA_2.n4598 GNDA_2.n4551 0.0682083
R14130 GNDA_2.n4600 GNDA_2.n4599 0.0682083
R14131 GNDA_2.n5215 GNDA_2.n144 0.0682083
R14132 GNDA_2.n5169 GNDA_2.n5158 0.0682083
R14133 GNDA_2.n5171 GNDA_2.n5170 0.0682083
R14134 GNDA_2.n5181 GNDA_2.n5180 0.0682083
R14135 GNDA_2.n5189 GNDA_2.n5154 0.0682083
R14136 GNDA_2.n5199 GNDA_2.n5152 0.0682083
R14137 GNDA_2.n5201 GNDA_2.n5200 0.0682083
R14138 GNDA_2.n4719 GNDA_2.n4715 0.0682083
R14139 GNDA_2.n4729 GNDA_2.n170 0.0682083
R14140 GNDA_2.n4731 GNDA_2.n4730 0.0682083
R14141 GNDA_2.n4741 GNDA_2.n4740 0.0682083
R14142 GNDA_2.n4749 GNDA_2.n166 0.0682083
R14143 GNDA_2.n4759 GNDA_2.n164 0.0682083
R14144 GNDA_2.n4761 GNDA_2.n4760 0.0682083
R14145 GNDA_2.n4704 GNDA_2.n4624 0.0682083
R14146 GNDA_2.n4650 GNDA_2.n4649 0.0682083
R14147 GNDA_2.n4652 GNDA_2.n4651 0.0682083
R14148 GNDA_2.n4656 GNDA_2.n4655 0.0682083
R14149 GNDA_2.n4658 GNDA_2.n4657 0.0682083
R14150 GNDA_2.n4662 GNDA_2.n4661 0.0682083
R14151 GNDA_2.n4664 GNDA_2.n4663 0.0682083
R14152 GNDA_2.n4482 GNDA_2.n4478 0.0682083
R14153 GNDA_2.n4492 GNDA_2.n210 0.0682083
R14154 GNDA_2.n4494 GNDA_2.n4493 0.0682083
R14155 GNDA_2.n4504 GNDA_2.n4503 0.0682083
R14156 GNDA_2.n4512 GNDA_2.n206 0.0682083
R14157 GNDA_2.n4522 GNDA_2.n204 0.0682083
R14158 GNDA_2.n4524 GNDA_2.n4523 0.0682083
R14159 GNDA_2.n4301 GNDA_2.n1093 0.0682083
R14160 GNDA_2.n4295 GNDA_2.n1098 0.0682083
R14161 GNDA_2.n4291 GNDA_2.n4290 0.0682083
R14162 GNDA_2.n4285 GNDA_2.n4284 0.0682083
R14163 GNDA_2.n4283 GNDA_2.n1108 0.0682083
R14164 GNDA_2.n4277 GNDA_2.n1113 0.0682083
R14165 GNDA_2.n4273 GNDA_2.n4272 0.0682083
R14166 GNDA_2.n4221 GNDA_2.n4217 0.0682083
R14167 GNDA_2.n4229 GNDA_2.n4202 0.0682083
R14168 GNDA_2.n4231 GNDA_2.n4230 0.0682083
R14169 GNDA_2.n4239 GNDA_2.n4238 0.0682083
R14170 GNDA_2.n4245 GNDA_2.n4194 0.0682083
R14171 GNDA_2.n4253 GNDA_2.n4190 0.0682083
R14172 GNDA_2.n4255 GNDA_2.n4254 0.0682083
R14173 GNDA_2.n4112 GNDA_2.n1089 0.0682083
R14174 GNDA_2.n4120 GNDA_2.n4105 0.0682083
R14175 GNDA_2.n4122 GNDA_2.n4121 0.0682083
R14176 GNDA_2.n4130 GNDA_2.n4129 0.0682083
R14177 GNDA_2.n4136 GNDA_2.n4097 0.0682083
R14178 GNDA_2.n4144 GNDA_2.n4093 0.0682083
R14179 GNDA_2.n4146 GNDA_2.n4145 0.0682083
R14180 GNDA_2.n4031 GNDA_2.n4027 0.0682083
R14181 GNDA_2.n4039 GNDA_2.n1153 0.0682083
R14182 GNDA_2.n4041 GNDA_2.n4040 0.0682083
R14183 GNDA_2.n4049 GNDA_2.n4048 0.0682083
R14184 GNDA_2.n4055 GNDA_2.n1145 0.0682083
R14185 GNDA_2.n4063 GNDA_2.n1141 0.0682083
R14186 GNDA_2.n4065 GNDA_2.n4064 0.0682083
R14187 GNDA_2.n1241 GNDA_2.n1161 0.0682083
R14188 GNDA_2.n1235 GNDA_2.n1167 0.0682083
R14189 GNDA_2.n1231 GNDA_2.n1230 0.0682083
R14190 GNDA_2.n1225 GNDA_2.n1224 0.0682083
R14191 GNDA_2.n1223 GNDA_2.n1183 0.0682083
R14192 GNDA_2.n1217 GNDA_2.n1191 0.0682083
R14193 GNDA_2.n1213 GNDA_2.n1212 0.0682083
R14194 GNDA_2.n3638 GNDA_2.n1245 0.0682083
R14195 GNDA_2.n3646 GNDA_2.n3631 0.0682083
R14196 GNDA_2.n3648 GNDA_2.n3647 0.0682083
R14197 GNDA_2.n3656 GNDA_2.n3655 0.0682083
R14198 GNDA_2.n3662 GNDA_2.n3623 0.0682083
R14199 GNDA_2.n3670 GNDA_2.n3619 0.0682083
R14200 GNDA_2.n3672 GNDA_2.n3671 0.0682083
R14201 GNDA_2.n3707 GNDA_2.n1252 0.0682083
R14202 GNDA_2.n3715 GNDA_2.n3700 0.0682083
R14203 GNDA_2.n3717 GNDA_2.n3716 0.0682083
R14204 GNDA_2.n3725 GNDA_2.n3724 0.0682083
R14205 GNDA_2.n3731 GNDA_2.n3692 0.0682083
R14206 GNDA_2.n3739 GNDA_2.n3688 0.0682083
R14207 GNDA_2.n3741 GNDA_2.n3740 0.0682083
R14208 GNDA_2.n3776 GNDA_2.n1256 0.0682083
R14209 GNDA_2.n3784 GNDA_2.n3769 0.0682083
R14210 GNDA_2.n3786 GNDA_2.n3785 0.0682083
R14211 GNDA_2.n3794 GNDA_2.n3793 0.0682083
R14212 GNDA_2.n3800 GNDA_2.n3761 0.0682083
R14213 GNDA_2.n3808 GNDA_2.n3757 0.0682083
R14214 GNDA_2.n3810 GNDA_2.n3809 0.0682083
R14215 GNDA_2.n3845 GNDA_2.n1260 0.0682083
R14216 GNDA_2.n3853 GNDA_2.n3838 0.0682083
R14217 GNDA_2.n3855 GNDA_2.n3854 0.0682083
R14218 GNDA_2.n3863 GNDA_2.n3862 0.0682083
R14219 GNDA_2.n3869 GNDA_2.n3830 0.0682083
R14220 GNDA_2.n3877 GNDA_2.n3826 0.0682083
R14221 GNDA_2.n3879 GNDA_2.n3878 0.0682083
R14222 GNDA_2.n3956 GNDA_2.n1264 0.0682083
R14223 GNDA_2.n3910 GNDA_2.n3899 0.0682083
R14224 GNDA_2.n3912 GNDA_2.n3911 0.0682083
R14225 GNDA_2.n3922 GNDA_2.n3921 0.0682083
R14226 GNDA_2.n3930 GNDA_2.n3895 0.0682083
R14227 GNDA_2.n3940 GNDA_2.n3893 0.0682083
R14228 GNDA_2.n3942 GNDA_2.n3941 0.0682083
R14229 GNDA_2.n3010 GNDA_2.n3009 0.0682083
R14230 GNDA_2.n3018 GNDA_2.n2993 0.0682083
R14231 GNDA_2.n3028 GNDA_2.n2989 0.0682083
R14232 GNDA_2.n3030 GNDA_2.n3029 0.0682083
R14233 GNDA_2.n3040 GNDA_2.n3039 0.0682083
R14234 GNDA_2.n3048 GNDA_2.n2981 0.0682083
R14235 GNDA_2.n3057 GNDA_2.n2977 0.0682083
R14236 GNDA_2.n294 GNDA_2.n215 0.0682083
R14237 GNDA_2.n288 GNDA_2.n220 0.0682083
R14238 GNDA_2.n284 GNDA_2.n283 0.0682083
R14239 GNDA_2.n278 GNDA_2.n277 0.0682083
R14240 GNDA_2.n276 GNDA_2.n236 0.0682083
R14241 GNDA_2.n270 GNDA_2.n244 0.0682083
R14242 GNDA_2.n266 GNDA_2.n265 0.0682083
R14243 GNDA_2.n655 GNDA_2.n651 0.0682083
R14244 GNDA_2.n663 GNDA_2.n647 0.0682083
R14245 GNDA_2.n665 GNDA_2.n664 0.0682083
R14246 GNDA_2.n673 GNDA_2.n672 0.0682083
R14247 GNDA_2.n679 GNDA_2.n639 0.0682083
R14248 GNDA_2.n687 GNDA_2.n635 0.0682083
R14249 GNDA_2.n689 GNDA_2.n688 0.0682083
R14250 GNDA_2.n971 GNDA_2.n967 0.0682083
R14251 GNDA_2.n979 GNDA_2.n461 0.0682083
R14252 GNDA_2.n981 GNDA_2.n980 0.0682083
R14253 GNDA_2.n989 GNDA_2.n988 0.0682083
R14254 GNDA_2.n995 GNDA_2.n453 0.0682083
R14255 GNDA_2.n1003 GNDA_2.n449 0.0682083
R14256 GNDA_2.n1005 GNDA_2.n1004 0.0682083
R14257 GNDA_2.n549 GNDA_2.n469 0.0682083
R14258 GNDA_2.n543 GNDA_2.n475 0.0682083
R14259 GNDA_2.n539 GNDA_2.n538 0.0682083
R14260 GNDA_2.n533 GNDA_2.n532 0.0682083
R14261 GNDA_2.n531 GNDA_2.n491 0.0682083
R14262 GNDA_2.n525 GNDA_2.n499 0.0682083
R14263 GNDA_2.n521 GNDA_2.n520 0.0682083
R14264 GNDA_2.n759 GNDA_2.n553 0.0682083
R14265 GNDA_2.n767 GNDA_2.n752 0.0682083
R14266 GNDA_2.n769 GNDA_2.n768 0.0682083
R14267 GNDA_2.n777 GNDA_2.n776 0.0682083
R14268 GNDA_2.n783 GNDA_2.n744 0.0682083
R14269 GNDA_2.n791 GNDA_2.n740 0.0682083
R14270 GNDA_2.n793 GNDA_2.n792 0.0682083
R14271 GNDA_2.n828 GNDA_2.n557 0.0682083
R14272 GNDA_2.n836 GNDA_2.n821 0.0682083
R14273 GNDA_2.n838 GNDA_2.n837 0.0682083
R14274 GNDA_2.n846 GNDA_2.n845 0.0682083
R14275 GNDA_2.n852 GNDA_2.n813 0.0682083
R14276 GNDA_2.n860 GNDA_2.n809 0.0682083
R14277 GNDA_2.n862 GNDA_2.n861 0.0682083
R14278 GNDA_2.n939 GNDA_2.n614 0.0682083
R14279 GNDA_2.n893 GNDA_2.n882 0.0682083
R14280 GNDA_2.n895 GNDA_2.n894 0.0682083
R14281 GNDA_2.n905 GNDA_2.n904 0.0682083
R14282 GNDA_2.n913 GNDA_2.n878 0.0682083
R14283 GNDA_2.n923 GNDA_2.n876 0.0682083
R14284 GNDA_2.n925 GNDA_2.n924 0.0682083
R14285 GNDA_2.n1034 GNDA_2.n1033 0.0672139
R14286 GNDA_2.n5061 GNDA_2.n5000 0.0672139
R14287 GNDA_2.n4985 GNDA_2.n4919 0.0672139
R14288 GNDA_2.n4855 GNDA_2.n4834 0.0672139
R14289 GNDA_2.n5145 GNDA_2.n4798 0.0672139
R14290 GNDA_2.n4609 GNDA_2.n4548 0.0672139
R14291 GNDA_2.n5210 GNDA_2.n5149 0.0672139
R14292 GNDA_2.n4770 GNDA_2.n161 0.0672139
R14293 GNDA_2.n4667 GNDA_2.n4646 0.0672139
R14294 GNDA_2.n4533 GNDA_2.n201 0.0672139
R14295 GNDA_2.n4268 GNDA_2.n4267 0.0672139
R14296 GNDA_2.n4262 GNDA_2.n4185 0.0672139
R14297 GNDA_2.n4153 GNDA_2.n4088 0.0672139
R14298 GNDA_2.n4072 GNDA_2.n1136 0.0672139
R14299 GNDA_2.n1208 GNDA_2.n1207 0.0672139
R14300 GNDA_2.n3679 GNDA_2.n3614 0.0672139
R14301 GNDA_2.n3748 GNDA_2.n3683 0.0672139
R14302 GNDA_2.n3817 GNDA_2.n3752 0.0672139
R14303 GNDA_2.n3886 GNDA_2.n3821 0.0672139
R14304 GNDA_2.n3951 GNDA_2.n3890 0.0672139
R14305 GNDA_2.n3001 GNDA_2.n3000 0.0672139
R14306 GNDA_2.n261 GNDA_2.n260 0.0672139
R14307 GNDA_2.n696 GNDA_2.n630 0.0672139
R14308 GNDA_2.n1012 GNDA_2.n444 0.0672139
R14309 GNDA_2.n516 GNDA_2.n515 0.0672139
R14310 GNDA_2.n800 GNDA_2.n735 0.0672139
R14311 GNDA_2.n869 GNDA_2.n804 0.0672139
R14312 GNDA_2.n934 GNDA_2.n873 0.0672139
R14313 GNDA_2.n1589 GNDA_2.n1588 0.0667303
R14314 GNDA_2.n4304 GNDA_2.n1091 0.0636702
R14315 GNDA_2.n1057 GNDA_2.n406 0.063
R14316 GNDA_2.n1050 GNDA_2.n1049 0.063
R14317 GNDA_2.n1039 GNDA_2.n421 0.063
R14318 GNDA_2.n5021 GNDA_2.n5020 0.063
R14319 GNDA_2.n5032 GNDA_2.n5005 0.063
R14320 GNDA_2.n5051 GNDA_2.n5050 0.063
R14321 GNDA_2.n4945 GNDA_2.n4944 0.063
R14322 GNDA_2.n4956 GNDA_2.n4924 0.063
R14323 GNDA_2.n4975 GNDA_2.n4974 0.063
R14324 GNDA_2.n4839 GNDA_2.n4838 0.063
R14325 GNDA_2.n4845 GNDA_2.n4844 0.063
R14326 GNDA_2.n4851 GNDA_2.n4850 0.063
R14327 GNDA_2.n5105 GNDA_2.n5104 0.063
R14328 GNDA_2.n5116 GNDA_2.n4803 0.063
R14329 GNDA_2.n5135 GNDA_2.n5134 0.063
R14330 GNDA_2.n4569 GNDA_2.n4568 0.063
R14331 GNDA_2.n4580 GNDA_2.n4553 0.063
R14332 GNDA_2.n4599 GNDA_2.n4598 0.063
R14333 GNDA_2.n5170 GNDA_2.n5169 0.063
R14334 GNDA_2.n5181 GNDA_2.n5154 0.063
R14335 GNDA_2.n5200 GNDA_2.n5199 0.063
R14336 GNDA_2.n4730 GNDA_2.n4729 0.063
R14337 GNDA_2.n4741 GNDA_2.n166 0.063
R14338 GNDA_2.n4760 GNDA_2.n4759 0.063
R14339 GNDA_2.n4651 GNDA_2.n4650 0.063
R14340 GNDA_2.n4657 GNDA_2.n4656 0.063
R14341 GNDA_2.n4663 GNDA_2.n4662 0.063
R14342 GNDA_2.n4493 GNDA_2.n4492 0.063
R14343 GNDA_2.n4504 GNDA_2.n206 0.063
R14344 GNDA_2.n4523 GNDA_2.n4522 0.063
R14345 GNDA_2.n4291 GNDA_2.n1098 0.063
R14346 GNDA_2.n4284 GNDA_2.n4283 0.063
R14347 GNDA_2.n4273 GNDA_2.n1113 0.063
R14348 GNDA_2.n4230 GNDA_2.n4229 0.063
R14349 GNDA_2.n4239 GNDA_2.n4194 0.063
R14350 GNDA_2.n4254 GNDA_2.n4253 0.063
R14351 GNDA_2.n4121 GNDA_2.n4120 0.063
R14352 GNDA_2.n4130 GNDA_2.n4097 0.063
R14353 GNDA_2.n4145 GNDA_2.n4144 0.063
R14354 GNDA_2.n4040 GNDA_2.n4039 0.063
R14355 GNDA_2.n4049 GNDA_2.n1145 0.063
R14356 GNDA_2.n4064 GNDA_2.n4063 0.063
R14357 GNDA_2.n1231 GNDA_2.n1167 0.063
R14358 GNDA_2.n1224 GNDA_2.n1223 0.063
R14359 GNDA_2.n1213 GNDA_2.n1191 0.063
R14360 GNDA_2.n3647 GNDA_2.n3646 0.063
R14361 GNDA_2.n3656 GNDA_2.n3623 0.063
R14362 GNDA_2.n3671 GNDA_2.n3670 0.063
R14363 GNDA_2.n3716 GNDA_2.n3715 0.063
R14364 GNDA_2.n3725 GNDA_2.n3692 0.063
R14365 GNDA_2.n3740 GNDA_2.n3739 0.063
R14366 GNDA_2.n3785 GNDA_2.n3784 0.063
R14367 GNDA_2.n3794 GNDA_2.n3761 0.063
R14368 GNDA_2.n3809 GNDA_2.n3808 0.063
R14369 GNDA_2.n3854 GNDA_2.n3853 0.063
R14370 GNDA_2.n3863 GNDA_2.n3830 0.063
R14371 GNDA_2.n3878 GNDA_2.n3877 0.063
R14372 GNDA_2.n3911 GNDA_2.n3910 0.063
R14373 GNDA_2.n3922 GNDA_2.n3895 0.063
R14374 GNDA_2.n3941 GNDA_2.n3940 0.063
R14375 GNDA_2.n3010 GNDA_2.n2993 0.063
R14376 GNDA_2.n3029 GNDA_2.n3028 0.063
R14377 GNDA_2.n3040 GNDA_2.n2981 0.063
R14378 GNDA_2.n3421 GNDA_2.n3420 0.063
R14379 GNDA_2.n3411 GNDA_2.n3410 0.063
R14380 GNDA_2.n284 GNDA_2.n220 0.063
R14381 GNDA_2.n277 GNDA_2.n276 0.063
R14382 GNDA_2.n266 GNDA_2.n244 0.063
R14383 GNDA_2.n601 GNDA_2.n595 0.063
R14384 GNDA_2.n570 GNDA_2.n386 0.063
R14385 GNDA_2.n664 GNDA_2.n663 0.063
R14386 GNDA_2.n673 GNDA_2.n639 0.063
R14387 GNDA_2.n688 GNDA_2.n687 0.063
R14388 GNDA_2.n980 GNDA_2.n979 0.063
R14389 GNDA_2.n989 GNDA_2.n453 0.063
R14390 GNDA_2.n1004 GNDA_2.n1003 0.063
R14391 GNDA_2.n539 GNDA_2.n475 0.063
R14392 GNDA_2.n532 GNDA_2.n531 0.063
R14393 GNDA_2.n521 GNDA_2.n499 0.063
R14394 GNDA_2.n768 GNDA_2.n767 0.063
R14395 GNDA_2.n777 GNDA_2.n744 0.063
R14396 GNDA_2.n792 GNDA_2.n791 0.063
R14397 GNDA_2.n837 GNDA_2.n836 0.063
R14398 GNDA_2.n846 GNDA_2.n813 0.063
R14399 GNDA_2.n861 GNDA_2.n860 0.063
R14400 GNDA_2.n894 GNDA_2.n893 0.063
R14401 GNDA_2.n905 GNDA_2.n878 0.063
R14402 GNDA_2.n924 GNDA_2.n923 0.063
R14403 GNDA_2.n4474 GNDA_2.n182 0.0629369
R14404 GNDA_2.n599 GNDA_2.n596 0.0626438
R14405 GNDA_2.n4340 GNDA_2.n4339 0.0626438
R14406 GNDA_2.n374 GNDA_2.n370 0.0626438
R14407 GNDA_2.n4358 GNDA_2.n4357 0.0626438
R14408 GNDA_2.n4401 GNDA_2.n337 0.0626438
R14409 GNDA_2.n4458 GNDA_2.n306 0.0626438
R14410 GNDA_2.n2670 GNDA_2.n2669 0.0626438
R14411 GNDA_2.n2695 GNDA_2.n2689 0.0626438
R14412 GNDA_2.n3067 GNDA_2.n2974 0.0626438
R14413 GNDA_2.n595 GNDA_2.n594 0.0577917
R14414 GNDA_2.n572 GNDA_2.n570 0.0577917
R14415 GNDA_2.n1016 GNDA_2.n404 0.0553333
R14416 GNDA_2.n413 GNDA_2.n412 0.0553333
R14417 GNDA_2.n1025 GNDA_2.n419 0.0553333
R14418 GNDA_2.n428 GNDA_2.n427 0.0553333
R14419 GNDA_2.n5014 GNDA_2.n5013 0.0553333
R14420 GNDA_2.n5028 GNDA_2.n5027 0.0553333
R14421 GNDA_2.n5044 GNDA_2.n5043 0.0553333
R14422 GNDA_2.n5058 GNDA_2.n5057 0.0553333
R14423 GNDA_2.n4938 GNDA_2.n4937 0.0553333
R14424 GNDA_2.n4952 GNDA_2.n4951 0.0553333
R14425 GNDA_2.n4968 GNDA_2.n4967 0.0553333
R14426 GNDA_2.n4982 GNDA_2.n4981 0.0553333
R14427 GNDA_2.n4887 GNDA_2.n4886 0.0553333
R14428 GNDA_2.n4878 GNDA_2.n4877 0.0553333
R14429 GNDA_2.n4869 GNDA_2.n4868 0.0553333
R14430 GNDA_2.n4860 GNDA_2.n4859 0.0553333
R14431 GNDA_2.n5098 GNDA_2.n5097 0.0553333
R14432 GNDA_2.n5112 GNDA_2.n5111 0.0553333
R14433 GNDA_2.n5128 GNDA_2.n5127 0.0553333
R14434 GNDA_2.n5142 GNDA_2.n5141 0.0553333
R14435 GNDA_2.n4562 GNDA_2.n4561 0.0553333
R14436 GNDA_2.n4576 GNDA_2.n4575 0.0553333
R14437 GNDA_2.n4592 GNDA_2.n4591 0.0553333
R14438 GNDA_2.n4606 GNDA_2.n4605 0.0553333
R14439 GNDA_2.n5163 GNDA_2.n5162 0.0553333
R14440 GNDA_2.n5177 GNDA_2.n5176 0.0553333
R14441 GNDA_2.n5193 GNDA_2.n5192 0.0553333
R14442 GNDA_2.n5207 GNDA_2.n5206 0.0553333
R14443 GNDA_2.n4723 GNDA_2.n4722 0.0553333
R14444 GNDA_2.n4737 GNDA_2.n4736 0.0553333
R14445 GNDA_2.n4753 GNDA_2.n4752 0.0553333
R14446 GNDA_2.n4767 GNDA_2.n4766 0.0553333
R14447 GNDA_2.n4699 GNDA_2.n4698 0.0553333
R14448 GNDA_2.n4690 GNDA_2.n4689 0.0553333
R14449 GNDA_2.n4681 GNDA_2.n4680 0.0553333
R14450 GNDA_2.n4672 GNDA_2.n4671 0.0553333
R14451 GNDA_2.n4486 GNDA_2.n4485 0.0553333
R14452 GNDA_2.n4500 GNDA_2.n4499 0.0553333
R14453 GNDA_2.n4516 GNDA_2.n4515 0.0553333
R14454 GNDA_2.n4530 GNDA_2.n4529 0.0553333
R14455 GNDA_2.n4157 GNDA_2.n1096 0.0553333
R14456 GNDA_2.n1105 GNDA_2.n1104 0.0553333
R14457 GNDA_2.n4166 GNDA_2.n1111 0.0553333
R14458 GNDA_2.n1120 GNDA_2.n1119 0.0553333
R14459 GNDA_2.n4205 GNDA_2.n4204 0.0553333
R14460 GNDA_2.n4235 GNDA_2.n4234 0.0553333
R14461 GNDA_2.n4193 GNDA_2.n4192 0.0553333
R14462 GNDA_2.n4259 GNDA_2.n4258 0.0553333
R14463 GNDA_2.n4108 GNDA_2.n4107 0.0553333
R14464 GNDA_2.n4126 GNDA_2.n4125 0.0553333
R14465 GNDA_2.n4096 GNDA_2.n4095 0.0553333
R14466 GNDA_2.n4150 GNDA_2.n4149 0.0553333
R14467 GNDA_2.n1156 GNDA_2.n1155 0.0553333
R14468 GNDA_2.n4045 GNDA_2.n4044 0.0553333
R14469 GNDA_2.n1144 GNDA_2.n1143 0.0553333
R14470 GNDA_2.n4069 GNDA_2.n4068 0.0553333
R14471 GNDA_2.n1168 GNDA_2.n1165 0.0553333
R14472 GNDA_2.n1179 GNDA_2.n1178 0.0553333
R14473 GNDA_2.n1192 GNDA_2.n1189 0.0553333
R14474 GNDA_2.n1203 GNDA_2.n1202 0.0553333
R14475 GNDA_2.n3634 GNDA_2.n3633 0.0553333
R14476 GNDA_2.n3652 GNDA_2.n3651 0.0553333
R14477 GNDA_2.n3622 GNDA_2.n3621 0.0553333
R14478 GNDA_2.n3676 GNDA_2.n3675 0.0553333
R14479 GNDA_2.n3703 GNDA_2.n3702 0.0553333
R14480 GNDA_2.n3721 GNDA_2.n3720 0.0553333
R14481 GNDA_2.n3691 GNDA_2.n3690 0.0553333
R14482 GNDA_2.n3745 GNDA_2.n3744 0.0553333
R14483 GNDA_2.n3772 GNDA_2.n3771 0.0553333
R14484 GNDA_2.n3790 GNDA_2.n3789 0.0553333
R14485 GNDA_2.n3760 GNDA_2.n3759 0.0553333
R14486 GNDA_2.n3814 GNDA_2.n3813 0.0553333
R14487 GNDA_2.n3841 GNDA_2.n3840 0.0553333
R14488 GNDA_2.n3859 GNDA_2.n3858 0.0553333
R14489 GNDA_2.n3829 GNDA_2.n3828 0.0553333
R14490 GNDA_2.n3883 GNDA_2.n3882 0.0553333
R14491 GNDA_2.n3904 GNDA_2.n3903 0.0553333
R14492 GNDA_2.n3918 GNDA_2.n3917 0.0553333
R14493 GNDA_2.n3934 GNDA_2.n3933 0.0553333
R14494 GNDA_2.n3948 GNDA_2.n3947 0.0553333
R14495 GNDA_2.n3006 GNDA_2.n3004 0.0553333
R14496 GNDA_2.n3022 GNDA_2.n2991 0.0553333
R14497 GNDA_2.n3036 GNDA_2.n3034 0.0553333
R14498 GNDA_2.n3052 GNDA_2.n2979 0.0553333
R14499 GNDA_2.n1593 GNDA_2.n1592 0.0553333
R14500 GNDA_2.n1607 GNDA_2.n1606 0.0553333
R14501 GNDA_2.n1623 GNDA_2.n1622 0.0553333
R14502 GNDA_2.n1637 GNDA_2.n1636 0.0553333
R14503 GNDA_2.n218 GNDA_2.n217 0.0553333
R14504 GNDA_2.n223 GNDA_2.n222 0.0553333
R14505 GNDA_2.n231 GNDA_2.n230 0.0553333
R14506 GNDA_2.n234 GNDA_2.n233 0.0553333
R14507 GNDA_2.n242 GNDA_2.n241 0.0553333
R14508 GNDA_2.n247 GNDA_2.n246 0.0553333
R14509 GNDA_2.n255 GNDA_2.n254 0.0553333
R14510 GNDA_2.n258 GNDA_2.n257 0.0553333
R14511 GNDA_2.n650 GNDA_2.n649 0.0553333
R14512 GNDA_2.n669 GNDA_2.n668 0.0553333
R14513 GNDA_2.n638 GNDA_2.n637 0.0553333
R14514 GNDA_2.n693 GNDA_2.n692 0.0553333
R14515 GNDA_2.n464 GNDA_2.n463 0.0553333
R14516 GNDA_2.n985 GNDA_2.n984 0.0553333
R14517 GNDA_2.n452 GNDA_2.n451 0.0553333
R14518 GNDA_2.n1009 GNDA_2.n1008 0.0553333
R14519 GNDA_2.n476 GNDA_2.n473 0.0553333
R14520 GNDA_2.n487 GNDA_2.n486 0.0553333
R14521 GNDA_2.n500 GNDA_2.n497 0.0553333
R14522 GNDA_2.n511 GNDA_2.n510 0.0553333
R14523 GNDA_2.n755 GNDA_2.n754 0.0553333
R14524 GNDA_2.n773 GNDA_2.n772 0.0553333
R14525 GNDA_2.n743 GNDA_2.n742 0.0553333
R14526 GNDA_2.n797 GNDA_2.n796 0.0553333
R14527 GNDA_2.n824 GNDA_2.n823 0.0553333
R14528 GNDA_2.n842 GNDA_2.n841 0.0553333
R14529 GNDA_2.n812 GNDA_2.n811 0.0553333
R14530 GNDA_2.n866 GNDA_2.n865 0.0553333
R14531 GNDA_2.n887 GNDA_2.n886 0.0553333
R14532 GNDA_2.n901 GNDA_2.n900 0.0553333
R14533 GNDA_2.n917 GNDA_2.n916 0.0553333
R14534 GNDA_2.n931 GNDA_2.n930 0.0553333
R14535 GNDA_2 GNDA_2.n5467 0.0517
R14536 GNDA_2 GNDA_2.n1898 0.0517
R14537 GNDA_2.n2843 GNDA_2 0.0517
R14538 GNDA_2.n2793 GNDA_2 0.0517
R14539 GNDA_2.n2117 GNDA_2 0.0517
R14540 GNDA_2.n5373 GNDA_2 0.0517
R14541 GNDA_2.n2246 GNDA_2 0.0517
R14542 GNDA_2.n3366 GNDA_2 0.0517
R14543 GNDA_2 GNDA_2.n0 0.0517
R14544 GNDA_2.n403 GNDA_2.n402 0.0514167
R14545 GNDA_2.n408 GNDA_2.n407 0.0514167
R14546 GNDA_2.n1019 GNDA_2.n409 0.0514167
R14547 GNDA_2.n1022 GNDA_2.n414 0.0514167
R14548 GNDA_2.n418 GNDA_2.n417 0.0514167
R14549 GNDA_2.n423 GNDA_2.n422 0.0514167
R14550 GNDA_2.n1028 GNDA_2.n424 0.0514167
R14551 GNDA_2.n1032 GNDA_2.n429 0.0514167
R14552 GNDA_2.n5064 GNDA_2.n4905 0.0514167
R14553 GNDA_2.n5018 GNDA_2.n5017 0.0514167
R14554 GNDA_2.n5024 GNDA_2.n5023 0.0514167
R14555 GNDA_2.n5034 GNDA_2.n5033 0.0514167
R14556 GNDA_2.n5038 GNDA_2.n5037 0.0514167
R14557 GNDA_2.n5048 GNDA_2.n5047 0.0514167
R14558 GNDA_2.n5054 GNDA_2.n5053 0.0514167
R14559 GNDA_2.n5062 GNDA_2.n4999 0.0514167
R14560 GNDA_2.n4932 GNDA_2.n4906 0.0514167
R14561 GNDA_2.n4942 GNDA_2.n4941 0.0514167
R14562 GNDA_2.n4948 GNDA_2.n4947 0.0514167
R14563 GNDA_2.n4958 GNDA_2.n4957 0.0514167
R14564 GNDA_2.n4962 GNDA_2.n4961 0.0514167
R14565 GNDA_2.n4972 GNDA_2.n4971 0.0514167
R14566 GNDA_2.n4978 GNDA_2.n4977 0.0514167
R14567 GNDA_2.n4986 GNDA_2.n4918 0.0514167
R14568 GNDA_2.n4890 GNDA_2.n4889 0.0514167
R14569 GNDA_2.n4884 GNDA_2.n4883 0.0514167
R14570 GNDA_2.n4881 GNDA_2.n4880 0.0514167
R14571 GNDA_2.n4875 GNDA_2.n4874 0.0514167
R14572 GNDA_2.n4872 GNDA_2.n4871 0.0514167
R14573 GNDA_2.n4866 GNDA_2.n4865 0.0514167
R14574 GNDA_2.n4863 GNDA_2.n4862 0.0514167
R14575 GNDA_2.n4857 GNDA_2.n4856 0.0514167
R14576 GNDA_2.n5092 GNDA_2.n4784 0.0514167
R14577 GNDA_2.n5102 GNDA_2.n5101 0.0514167
R14578 GNDA_2.n5108 GNDA_2.n5107 0.0514167
R14579 GNDA_2.n5118 GNDA_2.n5117 0.0514167
R14580 GNDA_2.n5122 GNDA_2.n5121 0.0514167
R14581 GNDA_2.n5132 GNDA_2.n5131 0.0514167
R14582 GNDA_2.n5138 GNDA_2.n5137 0.0514167
R14583 GNDA_2.n5146 GNDA_2.n4797 0.0514167
R14584 GNDA_2.n4612 GNDA_2.n186 0.0514167
R14585 GNDA_2.n4566 GNDA_2.n4565 0.0514167
R14586 GNDA_2.n4572 GNDA_2.n4571 0.0514167
R14587 GNDA_2.n4582 GNDA_2.n4581 0.0514167
R14588 GNDA_2.n4586 GNDA_2.n4585 0.0514167
R14589 GNDA_2.n4596 GNDA_2.n4595 0.0514167
R14590 GNDA_2.n4602 GNDA_2.n4601 0.0514167
R14591 GNDA_2.n4610 GNDA_2.n4547 0.0514167
R14592 GNDA_2.n5213 GNDA_2.n146 0.0514167
R14593 GNDA_2.n5167 GNDA_2.n5166 0.0514167
R14594 GNDA_2.n5173 GNDA_2.n5172 0.0514167
R14595 GNDA_2.n5183 GNDA_2.n5182 0.0514167
R14596 GNDA_2.n5187 GNDA_2.n5186 0.0514167
R14597 GNDA_2.n5197 GNDA_2.n5196 0.0514167
R14598 GNDA_2.n5203 GNDA_2.n5202 0.0514167
R14599 GNDA_2.n5211 GNDA_2.n5148 0.0514167
R14600 GNDA_2.n4717 GNDA_2.n148 0.0514167
R14601 GNDA_2.n4727 GNDA_2.n4726 0.0514167
R14602 GNDA_2.n4733 GNDA_2.n4732 0.0514167
R14603 GNDA_2.n4743 GNDA_2.n4742 0.0514167
R14604 GNDA_2.n4747 GNDA_2.n4746 0.0514167
R14605 GNDA_2.n4757 GNDA_2.n4756 0.0514167
R14606 GNDA_2.n4763 GNDA_2.n4762 0.0514167
R14607 GNDA_2.n4771 GNDA_2.n160 0.0514167
R14608 GNDA_2.n4702 GNDA_2.n4701 0.0514167
R14609 GNDA_2.n4696 GNDA_2.n4695 0.0514167
R14610 GNDA_2.n4693 GNDA_2.n4692 0.0514167
R14611 GNDA_2.n4687 GNDA_2.n4686 0.0514167
R14612 GNDA_2.n4684 GNDA_2.n4683 0.0514167
R14613 GNDA_2.n4678 GNDA_2.n4677 0.0514167
R14614 GNDA_2.n4675 GNDA_2.n4674 0.0514167
R14615 GNDA_2.n4669 GNDA_2.n4668 0.0514167
R14616 GNDA_2.n4480 GNDA_2.n188 0.0514167
R14617 GNDA_2.n4490 GNDA_2.n4489 0.0514167
R14618 GNDA_2.n4496 GNDA_2.n4495 0.0514167
R14619 GNDA_2.n4506 GNDA_2.n4505 0.0514167
R14620 GNDA_2.n4510 GNDA_2.n4509 0.0514167
R14621 GNDA_2.n4520 GNDA_2.n4519 0.0514167
R14622 GNDA_2.n4526 GNDA_2.n4525 0.0514167
R14623 GNDA_2.n4534 GNDA_2.n200 0.0514167
R14624 GNDA_2.n1095 GNDA_2.n1094 0.0514167
R14625 GNDA_2.n1100 GNDA_2.n1099 0.0514167
R14626 GNDA_2.n4160 GNDA_2.n1101 0.0514167
R14627 GNDA_2.n4163 GNDA_2.n1106 0.0514167
R14628 GNDA_2.n1110 GNDA_2.n1109 0.0514167
R14629 GNDA_2.n1115 GNDA_2.n1114 0.0514167
R14630 GNDA_2.n4169 GNDA_2.n1116 0.0514167
R14631 GNDA_2.n4266 GNDA_2.n1121 0.0514167
R14632 GNDA_2.n4219 GNDA_2.n4172 0.0514167
R14633 GNDA_2.n4227 GNDA_2.n4226 0.0514167
R14634 GNDA_2.n4201 GNDA_2.n4200 0.0514167
R14635 GNDA_2.n4197 GNDA_2.n4196 0.0514167
R14636 GNDA_2.n4243 GNDA_2.n4242 0.0514167
R14637 GNDA_2.n4251 GNDA_2.n4250 0.0514167
R14638 GNDA_2.n4189 GNDA_2.n4188 0.0514167
R14639 GNDA_2.n4263 GNDA_2.n4184 0.0514167
R14640 GNDA_2.n4110 GNDA_2.n4075 0.0514167
R14641 GNDA_2.n4118 GNDA_2.n4117 0.0514167
R14642 GNDA_2.n4104 GNDA_2.n4103 0.0514167
R14643 GNDA_2.n4100 GNDA_2.n4099 0.0514167
R14644 GNDA_2.n4134 GNDA_2.n4133 0.0514167
R14645 GNDA_2.n4142 GNDA_2.n4141 0.0514167
R14646 GNDA_2.n4092 GNDA_2.n4091 0.0514167
R14647 GNDA_2.n4154 GNDA_2.n4087 0.0514167
R14648 GNDA_2.n4029 GNDA_2.n1123 0.0514167
R14649 GNDA_2.n4037 GNDA_2.n4036 0.0514167
R14650 GNDA_2.n1152 GNDA_2.n1151 0.0514167
R14651 GNDA_2.n1148 GNDA_2.n1147 0.0514167
R14652 GNDA_2.n4053 GNDA_2.n4052 0.0514167
R14653 GNDA_2.n4061 GNDA_2.n4060 0.0514167
R14654 GNDA_2.n1140 GNDA_2.n1139 0.0514167
R14655 GNDA_2.n4073 GNDA_2.n1135 0.0514167
R14656 GNDA_2.n1163 GNDA_2.n1162 0.0514167
R14657 GNDA_2.n1171 GNDA_2.n1170 0.0514167
R14658 GNDA_2.n1176 GNDA_2.n1173 0.0514167
R14659 GNDA_2.n1184 GNDA_2.n1181 0.0514167
R14660 GNDA_2.n1187 GNDA_2.n1186 0.0514167
R14661 GNDA_2.n1195 GNDA_2.n1194 0.0514167
R14662 GNDA_2.n1200 GNDA_2.n1197 0.0514167
R14663 GNDA_2.n1206 GNDA_2.n1205 0.0514167
R14664 GNDA_2.n3636 GNDA_2.n3601 0.0514167
R14665 GNDA_2.n3644 GNDA_2.n3643 0.0514167
R14666 GNDA_2.n3630 GNDA_2.n3629 0.0514167
R14667 GNDA_2.n3626 GNDA_2.n3625 0.0514167
R14668 GNDA_2.n3660 GNDA_2.n3659 0.0514167
R14669 GNDA_2.n3668 GNDA_2.n3667 0.0514167
R14670 GNDA_2.n3618 GNDA_2.n3617 0.0514167
R14671 GNDA_2.n3680 GNDA_2.n3613 0.0514167
R14672 GNDA_2.n3705 GNDA_2.n3589 0.0514167
R14673 GNDA_2.n3713 GNDA_2.n3712 0.0514167
R14674 GNDA_2.n3699 GNDA_2.n3698 0.0514167
R14675 GNDA_2.n3695 GNDA_2.n3694 0.0514167
R14676 GNDA_2.n3729 GNDA_2.n3728 0.0514167
R14677 GNDA_2.n3737 GNDA_2.n3736 0.0514167
R14678 GNDA_2.n3687 GNDA_2.n3686 0.0514167
R14679 GNDA_2.n3749 GNDA_2.n3682 0.0514167
R14680 GNDA_2.n3774 GNDA_2.n3577 0.0514167
R14681 GNDA_2.n3782 GNDA_2.n3781 0.0514167
R14682 GNDA_2.n3768 GNDA_2.n3767 0.0514167
R14683 GNDA_2.n3764 GNDA_2.n3763 0.0514167
R14684 GNDA_2.n3798 GNDA_2.n3797 0.0514167
R14685 GNDA_2.n3806 GNDA_2.n3805 0.0514167
R14686 GNDA_2.n3756 GNDA_2.n3755 0.0514167
R14687 GNDA_2.n3818 GNDA_2.n3751 0.0514167
R14688 GNDA_2.n3843 GNDA_2.n3565 0.0514167
R14689 GNDA_2.n3851 GNDA_2.n3850 0.0514167
R14690 GNDA_2.n3837 GNDA_2.n3836 0.0514167
R14691 GNDA_2.n3833 GNDA_2.n3832 0.0514167
R14692 GNDA_2.n3867 GNDA_2.n3866 0.0514167
R14693 GNDA_2.n3875 GNDA_2.n3874 0.0514167
R14694 GNDA_2.n3825 GNDA_2.n3824 0.0514167
R14695 GNDA_2.n3887 GNDA_2.n3820 0.0514167
R14696 GNDA_2.n3954 GNDA_2.n1266 0.0514167
R14697 GNDA_2.n3908 GNDA_2.n3907 0.0514167
R14698 GNDA_2.n3914 GNDA_2.n3913 0.0514167
R14699 GNDA_2.n3924 GNDA_2.n3923 0.0514167
R14700 GNDA_2.n3928 GNDA_2.n3927 0.0514167
R14701 GNDA_2.n3938 GNDA_2.n3937 0.0514167
R14702 GNDA_2.n3944 GNDA_2.n3943 0.0514167
R14703 GNDA_2.n3952 GNDA_2.n3889 0.0514167
R14704 GNDA_2.n3002 GNDA_2.n2999 0.0514167
R14705 GNDA_2.n3012 GNDA_2.n2995 0.0514167
R14706 GNDA_2.n3016 GNDA_2.n3014 0.0514167
R14707 GNDA_2.n3026 GNDA_2.n3024 0.0514167
R14708 GNDA_2.n3032 GNDA_2.n2987 0.0514167
R14709 GNDA_2.n3042 GNDA_2.n2983 0.0514167
R14710 GNDA_2.n3046 GNDA_2.n3044 0.0514167
R14711 GNDA_2.n3055 GNDA_2.n3054 0.0514167
R14712 GNDA_2.n1587 GNDA_2.n1562 0.0514167
R14713 GNDA_2.n1597 GNDA_2.n1596 0.0514167
R14714 GNDA_2.n1603 GNDA_2.n1602 0.0514167
R14715 GNDA_2.n1613 GNDA_2.n1612 0.0514167
R14716 GNDA_2.n1617 GNDA_2.n1616 0.0514167
R14717 GNDA_2.n1627 GNDA_2.n1626 0.0514167
R14718 GNDA_2.n1633 GNDA_2.n1632 0.0514167
R14719 GNDA_2.n3436 GNDA_2.n1575 0.0514167
R14720 GNDA_2.n653 GNDA_2.n617 0.0514167
R14721 GNDA_2.n661 GNDA_2.n660 0.0514167
R14722 GNDA_2.n646 GNDA_2.n645 0.0514167
R14723 GNDA_2.n642 GNDA_2.n641 0.0514167
R14724 GNDA_2.n677 GNDA_2.n676 0.0514167
R14725 GNDA_2.n685 GNDA_2.n684 0.0514167
R14726 GNDA_2.n634 GNDA_2.n633 0.0514167
R14727 GNDA_2.n697 GNDA_2.n629 0.0514167
R14728 GNDA_2.n969 GNDA_2.n431 0.0514167
R14729 GNDA_2.n977 GNDA_2.n976 0.0514167
R14730 GNDA_2.n460 GNDA_2.n459 0.0514167
R14731 GNDA_2.n456 GNDA_2.n455 0.0514167
R14732 GNDA_2.n993 GNDA_2.n992 0.0514167
R14733 GNDA_2.n1001 GNDA_2.n1000 0.0514167
R14734 GNDA_2.n448 GNDA_2.n447 0.0514167
R14735 GNDA_2.n1013 GNDA_2.n443 0.0514167
R14736 GNDA_2.n471 GNDA_2.n470 0.0514167
R14737 GNDA_2.n479 GNDA_2.n478 0.0514167
R14738 GNDA_2.n484 GNDA_2.n481 0.0514167
R14739 GNDA_2.n492 GNDA_2.n489 0.0514167
R14740 GNDA_2.n495 GNDA_2.n494 0.0514167
R14741 GNDA_2.n503 GNDA_2.n502 0.0514167
R14742 GNDA_2.n508 GNDA_2.n505 0.0514167
R14743 GNDA_2.n514 GNDA_2.n513 0.0514167
R14744 GNDA_2.n757 GNDA_2.n722 0.0514167
R14745 GNDA_2.n765 GNDA_2.n764 0.0514167
R14746 GNDA_2.n751 GNDA_2.n750 0.0514167
R14747 GNDA_2.n747 GNDA_2.n746 0.0514167
R14748 GNDA_2.n781 GNDA_2.n780 0.0514167
R14749 GNDA_2.n789 GNDA_2.n788 0.0514167
R14750 GNDA_2.n739 GNDA_2.n738 0.0514167
R14751 GNDA_2.n801 GNDA_2.n734 0.0514167
R14752 GNDA_2.n826 GNDA_2.n710 0.0514167
R14753 GNDA_2.n834 GNDA_2.n833 0.0514167
R14754 GNDA_2.n820 GNDA_2.n819 0.0514167
R14755 GNDA_2.n816 GNDA_2.n815 0.0514167
R14756 GNDA_2.n850 GNDA_2.n849 0.0514167
R14757 GNDA_2.n858 GNDA_2.n857 0.0514167
R14758 GNDA_2.n808 GNDA_2.n807 0.0514167
R14759 GNDA_2.n870 GNDA_2.n803 0.0514167
R14760 GNDA_2.n937 GNDA_2.n616 0.0514167
R14761 GNDA_2.n891 GNDA_2.n890 0.0514167
R14762 GNDA_2.n897 GNDA_2.n896 0.0514167
R14763 GNDA_2.n907 GNDA_2.n906 0.0514167
R14764 GNDA_2.n911 GNDA_2.n910 0.0514167
R14765 GNDA_2.n921 GNDA_2.n920 0.0514167
R14766 GNDA_2.n927 GNDA_2.n926 0.0514167
R14767 GNDA_2.n935 GNDA_2.n872 0.0514167
R14768 GNDA_2.n226 GNDA_2.n225 0.0475
R14769 GNDA_2.n239 GNDA_2.n238 0.0475
R14770 GNDA_2.n250 GNDA_2.n249 0.0475
R14771 GNDA_2.n564 GNDA_2.n563 0.0421667
R14772 GNDA_2.n4477 GNDA_2.n4476 0.0421667
R14773 GNDA_2.n5249 GNDA_2.n5227 0.0421667
R14774 GNDA_2.n4418 GNDA_2.n325 0.0421667
R14775 GNDA_2.n4426 GNDA_2.n319 0.0421667
R14776 GNDA_2.n4443 GNDA_2.n316 0.0421667
R14777 GNDA_2.n4397 GNDA_2.n339 0.0421667
R14778 GNDA_2.n4378 GNDA_2.n4377 0.0421667
R14779 GNDA_2.n4413 GNDA_2.n329 0.0421667
R14780 GNDA_2.n4303 GNDA_2.n4302 0.0421667
R14781 GNDA_2.n3966 GNDA_2.n1257 0.0421667
R14782 GNDA_2.n3971 GNDA_2.n1253 0.0421667
R14783 GNDA_2.n3976 GNDA_2.n1249 0.0421667
R14784 GNDA_2.n4010 GNDA_2.n1246 0.0421667
R14785 GNDA_2.n4015 GNDA_2.n1242 0.0421667
R14786 GNDA_2.n4020 GNDA_2.n1158 0.0421667
R14787 GNDA_2.n4022 GNDA_2.n1085 0.0421667
R14788 GNDA_2.n4308 GNDA_2.n1090 0.0421667
R14789 GNDA_2.n4212 GNDA_2.n4207 0.0421667
R14790 GNDA_2.n2663 GNDA_2.n1683 0.0421667
R14791 GNDA_2.n299 GNDA_2.n212 0.0421667
R14792 GNDA_2.n4619 GNDA_2.n178 0.0421667
R14793 GNDA_2.n4709 GNDA_2.n175 0.0421667
R14794 GNDA_2.n173 GNDA_2.n142 0.0421667
R14795 GNDA_2.n5220 GNDA_2.n139 0.0421667
R14796 GNDA_2.n5223 GNDA_2.n138 0.0421667
R14797 GNDA_2.n5083 GNDA_2.n5082 0.0421667
R14798 GNDA_2.n5079 GNDA_2.n5078 0.0421667
R14799 GNDA_2.n5075 GNDA_2.n5074 0.0421667
R14800 GNDA_2.n5071 GNDA_2.n5070 0.0421667
R14801 GNDA_2.n394 GNDA_2.n392 0.0421667
R14802 GNDA_2.n950 GNDA_2.n554 0.0421667
R14803 GNDA_2.n955 GNDA_2.n550 0.0421667
R14804 GNDA_2.n960 GNDA_2.n466 0.0421667
R14805 GNDA_2.n962 GNDA_2.n400 0.0421667
R14806 GNDA_2.n1015 GNDA_2.n404 0.028198
R14807 GNDA_2.n1017 GNDA_2.n407 0.028198
R14808 GNDA_2.n1020 GNDA_2.n412 0.028198
R14809 GNDA_2.n1021 GNDA_2.n414 0.028198
R14810 GNDA_2.n1024 GNDA_2.n419 0.028198
R14811 GNDA_2.n1026 GNDA_2.n422 0.028198
R14812 GNDA_2.n1029 GNDA_2.n427 0.028198
R14813 GNDA_2.n1030 GNDA_2.n429 0.028198
R14814 GNDA_2.n5013 GNDA_2.n4988 0.028198
R14815 GNDA_2.n5017 GNDA_2.n4989 0.028198
R14816 GNDA_2.n5027 GNDA_2.n4991 0.028198
R14817 GNDA_2.n5033 GNDA_2.n4992 0.028198
R14818 GNDA_2.n5043 GNDA_2.n4994 0.028198
R14819 GNDA_2.n5047 GNDA_2.n4995 0.028198
R14820 GNDA_2.n5057 GNDA_2.n4997 0.028198
R14821 GNDA_2.n4999 GNDA_2.n4998 0.028198
R14822 GNDA_2.n4937 GNDA_2.n4907 0.028198
R14823 GNDA_2.n4941 GNDA_2.n4908 0.028198
R14824 GNDA_2.n4951 GNDA_2.n4910 0.028198
R14825 GNDA_2.n4957 GNDA_2.n4911 0.028198
R14826 GNDA_2.n4967 GNDA_2.n4913 0.028198
R14827 GNDA_2.n4971 GNDA_2.n4914 0.028198
R14828 GNDA_2.n4981 GNDA_2.n4916 0.028198
R14829 GNDA_2.n4918 GNDA_2.n4917 0.028198
R14830 GNDA_2.n4888 GNDA_2.n4887 0.028198
R14831 GNDA_2.n4885 GNDA_2.n4884 0.028198
R14832 GNDA_2.n4879 GNDA_2.n4878 0.028198
R14833 GNDA_2.n4876 GNDA_2.n4875 0.028198
R14834 GNDA_2.n4870 GNDA_2.n4869 0.028198
R14835 GNDA_2.n4867 GNDA_2.n4866 0.028198
R14836 GNDA_2.n4861 GNDA_2.n4860 0.028198
R14837 GNDA_2.n4858 GNDA_2.n4857 0.028198
R14838 GNDA_2.n5097 GNDA_2.n4785 0.028198
R14839 GNDA_2.n5101 GNDA_2.n4786 0.028198
R14840 GNDA_2.n5111 GNDA_2.n4788 0.028198
R14841 GNDA_2.n5117 GNDA_2.n4789 0.028198
R14842 GNDA_2.n5127 GNDA_2.n4791 0.028198
R14843 GNDA_2.n5131 GNDA_2.n4792 0.028198
R14844 GNDA_2.n5141 GNDA_2.n4794 0.028198
R14845 GNDA_2.n4797 GNDA_2.n4795 0.028198
R14846 GNDA_2.n4561 GNDA_2.n4536 0.028198
R14847 GNDA_2.n4565 GNDA_2.n4537 0.028198
R14848 GNDA_2.n4575 GNDA_2.n4539 0.028198
R14849 GNDA_2.n4581 GNDA_2.n4540 0.028198
R14850 GNDA_2.n4591 GNDA_2.n4542 0.028198
R14851 GNDA_2.n4595 GNDA_2.n4543 0.028198
R14852 GNDA_2.n4605 GNDA_2.n4545 0.028198
R14853 GNDA_2.n4547 GNDA_2.n4546 0.028198
R14854 GNDA_2.n5162 GNDA_2.n4773 0.028198
R14855 GNDA_2.n5166 GNDA_2.n4774 0.028198
R14856 GNDA_2.n5176 GNDA_2.n4776 0.028198
R14857 GNDA_2.n5182 GNDA_2.n4777 0.028198
R14858 GNDA_2.n5192 GNDA_2.n4779 0.028198
R14859 GNDA_2.n5196 GNDA_2.n4780 0.028198
R14860 GNDA_2.n5206 GNDA_2.n4782 0.028198
R14861 GNDA_2.n5148 GNDA_2.n4783 0.028198
R14862 GNDA_2.n4722 GNDA_2.n149 0.028198
R14863 GNDA_2.n4726 GNDA_2.n150 0.028198
R14864 GNDA_2.n4736 GNDA_2.n152 0.028198
R14865 GNDA_2.n4742 GNDA_2.n153 0.028198
R14866 GNDA_2.n4752 GNDA_2.n155 0.028198
R14867 GNDA_2.n4756 GNDA_2.n156 0.028198
R14868 GNDA_2.n4766 GNDA_2.n158 0.028198
R14869 GNDA_2.n160 GNDA_2.n159 0.028198
R14870 GNDA_2.n4700 GNDA_2.n4699 0.028198
R14871 GNDA_2.n4697 GNDA_2.n4696 0.028198
R14872 GNDA_2.n4691 GNDA_2.n4690 0.028198
R14873 GNDA_2.n4688 GNDA_2.n4687 0.028198
R14874 GNDA_2.n4682 GNDA_2.n4681 0.028198
R14875 GNDA_2.n4679 GNDA_2.n4678 0.028198
R14876 GNDA_2.n4673 GNDA_2.n4672 0.028198
R14877 GNDA_2.n4670 GNDA_2.n4669 0.028198
R14878 GNDA_2.n4485 GNDA_2.n189 0.028198
R14879 GNDA_2.n4489 GNDA_2.n190 0.028198
R14880 GNDA_2.n4499 GNDA_2.n192 0.028198
R14881 GNDA_2.n4505 GNDA_2.n193 0.028198
R14882 GNDA_2.n4515 GNDA_2.n195 0.028198
R14883 GNDA_2.n4519 GNDA_2.n196 0.028198
R14884 GNDA_2.n4529 GNDA_2.n198 0.028198
R14885 GNDA_2.n200 GNDA_2.n199 0.028198
R14886 GNDA_2.n4156 GNDA_2.n1096 0.028198
R14887 GNDA_2.n4158 GNDA_2.n1099 0.028198
R14888 GNDA_2.n4161 GNDA_2.n1104 0.028198
R14889 GNDA_2.n4162 GNDA_2.n1106 0.028198
R14890 GNDA_2.n4165 GNDA_2.n1111 0.028198
R14891 GNDA_2.n4167 GNDA_2.n1114 0.028198
R14892 GNDA_2.n4170 GNDA_2.n1119 0.028198
R14893 GNDA_2.n4171 GNDA_2.n1121 0.028198
R14894 GNDA_2.n4204 GNDA_2.n4173 0.028198
R14895 GNDA_2.n4226 GNDA_2.n4174 0.028198
R14896 GNDA_2.n4234 GNDA_2.n4176 0.028198
R14897 GNDA_2.n4196 GNDA_2.n4177 0.028198
R14898 GNDA_2.n4192 GNDA_2.n4179 0.028198
R14899 GNDA_2.n4250 GNDA_2.n4180 0.028198
R14900 GNDA_2.n4258 GNDA_2.n4182 0.028198
R14901 GNDA_2.n4184 GNDA_2.n4183 0.028198
R14902 GNDA_2.n4107 GNDA_2.n4076 0.028198
R14903 GNDA_2.n4117 GNDA_2.n4077 0.028198
R14904 GNDA_2.n4125 GNDA_2.n4079 0.028198
R14905 GNDA_2.n4099 GNDA_2.n4080 0.028198
R14906 GNDA_2.n4095 GNDA_2.n4082 0.028198
R14907 GNDA_2.n4141 GNDA_2.n4083 0.028198
R14908 GNDA_2.n4149 GNDA_2.n4085 0.028198
R14909 GNDA_2.n4087 GNDA_2.n4086 0.028198
R14910 GNDA_2.n1155 GNDA_2.n1124 0.028198
R14911 GNDA_2.n4036 GNDA_2.n1125 0.028198
R14912 GNDA_2.n4044 GNDA_2.n1127 0.028198
R14913 GNDA_2.n1147 GNDA_2.n1128 0.028198
R14914 GNDA_2.n1143 GNDA_2.n1130 0.028198
R14915 GNDA_2.n4060 GNDA_2.n1131 0.028198
R14916 GNDA_2.n4068 GNDA_2.n1133 0.028198
R14917 GNDA_2.n1135 GNDA_2.n1134 0.028198
R14918 GNDA_2.n1165 GNDA_2.n1164 0.028198
R14919 GNDA_2.n1170 GNDA_2.n1169 0.028198
R14920 GNDA_2.n1178 GNDA_2.n1177 0.028198
R14921 GNDA_2.n1181 GNDA_2.n1180 0.028198
R14922 GNDA_2.n1189 GNDA_2.n1188 0.028198
R14923 GNDA_2.n1194 GNDA_2.n1193 0.028198
R14924 GNDA_2.n1202 GNDA_2.n1201 0.028198
R14925 GNDA_2.n1205 GNDA_2.n1204 0.028198
R14926 GNDA_2.n3633 GNDA_2.n3602 0.028198
R14927 GNDA_2.n3643 GNDA_2.n3603 0.028198
R14928 GNDA_2.n3651 GNDA_2.n3605 0.028198
R14929 GNDA_2.n3625 GNDA_2.n3606 0.028198
R14930 GNDA_2.n3621 GNDA_2.n3608 0.028198
R14931 GNDA_2.n3667 GNDA_2.n3609 0.028198
R14932 GNDA_2.n3675 GNDA_2.n3611 0.028198
R14933 GNDA_2.n3613 GNDA_2.n3612 0.028198
R14934 GNDA_2.n3702 GNDA_2.n3590 0.028198
R14935 GNDA_2.n3712 GNDA_2.n3591 0.028198
R14936 GNDA_2.n3720 GNDA_2.n3593 0.028198
R14937 GNDA_2.n3694 GNDA_2.n3594 0.028198
R14938 GNDA_2.n3690 GNDA_2.n3596 0.028198
R14939 GNDA_2.n3736 GNDA_2.n3597 0.028198
R14940 GNDA_2.n3744 GNDA_2.n3599 0.028198
R14941 GNDA_2.n3682 GNDA_2.n3600 0.028198
R14942 GNDA_2.n3771 GNDA_2.n3578 0.028198
R14943 GNDA_2.n3781 GNDA_2.n3579 0.028198
R14944 GNDA_2.n3789 GNDA_2.n3581 0.028198
R14945 GNDA_2.n3763 GNDA_2.n3582 0.028198
R14946 GNDA_2.n3759 GNDA_2.n3584 0.028198
R14947 GNDA_2.n3805 GNDA_2.n3585 0.028198
R14948 GNDA_2.n3813 GNDA_2.n3587 0.028198
R14949 GNDA_2.n3751 GNDA_2.n3588 0.028198
R14950 GNDA_2.n3840 GNDA_2.n3566 0.028198
R14951 GNDA_2.n3850 GNDA_2.n3567 0.028198
R14952 GNDA_2.n3858 GNDA_2.n3569 0.028198
R14953 GNDA_2.n3832 GNDA_2.n3570 0.028198
R14954 GNDA_2.n3828 GNDA_2.n3572 0.028198
R14955 GNDA_2.n3874 GNDA_2.n3573 0.028198
R14956 GNDA_2.n3882 GNDA_2.n3575 0.028198
R14957 GNDA_2.n3820 GNDA_2.n3576 0.028198
R14958 GNDA_2.n3903 GNDA_2.n3554 0.028198
R14959 GNDA_2.n3907 GNDA_2.n3555 0.028198
R14960 GNDA_2.n3917 GNDA_2.n3557 0.028198
R14961 GNDA_2.n3923 GNDA_2.n3558 0.028198
R14962 GNDA_2.n3933 GNDA_2.n3560 0.028198
R14963 GNDA_2.n3937 GNDA_2.n3561 0.028198
R14964 GNDA_2.n3947 GNDA_2.n3563 0.028198
R14965 GNDA_2.n3889 GNDA_2.n3564 0.028198
R14966 GNDA_2.n3004 GNDA_2.n3003 0.028198
R14967 GNDA_2.n3005 GNDA_2.n2995 0.028198
R14968 GNDA_2.n3015 GNDA_2.n2991 0.028198
R14969 GNDA_2.n3024 GNDA_2.n3023 0.028198
R14970 GNDA_2.n3034 GNDA_2.n3033 0.028198
R14971 GNDA_2.n3035 GNDA_2.n2983 0.028198
R14972 GNDA_2.n3045 GNDA_2.n2979 0.028198
R14973 GNDA_2.n3054 GNDA_2.n3053 0.028198
R14974 GNDA_2.n1592 GNDA_2.n1563 0.028198
R14975 GNDA_2.n1596 GNDA_2.n1564 0.028198
R14976 GNDA_2.n1606 GNDA_2.n1566 0.028198
R14977 GNDA_2.n1612 GNDA_2.n1567 0.028198
R14978 GNDA_2.n1622 GNDA_2.n1569 0.028198
R14979 GNDA_2.n1626 GNDA_2.n1570 0.028198
R14980 GNDA_2.n1636 GNDA_2.n1572 0.028198
R14981 GNDA_2.n1575 GNDA_2.n1573 0.028198
R14982 GNDA_2.n1637 GNDA_2.n1573 0.028198
R14983 GNDA_2.n1633 GNDA_2.n1572 0.028198
R14984 GNDA_2.n1623 GNDA_2.n1570 0.028198
R14985 GNDA_2.n1617 GNDA_2.n1569 0.028198
R14986 GNDA_2.n1607 GNDA_2.n1567 0.028198
R14987 GNDA_2.n1603 GNDA_2.n1566 0.028198
R14988 GNDA_2.n1593 GNDA_2.n1564 0.028198
R14989 GNDA_2.n1587 GNDA_2.n1563 0.028198
R14990 GNDA_2.n3053 GNDA_2.n3052 0.028198
R14991 GNDA_2.n3046 GNDA_2.n3045 0.028198
R14992 GNDA_2.n3036 GNDA_2.n3035 0.028198
R14993 GNDA_2.n3033 GNDA_2.n3032 0.028198
R14994 GNDA_2.n3023 GNDA_2.n3022 0.028198
R14995 GNDA_2.n3016 GNDA_2.n3015 0.028198
R14996 GNDA_2.n3006 GNDA_2.n3005 0.028198
R14997 GNDA_2.n3003 GNDA_2.n3002 0.028198
R14998 GNDA_2.n3948 GNDA_2.n3564 0.028198
R14999 GNDA_2.n3944 GNDA_2.n3563 0.028198
R15000 GNDA_2.n3934 GNDA_2.n3561 0.028198
R15001 GNDA_2.n3928 GNDA_2.n3560 0.028198
R15002 GNDA_2.n3918 GNDA_2.n3558 0.028198
R15003 GNDA_2.n3914 GNDA_2.n3557 0.028198
R15004 GNDA_2.n3904 GNDA_2.n3555 0.028198
R15005 GNDA_2.n3554 GNDA_2.n1266 0.028198
R15006 GNDA_2.n3883 GNDA_2.n3576 0.028198
R15007 GNDA_2.n3825 GNDA_2.n3575 0.028198
R15008 GNDA_2.n3829 GNDA_2.n3573 0.028198
R15009 GNDA_2.n3867 GNDA_2.n3572 0.028198
R15010 GNDA_2.n3859 GNDA_2.n3570 0.028198
R15011 GNDA_2.n3837 GNDA_2.n3569 0.028198
R15012 GNDA_2.n3841 GNDA_2.n3567 0.028198
R15013 GNDA_2.n3843 GNDA_2.n3566 0.028198
R15014 GNDA_2.n3814 GNDA_2.n3588 0.028198
R15015 GNDA_2.n3756 GNDA_2.n3587 0.028198
R15016 GNDA_2.n3760 GNDA_2.n3585 0.028198
R15017 GNDA_2.n3798 GNDA_2.n3584 0.028198
R15018 GNDA_2.n3790 GNDA_2.n3582 0.028198
R15019 GNDA_2.n3768 GNDA_2.n3581 0.028198
R15020 GNDA_2.n3772 GNDA_2.n3579 0.028198
R15021 GNDA_2.n3774 GNDA_2.n3578 0.028198
R15022 GNDA_2.n3745 GNDA_2.n3600 0.028198
R15023 GNDA_2.n3687 GNDA_2.n3599 0.028198
R15024 GNDA_2.n3691 GNDA_2.n3597 0.028198
R15025 GNDA_2.n3729 GNDA_2.n3596 0.028198
R15026 GNDA_2.n3721 GNDA_2.n3594 0.028198
R15027 GNDA_2.n3699 GNDA_2.n3593 0.028198
R15028 GNDA_2.n3703 GNDA_2.n3591 0.028198
R15029 GNDA_2.n3705 GNDA_2.n3590 0.028198
R15030 GNDA_2.n3676 GNDA_2.n3612 0.028198
R15031 GNDA_2.n3618 GNDA_2.n3611 0.028198
R15032 GNDA_2.n3622 GNDA_2.n3609 0.028198
R15033 GNDA_2.n3660 GNDA_2.n3608 0.028198
R15034 GNDA_2.n3652 GNDA_2.n3606 0.028198
R15035 GNDA_2.n3630 GNDA_2.n3605 0.028198
R15036 GNDA_2.n3634 GNDA_2.n3603 0.028198
R15037 GNDA_2.n3636 GNDA_2.n3602 0.028198
R15038 GNDA_2.n1204 GNDA_2.n1203 0.028198
R15039 GNDA_2.n1201 GNDA_2.n1200 0.028198
R15040 GNDA_2.n1193 GNDA_2.n1192 0.028198
R15041 GNDA_2.n1188 GNDA_2.n1187 0.028198
R15042 GNDA_2.n1180 GNDA_2.n1179 0.028198
R15043 GNDA_2.n1177 GNDA_2.n1176 0.028198
R15044 GNDA_2.n1169 GNDA_2.n1168 0.028198
R15045 GNDA_2.n1164 GNDA_2.n1163 0.028198
R15046 GNDA_2.n4069 GNDA_2.n1134 0.028198
R15047 GNDA_2.n1140 GNDA_2.n1133 0.028198
R15048 GNDA_2.n1144 GNDA_2.n1131 0.028198
R15049 GNDA_2.n4053 GNDA_2.n1130 0.028198
R15050 GNDA_2.n4045 GNDA_2.n1128 0.028198
R15051 GNDA_2.n1152 GNDA_2.n1127 0.028198
R15052 GNDA_2.n1156 GNDA_2.n1125 0.028198
R15053 GNDA_2.n4029 GNDA_2.n1124 0.028198
R15054 GNDA_2.n4150 GNDA_2.n4086 0.028198
R15055 GNDA_2.n4092 GNDA_2.n4085 0.028198
R15056 GNDA_2.n4096 GNDA_2.n4083 0.028198
R15057 GNDA_2.n4134 GNDA_2.n4082 0.028198
R15058 GNDA_2.n4126 GNDA_2.n4080 0.028198
R15059 GNDA_2.n4104 GNDA_2.n4079 0.028198
R15060 GNDA_2.n4108 GNDA_2.n4077 0.028198
R15061 GNDA_2.n4110 GNDA_2.n4076 0.028198
R15062 GNDA_2.n4259 GNDA_2.n4183 0.028198
R15063 GNDA_2.n4189 GNDA_2.n4182 0.028198
R15064 GNDA_2.n4193 GNDA_2.n4180 0.028198
R15065 GNDA_2.n4243 GNDA_2.n4179 0.028198
R15066 GNDA_2.n4235 GNDA_2.n4177 0.028198
R15067 GNDA_2.n4201 GNDA_2.n4176 0.028198
R15068 GNDA_2.n4205 GNDA_2.n4174 0.028198
R15069 GNDA_2.n4219 GNDA_2.n4173 0.028198
R15070 GNDA_2.n4171 GNDA_2.n1120 0.028198
R15071 GNDA_2.n4170 GNDA_2.n4169 0.028198
R15072 GNDA_2.n4167 GNDA_2.n4166 0.028198
R15073 GNDA_2.n4165 GNDA_2.n1110 0.028198
R15074 GNDA_2.n4162 GNDA_2.n1105 0.028198
R15075 GNDA_2.n4161 GNDA_2.n4160 0.028198
R15076 GNDA_2.n4158 GNDA_2.n4157 0.028198
R15077 GNDA_2.n4156 GNDA_2.n1095 0.028198
R15078 GNDA_2.n4530 GNDA_2.n199 0.028198
R15079 GNDA_2.n4526 GNDA_2.n198 0.028198
R15080 GNDA_2.n4516 GNDA_2.n196 0.028198
R15081 GNDA_2.n4510 GNDA_2.n195 0.028198
R15082 GNDA_2.n4500 GNDA_2.n193 0.028198
R15083 GNDA_2.n4496 GNDA_2.n192 0.028198
R15084 GNDA_2.n4486 GNDA_2.n190 0.028198
R15085 GNDA_2.n4480 GNDA_2.n189 0.028198
R15086 GNDA_2.n4671 GNDA_2.n4670 0.028198
R15087 GNDA_2.n4674 GNDA_2.n4673 0.028198
R15088 GNDA_2.n4680 GNDA_2.n4679 0.028198
R15089 GNDA_2.n4683 GNDA_2.n4682 0.028198
R15090 GNDA_2.n4689 GNDA_2.n4688 0.028198
R15091 GNDA_2.n4692 GNDA_2.n4691 0.028198
R15092 GNDA_2.n4698 GNDA_2.n4697 0.028198
R15093 GNDA_2.n4701 GNDA_2.n4700 0.028198
R15094 GNDA_2.n4767 GNDA_2.n159 0.028198
R15095 GNDA_2.n4763 GNDA_2.n158 0.028198
R15096 GNDA_2.n4753 GNDA_2.n156 0.028198
R15097 GNDA_2.n4747 GNDA_2.n155 0.028198
R15098 GNDA_2.n4737 GNDA_2.n153 0.028198
R15099 GNDA_2.n4733 GNDA_2.n152 0.028198
R15100 GNDA_2.n4723 GNDA_2.n150 0.028198
R15101 GNDA_2.n4717 GNDA_2.n149 0.028198
R15102 GNDA_2.n5207 GNDA_2.n4783 0.028198
R15103 GNDA_2.n5203 GNDA_2.n4782 0.028198
R15104 GNDA_2.n5193 GNDA_2.n4780 0.028198
R15105 GNDA_2.n5187 GNDA_2.n4779 0.028198
R15106 GNDA_2.n5177 GNDA_2.n4777 0.028198
R15107 GNDA_2.n5173 GNDA_2.n4776 0.028198
R15108 GNDA_2.n5163 GNDA_2.n4774 0.028198
R15109 GNDA_2.n4773 GNDA_2.n146 0.028198
R15110 GNDA_2.n4606 GNDA_2.n4546 0.028198
R15111 GNDA_2.n4602 GNDA_2.n4545 0.028198
R15112 GNDA_2.n4592 GNDA_2.n4543 0.028198
R15113 GNDA_2.n4586 GNDA_2.n4542 0.028198
R15114 GNDA_2.n4576 GNDA_2.n4540 0.028198
R15115 GNDA_2.n4572 GNDA_2.n4539 0.028198
R15116 GNDA_2.n4562 GNDA_2.n4537 0.028198
R15117 GNDA_2.n4536 GNDA_2.n186 0.028198
R15118 GNDA_2.n5142 GNDA_2.n4795 0.028198
R15119 GNDA_2.n5138 GNDA_2.n4794 0.028198
R15120 GNDA_2.n5128 GNDA_2.n4792 0.028198
R15121 GNDA_2.n5122 GNDA_2.n4791 0.028198
R15122 GNDA_2.n5112 GNDA_2.n4789 0.028198
R15123 GNDA_2.n5108 GNDA_2.n4788 0.028198
R15124 GNDA_2.n5098 GNDA_2.n4786 0.028198
R15125 GNDA_2.n5092 GNDA_2.n4785 0.028198
R15126 GNDA_2.n4859 GNDA_2.n4858 0.028198
R15127 GNDA_2.n4862 GNDA_2.n4861 0.028198
R15128 GNDA_2.n4868 GNDA_2.n4867 0.028198
R15129 GNDA_2.n4871 GNDA_2.n4870 0.028198
R15130 GNDA_2.n4877 GNDA_2.n4876 0.028198
R15131 GNDA_2.n4880 GNDA_2.n4879 0.028198
R15132 GNDA_2.n4886 GNDA_2.n4885 0.028198
R15133 GNDA_2.n4889 GNDA_2.n4888 0.028198
R15134 GNDA_2.n4982 GNDA_2.n4917 0.028198
R15135 GNDA_2.n4978 GNDA_2.n4916 0.028198
R15136 GNDA_2.n4968 GNDA_2.n4914 0.028198
R15137 GNDA_2.n4962 GNDA_2.n4913 0.028198
R15138 GNDA_2.n4952 GNDA_2.n4911 0.028198
R15139 GNDA_2.n4948 GNDA_2.n4910 0.028198
R15140 GNDA_2.n4938 GNDA_2.n4908 0.028198
R15141 GNDA_2.n4932 GNDA_2.n4907 0.028198
R15142 GNDA_2.n5058 GNDA_2.n4998 0.028198
R15143 GNDA_2.n5054 GNDA_2.n4997 0.028198
R15144 GNDA_2.n5044 GNDA_2.n4995 0.028198
R15145 GNDA_2.n5038 GNDA_2.n4994 0.028198
R15146 GNDA_2.n5028 GNDA_2.n4992 0.028198
R15147 GNDA_2.n5024 GNDA_2.n4991 0.028198
R15148 GNDA_2.n5014 GNDA_2.n4989 0.028198
R15149 GNDA_2.n4988 GNDA_2.n4905 0.028198
R15150 GNDA_2.n649 GNDA_2.n618 0.028198
R15151 GNDA_2.n660 GNDA_2.n619 0.028198
R15152 GNDA_2.n668 GNDA_2.n621 0.028198
R15153 GNDA_2.n641 GNDA_2.n622 0.028198
R15154 GNDA_2.n637 GNDA_2.n624 0.028198
R15155 GNDA_2.n684 GNDA_2.n625 0.028198
R15156 GNDA_2.n692 GNDA_2.n627 0.028198
R15157 GNDA_2.n629 GNDA_2.n628 0.028198
R15158 GNDA_2.n463 GNDA_2.n432 0.028198
R15159 GNDA_2.n976 GNDA_2.n433 0.028198
R15160 GNDA_2.n984 GNDA_2.n435 0.028198
R15161 GNDA_2.n455 GNDA_2.n436 0.028198
R15162 GNDA_2.n451 GNDA_2.n438 0.028198
R15163 GNDA_2.n1000 GNDA_2.n439 0.028198
R15164 GNDA_2.n1008 GNDA_2.n441 0.028198
R15165 GNDA_2.n443 GNDA_2.n442 0.028198
R15166 GNDA_2.n473 GNDA_2.n472 0.028198
R15167 GNDA_2.n478 GNDA_2.n477 0.028198
R15168 GNDA_2.n486 GNDA_2.n485 0.028198
R15169 GNDA_2.n489 GNDA_2.n488 0.028198
R15170 GNDA_2.n497 GNDA_2.n496 0.028198
R15171 GNDA_2.n502 GNDA_2.n501 0.028198
R15172 GNDA_2.n510 GNDA_2.n509 0.028198
R15173 GNDA_2.n513 GNDA_2.n512 0.028198
R15174 GNDA_2.n754 GNDA_2.n723 0.028198
R15175 GNDA_2.n764 GNDA_2.n724 0.028198
R15176 GNDA_2.n772 GNDA_2.n726 0.028198
R15177 GNDA_2.n746 GNDA_2.n727 0.028198
R15178 GNDA_2.n742 GNDA_2.n729 0.028198
R15179 GNDA_2.n788 GNDA_2.n730 0.028198
R15180 GNDA_2.n796 GNDA_2.n732 0.028198
R15181 GNDA_2.n734 GNDA_2.n733 0.028198
R15182 GNDA_2.n823 GNDA_2.n711 0.028198
R15183 GNDA_2.n833 GNDA_2.n712 0.028198
R15184 GNDA_2.n841 GNDA_2.n714 0.028198
R15185 GNDA_2.n815 GNDA_2.n715 0.028198
R15186 GNDA_2.n811 GNDA_2.n717 0.028198
R15187 GNDA_2.n857 GNDA_2.n718 0.028198
R15188 GNDA_2.n865 GNDA_2.n720 0.028198
R15189 GNDA_2.n803 GNDA_2.n721 0.028198
R15190 GNDA_2.n886 GNDA_2.n699 0.028198
R15191 GNDA_2.n890 GNDA_2.n700 0.028198
R15192 GNDA_2.n900 GNDA_2.n702 0.028198
R15193 GNDA_2.n906 GNDA_2.n703 0.028198
R15194 GNDA_2.n916 GNDA_2.n705 0.028198
R15195 GNDA_2.n920 GNDA_2.n706 0.028198
R15196 GNDA_2.n930 GNDA_2.n708 0.028198
R15197 GNDA_2.n872 GNDA_2.n709 0.028198
R15198 GNDA_2.n931 GNDA_2.n709 0.028198
R15199 GNDA_2.n927 GNDA_2.n708 0.028198
R15200 GNDA_2.n917 GNDA_2.n706 0.028198
R15201 GNDA_2.n911 GNDA_2.n705 0.028198
R15202 GNDA_2.n901 GNDA_2.n703 0.028198
R15203 GNDA_2.n897 GNDA_2.n702 0.028198
R15204 GNDA_2.n887 GNDA_2.n700 0.028198
R15205 GNDA_2.n699 GNDA_2.n616 0.028198
R15206 GNDA_2.n866 GNDA_2.n721 0.028198
R15207 GNDA_2.n808 GNDA_2.n720 0.028198
R15208 GNDA_2.n812 GNDA_2.n718 0.028198
R15209 GNDA_2.n850 GNDA_2.n717 0.028198
R15210 GNDA_2.n842 GNDA_2.n715 0.028198
R15211 GNDA_2.n820 GNDA_2.n714 0.028198
R15212 GNDA_2.n824 GNDA_2.n712 0.028198
R15213 GNDA_2.n826 GNDA_2.n711 0.028198
R15214 GNDA_2.n797 GNDA_2.n733 0.028198
R15215 GNDA_2.n739 GNDA_2.n732 0.028198
R15216 GNDA_2.n743 GNDA_2.n730 0.028198
R15217 GNDA_2.n781 GNDA_2.n729 0.028198
R15218 GNDA_2.n773 GNDA_2.n727 0.028198
R15219 GNDA_2.n751 GNDA_2.n726 0.028198
R15220 GNDA_2.n755 GNDA_2.n724 0.028198
R15221 GNDA_2.n757 GNDA_2.n723 0.028198
R15222 GNDA_2.n512 GNDA_2.n511 0.028198
R15223 GNDA_2.n509 GNDA_2.n508 0.028198
R15224 GNDA_2.n501 GNDA_2.n500 0.028198
R15225 GNDA_2.n496 GNDA_2.n495 0.028198
R15226 GNDA_2.n488 GNDA_2.n487 0.028198
R15227 GNDA_2.n485 GNDA_2.n484 0.028198
R15228 GNDA_2.n477 GNDA_2.n476 0.028198
R15229 GNDA_2.n472 GNDA_2.n471 0.028198
R15230 GNDA_2.n1009 GNDA_2.n442 0.028198
R15231 GNDA_2.n448 GNDA_2.n441 0.028198
R15232 GNDA_2.n452 GNDA_2.n439 0.028198
R15233 GNDA_2.n993 GNDA_2.n438 0.028198
R15234 GNDA_2.n985 GNDA_2.n436 0.028198
R15235 GNDA_2.n460 GNDA_2.n435 0.028198
R15236 GNDA_2.n464 GNDA_2.n433 0.028198
R15237 GNDA_2.n969 GNDA_2.n432 0.028198
R15238 GNDA_2.n693 GNDA_2.n628 0.028198
R15239 GNDA_2.n634 GNDA_2.n627 0.028198
R15240 GNDA_2.n638 GNDA_2.n625 0.028198
R15241 GNDA_2.n677 GNDA_2.n624 0.028198
R15242 GNDA_2.n669 GNDA_2.n622 0.028198
R15243 GNDA_2.n646 GNDA_2.n621 0.028198
R15244 GNDA_2.n650 GNDA_2.n619 0.028198
R15245 GNDA_2.n653 GNDA_2.n618 0.028198
R15246 GNDA_2.n1030 GNDA_2.n428 0.028198
R15247 GNDA_2.n1029 GNDA_2.n1028 0.028198
R15248 GNDA_2.n1026 GNDA_2.n1025 0.028198
R15249 GNDA_2.n1024 GNDA_2.n418 0.028198
R15250 GNDA_2.n1021 GNDA_2.n413 0.028198
R15251 GNDA_2.n1020 GNDA_2.n1019 0.028198
R15252 GNDA_2.n1017 GNDA_2.n1016 0.028198
R15253 GNDA_2.n1015 GNDA_2.n403 0.028198
R15254 GNDA_2.n221 GNDA_2.n218 0.028198
R15255 GNDA_2.n232 GNDA_2.n231 0.028198
R15256 GNDA_2.n245 GNDA_2.n242 0.028198
R15257 GNDA_2.n256 GNDA_2.n255 0.028198
R15258 GNDA_2.n257 GNDA_2.n256 0.028198
R15259 GNDA_2.n246 GNDA_2.n245 0.028198
R15260 GNDA_2.n233 GNDA_2.n232 0.028198
R15261 GNDA_2.n222 GNDA_2.n221 0.028198
R15262 GNDA_2.n224 GNDA_2.n223 0.0262697
R15263 GNDA_2.n229 GNDA_2.n226 0.0262697
R15264 GNDA_2.n237 GNDA_2.n234 0.0262697
R15265 GNDA_2.n240 GNDA_2.n239 0.0262697
R15266 GNDA_2.n248 GNDA_2.n247 0.0262697
R15267 GNDA_2.n253 GNDA_2.n250 0.0262697
R15268 GNDA_2.n259 GNDA_2.n258 0.0262697
R15269 GNDA_2.n254 GNDA_2.n253 0.0262697
R15270 GNDA_2.n249 GNDA_2.n248 0.0262697
R15271 GNDA_2.n241 GNDA_2.n240 0.0262697
R15272 GNDA_2.n238 GNDA_2.n237 0.0262697
R15273 GNDA_2.n230 GNDA_2.n229 0.0262697
R15274 GNDA_2.n225 GNDA_2.n224 0.0262697
R15275 GNDA_2.n217 GNDA_2.n216 0.0262697
R15276 GNDA_2.n1018 GNDA_2.n409 0.0243392
R15277 GNDA_2.n1023 GNDA_2.n417 0.0243392
R15278 GNDA_2.n1027 GNDA_2.n424 0.0243392
R15279 GNDA_2.n5023 GNDA_2.n4990 0.0243392
R15280 GNDA_2.n5037 GNDA_2.n4993 0.0243392
R15281 GNDA_2.n5053 GNDA_2.n4996 0.0243392
R15282 GNDA_2.n4947 GNDA_2.n4909 0.0243392
R15283 GNDA_2.n4961 GNDA_2.n4912 0.0243392
R15284 GNDA_2.n4977 GNDA_2.n4915 0.0243392
R15285 GNDA_2.n4882 GNDA_2.n4881 0.0243392
R15286 GNDA_2.n4873 GNDA_2.n4872 0.0243392
R15287 GNDA_2.n4864 GNDA_2.n4863 0.0243392
R15288 GNDA_2.n5107 GNDA_2.n4787 0.0243392
R15289 GNDA_2.n5121 GNDA_2.n4790 0.0243392
R15290 GNDA_2.n5137 GNDA_2.n4793 0.0243392
R15291 GNDA_2.n4571 GNDA_2.n4538 0.0243392
R15292 GNDA_2.n4585 GNDA_2.n4541 0.0243392
R15293 GNDA_2.n4601 GNDA_2.n4544 0.0243392
R15294 GNDA_2.n5172 GNDA_2.n4775 0.0243392
R15295 GNDA_2.n5186 GNDA_2.n4778 0.0243392
R15296 GNDA_2.n5202 GNDA_2.n4781 0.0243392
R15297 GNDA_2.n4732 GNDA_2.n151 0.0243392
R15298 GNDA_2.n4746 GNDA_2.n154 0.0243392
R15299 GNDA_2.n4762 GNDA_2.n157 0.0243392
R15300 GNDA_2.n4694 GNDA_2.n4693 0.0243392
R15301 GNDA_2.n4685 GNDA_2.n4684 0.0243392
R15302 GNDA_2.n4676 GNDA_2.n4675 0.0243392
R15303 GNDA_2.n4495 GNDA_2.n191 0.0243392
R15304 GNDA_2.n4509 GNDA_2.n194 0.0243392
R15305 GNDA_2.n4525 GNDA_2.n197 0.0243392
R15306 GNDA_2.n4159 GNDA_2.n1101 0.0243392
R15307 GNDA_2.n4164 GNDA_2.n1109 0.0243392
R15308 GNDA_2.n4168 GNDA_2.n1116 0.0243392
R15309 GNDA_2.n4200 GNDA_2.n4175 0.0243392
R15310 GNDA_2.n4242 GNDA_2.n4178 0.0243392
R15311 GNDA_2.n4188 GNDA_2.n4181 0.0243392
R15312 GNDA_2.n4103 GNDA_2.n4078 0.0243392
R15313 GNDA_2.n4133 GNDA_2.n4081 0.0243392
R15314 GNDA_2.n4091 GNDA_2.n4084 0.0243392
R15315 GNDA_2.n1151 GNDA_2.n1126 0.0243392
R15316 GNDA_2.n4052 GNDA_2.n1129 0.0243392
R15317 GNDA_2.n1139 GNDA_2.n1132 0.0243392
R15318 GNDA_2.n1173 GNDA_2.n1172 0.0243392
R15319 GNDA_2.n1186 GNDA_2.n1185 0.0243392
R15320 GNDA_2.n1197 GNDA_2.n1196 0.0243392
R15321 GNDA_2.n3629 GNDA_2.n3604 0.0243392
R15322 GNDA_2.n3659 GNDA_2.n3607 0.0243392
R15323 GNDA_2.n3617 GNDA_2.n3610 0.0243392
R15324 GNDA_2.n3698 GNDA_2.n3592 0.0243392
R15325 GNDA_2.n3728 GNDA_2.n3595 0.0243392
R15326 GNDA_2.n3686 GNDA_2.n3598 0.0243392
R15327 GNDA_2.n3767 GNDA_2.n3580 0.0243392
R15328 GNDA_2.n3797 GNDA_2.n3583 0.0243392
R15329 GNDA_2.n3755 GNDA_2.n3586 0.0243392
R15330 GNDA_2.n3836 GNDA_2.n3568 0.0243392
R15331 GNDA_2.n3866 GNDA_2.n3571 0.0243392
R15332 GNDA_2.n3824 GNDA_2.n3574 0.0243392
R15333 GNDA_2.n3913 GNDA_2.n3556 0.0243392
R15334 GNDA_2.n3927 GNDA_2.n3559 0.0243392
R15335 GNDA_2.n3943 GNDA_2.n3562 0.0243392
R15336 GNDA_2.n3014 GNDA_2.n3013 0.0243392
R15337 GNDA_2.n3025 GNDA_2.n2987 0.0243392
R15338 GNDA_2.n3044 GNDA_2.n3043 0.0243392
R15339 GNDA_2.n1602 GNDA_2.n1565 0.0243392
R15340 GNDA_2.n1616 GNDA_2.n1568 0.0243392
R15341 GNDA_2.n1632 GNDA_2.n1571 0.0243392
R15342 GNDA_2.n1627 GNDA_2.n1571 0.0243392
R15343 GNDA_2.n1613 GNDA_2.n1568 0.0243392
R15344 GNDA_2.n1597 GNDA_2.n1565 0.0243392
R15345 GNDA_2.n3043 GNDA_2.n3042 0.0243392
R15346 GNDA_2.n3026 GNDA_2.n3025 0.0243392
R15347 GNDA_2.n3013 GNDA_2.n3012 0.0243392
R15348 GNDA_2.n3938 GNDA_2.n3562 0.0243392
R15349 GNDA_2.n3924 GNDA_2.n3559 0.0243392
R15350 GNDA_2.n3908 GNDA_2.n3556 0.0243392
R15351 GNDA_2.n3875 GNDA_2.n3574 0.0243392
R15352 GNDA_2.n3833 GNDA_2.n3571 0.0243392
R15353 GNDA_2.n3851 GNDA_2.n3568 0.0243392
R15354 GNDA_2.n3806 GNDA_2.n3586 0.0243392
R15355 GNDA_2.n3764 GNDA_2.n3583 0.0243392
R15356 GNDA_2.n3782 GNDA_2.n3580 0.0243392
R15357 GNDA_2.n3737 GNDA_2.n3598 0.0243392
R15358 GNDA_2.n3695 GNDA_2.n3595 0.0243392
R15359 GNDA_2.n3713 GNDA_2.n3592 0.0243392
R15360 GNDA_2.n3668 GNDA_2.n3610 0.0243392
R15361 GNDA_2.n3626 GNDA_2.n3607 0.0243392
R15362 GNDA_2.n3644 GNDA_2.n3604 0.0243392
R15363 GNDA_2.n1196 GNDA_2.n1195 0.0243392
R15364 GNDA_2.n1185 GNDA_2.n1184 0.0243392
R15365 GNDA_2.n1172 GNDA_2.n1171 0.0243392
R15366 GNDA_2.n4061 GNDA_2.n1132 0.0243392
R15367 GNDA_2.n1148 GNDA_2.n1129 0.0243392
R15368 GNDA_2.n4037 GNDA_2.n1126 0.0243392
R15369 GNDA_2.n4142 GNDA_2.n4084 0.0243392
R15370 GNDA_2.n4100 GNDA_2.n4081 0.0243392
R15371 GNDA_2.n4118 GNDA_2.n4078 0.0243392
R15372 GNDA_2.n4251 GNDA_2.n4181 0.0243392
R15373 GNDA_2.n4197 GNDA_2.n4178 0.0243392
R15374 GNDA_2.n4227 GNDA_2.n4175 0.0243392
R15375 GNDA_2.n4168 GNDA_2.n1115 0.0243392
R15376 GNDA_2.n4164 GNDA_2.n4163 0.0243392
R15377 GNDA_2.n4159 GNDA_2.n1100 0.0243392
R15378 GNDA_2.n4520 GNDA_2.n197 0.0243392
R15379 GNDA_2.n4506 GNDA_2.n194 0.0243392
R15380 GNDA_2.n4490 GNDA_2.n191 0.0243392
R15381 GNDA_2.n4677 GNDA_2.n4676 0.0243392
R15382 GNDA_2.n4686 GNDA_2.n4685 0.0243392
R15383 GNDA_2.n4695 GNDA_2.n4694 0.0243392
R15384 GNDA_2.n4757 GNDA_2.n157 0.0243392
R15385 GNDA_2.n4743 GNDA_2.n154 0.0243392
R15386 GNDA_2.n4727 GNDA_2.n151 0.0243392
R15387 GNDA_2.n5197 GNDA_2.n4781 0.0243392
R15388 GNDA_2.n5183 GNDA_2.n4778 0.0243392
R15389 GNDA_2.n5167 GNDA_2.n4775 0.0243392
R15390 GNDA_2.n4596 GNDA_2.n4544 0.0243392
R15391 GNDA_2.n4582 GNDA_2.n4541 0.0243392
R15392 GNDA_2.n4566 GNDA_2.n4538 0.0243392
R15393 GNDA_2.n5132 GNDA_2.n4793 0.0243392
R15394 GNDA_2.n5118 GNDA_2.n4790 0.0243392
R15395 GNDA_2.n5102 GNDA_2.n4787 0.0243392
R15396 GNDA_2.n4865 GNDA_2.n4864 0.0243392
R15397 GNDA_2.n4874 GNDA_2.n4873 0.0243392
R15398 GNDA_2.n4883 GNDA_2.n4882 0.0243392
R15399 GNDA_2.n4972 GNDA_2.n4915 0.0243392
R15400 GNDA_2.n4958 GNDA_2.n4912 0.0243392
R15401 GNDA_2.n4942 GNDA_2.n4909 0.0243392
R15402 GNDA_2.n5048 GNDA_2.n4996 0.0243392
R15403 GNDA_2.n5034 GNDA_2.n4993 0.0243392
R15404 GNDA_2.n5018 GNDA_2.n4990 0.0243392
R15405 GNDA_2.n645 GNDA_2.n620 0.0243392
R15406 GNDA_2.n676 GNDA_2.n623 0.0243392
R15407 GNDA_2.n633 GNDA_2.n626 0.0243392
R15408 GNDA_2.n459 GNDA_2.n434 0.0243392
R15409 GNDA_2.n992 GNDA_2.n437 0.0243392
R15410 GNDA_2.n447 GNDA_2.n440 0.0243392
R15411 GNDA_2.n481 GNDA_2.n480 0.0243392
R15412 GNDA_2.n494 GNDA_2.n493 0.0243392
R15413 GNDA_2.n505 GNDA_2.n504 0.0243392
R15414 GNDA_2.n750 GNDA_2.n725 0.0243392
R15415 GNDA_2.n780 GNDA_2.n728 0.0243392
R15416 GNDA_2.n738 GNDA_2.n731 0.0243392
R15417 GNDA_2.n819 GNDA_2.n713 0.0243392
R15418 GNDA_2.n849 GNDA_2.n716 0.0243392
R15419 GNDA_2.n807 GNDA_2.n719 0.0243392
R15420 GNDA_2.n896 GNDA_2.n701 0.0243392
R15421 GNDA_2.n910 GNDA_2.n704 0.0243392
R15422 GNDA_2.n926 GNDA_2.n707 0.0243392
R15423 GNDA_2.n921 GNDA_2.n707 0.0243392
R15424 GNDA_2.n907 GNDA_2.n704 0.0243392
R15425 GNDA_2.n891 GNDA_2.n701 0.0243392
R15426 GNDA_2.n858 GNDA_2.n719 0.0243392
R15427 GNDA_2.n816 GNDA_2.n716 0.0243392
R15428 GNDA_2.n834 GNDA_2.n713 0.0243392
R15429 GNDA_2.n789 GNDA_2.n731 0.0243392
R15430 GNDA_2.n747 GNDA_2.n728 0.0243392
R15431 GNDA_2.n765 GNDA_2.n725 0.0243392
R15432 GNDA_2.n504 GNDA_2.n503 0.0243392
R15433 GNDA_2.n493 GNDA_2.n492 0.0243392
R15434 GNDA_2.n480 GNDA_2.n479 0.0243392
R15435 GNDA_2.n1001 GNDA_2.n440 0.0243392
R15436 GNDA_2.n456 GNDA_2.n437 0.0243392
R15437 GNDA_2.n977 GNDA_2.n434 0.0243392
R15438 GNDA_2.n685 GNDA_2.n626 0.0243392
R15439 GNDA_2.n642 GNDA_2.n623 0.0243392
R15440 GNDA_2.n661 GNDA_2.n620 0.0243392
R15441 GNDA_2.n1027 GNDA_2.n423 0.0243392
R15442 GNDA_2.n1023 GNDA_2.n1022 0.0243392
R15443 GNDA_2.n1018 GNDA_2.n408 0.0243392
R15444 GNDA_2.n564 GNDA_2.n561 0.0217373
R15445 GNDA_2.n5068 GNDA_2.n4901 0.0217373
R15446 GNDA_2.n5069 GNDA_2.n4901 0.0217373
R15447 GNDA_2.n4899 GNDA_2.n4896 0.0217373
R15448 GNDA_2.n4900 GNDA_2.n4896 0.0217373
R15449 GNDA_2.n4894 GNDA_2.n4810 0.0217373
R15450 GNDA_2.n4895 GNDA_2.n4810 0.0217373
R15451 GNDA_2.n5087 GNDA_2.n5084 0.0217373
R15452 GNDA_2.n5088 GNDA_2.n5087 0.0217373
R15453 GNDA_2.n143 GNDA_2.n141 0.0217373
R15454 GNDA_2.n143 GNDA_2.n140 0.0217373
R15455 GNDA_2.n4712 GNDA_2.n174 0.0217373
R15456 GNDA_2.n4713 GNDA_2.n4712 0.0217373
R15457 GNDA_2.n4623 GNDA_2.n177 0.0217373
R15458 GNDA_2.n4623 GNDA_2.n176 0.0217373
R15459 GNDA_2.n5245 GNDA_2.n5244 0.0217373
R15460 GNDA_2.n5248 GNDA_2.n5247 0.0217373
R15461 GNDA_2.n5250 GNDA_2.n136 0.0217373
R15462 GNDA_2.n5221 GNDA_2.n137 0.0217373
R15463 GNDA_2.n5222 GNDA_2.n5221 0.0217373
R15464 GNDA_2.n5243 GNDA_2.n5228 0.0217373
R15465 GNDA_2.n5246 GNDA_2.n5245 0.0217373
R15466 GNDA_2.n359 GNDA_2.n358 0.0217373
R15467 GNDA_2.n5248 GNDA_2.n134 0.0217373
R15468 GNDA_2.n136 GNDA_2.n134 0.0217373
R15469 GNDA_2.n4419 GNDA_2.n4418 0.0217373
R15470 GNDA_2.n4432 GNDA_2.n4428 0.0217373
R15471 GNDA_2.n4437 GNDA_2.n4436 0.0217373
R15472 GNDA_2.n4439 GNDA_2.n317 0.0217373
R15473 GNDA_2.n4442 GNDA_2.n318 0.0217373
R15474 GNDA_2.n4435 GNDA_2.n4428 0.0217373
R15475 GNDA_2.n4438 GNDA_2.n4437 0.0217373
R15476 GNDA_2.n4423 GNDA_2.n319 0.0217373
R15477 GNDA_2.n4427 GNDA_2.n317 0.0217373
R15478 GNDA_2.n4427 GNDA_2.n318 0.0217373
R15479 GNDA_2.n4394 GNDA_2.n339 0.0217373
R15480 GNDA_2.n4376 GNDA_2.n310 0.0217373
R15481 GNDA_2.n311 GNDA_2.n308 0.0217373
R15482 GNDA_2.n4445 GNDA_2.n313 0.0217373
R15483 GNDA_2.n353 GNDA_2.n352 0.0217373
R15484 GNDA_2.n357 GNDA_2.n355 0.0217373
R15485 GNDA_2.n4451 GNDA_2.n309 0.0217373
R15486 GNDA_2.n4450 GNDA_2.n308 0.0217373
R15487 GNDA_2.n4447 GNDA_2.n314 0.0217373
R15488 GNDA_2.n4446 GNDA_2.n4445 0.0217373
R15489 GNDA_2.n365 GNDA_2.n364 0.0217373
R15490 GNDA_2.n362 GNDA_2.n352 0.0217373
R15491 GNDA_2.n358 GNDA_2.n356 0.0217373
R15492 GNDA_2.n4386 GNDA_2.n341 0.0217373
R15493 GNDA_2.n4379 GNDA_2.n4375 0.0217373
R15494 GNDA_2.n4376 GNDA_2.n4375 0.0217373
R15495 GNDA_2.n4390 GNDA_2.n4389 0.0217373
R15496 GNDA_2.n4393 GNDA_2.n4392 0.0217373
R15497 GNDA_2.n4393 GNDA_2.n340 0.0217373
R15498 GNDA_2.n323 GNDA_2.n322 0.0217373
R15499 GNDA_2.n323 GNDA_2.n320 0.0217373
R15500 GNDA_2.n326 GNDA_2.n324 0.0217373
R15501 GNDA_2.n4416 GNDA_2.n326 0.0217373
R15502 GNDA_2.n4415 GNDA_2.n4414 0.0217373
R15503 GNDA_2.n4412 GNDA_2.n330 0.0217373
R15504 GNDA_2.n4388 GNDA_2.n341 0.0217373
R15505 GNDA_2.n4391 GNDA_2.n4390 0.0217373
R15506 GNDA_2.n4396 GNDA_2.n4392 0.0217373
R15507 GNDA_2.n340 GNDA_2.n321 0.0217373
R15508 GNDA_2.n4395 GNDA_2.n4394 0.0217373
R15509 GNDA_2.n4425 GNDA_2.n322 0.0217373
R15510 GNDA_2.n4422 GNDA_2.n320 0.0217373
R15511 GNDA_2.n4424 GNDA_2.n4423 0.0217373
R15512 GNDA_2.n4421 GNDA_2.n324 0.0217373
R15513 GNDA_2.n4417 GNDA_2.n4416 0.0217373
R15514 GNDA_2.n4420 GNDA_2.n4419 0.0217373
R15515 GNDA_2.n4000 GNDA_2.n3978 0.0217373
R15516 GNDA_2.n4414 GNDA_2.n328 0.0217373
R15517 GNDA_2.n330 GNDA_2.n328 0.0217373
R15518 GNDA_2.n3993 GNDA_2.n3980 0.0217373
R15519 GNDA_2.n3997 GNDA_2.n3996 0.0217373
R15520 GNDA_2.n4004 GNDA_2.n4003 0.0217373
R15521 GNDA_2.n4006 GNDA_2.n1247 0.0217373
R15522 GNDA_2.n4009 GNDA_2.n1248 0.0217373
R15523 GNDA_2.n3995 GNDA_2.n3980 0.0217373
R15524 GNDA_2.n3998 GNDA_2.n3997 0.0217373
R15525 GNDA_2.n4002 GNDA_2.n3978 0.0217373
R15526 GNDA_2.n4005 GNDA_2.n4004 0.0217373
R15527 GNDA_2.n4216 GNDA_2.n4206 0.0217373
R15528 GNDA_2.n4026 GNDA_2.n1157 0.0217373
R15529 GNDA_2.n4019 GNDA_2.n1160 0.0217373
R15530 GNDA_2.n4014 GNDA_2.n1244 0.0217373
R15531 GNDA_2.n3975 GNDA_2.n1251 0.0217373
R15532 GNDA_2.n3970 GNDA_2.n1255 0.0217373
R15533 GNDA_2.n3965 GNDA_2.n1259 0.0217373
R15534 GNDA_2.n3961 GNDA_2.n1261 0.0217373
R15535 GNDA_2.n3962 GNDA_2.n1258 0.0217373
R15536 GNDA_2.n3962 GNDA_2.n1259 0.0217373
R15537 GNDA_2.n3967 GNDA_2.n1254 0.0217373
R15538 GNDA_2.n3967 GNDA_2.n1255 0.0217373
R15539 GNDA_2.n3972 GNDA_2.n1250 0.0217373
R15540 GNDA_2.n3972 GNDA_2.n1251 0.0217373
R15541 GNDA_2.n4011 GNDA_2.n1243 0.0217373
R15542 GNDA_2.n4011 GNDA_2.n1244 0.0217373
R15543 GNDA_2.n4016 GNDA_2.n1159 0.0217373
R15544 GNDA_2.n4016 GNDA_2.n1160 0.0217373
R15545 GNDA_2.n4023 GNDA_2.n4021 0.0217373
R15546 GNDA_2.n4021 GNDA_2.n1157 0.0217373
R15547 GNDA_2.n4213 GNDA_2.n4211 0.0217373
R15548 GNDA_2.n4211 GNDA_2.n4206 0.0217373
R15549 GNDA_2.n3977 GNDA_2.n1247 0.0217373
R15550 GNDA_2.n3977 GNDA_2.n1248 0.0217373
R15551 GNDA_2.n3958 GNDA_2.n1262 0.0217373
R15552 GNDA_2.n1263 GNDA_2.n1261 0.0217373
R15553 GNDA_2.n3958 GNDA_2.n3957 0.0217373
R15554 GNDA_2.n2823 GNDA_2.n2668 0.0217373
R15555 GNDA_2.n2826 GNDA_2.n2664 0.0217373
R15556 GNDA_2.n2691 GNDA_2.n2666 0.0217373
R15557 GNDA_2.n2668 GNDA_2.n2667 0.0217373
R15558 GNDA_2.n2661 GNDA_2.n2660 0.0217373
R15559 GNDA_2.n2664 GNDA_2.n2660 0.0217373
R15560 GNDA_2.n3058 GNDA_2.n2975 0.0217373
R15561 GNDA_2.n3384 GNDA_2.n1681 0.0217373
R15562 GNDA_2.n3059 GNDA_2.n2976 0.0217373
R15563 GNDA_2.n2975 GNDA_2.n1679 0.0217373
R15564 GNDA_2.n3385 GNDA_2.n1682 0.0217373
R15565 GNDA_2.n3424 GNDA_2.n1648 0.0217373
R15566 GNDA_2.n3431 GNDA_2.n3429 0.0217373
R15567 GNDA_2.n3427 GNDA_2.n1642 0.0217373
R15568 GNDA_2.n1647 GNDA_2.n1645 0.0217373
R15569 GNDA_2.n3429 GNDA_2.n1643 0.0217373
R15570 GNDA_2.n3428 GNDA_2.n3427 0.0217373
R15571 GNDA_2.n1648 GNDA_2.n1646 0.0217373
R15572 GNDA_2.n298 GNDA_2.n214 0.0217373
R15573 GNDA_2.n4616 GNDA_2.n178 0.0217373
R15574 GNDA_2.n4706 GNDA_2.n175 0.0217373
R15575 GNDA_2.n173 GNDA_2.n172 0.0217373
R15576 GNDA_2.n5217 GNDA_2.n139 0.0217373
R15577 GNDA_2.n5224 GNDA_2.n5223 0.0217373
R15578 GNDA_2.n5083 GNDA_2.n4809 0.0217373
R15579 GNDA_2.n5080 GNDA_2.n5079 0.0217373
R15580 GNDA_2.n5076 GNDA_2.n5075 0.0217373
R15581 GNDA_2.n5072 GNDA_2.n5071 0.0217373
R15582 GNDA_2.n295 GNDA_2.n213 0.0217373
R15583 GNDA_2.n295 GNDA_2.n214 0.0217373
R15584 GNDA_2.n4708 GNDA_2.n177 0.0217373
R15585 GNDA_2.n4705 GNDA_2.n176 0.0217373
R15586 GNDA_2.n4707 GNDA_2.n4706 0.0217373
R15587 GNDA_2.n4710 GNDA_2.n174 0.0217373
R15588 GNDA_2.n4714 GNDA_2.n4713 0.0217373
R15589 GNDA_2.n4711 GNDA_2.n172 0.0217373
R15590 GNDA_2.n5219 GNDA_2.n141 0.0217373
R15591 GNDA_2.n5216 GNDA_2.n140 0.0217373
R15592 GNDA_2.n5218 GNDA_2.n5217 0.0217373
R15593 GNDA_2.n4617 GNDA_2.n4616 0.0217373
R15594 GNDA_2.n5085 GNDA_2.n5084 0.0217373
R15595 GNDA_2.n5089 GNDA_2.n5088 0.0217373
R15596 GNDA_2.n5086 GNDA_2.n4809 0.0217373
R15597 GNDA_2.n4894 GNDA_2.n4811 0.0217373
R15598 GNDA_2.n4895 GNDA_2.n4893 0.0217373
R15599 GNDA_2.n5081 GNDA_2.n5080 0.0217373
R15600 GNDA_2.n4899 GNDA_2.n4897 0.0217373
R15601 GNDA_2.n4900 GNDA_2.n4898 0.0217373
R15602 GNDA_2.n5077 GNDA_2.n5076 0.0217373
R15603 GNDA_2.n5068 GNDA_2.n4902 0.0217373
R15604 GNDA_2.n5069 GNDA_2.n5067 0.0217373
R15605 GNDA_2.n5073 GNDA_2.n5072 0.0217373
R15606 GNDA_2.n5226 GNDA_2.n137 0.0217373
R15607 GNDA_2.n5225 GNDA_2.n5224 0.0217373
R15608 GNDA_2.n398 GNDA_2.n391 0.0217373
R15609 GNDA_2.n399 GNDA_2.n389 0.0217373
R15610 GNDA_2.n1070 GNDA_2.n390 0.0217373
R15611 GNDA_2.n1069 GNDA_2.n389 0.0217373
R15612 GNDA_2.n602 GNDA_2.n566 0.0217373
R15613 GNDA_2.n395 GNDA_2.n393 0.0217373
R15614 GNDA_2.n393 GNDA_2.n391 0.0217373
R15615 GNDA_2.n606 GNDA_2.n605 0.0217373
R15616 GNDA_2.n610 GNDA_2.n565 0.0217373
R15617 GNDA_2.n611 GNDA_2.n610 0.0217373
R15618 GNDA_2.n604 GNDA_2.n566 0.0217373
R15619 GNDA_2.n607 GNDA_2.n606 0.0217373
R15620 GNDA_2.n608 GNDA_2.n565 0.0217373
R15621 GNDA_2.n612 GNDA_2.n611 0.0217373
R15622 GNDA_2.n609 GNDA_2.n561 0.0217373
R15623 GNDA_2.n966 GNDA_2.n465 0.0217373
R15624 GNDA_2.n959 GNDA_2.n468 0.0217373
R15625 GNDA_2.n954 GNDA_2.n552 0.0217373
R15626 GNDA_2.n949 GNDA_2.n556 0.0217373
R15627 GNDA_2.n945 GNDA_2.n558 0.0217373
R15628 GNDA_2.n946 GNDA_2.n555 0.0217373
R15629 GNDA_2.n946 GNDA_2.n556 0.0217373
R15630 GNDA_2.n951 GNDA_2.n551 0.0217373
R15631 GNDA_2.n951 GNDA_2.n552 0.0217373
R15632 GNDA_2.n956 GNDA_2.n467 0.0217373
R15633 GNDA_2.n956 GNDA_2.n468 0.0217373
R15634 GNDA_2.n963 GNDA_2.n961 0.0217373
R15635 GNDA_2.n961 GNDA_2.n465 0.0217373
R15636 GNDA_2.n941 GNDA_2.n559 0.0217373
R15637 GNDA_2.n560 GNDA_2.n558 0.0217373
R15638 GNDA_2.n941 GNDA_2.n940 0.0217373
R15639 GNDA_2.n5243 GNDA_2.n5242 0.0217373
R15640 GNDA_2.n5244 GNDA_2.n5241 0.0217373
R15641 GNDA_2.n5242 GNDA_2.n5240 0.0217373
R15642 GNDA_2.n356 GNDA_2.n354 0.0217373
R15643 GNDA_2.n5251 GNDA_2.n135 0.0217373
R15644 GNDA_2.n5227 GNDA_2.n135 0.0217373
R15645 GNDA_2.n366 GNDA_2.n365 0.0217373
R15646 GNDA_2.n4435 GNDA_2.n4434 0.0217373
R15647 GNDA_2.n4436 GNDA_2.n4433 0.0217373
R15648 GNDA_2.n4434 GNDA_2.n4430 0.0217373
R15649 GNDA_2.n4441 GNDA_2.n4440 0.0217373
R15650 GNDA_2.n314 GNDA_2.n312 0.0217373
R15651 GNDA_2.n4440 GNDA_2.n316 0.0217373
R15652 GNDA_2.n4454 GNDA_2.n309 0.0217373
R15653 GNDA_2.n4452 GNDA_2.n311 0.0217373
R15654 GNDA_2.n4448 GNDA_2.n313 0.0217373
R15655 GNDA_2.n363 GNDA_2.n353 0.0217373
R15656 GNDA_2.n360 GNDA_2.n355 0.0217373
R15657 GNDA_2.n4453 GNDA_2.n4452 0.0217373
R15658 GNDA_2.n4455 GNDA_2.n4454 0.0217373
R15659 GNDA_2.n4449 GNDA_2.n4448 0.0217373
R15660 GNDA_2.n4444 GNDA_2.n312 0.0217373
R15661 GNDA_2.n363 GNDA_2.n315 0.0217373
R15662 GNDA_2.n367 GNDA_2.n366 0.0217373
R15663 GNDA_2.n361 GNDA_2.n360 0.0217373
R15664 GNDA_2.n4388 GNDA_2.n342 0.0217373
R15665 GNDA_2.n4381 GNDA_2.n4380 0.0217373
R15666 GNDA_2.n4380 GNDA_2.n4377 0.0217373
R15667 GNDA_2.n4389 GNDA_2.n4387 0.0217373
R15668 GNDA_2.n4002 GNDA_2.n3979 0.0217373
R15669 GNDA_2.n4411 GNDA_2.n327 0.0217373
R15670 GNDA_2.n329 GNDA_2.n327 0.0217373
R15671 GNDA_2.n3995 GNDA_2.n3981 0.0217373
R15672 GNDA_2.n3996 GNDA_2.n3994 0.0217373
R15673 GNDA_2.n4003 GNDA_2.n4001 0.0217373
R15674 GNDA_2.n4001 GNDA_2.n3999 0.0217373
R15675 GNDA_2.n3959 GNDA_2.n1263 0.0217373
R15676 GNDA_2.n3964 GNDA_2.n3963 0.0217373
R15677 GNDA_2.n3969 GNDA_2.n3968 0.0217373
R15678 GNDA_2.n3974 GNDA_2.n3973 0.0217373
R15679 GNDA_2.n4008 GNDA_2.n4007 0.0217373
R15680 GNDA_2.n4013 GNDA_2.n4012 0.0217373
R15681 GNDA_2.n4018 GNDA_2.n4017 0.0217373
R15682 GNDA_2.n4025 GNDA_2.n4024 0.0217373
R15683 GNDA_2.n4310 GNDA_2.n1087 0.0217373
R15684 GNDA_2.n4215 GNDA_2.n4214 0.0217373
R15685 GNDA_2.n3963 GNDA_2.n1257 0.0217373
R15686 GNDA_2.n3968 GNDA_2.n1253 0.0217373
R15687 GNDA_2.n3973 GNDA_2.n1249 0.0217373
R15688 GNDA_2.n4012 GNDA_2.n1242 0.0217373
R15689 GNDA_2.n4017 GNDA_2.n1158 0.0217373
R15690 GNDA_2.n4024 GNDA_2.n4022 0.0217373
R15691 GNDA_2.n1090 GNDA_2.n1087 0.0217373
R15692 GNDA_2.n4214 GNDA_2.n4212 0.0217373
R15693 GNDA_2.n4007 GNDA_2.n1246 0.0217373
R15694 GNDA_2.n3960 GNDA_2.n1262 0.0217373
R15695 GNDA_2.n2667 GNDA_2.n2665 0.0217373
R15696 GNDA_2.n2824 GNDA_2.n2666 0.0217373
R15697 GNDA_2.n2825 GNDA_2.n2824 0.0217373
R15698 GNDA_2.n2692 GNDA_2.n2665 0.0217373
R15699 GNDA_2.n2827 GNDA_2.n2662 0.0217373
R15700 GNDA_2.n1682 GNDA_2.n1680 0.0217373
R15701 GNDA_2.n2663 GNDA_2.n2662 0.0217373
R15702 GNDA_2.n3062 GNDA_2.n2976 0.0217373
R15703 GNDA_2.n3060 GNDA_2.n3058 0.0217373
R15704 GNDA_2.n3386 GNDA_2.n1681 0.0217373
R15705 GNDA_2.n3061 GNDA_2.n3060 0.0217373
R15706 GNDA_2.n3063 GNDA_2.n3062 0.0217373
R15707 GNDA_2.n3387 GNDA_2.n3386 0.0217373
R15708 GNDA_2.n3383 GNDA_2.n1680 0.0217373
R15709 GNDA_2.n1646 GNDA_2.n1644 0.0217373
R15710 GNDA_2.n1643 GNDA_2.n1641 0.0217373
R15711 GNDA_2.n3432 GNDA_2.n1642 0.0217373
R15712 GNDA_2.n3425 GNDA_2.n1645 0.0217373
R15713 GNDA_2.n3433 GNDA_2.n3432 0.0217373
R15714 GNDA_2.n3426 GNDA_2.n3425 0.0217373
R15715 GNDA_2.n297 GNDA_2.n296 0.0217373
R15716 GNDA_2.n296 GNDA_2.n212 0.0217373
R15717 GNDA_2.n1073 GNDA_2.n390 0.0217373
R15718 GNDA_2.n1071 GNDA_2.n399 0.0217373
R15719 GNDA_2.n1072 GNDA_2.n1071 0.0217373
R15720 GNDA_2.n1074 GNDA_2.n1073 0.0217373
R15721 GNDA_2.n604 GNDA_2.n567 0.0217373
R15722 GNDA_2.n397 GNDA_2.n396 0.0217373
R15723 GNDA_2.n396 GNDA_2.n394 0.0217373
R15724 GNDA_2.n605 GNDA_2.n603 0.0217373
R15725 GNDA_2.n943 GNDA_2.n560 0.0217373
R15726 GNDA_2.n948 GNDA_2.n947 0.0217373
R15727 GNDA_2.n953 GNDA_2.n952 0.0217373
R15728 GNDA_2.n958 GNDA_2.n957 0.0217373
R15729 GNDA_2.n965 GNDA_2.n964 0.0217373
R15730 GNDA_2.n947 GNDA_2.n554 0.0217373
R15731 GNDA_2.n952 GNDA_2.n550 0.0217373
R15732 GNDA_2.n957 GNDA_2.n466 0.0217373
R15733 GNDA_2.n964 GNDA_2.n962 0.0217373
R15734 GNDA_2.n944 GNDA_2.n559 0.0217373
R15735 GNDA_2.n943 GNDA_2.n942 0.0217373
R15736 GNDA_2.n183 GNDA_2.n181 0.0181756
R15737 GNDA_2.n183 GNDA_2.n179 0.0181756
R15738 GNDA_2.n4307 GNDA_2.n4306 0.0181756
R15739 GNDA_2.n4309 GNDA_2.n1088 0.0181756
R15740 GNDA_2.n4307 GNDA_2.n1086 0.0181756
R15741 GNDA_2.n1088 GNDA_2.n1086 0.0181756
R15742 GNDA_2.n4618 GNDA_2.n181 0.0181756
R15743 GNDA_2.n4615 GNDA_2.n179 0.0181756
R15744 GNDA_2.n3953 GNDA_2.n3888 0.0107812
R15745 GNDA_2.n3888 GNDA_2.n3819 0.0107812
R15746 GNDA_2.n3819 GNDA_2.n3750 0.0107812
R15747 GNDA_2.n3750 GNDA_2.n3681 0.0107812
R15748 GNDA_2.n3681 GNDA_2.n1122 0.0107812
R15749 GNDA_2.n4074 GNDA_2.n1122 0.0107812
R15750 GNDA_2.n4155 GNDA_2.n4074 0.0107812
R15751 GNDA_2.n4265 GNDA_2.n4155 0.0107812
R15752 GNDA_2.n4265 GNDA_2.n4264 0.0107812
R15753 GNDA_2.n4535 GNDA_2.n187 0.0107812
R15754 GNDA_2.n4611 GNDA_2.n4535 0.0107812
R15755 GNDA_2.n4611 GNDA_2.n147 0.0107812
R15756 GNDA_2.n4772 GNDA_2.n147 0.0107812
R15757 GNDA_2.n5212 GNDA_2.n4772 0.0107812
R15758 GNDA_2.n5212 GNDA_2.n5147 0.0107812
R15759 GNDA_2.n5147 GNDA_2.n4796 0.0107812
R15760 GNDA_2.n4987 GNDA_2.n4796 0.0107812
R15761 GNDA_2.n5063 GNDA_2.n4987 0.0107812
R15762 GNDA_2.n936 GNDA_2.n698 0.0107812
R15763 GNDA_2.n936 GNDA_2.n871 0.0107812
R15764 GNDA_2.n871 GNDA_2.n802 0.0107812
R15765 GNDA_2.n802 GNDA_2.n430 0.0107812
R15766 GNDA_2.n1014 GNDA_2.n430 0.0107812
R15767 GNDA_2.n1031 GNDA_2.n1014 0.0107812
R15768 GNDA_2.n3512 GNDA_2.n1429 0.00182188
R15769 GNDA_2.n3441 GNDA_2.n1495 0.00182188
R15770 GNDA_2.n3547 GNDA_2.n1347 0.00182188
R15771 GNDA_2.n3443 GNDA_2.n1429 0.00166081
R15772 GNDA_2.n1413 GNDA_2.n1365 0.00166081
R15773 GNDA_2.n3444 GNDA_2.n1365 0.00166081
R15774 GNDA_2.n1414 GNDA_2.n1366 0.00166081
R15775 GNDA_2.n3445 GNDA_2.n1366 0.00166081
R15776 GNDA_2.n1415 GNDA_2.n1367 0.00166081
R15777 GNDA_2.n3446 GNDA_2.n1367 0.00166081
R15778 GNDA_2.n1416 GNDA_2.n1368 0.00166081
R15779 GNDA_2.n3447 GNDA_2.n1368 0.00166081
R15780 GNDA_2.n1417 GNDA_2.n1369 0.00166081
R15781 GNDA_2.n3448 GNDA_2.n1369 0.00166081
R15782 GNDA_2.n1418 GNDA_2.n1370 0.00166081
R15783 GNDA_2.n3449 GNDA_2.n1370 0.00166081
R15784 GNDA_2.n1419 GNDA_2.n1371 0.00166081
R15785 GNDA_2.n3450 GNDA_2.n1371 0.00166081
R15786 GNDA_2.n1420 GNDA_2.n1372 0.00166081
R15787 GNDA_2.n3451 GNDA_2.n1372 0.00166081
R15788 GNDA_2.n1421 GNDA_2.n1373 0.00166081
R15789 GNDA_2.n3452 GNDA_2.n1373 0.00166081
R15790 GNDA_2.n1422 GNDA_2.n1374 0.00166081
R15791 GNDA_2.n3453 GNDA_2.n1374 0.00166081
R15792 GNDA_2.n1423 GNDA_2.n1375 0.00166081
R15793 GNDA_2.n3454 GNDA_2.n1375 0.00166081
R15794 GNDA_2.n1424 GNDA_2.n1376 0.00166081
R15795 GNDA_2.n3455 GNDA_2.n1376 0.00166081
R15796 GNDA_2.n1425 GNDA_2.n1377 0.00166081
R15797 GNDA_2.n3456 GNDA_2.n1377 0.00166081
R15798 GNDA_2.n1426 GNDA_2.n1378 0.00166081
R15799 GNDA_2.n3457 GNDA_2.n1378 0.00166081
R15800 GNDA_2.n1427 GNDA_2.n1379 0.00166081
R15801 GNDA_2.n3458 GNDA_2.n1379 0.00166081
R15802 GNDA_2.n3492 GNDA_2.n3491 0.00166081
R15803 GNDA_2.n3509 GNDA_2.n1380 0.00166081
R15804 GNDA_2.n1496 GNDA_2.n1495 0.00166081
R15805 GNDA_2.n1479 GNDA_2.n1431 0.00166081
R15806 GNDA_2.n1497 GNDA_2.n1431 0.00166081
R15807 GNDA_2.n1480 GNDA_2.n1432 0.00166081
R15808 GNDA_2.n1498 GNDA_2.n1432 0.00166081
R15809 GNDA_2.n1481 GNDA_2.n1433 0.00166081
R15810 GNDA_2.n1499 GNDA_2.n1433 0.00166081
R15811 GNDA_2.n1482 GNDA_2.n1434 0.00166081
R15812 GNDA_2.n1500 GNDA_2.n1434 0.00166081
R15813 GNDA_2.n1483 GNDA_2.n1435 0.00166081
R15814 GNDA_2.n1501 GNDA_2.n1435 0.00166081
R15815 GNDA_2.n1484 GNDA_2.n1436 0.00166081
R15816 GNDA_2.n1502 GNDA_2.n1436 0.00166081
R15817 GNDA_2.n1485 GNDA_2.n1437 0.00166081
R15818 GNDA_2.n1503 GNDA_2.n1437 0.00166081
R15819 GNDA_2.n1486 GNDA_2.n1438 0.00166081
R15820 GNDA_2.n1504 GNDA_2.n1438 0.00166081
R15821 GNDA_2.n1487 GNDA_2.n1439 0.00166081
R15822 GNDA_2.n1505 GNDA_2.n1439 0.00166081
R15823 GNDA_2.n1488 GNDA_2.n1440 0.00166081
R15824 GNDA_2.n1506 GNDA_2.n1440 0.00166081
R15825 GNDA_2.n1489 GNDA_2.n1441 0.00166081
R15826 GNDA_2.n1507 GNDA_2.n1441 0.00166081
R15827 GNDA_2.n1490 GNDA_2.n1442 0.00166081
R15828 GNDA_2.n1508 GNDA_2.n1442 0.00166081
R15829 GNDA_2.n1491 GNDA_2.n1443 0.00166081
R15830 GNDA_2.n1509 GNDA_2.n1443 0.00166081
R15831 GNDA_2.n1492 GNDA_2.n1444 0.00166081
R15832 GNDA_2.n1510 GNDA_2.n1444 0.00166081
R15833 GNDA_2.n1493 GNDA_2.n1445 0.00166081
R15834 GNDA_2.n1511 GNDA_2.n1445 0.00166081
R15835 GNDA_2.n1545 GNDA_2.n1544 0.00166081
R15836 GNDA_2.n3438 GNDA_2.n1446 0.00166081
R15837 GNDA_2.n1561 GNDA_2.n1494 0.00166081
R15838 GNDA_2.n1514 GNDA_2.n1513 0.00166081
R15839 GNDA_2.n1560 GNDA_2.n1478 0.00166081
R15840 GNDA_2.n1516 GNDA_2.n1515 0.00166081
R15841 GNDA_2.n1559 GNDA_2.n1477 0.00166081
R15842 GNDA_2.n1518 GNDA_2.n1517 0.00166081
R15843 GNDA_2.n1558 GNDA_2.n1476 0.00166081
R15844 GNDA_2.n1520 GNDA_2.n1519 0.00166081
R15845 GNDA_2.n1557 GNDA_2.n1475 0.00166081
R15846 GNDA_2.n1522 GNDA_2.n1521 0.00166081
R15847 GNDA_2.n1556 GNDA_2.n1474 0.00166081
R15848 GNDA_2.n1524 GNDA_2.n1523 0.00166081
R15849 GNDA_2.n1555 GNDA_2.n1473 0.00166081
R15850 GNDA_2.n1526 GNDA_2.n1525 0.00166081
R15851 GNDA_2.n1554 GNDA_2.n1472 0.00166081
R15852 GNDA_2.n1528 GNDA_2.n1527 0.00166081
R15853 GNDA_2.n1553 GNDA_2.n1471 0.00166081
R15854 GNDA_2.n1530 GNDA_2.n1529 0.00166081
R15855 GNDA_2.n1552 GNDA_2.n1470 0.00166081
R15856 GNDA_2.n1532 GNDA_2.n1531 0.00166081
R15857 GNDA_2.n1551 GNDA_2.n1469 0.00166081
R15858 GNDA_2.n1534 GNDA_2.n1533 0.00166081
R15859 GNDA_2.n1550 GNDA_2.n1468 0.00166081
R15860 GNDA_2.n1536 GNDA_2.n1535 0.00166081
R15861 GNDA_2.n1549 GNDA_2.n1467 0.00166081
R15862 GNDA_2.n1538 GNDA_2.n1537 0.00166081
R15863 GNDA_2.n1548 GNDA_2.n1466 0.00166081
R15864 GNDA_2.n1540 GNDA_2.n1539 0.00166081
R15865 GNDA_2.n1547 GNDA_2.n1465 0.00166081
R15866 GNDA_2.n1542 GNDA_2.n1541 0.00166081
R15867 GNDA_2.n1546 GNDA_2.n1464 0.00166081
R15868 GNDA_2.n3440 GNDA_2.n1543 0.00166081
R15869 GNDA_2.n3439 GNDA_2.n1463 0.00166081
R15870 GNDA_2.n3442 GNDA_2.n1430 0.00166081
R15871 GNDA_2.n3508 GNDA_2.n1428 0.00166081
R15872 GNDA_2.n3461 GNDA_2.n3460 0.00166081
R15873 GNDA_2.n3507 GNDA_2.n1412 0.00166081
R15874 GNDA_2.n3463 GNDA_2.n3462 0.00166081
R15875 GNDA_2.n3506 GNDA_2.n1411 0.00166081
R15876 GNDA_2.n3465 GNDA_2.n3464 0.00166081
R15877 GNDA_2.n3505 GNDA_2.n1410 0.00166081
R15878 GNDA_2.n3467 GNDA_2.n3466 0.00166081
R15879 GNDA_2.n3504 GNDA_2.n1409 0.00166081
R15880 GNDA_2.n3469 GNDA_2.n3468 0.00166081
R15881 GNDA_2.n3503 GNDA_2.n1408 0.00166081
R15882 GNDA_2.n3471 GNDA_2.n3470 0.00166081
R15883 GNDA_2.n3502 GNDA_2.n1407 0.00166081
R15884 GNDA_2.n3473 GNDA_2.n3472 0.00166081
R15885 GNDA_2.n3501 GNDA_2.n1406 0.00166081
R15886 GNDA_2.n3475 GNDA_2.n3474 0.00166081
R15887 GNDA_2.n3500 GNDA_2.n1405 0.00166081
R15888 GNDA_2.n3477 GNDA_2.n3476 0.00166081
R15889 GNDA_2.n3499 GNDA_2.n1404 0.00166081
R15890 GNDA_2.n3479 GNDA_2.n3478 0.00166081
R15891 GNDA_2.n3498 GNDA_2.n1403 0.00166081
R15892 GNDA_2.n3481 GNDA_2.n3480 0.00166081
R15893 GNDA_2.n3497 GNDA_2.n1402 0.00166081
R15894 GNDA_2.n3483 GNDA_2.n3482 0.00166081
R15895 GNDA_2.n3496 GNDA_2.n1401 0.00166081
R15896 GNDA_2.n3485 GNDA_2.n3484 0.00166081
R15897 GNDA_2.n3495 GNDA_2.n1400 0.00166081
R15898 GNDA_2.n3487 GNDA_2.n3486 0.00166081
R15899 GNDA_2.n3494 GNDA_2.n1399 0.00166081
R15900 GNDA_2.n3489 GNDA_2.n3488 0.00166081
R15901 GNDA_2.n3493 GNDA_2.n1398 0.00166081
R15902 GNDA_2.n3511 GNDA_2.n3490 0.00166081
R15903 GNDA_2.n3510 GNDA_2.n1397 0.00166081
R15904 GNDA_2.n3513 GNDA_2.n1364 0.00166081
R15905 GNDA_2.n3530 GNDA_2.n1283 0.00166081
R15906 GNDA_2.n3550 GNDA_2.n3548 0.00166081
R15907 GNDA_2.n3549 GNDA_2.n1282 0.00166081
R15908 GNDA_2.n3532 GNDA_2.n1285 0.00166081
R15909 GNDA_2.n1315 GNDA_2.n1281 0.00166081
R15910 GNDA_2.n3533 GNDA_2.n1286 0.00166081
R15911 GNDA_2.n1314 GNDA_2.n1280 0.00166081
R15912 GNDA_2.n3534 GNDA_2.n1287 0.00166081
R15913 GNDA_2.n1313 GNDA_2.n1279 0.00166081
R15914 GNDA_2.n3535 GNDA_2.n1288 0.00166081
R15915 GNDA_2.n1312 GNDA_2.n1278 0.00166081
R15916 GNDA_2.n3536 GNDA_2.n1289 0.00166081
R15917 GNDA_2.n1311 GNDA_2.n1277 0.00166081
R15918 GNDA_2.n3537 GNDA_2.n1290 0.00166081
R15919 GNDA_2.n1310 GNDA_2.n1276 0.00166081
R15920 GNDA_2.n3538 GNDA_2.n1291 0.00166081
R15921 GNDA_2.n1309 GNDA_2.n1275 0.00166081
R15922 GNDA_2.n3539 GNDA_2.n1292 0.00166081
R15923 GNDA_2.n1308 GNDA_2.n1274 0.00166081
R15924 GNDA_2.n3540 GNDA_2.n1293 0.00166081
R15925 GNDA_2.n1307 GNDA_2.n1273 0.00166081
R15926 GNDA_2.n3541 GNDA_2.n1294 0.00166081
R15927 GNDA_2.n1306 GNDA_2.n1272 0.00166081
R15928 GNDA_2.n3542 GNDA_2.n1295 0.00166081
R15929 GNDA_2.n1305 GNDA_2.n1271 0.00166081
R15930 GNDA_2.n3543 GNDA_2.n1296 0.00166081
R15931 GNDA_2.n1304 GNDA_2.n1270 0.00166081
R15932 GNDA_2.n3544 GNDA_2.n1297 0.00166081
R15933 GNDA_2.n1303 GNDA_2.n1269 0.00166081
R15934 GNDA_2.n3545 GNDA_2.n1298 0.00166081
R15935 GNDA_2.n1302 GNDA_2.n1268 0.00166081
R15936 GNDA_2.n3546 GNDA_2.n1299 0.00166081
R15937 GNDA_2.n1301 GNDA_2.n1267 0.00166081
R15938 GNDA_2.n3552 GNDA_2.n1300 0.00166081
R15939 GNDA_2.n1561 GNDA_2.n1512 0.00166081
R15940 GNDA_2.n1511 GNDA_2.n1447 0.00166081
R15941 GNDA_2.n1510 GNDA_2.n1448 0.00166081
R15942 GNDA_2.n1509 GNDA_2.n1449 0.00166081
R15943 GNDA_2.n1508 GNDA_2.n1450 0.00166081
R15944 GNDA_2.n1507 GNDA_2.n1451 0.00166081
R15945 GNDA_2.n1506 GNDA_2.n1452 0.00166081
R15946 GNDA_2.n1505 GNDA_2.n1453 0.00166081
R15947 GNDA_2.n1504 GNDA_2.n1454 0.00166081
R15948 GNDA_2.n1503 GNDA_2.n1455 0.00166081
R15949 GNDA_2.n1502 GNDA_2.n1456 0.00166081
R15950 GNDA_2.n1501 GNDA_2.n1457 0.00166081
R15951 GNDA_2.n1500 GNDA_2.n1458 0.00166081
R15952 GNDA_2.n1499 GNDA_2.n1459 0.00166081
R15953 GNDA_2.n1498 GNDA_2.n1460 0.00166081
R15954 GNDA_2.n1497 GNDA_2.n1461 0.00166081
R15955 GNDA_2.n1496 GNDA_2.n1462 0.00166081
R15956 GNDA_2.n1544 GNDA_2.n1447 0.00166081
R15957 GNDA_2.n1493 GNDA_2.n1448 0.00166081
R15958 GNDA_2.n1492 GNDA_2.n1449 0.00166081
R15959 GNDA_2.n1491 GNDA_2.n1450 0.00166081
R15960 GNDA_2.n1490 GNDA_2.n1451 0.00166081
R15961 GNDA_2.n1489 GNDA_2.n1452 0.00166081
R15962 GNDA_2.n1488 GNDA_2.n1453 0.00166081
R15963 GNDA_2.n1487 GNDA_2.n1454 0.00166081
R15964 GNDA_2.n1486 GNDA_2.n1455 0.00166081
R15965 GNDA_2.n1485 GNDA_2.n1456 0.00166081
R15966 GNDA_2.n1484 GNDA_2.n1457 0.00166081
R15967 GNDA_2.n1483 GNDA_2.n1458 0.00166081
R15968 GNDA_2.n1482 GNDA_2.n1459 0.00166081
R15969 GNDA_2.n1481 GNDA_2.n1460 0.00166081
R15970 GNDA_2.n1480 GNDA_2.n1461 0.00166081
R15971 GNDA_2.n1479 GNDA_2.n1462 0.00166081
R15972 GNDA_2.n1513 GNDA_2.n1494 0.00166081
R15973 GNDA_2.n1560 GNDA_2.n1514 0.00166081
R15974 GNDA_2.n1515 GNDA_2.n1478 0.00166081
R15975 GNDA_2.n1559 GNDA_2.n1516 0.00166081
R15976 GNDA_2.n1517 GNDA_2.n1477 0.00166081
R15977 GNDA_2.n1558 GNDA_2.n1518 0.00166081
R15978 GNDA_2.n1519 GNDA_2.n1476 0.00166081
R15979 GNDA_2.n1557 GNDA_2.n1520 0.00166081
R15980 GNDA_2.n1521 GNDA_2.n1475 0.00166081
R15981 GNDA_2.n1556 GNDA_2.n1522 0.00166081
R15982 GNDA_2.n1523 GNDA_2.n1474 0.00166081
R15983 GNDA_2.n1555 GNDA_2.n1524 0.00166081
R15984 GNDA_2.n1525 GNDA_2.n1473 0.00166081
R15985 GNDA_2.n1554 GNDA_2.n1526 0.00166081
R15986 GNDA_2.n1527 GNDA_2.n1472 0.00166081
R15987 GNDA_2.n1553 GNDA_2.n1528 0.00166081
R15988 GNDA_2.n1529 GNDA_2.n1471 0.00166081
R15989 GNDA_2.n1552 GNDA_2.n1530 0.00166081
R15990 GNDA_2.n1531 GNDA_2.n1470 0.00166081
R15991 GNDA_2.n1551 GNDA_2.n1532 0.00166081
R15992 GNDA_2.n1533 GNDA_2.n1469 0.00166081
R15993 GNDA_2.n1550 GNDA_2.n1534 0.00166081
R15994 GNDA_2.n1535 GNDA_2.n1468 0.00166081
R15995 GNDA_2.n1549 GNDA_2.n1536 0.00166081
R15996 GNDA_2.n1537 GNDA_2.n1467 0.00166081
R15997 GNDA_2.n1548 GNDA_2.n1538 0.00166081
R15998 GNDA_2.n1539 GNDA_2.n1466 0.00166081
R15999 GNDA_2.n1547 GNDA_2.n1540 0.00166081
R16000 GNDA_2.n1541 GNDA_2.n1465 0.00166081
R16001 GNDA_2.n1546 GNDA_2.n1542 0.00166081
R16002 GNDA_2.n1543 GNDA_2.n1464 0.00166081
R16003 GNDA_2.n3440 GNDA_2.n3439 0.00166081
R16004 GNDA_2.n1463 GNDA_2.n1430 0.00166081
R16005 GNDA_2.n1545 GNDA_2.n1446 0.00166081
R16006 GNDA_2.n3508 GNDA_2.n3459 0.00166081
R16007 GNDA_2.n3458 GNDA_2.n1381 0.00166081
R16008 GNDA_2.n3457 GNDA_2.n1382 0.00166081
R16009 GNDA_2.n3456 GNDA_2.n1383 0.00166081
R16010 GNDA_2.n3455 GNDA_2.n1384 0.00166081
R16011 GNDA_2.n3454 GNDA_2.n1385 0.00166081
R16012 GNDA_2.n3453 GNDA_2.n1386 0.00166081
R16013 GNDA_2.n3452 GNDA_2.n1387 0.00166081
R16014 GNDA_2.n3451 GNDA_2.n1388 0.00166081
R16015 GNDA_2.n3450 GNDA_2.n1389 0.00166081
R16016 GNDA_2.n3449 GNDA_2.n1390 0.00166081
R16017 GNDA_2.n3448 GNDA_2.n1391 0.00166081
R16018 GNDA_2.n3447 GNDA_2.n1392 0.00166081
R16019 GNDA_2.n3446 GNDA_2.n1393 0.00166081
R16020 GNDA_2.n3445 GNDA_2.n1394 0.00166081
R16021 GNDA_2.n3444 GNDA_2.n1395 0.00166081
R16022 GNDA_2.n3443 GNDA_2.n1396 0.00166081
R16023 GNDA_2.n3491 GNDA_2.n1381 0.00166081
R16024 GNDA_2.n1427 GNDA_2.n1382 0.00166081
R16025 GNDA_2.n1426 GNDA_2.n1383 0.00166081
R16026 GNDA_2.n1425 GNDA_2.n1384 0.00166081
R16027 GNDA_2.n1424 GNDA_2.n1385 0.00166081
R16028 GNDA_2.n1423 GNDA_2.n1386 0.00166081
R16029 GNDA_2.n1422 GNDA_2.n1387 0.00166081
R16030 GNDA_2.n1421 GNDA_2.n1388 0.00166081
R16031 GNDA_2.n1420 GNDA_2.n1389 0.00166081
R16032 GNDA_2.n1419 GNDA_2.n1390 0.00166081
R16033 GNDA_2.n1418 GNDA_2.n1391 0.00166081
R16034 GNDA_2.n1417 GNDA_2.n1392 0.00166081
R16035 GNDA_2.n1416 GNDA_2.n1393 0.00166081
R16036 GNDA_2.n1415 GNDA_2.n1394 0.00166081
R16037 GNDA_2.n1414 GNDA_2.n1395 0.00166081
R16038 GNDA_2.n1413 GNDA_2.n1396 0.00166081
R16039 GNDA_2.n3460 GNDA_2.n1428 0.00166081
R16040 GNDA_2.n3507 GNDA_2.n3461 0.00166081
R16041 GNDA_2.n3462 GNDA_2.n1412 0.00166081
R16042 GNDA_2.n3506 GNDA_2.n3463 0.00166081
R16043 GNDA_2.n3464 GNDA_2.n1411 0.00166081
R16044 GNDA_2.n3505 GNDA_2.n3465 0.00166081
R16045 GNDA_2.n3466 GNDA_2.n1410 0.00166081
R16046 GNDA_2.n3504 GNDA_2.n3467 0.00166081
R16047 GNDA_2.n3468 GNDA_2.n1409 0.00166081
R16048 GNDA_2.n3503 GNDA_2.n3469 0.00166081
R16049 GNDA_2.n3470 GNDA_2.n1408 0.00166081
R16050 GNDA_2.n3502 GNDA_2.n3471 0.00166081
R16051 GNDA_2.n3472 GNDA_2.n1407 0.00166081
R16052 GNDA_2.n3501 GNDA_2.n3473 0.00166081
R16053 GNDA_2.n3474 GNDA_2.n1406 0.00166081
R16054 GNDA_2.n3500 GNDA_2.n3475 0.00166081
R16055 GNDA_2.n3476 GNDA_2.n1405 0.00166081
R16056 GNDA_2.n3499 GNDA_2.n3477 0.00166081
R16057 GNDA_2.n3478 GNDA_2.n1404 0.00166081
R16058 GNDA_2.n3498 GNDA_2.n3479 0.00166081
R16059 GNDA_2.n3480 GNDA_2.n1403 0.00166081
R16060 GNDA_2.n3497 GNDA_2.n3481 0.00166081
R16061 GNDA_2.n3482 GNDA_2.n1402 0.00166081
R16062 GNDA_2.n3496 GNDA_2.n3483 0.00166081
R16063 GNDA_2.n3484 GNDA_2.n1401 0.00166081
R16064 GNDA_2.n3495 GNDA_2.n3485 0.00166081
R16065 GNDA_2.n3486 GNDA_2.n1400 0.00166081
R16066 GNDA_2.n3494 GNDA_2.n3487 0.00166081
R16067 GNDA_2.n3488 GNDA_2.n1399 0.00166081
R16068 GNDA_2.n3493 GNDA_2.n3489 0.00166081
R16069 GNDA_2.n3490 GNDA_2.n1398 0.00166081
R16070 GNDA_2.n3511 GNDA_2.n3510 0.00166081
R16071 GNDA_2.n1397 GNDA_2.n1364 0.00166081
R16072 GNDA_2.n3492 GNDA_2.n1380 0.00166081
R16073 GNDA_2.n3551 GNDA_2.n3531 0.00166081
R16074 GNDA_2.n3514 GNDA_2.n1347 0.00166081
R16075 GNDA_2.n1348 GNDA_2.n1316 0.00166081
R16076 GNDA_2.n3515 GNDA_2.n1346 0.00166081
R16077 GNDA_2.n1349 GNDA_2.n1317 0.00166081
R16078 GNDA_2.n3516 GNDA_2.n1345 0.00166081
R16079 GNDA_2.n1350 GNDA_2.n1318 0.00166081
R16080 GNDA_2.n3517 GNDA_2.n1344 0.00166081
R16081 GNDA_2.n1351 GNDA_2.n1319 0.00166081
R16082 GNDA_2.n3518 GNDA_2.n1343 0.00166081
R16083 GNDA_2.n1352 GNDA_2.n1320 0.00166081
R16084 GNDA_2.n3519 GNDA_2.n1342 0.00166081
R16085 GNDA_2.n1353 GNDA_2.n1321 0.00166081
R16086 GNDA_2.n3520 GNDA_2.n1341 0.00166081
R16087 GNDA_2.n1354 GNDA_2.n1322 0.00166081
R16088 GNDA_2.n3521 GNDA_2.n1340 0.00166081
R16089 GNDA_2.n1355 GNDA_2.n1323 0.00166081
R16090 GNDA_2.n3522 GNDA_2.n1339 0.00166081
R16091 GNDA_2.n1356 GNDA_2.n1324 0.00166081
R16092 GNDA_2.n3523 GNDA_2.n1338 0.00166081
R16093 GNDA_2.n1357 GNDA_2.n1325 0.00166081
R16094 GNDA_2.n3524 GNDA_2.n1337 0.00166081
R16095 GNDA_2.n1358 GNDA_2.n1326 0.00166081
R16096 GNDA_2.n3525 GNDA_2.n1336 0.00166081
R16097 GNDA_2.n1359 GNDA_2.n1327 0.00166081
R16098 GNDA_2.n3526 GNDA_2.n1335 0.00166081
R16099 GNDA_2.n1360 GNDA_2.n1328 0.00166081
R16100 GNDA_2.n3527 GNDA_2.n1334 0.00166081
R16101 GNDA_2.n1361 GNDA_2.n1329 0.00166081
R16102 GNDA_2.n3528 GNDA_2.n1333 0.00166081
R16103 GNDA_2.n1362 GNDA_2.n1330 0.00166081
R16104 GNDA_2.n3529 GNDA_2.n1332 0.00166081
R16105 GNDA_2.n1331 GNDA_2.n1284 0.00166081
R16106 GNDA_2.n3529 GNDA_2.n1331 0.00166081
R16107 GNDA_2.n3528 GNDA_2.n1330 0.00166081
R16108 GNDA_2.n3527 GNDA_2.n1329 0.00166081
R16109 GNDA_2.n3526 GNDA_2.n1328 0.00166081
R16110 GNDA_2.n3525 GNDA_2.n1327 0.00166081
R16111 GNDA_2.n3524 GNDA_2.n1326 0.00166081
R16112 GNDA_2.n3523 GNDA_2.n1325 0.00166081
R16113 GNDA_2.n3522 GNDA_2.n1324 0.00166081
R16114 GNDA_2.n3521 GNDA_2.n1323 0.00166081
R16115 GNDA_2.n3520 GNDA_2.n1322 0.00166081
R16116 GNDA_2.n3519 GNDA_2.n1321 0.00166081
R16117 GNDA_2.n3518 GNDA_2.n1320 0.00166081
R16118 GNDA_2.n3517 GNDA_2.n1319 0.00166081
R16119 GNDA_2.n3516 GNDA_2.n1318 0.00166081
R16120 GNDA_2.n3515 GNDA_2.n1317 0.00166081
R16121 GNDA_2.n3514 GNDA_2.n1316 0.00166081
R16122 GNDA_2.n3547 GNDA_2.n3531 0.00166081
R16123 GNDA_2.n1363 GNDA_2.n1283 0.00166081
R16124 GNDA_2.n1362 GNDA_2.n1332 0.00166081
R16125 GNDA_2.n1361 GNDA_2.n1333 0.00166081
R16126 GNDA_2.n1360 GNDA_2.n1334 0.00166081
R16127 GNDA_2.n1359 GNDA_2.n1335 0.00166081
R16128 GNDA_2.n1358 GNDA_2.n1336 0.00166081
R16129 GNDA_2.n1357 GNDA_2.n1337 0.00166081
R16130 GNDA_2.n1356 GNDA_2.n1338 0.00166081
R16131 GNDA_2.n1355 GNDA_2.n1339 0.00166081
R16132 GNDA_2.n1354 GNDA_2.n1340 0.00166081
R16133 GNDA_2.n1353 GNDA_2.n1341 0.00166081
R16134 GNDA_2.n1352 GNDA_2.n1342 0.00166081
R16135 GNDA_2.n1351 GNDA_2.n1343 0.00166081
R16136 GNDA_2.n1350 GNDA_2.n1344 0.00166081
R16137 GNDA_2.n1349 GNDA_2.n1345 0.00166081
R16138 GNDA_2.n1348 GNDA_2.n1346 0.00166081
R16139 GNDA_2.n3548 GNDA_2.n1363 0.00166081
R16140 GNDA_2.n3553 GNDA_2.n1284 0.00166081
R16141 GNDA_2.n3550 GNDA_2.n3549 0.00166081
R16142 GNDA_2.n3532 GNDA_2.n1282 0.00166081
R16143 GNDA_2.n1315 GNDA_2.n1285 0.00166081
R16144 GNDA_2.n3533 GNDA_2.n1281 0.00166081
R16145 GNDA_2.n1314 GNDA_2.n1286 0.00166081
R16146 GNDA_2.n3534 GNDA_2.n1280 0.00166081
R16147 GNDA_2.n1313 GNDA_2.n1287 0.00166081
R16148 GNDA_2.n3535 GNDA_2.n1279 0.00166081
R16149 GNDA_2.n1312 GNDA_2.n1288 0.00166081
R16150 GNDA_2.n3536 GNDA_2.n1278 0.00166081
R16151 GNDA_2.n1311 GNDA_2.n1289 0.00166081
R16152 GNDA_2.n3537 GNDA_2.n1277 0.00166081
R16153 GNDA_2.n1310 GNDA_2.n1290 0.00166081
R16154 GNDA_2.n3538 GNDA_2.n1276 0.00166081
R16155 GNDA_2.n1309 GNDA_2.n1291 0.00166081
R16156 GNDA_2.n3539 GNDA_2.n1275 0.00166081
R16157 GNDA_2.n1308 GNDA_2.n1292 0.00166081
R16158 GNDA_2.n3540 GNDA_2.n1274 0.00166081
R16159 GNDA_2.n1307 GNDA_2.n1293 0.00166081
R16160 GNDA_2.n3541 GNDA_2.n1273 0.00166081
R16161 GNDA_2.n1306 GNDA_2.n1294 0.00166081
R16162 GNDA_2.n3542 GNDA_2.n1272 0.00166081
R16163 GNDA_2.n1305 GNDA_2.n1295 0.00166081
R16164 GNDA_2.n3543 GNDA_2.n1271 0.00166081
R16165 GNDA_2.n1304 GNDA_2.n1296 0.00166081
R16166 GNDA_2.n3544 GNDA_2.n1270 0.00166081
R16167 GNDA_2.n1303 GNDA_2.n1297 0.00166081
R16168 GNDA_2.n3545 GNDA_2.n1269 0.00166081
R16169 GNDA_2.n1302 GNDA_2.n1298 0.00166081
R16170 GNDA_2.n3546 GNDA_2.n1268 0.00166081
R16171 GNDA_2.n1301 GNDA_2.n1299 0.00166081
R16172 GNDA_2.n1300 GNDA_2.n1267 0.00166081
R16173 two_stage_opamp_dummy_magic_29_0.Vb2.n2 two_stage_opamp_dummy_magic_29_0.Vb2.t22 752.422
R16174 two_stage_opamp_dummy_magic_29_0.Vb2.n0 two_stage_opamp_dummy_magic_29_0.Vb2.t15 752.422
R16175 two_stage_opamp_dummy_magic_29_0.Vb2.n2 two_stage_opamp_dummy_magic_29_0.Vb2.t28 752.234
R16176 two_stage_opamp_dummy_magic_29_0.Vb2.n2 two_stage_opamp_dummy_magic_29_0.Vb2.t25 752.234
R16177 two_stage_opamp_dummy_magic_29_0.Vb2.n3 two_stage_opamp_dummy_magic_29_0.Vb2.t32 752.234
R16178 two_stage_opamp_dummy_magic_29_0.Vb2.n3 two_stage_opamp_dummy_magic_29_0.Vb2.t18 752.234
R16179 two_stage_opamp_dummy_magic_29_0.Vb2.n3 two_stage_opamp_dummy_magic_29_0.Vb2.t20 752.234
R16180 two_stage_opamp_dummy_magic_29_0.Vb2.n3 two_stage_opamp_dummy_magic_29_0.Vb2.t24 752.234
R16181 two_stage_opamp_dummy_magic_29_0.Vb2.n4 two_stage_opamp_dummy_magic_29_0.Vb2.t21 752.234
R16182 two_stage_opamp_dummy_magic_29_0.Vb2.n4 two_stage_opamp_dummy_magic_29_0.Vb2.t26 752.234
R16183 two_stage_opamp_dummy_magic_29_0.Vb2.n4 two_stage_opamp_dummy_magic_29_0.Vb2.t11 752.234
R16184 two_stage_opamp_dummy_magic_29_0.Vb2.n5 two_stage_opamp_dummy_magic_29_0.Vb2.t31 752.234
R16185 two_stage_opamp_dummy_magic_29_0.Vb2.n5 two_stage_opamp_dummy_magic_29_0.Vb2.t27 752.234
R16186 two_stage_opamp_dummy_magic_29_0.Vb2.n1 two_stage_opamp_dummy_magic_29_0.Vb2.t12 752.234
R16187 two_stage_opamp_dummy_magic_29_0.Vb2.n1 two_stage_opamp_dummy_magic_29_0.Vb2.t14 752.234
R16188 two_stage_opamp_dummy_magic_29_0.Vb2.n1 two_stage_opamp_dummy_magic_29_0.Vb2.t16 752.234
R16189 two_stage_opamp_dummy_magic_29_0.Vb2.n1 two_stage_opamp_dummy_magic_29_0.Vb2.t19 752.234
R16190 two_stage_opamp_dummy_magic_29_0.Vb2.n0 two_stage_opamp_dummy_magic_29_0.Vb2.t23 752.234
R16191 two_stage_opamp_dummy_magic_29_0.Vb2.n0 two_stage_opamp_dummy_magic_29_0.Vb2.t29 752.234
R16192 two_stage_opamp_dummy_magic_29_0.Vb2.n0 two_stage_opamp_dummy_magic_29_0.Vb2.t13 752.234
R16193 two_stage_opamp_dummy_magic_29_0.Vb2.n17 two_stage_opamp_dummy_magic_29_0.Vb2.t17 746.673
R16194 two_stage_opamp_dummy_magic_29_0.Vb2.n14 two_stage_opamp_dummy_magic_29_0.Vb2.t8 745.726
R16195 two_stage_opamp_dummy_magic_29_0.Vb2.n16 two_stage_opamp_dummy_magic_29_0.Vb2.t30 587.551
R16196 two_stage_opamp_dummy_magic_29_0.Vb2.n8 two_stage_opamp_dummy_magic_29_0.Vb2.n6 140.546
R16197 two_stage_opamp_dummy_magic_29_0.Vb2.n12 two_stage_opamp_dummy_magic_29_0.Vb2.n11 139.297
R16198 two_stage_opamp_dummy_magic_29_0.Vb2.n10 two_stage_opamp_dummy_magic_29_0.Vb2.n9 139.297
R16199 two_stage_opamp_dummy_magic_29_0.Vb2.n8 two_stage_opamp_dummy_magic_29_0.Vb2.n7 139.297
R16200 two_stage_opamp_dummy_magic_29_0.Vb2.n14 two_stage_opamp_dummy_magic_29_0.Vb2.n13 67.0547
R16201 bgr_11_0.VB2_CUR_BIAS two_stage_opamp_dummy_magic_29_0.Vb2.n18 41.0474
R16202 two_stage_opamp_dummy_magic_29_0.Vb2.n11 two_stage_opamp_dummy_magic_29_0.Vb2.t3 24.0005
R16203 two_stage_opamp_dummy_magic_29_0.Vb2.n11 two_stage_opamp_dummy_magic_29_0.Vb2.t7 24.0005
R16204 two_stage_opamp_dummy_magic_29_0.Vb2.n9 two_stage_opamp_dummy_magic_29_0.Vb2.t4 24.0005
R16205 two_stage_opamp_dummy_magic_29_0.Vb2.n9 two_stage_opamp_dummy_magic_29_0.Vb2.t6 24.0005
R16206 two_stage_opamp_dummy_magic_29_0.Vb2.n7 two_stage_opamp_dummy_magic_29_0.Vb2.t0 24.0005
R16207 two_stage_opamp_dummy_magic_29_0.Vb2.n7 two_stage_opamp_dummy_magic_29_0.Vb2.t5 24.0005
R16208 two_stage_opamp_dummy_magic_29_0.Vb2.n6 two_stage_opamp_dummy_magic_29_0.Vb2.t1 24.0005
R16209 two_stage_opamp_dummy_magic_29_0.Vb2.n6 two_stage_opamp_dummy_magic_29_0.Vb2.t2 24.0005
R16210 bgr_11_0.VB2_CUR_BIAS two_stage_opamp_dummy_magic_29_0.Vb2.n12 21.5317
R16211 two_stage_opamp_dummy_magic_29_0.Vb2.n15 two_stage_opamp_dummy_magic_29_0.Vb2.n4 13.5005
R16212 two_stage_opamp_dummy_magic_29_0.Vb2.n18 two_stage_opamp_dummy_magic_29_0.Vb2.n5 12.5005
R16213 two_stage_opamp_dummy_magic_29_0.Vb2.n13 two_stage_opamp_dummy_magic_29_0.Vb2.t9 11.2576
R16214 two_stage_opamp_dummy_magic_29_0.Vb2.n13 two_stage_opamp_dummy_magic_29_0.Vb2.t10 11.2576
R16215 two_stage_opamp_dummy_magic_29_0.Vb2.n10 two_stage_opamp_dummy_magic_29_0.Vb2.n8 6.21925
R16216 two_stage_opamp_dummy_magic_29_0.Vb2.n15 two_stage_opamp_dummy_magic_29_0.Vb2.n14 4.5005
R16217 two_stage_opamp_dummy_magic_29_0.Vb2.n17 two_stage_opamp_dummy_magic_29_0.Vb2.n16 3.58175
R16218 two_stage_opamp_dummy_magic_29_0.Vb2.n16 two_stage_opamp_dummy_magic_29_0.Vb2.n15 1.48488
R16219 two_stage_opamp_dummy_magic_29_0.Vb2.n12 two_stage_opamp_dummy_magic_29_0.Vb2.n10 1.2505
R16220 two_stage_opamp_dummy_magic_29_0.Vb2.n18 two_stage_opamp_dummy_magic_29_0.Vb2.n17 1.12238
R16221 two_stage_opamp_dummy_magic_29_0.Vb2.n4 two_stage_opamp_dummy_magic_29_0.Vb2.n3 0.7505
R16222 two_stage_opamp_dummy_magic_29_0.Vb2.n3 two_stage_opamp_dummy_magic_29_0.Vb2.n2 0.7505
R16223 two_stage_opamp_dummy_magic_29_0.Vb2.n1 two_stage_opamp_dummy_magic_29_0.Vb2.n0 0.7505
R16224 two_stage_opamp_dummy_magic_29_0.Vb2.n5 two_stage_opamp_dummy_magic_29_0.Vb2.n1 0.7505
R16225 two_stage_opamp_dummy_magic_29_0.Y.n53 two_stage_opamp_dummy_magic_29_0.Y.t34 1172.87
R16226 two_stage_opamp_dummy_magic_29_0.Y.n49 two_stage_opamp_dummy_magic_29_0.Y.t25 1172.87
R16227 two_stage_opamp_dummy_magic_29_0.Y.n53 two_stage_opamp_dummy_magic_29_0.Y.t26 996.134
R16228 two_stage_opamp_dummy_magic_29_0.Y.n54 two_stage_opamp_dummy_magic_29_0.Y.t44 996.134
R16229 two_stage_opamp_dummy_magic_29_0.Y.n55 two_stage_opamp_dummy_magic_29_0.Y.t29 996.134
R16230 two_stage_opamp_dummy_magic_29_0.Y.n56 two_stage_opamp_dummy_magic_29_0.Y.t46 996.134
R16231 two_stage_opamp_dummy_magic_29_0.Y.n52 two_stage_opamp_dummy_magic_29_0.Y.t32 996.134
R16232 two_stage_opamp_dummy_magic_29_0.Y.n51 two_stage_opamp_dummy_magic_29_0.Y.t38 996.134
R16233 two_stage_opamp_dummy_magic_29_0.Y.n50 two_stage_opamp_dummy_magic_29_0.Y.t51 996.134
R16234 two_stage_opamp_dummy_magic_29_0.Y.n49 two_stage_opamp_dummy_magic_29_0.Y.t41 996.134
R16235 two_stage_opamp_dummy_magic_29_0.Y.n71 two_stage_opamp_dummy_magic_29_0.Y.t30 690.867
R16236 two_stage_opamp_dummy_magic_29_0.Y.n64 two_stage_opamp_dummy_magic_29_0.Y.t49 690.867
R16237 two_stage_opamp_dummy_magic_29_0.Y.n80 two_stage_opamp_dummy_magic_29_0.Y.t33 530.201
R16238 two_stage_opamp_dummy_magic_29_0.Y.n73 two_stage_opamp_dummy_magic_29_0.Y.t52 530.201
R16239 two_stage_opamp_dummy_magic_29_0.Y.n71 two_stage_opamp_dummy_magic_29_0.Y.t50 514.134
R16240 two_stage_opamp_dummy_magic_29_0.Y.n64 two_stage_opamp_dummy_magic_29_0.Y.t37 514.134
R16241 two_stage_opamp_dummy_magic_29_0.Y.n65 two_stage_opamp_dummy_magic_29_0.Y.t47 514.134
R16242 two_stage_opamp_dummy_magic_29_0.Y.n66 two_stage_opamp_dummy_magic_29_0.Y.t35 514.134
R16243 two_stage_opamp_dummy_magic_29_0.Y.n67 two_stage_opamp_dummy_magic_29_0.Y.t28 514.134
R16244 two_stage_opamp_dummy_magic_29_0.Y.n68 two_stage_opamp_dummy_magic_29_0.Y.t43 514.134
R16245 two_stage_opamp_dummy_magic_29_0.Y.n69 two_stage_opamp_dummy_magic_29_0.Y.t54 514.134
R16246 two_stage_opamp_dummy_magic_29_0.Y.n70 two_stage_opamp_dummy_magic_29_0.Y.t40 514.134
R16247 two_stage_opamp_dummy_magic_29_0.Y.n80 two_stage_opamp_dummy_magic_29_0.Y.t53 353.467
R16248 two_stage_opamp_dummy_magic_29_0.Y.n79 two_stage_opamp_dummy_magic_29_0.Y.t42 353.467
R16249 two_stage_opamp_dummy_magic_29_0.Y.n78 two_stage_opamp_dummy_magic_29_0.Y.t27 353.467
R16250 two_stage_opamp_dummy_magic_29_0.Y.n77 two_stage_opamp_dummy_magic_29_0.Y.t45 353.467
R16251 two_stage_opamp_dummy_magic_29_0.Y.n76 two_stage_opamp_dummy_magic_29_0.Y.t31 353.467
R16252 two_stage_opamp_dummy_magic_29_0.Y.n75 two_stage_opamp_dummy_magic_29_0.Y.t36 353.467
R16253 two_stage_opamp_dummy_magic_29_0.Y.n74 two_stage_opamp_dummy_magic_29_0.Y.t48 353.467
R16254 two_stage_opamp_dummy_magic_29_0.Y.n73 two_stage_opamp_dummy_magic_29_0.Y.t39 353.467
R16255 two_stage_opamp_dummy_magic_29_0.Y.n52 two_stage_opamp_dummy_magic_29_0.Y.n51 176.733
R16256 two_stage_opamp_dummy_magic_29_0.Y.n51 two_stage_opamp_dummy_magic_29_0.Y.n50 176.733
R16257 two_stage_opamp_dummy_magic_29_0.Y.n50 two_stage_opamp_dummy_magic_29_0.Y.n49 176.733
R16258 two_stage_opamp_dummy_magic_29_0.Y.n54 two_stage_opamp_dummy_magic_29_0.Y.n53 176.733
R16259 two_stage_opamp_dummy_magic_29_0.Y.n55 two_stage_opamp_dummy_magic_29_0.Y.n54 176.733
R16260 two_stage_opamp_dummy_magic_29_0.Y.n56 two_stage_opamp_dummy_magic_29_0.Y.n55 176.733
R16261 two_stage_opamp_dummy_magic_29_0.Y.n79 two_stage_opamp_dummy_magic_29_0.Y.n78 176.733
R16262 two_stage_opamp_dummy_magic_29_0.Y.n78 two_stage_opamp_dummy_magic_29_0.Y.n77 176.733
R16263 two_stage_opamp_dummy_magic_29_0.Y.n77 two_stage_opamp_dummy_magic_29_0.Y.n76 176.733
R16264 two_stage_opamp_dummy_magic_29_0.Y.n76 two_stage_opamp_dummy_magic_29_0.Y.n75 176.733
R16265 two_stage_opamp_dummy_magic_29_0.Y.n75 two_stage_opamp_dummy_magic_29_0.Y.n74 176.733
R16266 two_stage_opamp_dummy_magic_29_0.Y.n74 two_stage_opamp_dummy_magic_29_0.Y.n73 176.733
R16267 two_stage_opamp_dummy_magic_29_0.Y.n70 two_stage_opamp_dummy_magic_29_0.Y.n69 176.733
R16268 two_stage_opamp_dummy_magic_29_0.Y.n69 two_stage_opamp_dummy_magic_29_0.Y.n68 176.733
R16269 two_stage_opamp_dummy_magic_29_0.Y.n68 two_stage_opamp_dummy_magic_29_0.Y.n67 176.733
R16270 two_stage_opamp_dummy_magic_29_0.Y.n67 two_stage_opamp_dummy_magic_29_0.Y.n66 176.733
R16271 two_stage_opamp_dummy_magic_29_0.Y.n66 two_stage_opamp_dummy_magic_29_0.Y.n65 176.733
R16272 two_stage_opamp_dummy_magic_29_0.Y.n65 two_stage_opamp_dummy_magic_29_0.Y.n64 176.733
R16273 two_stage_opamp_dummy_magic_29_0.Y.n82 two_stage_opamp_dummy_magic_29_0.Y.n81 165.472
R16274 two_stage_opamp_dummy_magic_29_0.Y.n82 two_stage_opamp_dummy_magic_29_0.Y.n72 165.472
R16275 two_stage_opamp_dummy_magic_29_0.Y.n59 two_stage_opamp_dummy_magic_29_0.Y.n58 152
R16276 two_stage_opamp_dummy_magic_29_0.Y.n60 two_stage_opamp_dummy_magic_29_0.Y.n59 131.571
R16277 two_stage_opamp_dummy_magic_29_0.Y.n59 two_stage_opamp_dummy_magic_29_0.Y.n57 124.517
R16278 two_stage_opamp_dummy_magic_29_0.Y.n84 two_stage_opamp_dummy_magic_29_0.Y.n82 74.5372
R16279 two_stage_opamp_dummy_magic_29_0.Y.n110 two_stage_opamp_dummy_magic_29_0.Y.n109 66.0338
R16280 two_stage_opamp_dummy_magic_29_0.Y.n94 two_stage_opamp_dummy_magic_29_0.Y.n93 66.0338
R16281 two_stage_opamp_dummy_magic_29_0.Y.n97 two_stage_opamp_dummy_magic_29_0.Y.n96 66.0338
R16282 two_stage_opamp_dummy_magic_29_0.Y.n100 two_stage_opamp_dummy_magic_29_0.Y.n99 66.0338
R16283 two_stage_opamp_dummy_magic_29_0.Y.n104 two_stage_opamp_dummy_magic_29_0.Y.n103 66.0338
R16284 two_stage_opamp_dummy_magic_29_0.Y.n107 two_stage_opamp_dummy_magic_29_0.Y.n106 66.0338
R16285 two_stage_opamp_dummy_magic_29_0.Y.n8 two_stage_opamp_dummy_magic_29_0.Y.n6 54.7984
R16286 two_stage_opamp_dummy_magic_29_0.Y.n8 two_stage_opamp_dummy_magic_29_0.Y.n7 54.4547
R16287 two_stage_opamp_dummy_magic_29_0.Y.n10 two_stage_opamp_dummy_magic_29_0.Y.n9 54.4547
R16288 two_stage_opamp_dummy_magic_29_0.Y.n12 two_stage_opamp_dummy_magic_29_0.Y.n11 54.4547
R16289 two_stage_opamp_dummy_magic_29_0.Y.n14 two_stage_opamp_dummy_magic_29_0.Y.n13 54.4547
R16290 two_stage_opamp_dummy_magic_29_0.Y.n16 two_stage_opamp_dummy_magic_29_0.Y.n15 54.4547
R16291 two_stage_opamp_dummy_magic_29_0.Y.n43 two_stage_opamp_dummy_magic_29_0.Y.t2 41.0384
R16292 two_stage_opamp_dummy_magic_29_0.Y.n57 two_stage_opamp_dummy_magic_29_0.Y.n52 40.1672
R16293 two_stage_opamp_dummy_magic_29_0.Y.n57 two_stage_opamp_dummy_magic_29_0.Y.n56 40.1672
R16294 two_stage_opamp_dummy_magic_29_0.Y.n81 two_stage_opamp_dummy_magic_29_0.Y.n79 40.1672
R16295 two_stage_opamp_dummy_magic_29_0.Y.n81 two_stage_opamp_dummy_magic_29_0.Y.n80 40.1672
R16296 two_stage_opamp_dummy_magic_29_0.Y.n72 two_stage_opamp_dummy_magic_29_0.Y.n70 40.1672
R16297 two_stage_opamp_dummy_magic_29_0.Y.n72 two_stage_opamp_dummy_magic_29_0.Y.n71 40.1672
R16298 two_stage_opamp_dummy_magic_29_0.Y.n61 two_stage_opamp_dummy_magic_29_0.Y.n60 16.3217
R16299 two_stage_opamp_dummy_magic_29_0.Y.n6 two_stage_opamp_dummy_magic_29_0.Y.t5 16.0005
R16300 two_stage_opamp_dummy_magic_29_0.Y.n6 two_stage_opamp_dummy_magic_29_0.Y.t4 16.0005
R16301 two_stage_opamp_dummy_magic_29_0.Y.n7 two_stage_opamp_dummy_magic_29_0.Y.t1 16.0005
R16302 two_stage_opamp_dummy_magic_29_0.Y.n7 two_stage_opamp_dummy_magic_29_0.Y.t6 16.0005
R16303 two_stage_opamp_dummy_magic_29_0.Y.n9 two_stage_opamp_dummy_magic_29_0.Y.t7 16.0005
R16304 two_stage_opamp_dummy_magic_29_0.Y.n9 two_stage_opamp_dummy_magic_29_0.Y.t12 16.0005
R16305 two_stage_opamp_dummy_magic_29_0.Y.n11 two_stage_opamp_dummy_magic_29_0.Y.t10 16.0005
R16306 two_stage_opamp_dummy_magic_29_0.Y.n11 two_stage_opamp_dummy_magic_29_0.Y.t8 16.0005
R16307 two_stage_opamp_dummy_magic_29_0.Y.n13 two_stage_opamp_dummy_magic_29_0.Y.t23 16.0005
R16308 two_stage_opamp_dummy_magic_29_0.Y.n13 two_stage_opamp_dummy_magic_29_0.Y.t11 16.0005
R16309 two_stage_opamp_dummy_magic_29_0.Y.n15 two_stage_opamp_dummy_magic_29_0.Y.t3 16.0005
R16310 two_stage_opamp_dummy_magic_29_0.Y.n15 two_stage_opamp_dummy_magic_29_0.Y.t9 16.0005
R16311 two_stage_opamp_dummy_magic_29_0.Y.n58 two_stage_opamp_dummy_magic_29_0.Y.n48 12.8005
R16312 two_stage_opamp_dummy_magic_29_0.Y.n109 two_stage_opamp_dummy_magic_29_0.Y.t24 11.2576
R16313 two_stage_opamp_dummy_magic_29_0.Y.n109 two_stage_opamp_dummy_magic_29_0.Y.t17 11.2576
R16314 two_stage_opamp_dummy_magic_29_0.Y.n93 two_stage_opamp_dummy_magic_29_0.Y.t13 11.2576
R16315 two_stage_opamp_dummy_magic_29_0.Y.n93 two_stage_opamp_dummy_magic_29_0.Y.t0 11.2576
R16316 two_stage_opamp_dummy_magic_29_0.Y.n96 two_stage_opamp_dummy_magic_29_0.Y.t19 11.2576
R16317 two_stage_opamp_dummy_magic_29_0.Y.n96 two_stage_opamp_dummy_magic_29_0.Y.t21 11.2576
R16318 two_stage_opamp_dummy_magic_29_0.Y.n99 two_stage_opamp_dummy_magic_29_0.Y.t16 11.2576
R16319 two_stage_opamp_dummy_magic_29_0.Y.n99 two_stage_opamp_dummy_magic_29_0.Y.t14 11.2576
R16320 two_stage_opamp_dummy_magic_29_0.Y.n103 two_stage_opamp_dummy_magic_29_0.Y.t20 11.2576
R16321 two_stage_opamp_dummy_magic_29_0.Y.n103 two_stage_opamp_dummy_magic_29_0.Y.t18 11.2576
R16322 two_stage_opamp_dummy_magic_29_0.Y.n106 two_stage_opamp_dummy_magic_29_0.Y.t22 11.2576
R16323 two_stage_opamp_dummy_magic_29_0.Y.n106 two_stage_opamp_dummy_magic_29_0.Y.t15 11.2576
R16324 two_stage_opamp_dummy_magic_29_0.Y.n17 two_stage_opamp_dummy_magic_29_0.Y.n16 11.1099
R16325 two_stage_opamp_dummy_magic_29_0.Y.n58 two_stage_opamp_dummy_magic_29_0.Y.n46 9.36264
R16326 two_stage_opamp_dummy_magic_29_0.Y.n48 two_stage_opamp_dummy_magic_29_0.Y.n47 9.3005
R16327 two_stage_opamp_dummy_magic_29_0.Y.n119 two_stage_opamp_dummy_magic_29_0.Y.n25 5.78175
R16328 two_stage_opamp_dummy_magic_29_0.Y.n98 two_stage_opamp_dummy_magic_29_0.Y.n94 5.66717
R16329 two_stage_opamp_dummy_magic_29_0.Y.n95 two_stage_opamp_dummy_magic_29_0.Y.n94 5.66717
R16330 two_stage_opamp_dummy_magic_29_0.Y.n110 two_stage_opamp_dummy_magic_29_0.Y.n108 5.66717
R16331 two_stage_opamp_dummy_magic_29_0.Y.n18 two_stage_opamp_dummy_magic_29_0.Y.n17 5.46373
R16332 two_stage_opamp_dummy_magic_29_0.Y.n19 two_stage_opamp_dummy_magic_29_0.Y.n5 5.438
R16333 two_stage_opamp_dummy_magic_29_0.Y.n21 two_stage_opamp_dummy_magic_29_0.Y.n4 5.438
R16334 two_stage_opamp_dummy_magic_29_0.Y.n125 two_stage_opamp_dummy_magic_29_0.Y.n1 5.438
R16335 two_stage_opamp_dummy_magic_29_0.Y.n121 two_stage_opamp_dummy_magic_29_0.Y.n25 5.438
R16336 two_stage_opamp_dummy_magic_29_0.Y.n60 two_stage_opamp_dummy_magic_29_0.Y.n48 5.33141
R16337 two_stage_opamp_dummy_magic_29_0.Y.n98 two_stage_opamp_dummy_magic_29_0.Y.n97 5.29217
R16338 two_stage_opamp_dummy_magic_29_0.Y.n97 two_stage_opamp_dummy_magic_29_0.Y.n95 5.29217
R16339 two_stage_opamp_dummy_magic_29_0.Y.n101 two_stage_opamp_dummy_magic_29_0.Y.n100 5.29217
R16340 two_stage_opamp_dummy_magic_29_0.Y.n100 two_stage_opamp_dummy_magic_29_0.Y.n92 5.29217
R16341 two_stage_opamp_dummy_magic_29_0.Y.n104 two_stage_opamp_dummy_magic_29_0.Y.n102 5.29217
R16342 two_stage_opamp_dummy_magic_29_0.Y.n105 two_stage_opamp_dummy_magic_29_0.Y.n104 5.29217
R16343 two_stage_opamp_dummy_magic_29_0.Y.n107 two_stage_opamp_dummy_magic_29_0.Y.n91 5.29217
R16344 two_stage_opamp_dummy_magic_29_0.Y.n108 two_stage_opamp_dummy_magic_29_0.Y.n107 5.29217
R16345 two_stage_opamp_dummy_magic_29_0.Y.n111 two_stage_opamp_dummy_magic_29_0.Y.n110 5.29217
R16346 two_stage_opamp_dummy_magic_29_0.Y.n117 two_stage_opamp_dummy_magic_29_0.Y.n28 4.5005
R16347 two_stage_opamp_dummy_magic_29_0.Y.n117 two_stage_opamp_dummy_magic_29_0.Y.n30 4.5005
R16348 two_stage_opamp_dummy_magic_29_0.Y.n117 two_stage_opamp_dummy_magic_29_0.Y.n27 4.5005
R16349 two_stage_opamp_dummy_magic_29_0.Y.n117 two_stage_opamp_dummy_magic_29_0.Y.n116 4.5005
R16350 two_stage_opamp_dummy_magic_29_0.Y.n34 two_stage_opamp_dummy_magic_29_0.Y.n32 4.5005
R16351 two_stage_opamp_dummy_magic_29_0.Y.n83 two_stage_opamp_dummy_magic_29_0.Y.n36 4.5005
R16352 two_stage_opamp_dummy_magic_29_0.Y.n85 two_stage_opamp_dummy_magic_29_0.Y.n84 4.5005
R16353 two_stage_opamp_dummy_magic_29_0.Y.n84 two_stage_opamp_dummy_magic_29_0.Y.n83 4.5005
R16354 two_stage_opamp_dummy_magic_29_0.Y.n62 two_stage_opamp_dummy_magic_29_0.Y.n61 4.5005
R16355 two_stage_opamp_dummy_magic_29_0.Y.n40 two_stage_opamp_dummy_magic_29_0.Y.n39 4.5005
R16356 two_stage_opamp_dummy_magic_29_0.Y.n112 two_stage_opamp_dummy_magic_29_0.Y.n111 2.35543
R16357 two_stage_opamp_dummy_magic_29_0.Y.n41 two_stage_opamp_dummy_magic_29_0.Y.n38 2.26187
R16358 two_stage_opamp_dummy_magic_29_0.Y.n42 two_stage_opamp_dummy_magic_29_0.Y.n41 2.26187
R16359 two_stage_opamp_dummy_magic_29_0.Y.n112 two_stage_opamp_dummy_magic_29_0.Y.n29 2.24654
R16360 two_stage_opamp_dummy_magic_29_0.Y.n89 two_stage_opamp_dummy_magic_29_0.Y.n88 2.24654
R16361 two_stage_opamp_dummy_magic_29_0.Y.n34 two_stage_opamp_dummy_magic_29_0.Y.n33 2.24063
R16362 two_stage_opamp_dummy_magic_29_0.Y.n34 two_stage_opamp_dummy_magic_29_0.Y.n31 2.24063
R16363 two_stage_opamp_dummy_magic_29_0.Y.n117 two_stage_opamp_dummy_magic_29_0.Y.n26 2.24063
R16364 two_stage_opamp_dummy_magic_29_0.Y.n86 two_stage_opamp_dummy_magic_29_0.Y.n85 2.24063
R16365 two_stage_opamp_dummy_magic_29_0.Y.n63 two_stage_opamp_dummy_magic_29_0.Y.n37 2.24063
R16366 two_stage_opamp_dummy_magic_29_0.Y.n45 two_stage_opamp_dummy_magic_29_0.Y.n38 2.24063
R16367 two_stage_opamp_dummy_magic_29_0.Y.n114 two_stage_opamp_dummy_magic_29_0.Y.n113 2.24063
R16368 two_stage_opamp_dummy_magic_29_0.Y.n114 two_stage_opamp_dummy_magic_29_0.Y.n90 2.24063
R16369 two_stage_opamp_dummy_magic_29_0.Y.n115 two_stage_opamp_dummy_magic_29_0.Y.n114 2.24063
R16370 two_stage_opamp_dummy_magic_29_0.Y.n87 two_stage_opamp_dummy_magic_29_0.Y.n35 2.24063
R16371 two_stage_opamp_dummy_magic_29_0.Y.n44 two_stage_opamp_dummy_magic_29_0.Y.n43 2.24063
R16372 two_stage_opamp_dummy_magic_29_0.Y.n62 two_stage_opamp_dummy_magic_29_0.Y.n46 2.22018
R16373 two_stage_opamp_dummy_magic_29_0.Y.n62 two_stage_opamp_dummy_magic_29_0.Y.n45 0.682792
R16374 two_stage_opamp_dummy_magic_29_0.Y.n119 two_stage_opamp_dummy_magic_29_0.Y.n118 0.643357
R16375 two_stage_opamp_dummy_magic_29_0.Y.n120 two_stage_opamp_dummy_magic_29_0.Y.n24 0.643357
R16376 two_stage_opamp_dummy_magic_29_0.Y.n122 two_stage_opamp_dummy_magic_29_0.Y.n121 0.643357
R16377 two_stage_opamp_dummy_magic_29_0.Y.n123 two_stage_opamp_dummy_magic_29_0.Y.n2 0.643357
R16378 two_stage_opamp_dummy_magic_29_0.Y.n125 two_stage_opamp_dummy_magic_29_0.Y.n124 0.643357
R16379 two_stage_opamp_dummy_magic_29_0.Y.n23 two_stage_opamp_dummy_magic_29_0.Y.n0 0.643357
R16380 two_stage_opamp_dummy_magic_29_0.Y.n22 two_stage_opamp_dummy_magic_29_0.Y.n21 0.643357
R16381 two_stage_opamp_dummy_magic_29_0.Y.n20 two_stage_opamp_dummy_magic_29_0.Y.n3 0.643357
R16382 two_stage_opamp_dummy_magic_29_0.Y.n88 two_stage_opamp_dummy_magic_29_0.Y.n87 0.479667
R16383 two_stage_opamp_dummy_magic_29_0.Y.n85 two_stage_opamp_dummy_magic_29_0.Y.n62 0.46925
R16384 two_stage_opamp_dummy_magic_29_0.Y.n108 two_stage_opamp_dummy_magic_29_0.Y.n105 0.3755
R16385 two_stage_opamp_dummy_magic_29_0.Y.n105 two_stage_opamp_dummy_magic_29_0.Y.n92 0.3755
R16386 two_stage_opamp_dummy_magic_29_0.Y.n95 two_stage_opamp_dummy_magic_29_0.Y.n92 0.3755
R16387 two_stage_opamp_dummy_magic_29_0.Y.n111 two_stage_opamp_dummy_magic_29_0.Y.n91 0.3755
R16388 two_stage_opamp_dummy_magic_29_0.Y.n102 two_stage_opamp_dummy_magic_29_0.Y.n91 0.3755
R16389 two_stage_opamp_dummy_magic_29_0.Y.n102 two_stage_opamp_dummy_magic_29_0.Y.n101 0.3755
R16390 two_stage_opamp_dummy_magic_29_0.Y.n101 two_stage_opamp_dummy_magic_29_0.Y.n98 0.3755
R16391 two_stage_opamp_dummy_magic_29_0.Y.n16 two_stage_opamp_dummy_magic_29_0.Y.n14 0.34425
R16392 two_stage_opamp_dummy_magic_29_0.Y.n14 two_stage_opamp_dummy_magic_29_0.Y.n12 0.34425
R16393 two_stage_opamp_dummy_magic_29_0.Y.n12 two_stage_opamp_dummy_magic_29_0.Y.n10 0.34425
R16394 two_stage_opamp_dummy_magic_29_0.Y.n10 two_stage_opamp_dummy_magic_29_0.Y.n8 0.34425
R16395 two_stage_opamp_dummy_magic_29_0.Y.n17 two_stage_opamp_dummy_magic_29_0.Y.n5 0.34425
R16396 two_stage_opamp_dummy_magic_29_0.Y.n5 two_stage_opamp_dummy_magic_29_0.Y.n4 0.34425
R16397 two_stage_opamp_dummy_magic_29_0.Y.n4 two_stage_opamp_dummy_magic_29_0.Y.n1 0.34425
R16398 two_stage_opamp_dummy_magic_29_0.Y.n25 two_stage_opamp_dummy_magic_29_0.Y.n1 0.34425
R16399 two_stage_opamp_dummy_magic_29_0.Y.n118 two_stage_opamp_dummy_magic_29_0.Y.n117 0.270589
R16400 two_stage_opamp_dummy_magic_29_0.Y.n18 two_stage_opamp_dummy_magic_29_0.Y.n3 0.242602
R16401 two_stage_opamp_dummy_magic_29_0.Y.n61 two_stage_opamp_dummy_magic_29_0.Y.n47 0.1255
R16402 two_stage_opamp_dummy_magic_29_0.Y.n47 two_stage_opamp_dummy_magic_29_0.Y.n46 0.0626438
R16403 two_stage_opamp_dummy_magic_29_0.Y.n85 two_stage_opamp_dummy_magic_29_0.Y.n37 0.0421667
R16404 two_stage_opamp_dummy_magic_29_0.Y.n20 two_stage_opamp_dummy_magic_29_0.Y.n19 0.0250536
R16405 two_stage_opamp_dummy_magic_29_0.Y.n21 two_stage_opamp_dummy_magic_29_0.Y.n20 0.0250536
R16406 two_stage_opamp_dummy_magic_29_0.Y.n21 two_stage_opamp_dummy_magic_29_0.Y.n0 0.0250536
R16407 two_stage_opamp_dummy_magic_29_0.Y.n125 two_stage_opamp_dummy_magic_29_0.Y.n2 0.0250536
R16408 two_stage_opamp_dummy_magic_29_0.Y.n121 two_stage_opamp_dummy_magic_29_0.Y.n2 0.0250536
R16409 two_stage_opamp_dummy_magic_29_0.Y.n121 two_stage_opamp_dummy_magic_29_0.Y.n120 0.0250536
R16410 two_stage_opamp_dummy_magic_29_0.Y.n120 two_stage_opamp_dummy_magic_29_0.Y.n119 0.0250536
R16411 two_stage_opamp_dummy_magic_29_0.Y.n22 two_stage_opamp_dummy_magic_29_0.Y.n3 0.0250536
R16412 two_stage_opamp_dummy_magic_29_0.Y.n23 two_stage_opamp_dummy_magic_29_0.Y.n22 0.0250536
R16413 two_stage_opamp_dummy_magic_29_0.Y.n124 two_stage_opamp_dummy_magic_29_0.Y.n23 0.0250536
R16414 two_stage_opamp_dummy_magic_29_0.Y.n124 two_stage_opamp_dummy_magic_29_0.Y.n123 0.0250536
R16415 two_stage_opamp_dummy_magic_29_0.Y.n123 two_stage_opamp_dummy_magic_29_0.Y.n122 0.0250536
R16416 two_stage_opamp_dummy_magic_29_0.Y.n122 two_stage_opamp_dummy_magic_29_0.Y.n24 0.0250536
R16417 two_stage_opamp_dummy_magic_29_0.Y.n118 two_stage_opamp_dummy_magic_29_0.Y.n24 0.0250536
R16418 two_stage_opamp_dummy_magic_29_0.Y.n19 two_stage_opamp_dummy_magic_29_0.Y.n18 0.024102
R16419 two_stage_opamp_dummy_magic_29_0.Y.n33 two_stage_opamp_dummy_magic_29_0.Y.n30 0.0217373
R16420 two_stage_opamp_dummy_magic_29_0.Y.n116 two_stage_opamp_dummy_magic_29_0.Y.n31 0.0217373
R16421 two_stage_opamp_dummy_magic_29_0.Y.n32 two_stage_opamp_dummy_magic_29_0.Y.n26 0.0217373
R16422 two_stage_opamp_dummy_magic_29_0.Y.n87 two_stage_opamp_dummy_magic_29_0.Y.n86 0.0217373
R16423 two_stage_opamp_dummy_magic_29_0.Y.n84 two_stage_opamp_dummy_magic_29_0.Y.n63 0.0217373
R16424 two_stage_opamp_dummy_magic_29_0.Y.n33 two_stage_opamp_dummy_magic_29_0.Y.n28 0.0217373
R16425 two_stage_opamp_dummy_magic_29_0.Y.n31 two_stage_opamp_dummy_magic_29_0.Y.n27 0.0217373
R16426 two_stage_opamp_dummy_magic_29_0.Y.n88 two_stage_opamp_dummy_magic_29_0.Y.n26 0.0217373
R16427 two_stage_opamp_dummy_magic_29_0.Y.n86 two_stage_opamp_dummy_magic_29_0.Y.n36 0.0217373
R16428 two_stage_opamp_dummy_magic_29_0.Y.n63 two_stage_opamp_dummy_magic_29_0.Y.n36 0.0217373
R16429 two_stage_opamp_dummy_magic_29_0.Y.n40 two_stage_opamp_dummy_magic_29_0.Y.n38 0.0217373
R16430 two_stage_opamp_dummy_magic_29_0.Y.n41 two_stage_opamp_dummy_magic_29_0.Y.n39 0.0217373
R16431 two_stage_opamp_dummy_magic_29_0.Y.n113 two_stage_opamp_dummy_magic_29_0.Y.n28 0.0217373
R16432 two_stage_opamp_dummy_magic_29_0.Y.n90 two_stage_opamp_dummy_magic_29_0.Y.n27 0.0217373
R16433 two_stage_opamp_dummy_magic_29_0.Y.n115 two_stage_opamp_dummy_magic_29_0.Y.n32 0.0217373
R16434 two_stage_opamp_dummy_magic_29_0.Y.n113 two_stage_opamp_dummy_magic_29_0.Y.n112 0.0217373
R16435 two_stage_opamp_dummy_magic_29_0.Y.n90 two_stage_opamp_dummy_magic_29_0.Y.n30 0.0217373
R16436 two_stage_opamp_dummy_magic_29_0.Y.n116 two_stage_opamp_dummy_magic_29_0.Y.n115 0.0217373
R16437 two_stage_opamp_dummy_magic_29_0.Y.n83 two_stage_opamp_dummy_magic_29_0.Y.n35 0.0217373
R16438 two_stage_opamp_dummy_magic_29_0.Y.n44 two_stage_opamp_dummy_magic_29_0.Y.n39 0.0217373
R16439 two_stage_opamp_dummy_magic_29_0.Y.n37 two_stage_opamp_dummy_magic_29_0.Y.n35 0.0217373
R16440 two_stage_opamp_dummy_magic_29_0.Y.n42 two_stage_opamp_dummy_magic_29_0.Y.n40 0.0217373
R16441 two_stage_opamp_dummy_magic_29_0.Y.n43 two_stage_opamp_dummy_magic_29_0.Y.n42 0.0217373
R16442 two_stage_opamp_dummy_magic_29_0.Y.n45 two_stage_opamp_dummy_magic_29_0.Y.n44 0.0217373
R16443 two_stage_opamp_dummy_magic_29_0.Y two_stage_opamp_dummy_magic_29_0.Y.n0 0.016125
R16444 two_stage_opamp_dummy_magic_29_0.Y.n34 two_stage_opamp_dummy_magic_29_0.Y.n29 0.00991089
R16445 two_stage_opamp_dummy_magic_29_0.Y.n114 two_stage_opamp_dummy_magic_29_0.Y.n89 0.00991089
R16446 two_stage_opamp_dummy_magic_29_0.Y.n117 two_stage_opamp_dummy_magic_29_0.Y.n29 0.00991089
R16447 two_stage_opamp_dummy_magic_29_0.Y.n89 two_stage_opamp_dummy_magic_29_0.Y.n34 0.00991089
R16448 two_stage_opamp_dummy_magic_29_0.Y two_stage_opamp_dummy_magic_29_0.Y.n125 0.00942857
R16449 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.n0 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.t5 447.279
R16450 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.n0 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.t7 446.967
R16451 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.n1 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.t2 446.967
R16452 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.n2 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.t3 446.967
R16453 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.n5 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.t8 344.772
R16454 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.n8 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.t9 281.168
R16455 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.n7 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.t4 281.168
R16456 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.n6 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.t6 281.168
R16457 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.n8 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.n7 205.946
R16458 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.n7 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.n6 205.946
R16459 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.n7 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.n4 165.8
R16460 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.n9 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.n8 165.8
R16461 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.n3 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.t1 108.615
R16462 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.n10 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.t0 108.615
R16463 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.n6 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.n5 63.4857
R16464 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.n5 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.n4 51.5193
R16465 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.n10 15.6567
R16466 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.n3 10.5317
R16467 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.n3 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.n2 6.0005
R16468 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.n10 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.n9 6.0005
R16469 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.n2 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.n1 0.313
R16470 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.n1 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.n0 0.313
R16471 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.n9 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.n4 0.313
R16472 VOUT-.n179 VOUT-.t10 110.386
R16473 VOUT-.n39 VOUT-.n38 34.9935
R16474 VOUT-.n28 VOUT-.n27 34.9935
R16475 VOUT-.n30 VOUT-.n29 34.9935
R16476 VOUT-.n33 VOUT-.n32 34.9935
R16477 VOUT-.n36 VOUT-.n35 34.9935
R16478 VOUT-.n42 VOUT-.n41 34.9935
R16479 VOUT-.n186 VOUT-.n185 9.73997
R16480 VOUT-.n182 VOUT-.n181 9.73997
R16481 VOUT-.n189 VOUT-.n188 9.73997
R16482 VOUT-.n187 VOUT-.n182 6.64633
R16483 VOUT-.n187 VOUT-.n186 6.64633
R16484 VOUT-.n38 VOUT-.t11 6.56717
R16485 VOUT-.n38 VOUT-.t18 6.56717
R16486 VOUT-.n27 VOUT-.t17 6.56717
R16487 VOUT-.n27 VOUT-.t14 6.56717
R16488 VOUT-.n29 VOUT-.t0 6.56717
R16489 VOUT-.n29 VOUT-.t3 6.56717
R16490 VOUT-.n32 VOUT-.t12 6.56717
R16491 VOUT-.n32 VOUT-.t15 6.56717
R16492 VOUT-.n35 VOUT-.t1 6.56717
R16493 VOUT-.n35 VOUT-.t13 6.56717
R16494 VOUT-.n41 VOUT-.t2 6.56717
R16495 VOUT-.n41 VOUT-.t16 6.56717
R16496 VOUT-.n31 VOUT-.n28 6.3755
R16497 VOUT-.n40 VOUT-.n39 6.3755
R16498 VOUT-.n189 VOUT-.n187 6.02133
R16499 VOUT-.n31 VOUT-.n30 5.813
R16500 VOUT-.n34 VOUT-.n33 5.813
R16501 VOUT-.n37 VOUT-.n36 5.813
R16502 VOUT-.n42 VOUT-.n40 5.813
R16503 VOUT-.n46 VOUT-.n26 5.063
R16504 VOUT-.n43 VOUT-.n19 5.063
R16505 VOUT-.n111 VOUT-.t131 4.8295
R16506 VOUT-.n110 VOUT-.t39 4.8295
R16507 VOUT-.n109 VOUT-.t75 4.8295
R16508 VOUT-.n108 VOUT-.t64 4.8295
R16509 VOUT-.n125 VOUT-.t98 4.8295
R16510 VOUT-.n126 VOUT-.t69 4.8295
R16511 VOUT-.n128 VOUT-.t141 4.8295
R16512 VOUT-.n129 VOUT-.t109 4.8295
R16513 VOUT-.n131 VOUT-.t101 4.8295
R16514 VOUT-.n132 VOUT-.t72 4.8295
R16515 VOUT-.n134 VOUT-.t138 4.8295
R16516 VOUT-.n135 VOUT-.t103 4.8295
R16517 VOUT-.n137 VOUT-.t96 4.8295
R16518 VOUT-.n138 VOUT-.t65 4.8295
R16519 VOUT-.n140 VOUT-.t56 4.8295
R16520 VOUT-.n141 VOUT-.t26 4.8295
R16521 VOUT-.n143 VOUT-.t90 4.8295
R16522 VOUT-.n144 VOUT-.t58 4.8295
R16523 VOUT-.n146 VOUT-.t53 4.8295
R16524 VOUT-.n147 VOUT-.t19 4.8295
R16525 VOUT-.n149 VOUT-.t154 4.8295
R16526 VOUT-.n150 VOUT-.t121 4.8295
R16527 VOUT-.n71 VOUT-.t83 4.8295
R16528 VOUT-.n73 VOUT-.t43 4.8295
R16529 VOUT-.n87 VOUT-.t37 4.8295
R16530 VOUT-.n88 VOUT-.t147 4.8295
R16531 VOUT-.n90 VOUT-.t74 4.8295
R16532 VOUT-.n91 VOUT-.t41 4.8295
R16533 VOUT-.n93 VOUT-.t87 4.8295
R16534 VOUT-.n94 VOUT-.t104 4.8295
R16535 VOUT-.n96 VOUT-.t102 4.8295
R16536 VOUT-.n97 VOUT-.t71 4.8295
R16537 VOUT-.n99 VOUT-.t68 4.8295
R16538 VOUT-.n100 VOUT-.t36 4.8295
R16539 VOUT-.n102 VOUT-.t107 4.8295
R16540 VOUT-.n103 VOUT-.t76 4.8295
R16541 VOUT-.n105 VOUT-.t148 4.8295
R16542 VOUT-.n106 VOUT-.t116 4.8295
R16543 VOUT-.n152 VOUT-.t113 4.8295
R16544 VOUT-.n112 VOUT-.t30 4.8154
R16545 VOUT-.n115 VOUT-.t62 4.8154
R16546 VOUT-.n113 VOUT-.t143 4.81305
R16547 VOUT-.n116 VOUT-.t38 4.81305
R16548 VOUT-.n114 VOUT-.t24 4.806
R16549 VOUT-.n117 VOUT-.t79 4.806
R16550 VOUT-.n118 VOUT-.t117 4.806
R16551 VOUT-.n74 VOUT-.t155 4.806
R16552 VOUT-.n75 VOUT-.t133 4.806
R16553 VOUT-.n76 VOUT-.t150 4.806
R16554 VOUT-.n77 VOUT-.t47 4.806
R16555 VOUT-.n78 VOUT-.t25 4.806
R16556 VOUT-.n79 VOUT-.t63 4.806
R16557 VOUT-.n80 VOUT-.t99 4.806
R16558 VOUT-.n81 VOUT-.t139 4.806
R16559 VOUT-.n82 VOUT-.t119 4.806
R16560 VOUT-.n83 VOUT-.t157 4.806
R16561 VOUT-.n84 VOUT-.t52 4.806
R16562 VOUT-.n85 VOUT-.t33 4.806
R16563 VOUT-.n111 VOUT-.t156 4.5005
R16564 VOUT-.n110 VOUT-.t135 4.5005
R16565 VOUT-.n109 VOUT-.t32 4.5005
R16566 VOUT-.n108 VOUT-.t86 4.5005
R16567 VOUT-.n124 VOUT-.t48 4.5005
R16568 VOUT-.n123 VOUT-.t151 4.5005
R16569 VOUT-.n122 VOUT-.t35 4.5005
R16570 VOUT-.n121 VOUT-.t137 4.5005
R16571 VOUT-.n120 VOUT-.t94 4.5005
R16572 VOUT-.n119 VOUT-.t120 4.5005
R16573 VOUT-.n118 VOUT-.t81 4.5005
R16574 VOUT-.n117 VOUT-.t42 4.5005
R16575 VOUT-.n116 VOUT-.t142 4.5005
R16576 VOUT-.n115 VOUT-.t29 4.5005
R16577 VOUT-.n114 VOUT-.t130 4.5005
R16578 VOUT-.n113 VOUT-.t111 4.5005
R16579 VOUT-.n112 VOUT-.t136 4.5005
R16580 VOUT-.n125 VOUT-.t124 4.5005
R16581 VOUT-.n127 VOUT-.t82 4.5005
R16582 VOUT-.n126 VOUT-.t44 4.5005
R16583 VOUT-.n128 VOUT-.t89 4.5005
R16584 VOUT-.n130 VOUT-.t54 4.5005
R16585 VOUT-.n129 VOUT-.t20 4.5005
R16586 VOUT-.n131 VOUT-.t51 4.5005
R16587 VOUT-.n133 VOUT-.t160 4.5005
R16588 VOUT-.n132 VOUT-.t123 4.5005
R16589 VOUT-.n134 VOUT-.t84 4.5005
R16590 VOUT-.n136 VOUT-.t49 4.5005
R16591 VOUT-.n135 VOUT-.t159 4.5005
R16592 VOUT-.n137 VOUT-.t45 4.5005
R16593 VOUT-.n139 VOUT-.t152 4.5005
R16594 VOUT-.n138 VOUT-.t118 4.5005
R16595 VOUT-.n140 VOUT-.t145 4.5005
R16596 VOUT-.n142 VOUT-.t112 4.5005
R16597 VOUT-.n141 VOUT-.t77 4.5005
R16598 VOUT-.n143 VOUT-.t40 4.5005
R16599 VOUT-.n145 VOUT-.t144 4.5005
R16600 VOUT-.n144 VOUT-.t110 4.5005
R16601 VOUT-.n146 VOUT-.t140 4.5005
R16602 VOUT-.n148 VOUT-.t106 4.5005
R16603 VOUT-.n147 VOUT-.t73 4.5005
R16604 VOUT-.n149 VOUT-.t100 4.5005
R16605 VOUT-.n151 VOUT-.t67 4.5005
R16606 VOUT-.n150 VOUT-.t34 4.5005
R16607 VOUT-.n71 VOUT-.t105 4.5005
R16608 VOUT-.n72 VOUT-.t70 4.5005
R16609 VOUT-.n73 VOUT-.t66 4.5005
R16610 VOUT-.n86 VOUT-.t31 4.5005
R16611 VOUT-.n85 VOUT-.t132 4.5005
R16612 VOUT-.n84 VOUT-.t153 4.5005
R16613 VOUT-.n83 VOUT-.t115 4.5005
R16614 VOUT-.n82 VOUT-.t78 4.5005
R16615 VOUT-.n81 VOUT-.t97 4.5005
R16616 VOUT-.n80 VOUT-.t59 4.5005
R16617 VOUT-.n79 VOUT-.t22 4.5005
R16618 VOUT-.n78 VOUT-.t126 4.5005
R16619 VOUT-.n77 VOUT-.t146 4.5005
R16620 VOUT-.n76 VOUT-.t108 4.5005
R16621 VOUT-.n75 VOUT-.t88 4.5005
R16622 VOUT-.n74 VOUT-.t114 4.5005
R16623 VOUT-.n87 VOUT-.t129 4.5005
R16624 VOUT-.n89 VOUT-.t92 4.5005
R16625 VOUT-.n88 VOUT-.t57 4.5005
R16626 VOUT-.n90 VOUT-.t23 4.5005
R16627 VOUT-.n92 VOUT-.t128 4.5005
R16628 VOUT-.n91 VOUT-.t91 4.5005
R16629 VOUT-.n93 VOUT-.t46 4.5005
R16630 VOUT-.n95 VOUT-.t95 4.5005
R16631 VOUT-.n94 VOUT-.t149 4.5005
R16632 VOUT-.n96 VOUT-.t50 4.5005
R16633 VOUT-.n98 VOUT-.t158 4.5005
R16634 VOUT-.n97 VOUT-.t122 4.5005
R16635 VOUT-.n99 VOUT-.t161 4.5005
R16636 VOUT-.n101 VOUT-.t125 4.5005
R16637 VOUT-.n100 VOUT-.t85 4.5005
R16638 VOUT-.n102 VOUT-.t55 4.5005
R16639 VOUT-.n104 VOUT-.t21 4.5005
R16640 VOUT-.n103 VOUT-.t127 4.5005
R16641 VOUT-.n105 VOUT-.t93 4.5005
R16642 VOUT-.n107 VOUT-.t60 4.5005
R16643 VOUT-.n106 VOUT-.t27 4.5005
R16644 VOUT-.n152 VOUT-.t61 4.5005
R16645 VOUT-.n153 VOUT-.t28 4.5005
R16646 VOUT-.n154 VOUT-.t134 4.5005
R16647 VOUT-.n155 VOUT-.t80 4.5005
R16648 VOUT-.n47 VOUT-.n46 4.5005
R16649 VOUT-.n45 VOUT-.n24 4.5005
R16650 VOUT-.n44 VOUT-.n23 4.5005
R16651 VOUT-.n43 VOUT-.n20 4.5005
R16652 VOUT-.n65 VOUT-.n64 4.5005
R16653 VOUT-.n16 VOUT-.n13 4.5005
R16654 VOUT-.n65 VOUT-.n13 4.5005
R16655 VOUT-.n66 VOUT-.n9 4.5005
R16656 VOUT-.n66 VOUT-.n11 4.5005
R16657 VOUT-.n66 VOUT-.n65 4.5005
R16658 VOUT-.n164 VOUT-.n69 4.5005
R16659 VOUT-.n165 VOUT-.n164 4.5005
R16660 VOUT-.n165 VOUT-.n5 4.5005
R16661 VOUT-.n166 VOUT-.n4 4.5005
R16662 VOUT-.n166 VOUT-.n165 4.5005
R16663 VOUT-.n178 VOUT-.n177 4.5005
R16664 VOUT-.n178 VOUT-.n1 4.5005
R16665 VOUT-.n174 VOUT-.n1 4.5005
R16666 VOUT-.n171 VOUT-.n1 4.5005
R16667 VOUT-.n172 VOUT-.n1 4.5005
R16668 VOUT-.n174 VOUT-.n173 4.5005
R16669 VOUT-.n173 VOUT-.n171 4.5005
R16670 VOUT-.n173 VOUT-.n172 4.5005
R16671 VOUT-.n185 VOUT-.t7 3.42907
R16672 VOUT-.n185 VOUT-.t4 3.42907
R16673 VOUT-.n181 VOUT-.t5 3.42907
R16674 VOUT-.n181 VOUT-.t8 3.42907
R16675 VOUT-.n188 VOUT-.t9 3.42907
R16676 VOUT-.n188 VOUT-.t6 3.42907
R16677 VOUT-.n63 VOUT-.n62 2.24601
R16678 VOUT-.n14 VOUT-.n8 2.24601
R16679 VOUT-.n176 VOUT-.n175 2.24601
R16680 VOUT-.n170 VOUT-.n169 2.24601
R16681 VOUT-.n163 VOUT-.n162 2.24477
R16682 VOUT-.n7 VOUT-.n2 2.24477
R16683 VOUT-.n66 VOUT-.n10 2.24063
R16684 VOUT-.n166 VOUT-.n3 2.24063
R16685 VOUT-.n173 VOUT-.n0 2.24063
R16686 VOUT-.n13 VOUT-.n12 2.24063
R16687 VOUT-.n164 VOUT-.n67 2.24063
R16688 VOUT-.n68 VOUT-.n5 2.24063
R16689 VOUT-.n177 VOUT-.n168 2.24063
R16690 VOUT-.n177 VOUT-.n167 2.24063
R16691 VOUT-.n64 VOUT-.n17 2.23934
R16692 VOUT-.n64 VOUT-.n15 2.23934
R16693 VOUT-.n186 VOUT-.n184 1.83719
R16694 VOUT-.n197 VOUT-.n182 1.72967
R16695 VOUT-.n190 VOUT-.n189 1.72967
R16696 VOUT-.n50 VOUT-.n25 1.5005
R16697 VOUT-.n52 VOUT-.n51 1.5005
R16698 VOUT-.n53 VOUT-.n22 1.5005
R16699 VOUT-.n55 VOUT-.n54 1.5005
R16700 VOUT-.n56 VOUT-.n21 1.5005
R16701 VOUT-.n58 VOUT-.n57 1.5005
R16702 VOUT-.n59 VOUT-.n18 1.5005
R16703 VOUT-.n61 VOUT-.n60 1.5005
R16704 VOUT-.n192 VOUT-.n191 1.5005
R16705 VOUT-.n193 VOUT-.n183 1.5005
R16706 VOUT-.n195 VOUT-.n194 1.5005
R16707 VOUT-.n196 VOUT-.n180 1.5005
R16708 VOUT-.n198 VOUT-.n197 1.5005
R16709 VOUT-.n30 VOUT-.n20 1.313
R16710 VOUT-.n33 VOUT-.n23 1.313
R16711 VOUT-.n36 VOUT-.n24 1.313
R16712 VOUT-.n47 VOUT-.n42 1.313
R16713 VOUT-.n28 VOUT-.n19 1.313
R16714 VOUT-.n39 VOUT-.n26 1.313
R16715 VOUT-.n162 VOUT-.n161 1.1455
R16716 VOUT-.n156 VOUT-.n6 1.13717
R16717 VOUT-.n158 VOUT-.n157 1.13717
R16718 VOUT-.n160 VOUT-.n159 1.13717
R16719 VOUT-.n165 VOUT-.n6 1.13717
R16720 VOUT-.n158 VOUT-.n7 1.13717
R16721 VOUT-.n159 VOUT-.n4 1.13717
R16722 VOUT-.n70 VOUT-.n69 1.13717
R16723 VOUT-.n62 VOUT-.n61 0.859875
R16724 VOUT-.n49 VOUT-.n26 0.715216
R16725 VOUT-.n58 VOUT-.n20 0.65675
R16726 VOUT-.n54 VOUT-.n23 0.65675
R16727 VOUT-.n52 VOUT-.n24 0.65675
R16728 VOUT-.n48 VOUT-.n47 0.65675
R16729 VOUT-.n60 VOUT-.n19 0.65675
R16730 VOUT-.n161 VOUT-.n160 0.585
R16731 VOUT-.n50 VOUT-.n49 0.564601
R16732 VOUT-.n46 VOUT-.n45 0.563
R16733 VOUT-.n45 VOUT-.n44 0.563
R16734 VOUT-.n44 VOUT-.n43 0.563
R16735 VOUT-.n34 VOUT-.n31 0.563
R16736 VOUT-.n37 VOUT-.n34 0.563
R16737 VOUT-.n40 VOUT-.n37 0.563
R16738 VOUT-.n179 VOUT-.n178 0.557792
R16739 VOUT-.n177 VOUT-.n166 0.5455
R16740 VOUT-.n124 VOUT-.n108 0.3295
R16741 VOUT-.n124 VOUT-.n123 0.3295
R16742 VOUT-.n123 VOUT-.n122 0.3295
R16743 VOUT-.n122 VOUT-.n121 0.3295
R16744 VOUT-.n121 VOUT-.n120 0.3295
R16745 VOUT-.n120 VOUT-.n119 0.3295
R16746 VOUT-.n119 VOUT-.n118 0.3295
R16747 VOUT-.n118 VOUT-.n117 0.3295
R16748 VOUT-.n117 VOUT-.n116 0.3295
R16749 VOUT-.n116 VOUT-.n115 0.3295
R16750 VOUT-.n115 VOUT-.n114 0.3295
R16751 VOUT-.n114 VOUT-.n113 0.3295
R16752 VOUT-.n113 VOUT-.n112 0.3295
R16753 VOUT-.n127 VOUT-.n125 0.3295
R16754 VOUT-.n127 VOUT-.n126 0.3295
R16755 VOUT-.n130 VOUT-.n128 0.3295
R16756 VOUT-.n130 VOUT-.n129 0.3295
R16757 VOUT-.n133 VOUT-.n131 0.3295
R16758 VOUT-.n133 VOUT-.n132 0.3295
R16759 VOUT-.n136 VOUT-.n134 0.3295
R16760 VOUT-.n136 VOUT-.n135 0.3295
R16761 VOUT-.n139 VOUT-.n137 0.3295
R16762 VOUT-.n139 VOUT-.n138 0.3295
R16763 VOUT-.n142 VOUT-.n140 0.3295
R16764 VOUT-.n142 VOUT-.n141 0.3295
R16765 VOUT-.n145 VOUT-.n143 0.3295
R16766 VOUT-.n145 VOUT-.n144 0.3295
R16767 VOUT-.n148 VOUT-.n146 0.3295
R16768 VOUT-.n148 VOUT-.n147 0.3295
R16769 VOUT-.n151 VOUT-.n149 0.3295
R16770 VOUT-.n151 VOUT-.n150 0.3295
R16771 VOUT-.n72 VOUT-.n71 0.3295
R16772 VOUT-.n86 VOUT-.n73 0.3295
R16773 VOUT-.n86 VOUT-.n85 0.3295
R16774 VOUT-.n85 VOUT-.n84 0.3295
R16775 VOUT-.n84 VOUT-.n83 0.3295
R16776 VOUT-.n83 VOUT-.n82 0.3295
R16777 VOUT-.n82 VOUT-.n81 0.3295
R16778 VOUT-.n81 VOUT-.n80 0.3295
R16779 VOUT-.n80 VOUT-.n79 0.3295
R16780 VOUT-.n79 VOUT-.n78 0.3295
R16781 VOUT-.n78 VOUT-.n77 0.3295
R16782 VOUT-.n77 VOUT-.n76 0.3295
R16783 VOUT-.n76 VOUT-.n75 0.3295
R16784 VOUT-.n75 VOUT-.n74 0.3295
R16785 VOUT-.n89 VOUT-.n87 0.3295
R16786 VOUT-.n89 VOUT-.n88 0.3295
R16787 VOUT-.n92 VOUT-.n90 0.3295
R16788 VOUT-.n92 VOUT-.n91 0.3295
R16789 VOUT-.n95 VOUT-.n93 0.3295
R16790 VOUT-.n95 VOUT-.n94 0.3295
R16791 VOUT-.n98 VOUT-.n96 0.3295
R16792 VOUT-.n98 VOUT-.n97 0.3295
R16793 VOUT-.n101 VOUT-.n99 0.3295
R16794 VOUT-.n101 VOUT-.n100 0.3295
R16795 VOUT-.n104 VOUT-.n102 0.3295
R16796 VOUT-.n104 VOUT-.n103 0.3295
R16797 VOUT-.n107 VOUT-.n105 0.3295
R16798 VOUT-.n107 VOUT-.n106 0.3295
R16799 VOUT-.n153 VOUT-.n152 0.3295
R16800 VOUT-.n154 VOUT-.n153 0.3295
R16801 VOUT-.n192 VOUT-.n184 0.314966
R16802 VOUT-.n155 VOUT-.n154 0.3107
R16803 VOUT-.n119 VOUT-.n111 0.306
R16804 VOUT-.n120 VOUT-.n110 0.306
R16805 VOUT-.n121 VOUT-.n109 0.306
R16806 VOUT-.n127 VOUT-.n124 0.2825
R16807 VOUT-.n130 VOUT-.n127 0.2825
R16808 VOUT-.n133 VOUT-.n130 0.2825
R16809 VOUT-.n136 VOUT-.n133 0.2825
R16810 VOUT-.n139 VOUT-.n136 0.2825
R16811 VOUT-.n142 VOUT-.n139 0.2825
R16812 VOUT-.n145 VOUT-.n142 0.2825
R16813 VOUT-.n148 VOUT-.n145 0.2825
R16814 VOUT-.n151 VOUT-.n148 0.2825
R16815 VOUT-.n86 VOUT-.n72 0.2825
R16816 VOUT-.n89 VOUT-.n86 0.2825
R16817 VOUT-.n92 VOUT-.n89 0.2825
R16818 VOUT-.n95 VOUT-.n92 0.2825
R16819 VOUT-.n98 VOUT-.n95 0.2825
R16820 VOUT-.n101 VOUT-.n98 0.2825
R16821 VOUT-.n104 VOUT-.n101 0.2825
R16822 VOUT-.n107 VOUT-.n104 0.2825
R16823 VOUT-.n153 VOUT-.n107 0.2825
R16824 VOUT-.n153 VOUT-.n151 0.2825
R16825 VOUT-.n164 VOUT-.n66 0.2455
R16826 VOUT- VOUT-.n179 0.198417
R16827 VOUT- VOUT-.n198 0.182792
R16828 VOUT-.n156 VOUT-.n155 0.138367
R16829 VOUT-.n190 VOUT-.n184 0.0891864
R16830 VOUT-.n60 VOUT-.n59 0.0577917
R16831 VOUT-.n59 VOUT-.n58 0.0577917
R16832 VOUT-.n58 VOUT-.n21 0.0577917
R16833 VOUT-.n54 VOUT-.n21 0.0577917
R16834 VOUT-.n54 VOUT-.n53 0.0577917
R16835 VOUT-.n53 VOUT-.n52 0.0577917
R16836 VOUT-.n52 VOUT-.n25 0.0577917
R16837 VOUT-.n48 VOUT-.n25 0.0577917
R16838 VOUT-.n61 VOUT-.n18 0.0577917
R16839 VOUT-.n57 VOUT-.n18 0.0577917
R16840 VOUT-.n57 VOUT-.n56 0.0577917
R16841 VOUT-.n56 VOUT-.n55 0.0577917
R16842 VOUT-.n55 VOUT-.n22 0.0577917
R16843 VOUT-.n51 VOUT-.n22 0.0577917
R16844 VOUT-.n51 VOUT-.n50 0.0577917
R16845 VOUT-.n49 VOUT-.n48 0.054517
R16846 VOUT-.n171 VOUT-.n170 0.047375
R16847 VOUT-.n175 VOUT-.n174 0.047375
R16848 VOUT-.n165 VOUT-.n7 0.0421667
R16849 VOUT-.n65 VOUT-.n14 0.0421667
R16850 VOUT-.n197 VOUT-.n196 0.0421667
R16851 VOUT-.n196 VOUT-.n195 0.0421667
R16852 VOUT-.n195 VOUT-.n183 0.0421667
R16853 VOUT-.n191 VOUT-.n183 0.0421667
R16854 VOUT-.n191 VOUT-.n190 0.0421667
R16855 VOUT-.n198 VOUT-.n180 0.0421667
R16856 VOUT-.n194 VOUT-.n180 0.0421667
R16857 VOUT-.n194 VOUT-.n193 0.0421667
R16858 VOUT-.n193 VOUT-.n192 0.0421667
R16859 VOUT-.n15 VOUT-.n14 0.0243161
R16860 VOUT-.n17 VOUT-.n9 0.0243161
R16861 VOUT-.n17 VOUT-.n16 0.0243161
R16862 VOUT-.n15 VOUT-.n11 0.0243161
R16863 VOUT-.n162 VOUT-.n3 0.0217373
R16864 VOUT-.n62 VOUT-.n10 0.0217373
R16865 VOUT-.n16 VOUT-.n10 0.0217373
R16866 VOUT-.n69 VOUT-.n3 0.0217373
R16867 VOUT-.n178 VOUT-.n0 0.0217373
R16868 VOUT-.n175 VOUT-.n0 0.0217373
R16869 VOUT-.n67 VOUT-.n7 0.0217373
R16870 VOUT-.n69 VOUT-.n68 0.0217373
R16871 VOUT-.n12 VOUT-.n9 0.0217373
R16872 VOUT-.n12 VOUT-.n11 0.0217373
R16873 VOUT-.n67 VOUT-.n4 0.0217373
R16874 VOUT-.n68 VOUT-.n4 0.0217373
R16875 VOUT-.n172 VOUT-.n167 0.0217373
R16876 VOUT-.n171 VOUT-.n168 0.0217373
R16877 VOUT-.n174 VOUT-.n168 0.0217373
R16878 VOUT-.n170 VOUT-.n167 0.0217373
R16879 VOUT-.n157 VOUT-.n156 0.0161667
R16880 VOUT-.n160 VOUT-.n157 0.0161667
R16881 VOUT-.n158 VOUT-.n6 0.0161667
R16882 VOUT-.n159 VOUT-.n158 0.0161667
R16883 VOUT-.n159 VOUT-.n70 0.0161667
R16884 VOUT-.n163 VOUT-.n5 0.0134654
R16885 VOUT-.n166 VOUT-.n2 0.0134654
R16886 VOUT-.n164 VOUT-.n163 0.0134654
R16887 VOUT-.n5 VOUT-.n2 0.0134654
R16888 VOUT-.n63 VOUT-.n13 0.0109778
R16889 VOUT-.n66 VOUT-.n8 0.0109778
R16890 VOUT-.n176 VOUT-.n1 0.0109778
R16891 VOUT-.n173 VOUT-.n169 0.0109778
R16892 VOUT-.n64 VOUT-.n63 0.0109778
R16893 VOUT-.n13 VOUT-.n8 0.0109778
R16894 VOUT-.n177 VOUT-.n176 0.0109778
R16895 VOUT-.n169 VOUT-.n1 0.0109778
R16896 VOUT-.n161 VOUT-.n70 0.00872683
R16897 two_stage_opamp_dummy_magic_29_0.Vb2_2.n2 two_stage_opamp_dummy_magic_29_0.Vb2_2.t3 661.375
R16898 two_stage_opamp_dummy_magic_29_0.Vb2_2.n4 two_stage_opamp_dummy_magic_29_0.Vb2_2.t0 661.375
R16899 two_stage_opamp_dummy_magic_29_0.Vb2_2.t4 two_stage_opamp_dummy_magic_29_0.Vb2_2.n0 213.131
R16900 two_stage_opamp_dummy_magic_29_0.Vb2_2.n3 two_stage_opamp_dummy_magic_29_0.Vb2_2.t1 213.131
R16901 two_stage_opamp_dummy_magic_29_0.Vb2_2.n6 two_stage_opamp_dummy_magic_29_0.Vb2_2.n1 154.851
R16902 two_stage_opamp_dummy_magic_29_0.Vb2_2.t8 two_stage_opamp_dummy_magic_29_0.Vb2_2.t4 146.155
R16903 two_stage_opamp_dummy_magic_29_0.Vb2_2.t1 two_stage_opamp_dummy_magic_29_0.Vb2_2.t8 146.155
R16904 two_stage_opamp_dummy_magic_29_0.Vb2_2.t5 two_stage_opamp_dummy_magic_29_0.Vb2_2.n0 76.2576
R16905 two_stage_opamp_dummy_magic_29_0.Vb2_2.n3 two_stage_opamp_dummy_magic_29_0.Vb2_2.t2 76.2576
R16906 two_stage_opamp_dummy_magic_29_0.Vb2_2.n7 two_stage_opamp_dummy_magic_29_0.Vb2_2.n6 66.4503
R16907 two_stage_opamp_dummy_magic_29_0.Vb2_2.n1 two_stage_opamp_dummy_magic_29_0.Vb2_2.t6 21.8894
R16908 two_stage_opamp_dummy_magic_29_0.Vb2_2.n1 two_stage_opamp_dummy_magic_29_0.Vb2_2.t7 21.8894
R16909 two_stage_opamp_dummy_magic_29_0.Vb2_2.t5 two_stage_opamp_dummy_magic_29_0.Vb2_2.n7 11.2576
R16910 two_stage_opamp_dummy_magic_29_0.Vb2_2.n7 two_stage_opamp_dummy_magic_29_0.Vb2_2.t9 11.2576
R16911 two_stage_opamp_dummy_magic_29_0.Vb2_2.n5 two_stage_opamp_dummy_magic_29_0.Vb2_2.n4 5.1255
R16912 two_stage_opamp_dummy_magic_29_0.Vb2_2.n6 two_stage_opamp_dummy_magic_29_0.Vb2_2.n5 4.91195
R16913 two_stage_opamp_dummy_magic_29_0.Vb2_2.n5 two_stage_opamp_dummy_magic_29_0.Vb2_2.n2 4.7505
R16914 two_stage_opamp_dummy_magic_29_0.Vb2_2.n4 two_stage_opamp_dummy_magic_29_0.Vb2_2.n3 1.888
R16915 two_stage_opamp_dummy_magic_29_0.Vb2_2.n2 two_stage_opamp_dummy_magic_29_0.Vb2_2.n0 1.888
R16916 bgr_11_0.V_TOP.n23 bgr_11_0.V_TOP.n21 344.178
R16917 bgr_11_0.V_TOP.n23 bgr_11_0.V_TOP.n22 334.772
R16918 bgr_11_0.V_TOP.n1 bgr_11_0.V_TOP.t37 312.798
R16919 bgr_11_0.V_TOP bgr_11_0.V_TOP.t21 312.639
R16920 bgr_11_0.V_TOP.n36 bgr_11_0.V_TOP.t45 312.5
R16921 bgr_11_0.V_TOP.n42 bgr_11_0.V_TOP.t33 310.401
R16922 bgr_11_0.V_TOP.n41 bgr_11_0.V_TOP.t42 310.401
R16923 bgr_11_0.V_TOP.n40 bgr_11_0.V_TOP.t49 310.401
R16924 bgr_11_0.V_TOP.n39 bgr_11_0.V_TOP.t26 310.401
R16925 bgr_11_0.V_TOP.n38 bgr_11_0.V_TOP.t25 310.401
R16926 bgr_11_0.V_TOP.n37 bgr_11_0.V_TOP.t36 310.401
R16927 bgr_11_0.V_TOP.n5 bgr_11_0.V_TOP.t27 310.401
R16928 bgr_11_0.V_TOP.n4 bgr_11_0.V_TOP.t39 310.401
R16929 bgr_11_0.V_TOP.n3 bgr_11_0.V_TOP.t48 310.401
R16930 bgr_11_0.V_TOP.n2 bgr_11_0.V_TOP.t23 310.401
R16931 bgr_11_0.V_TOP.n1 bgr_11_0.V_TOP.t38 310.401
R16932 bgr_11_0.V_TOP.n34 bgr_11_0.V_TOP.t14 308
R16933 bgr_11_0.V_TOP.n7 bgr_11_0.V_TOP.t29 305.901
R16934 bgr_11_0.V_TOP.n31 bgr_11_0.V_TOP.n30 301.933
R16935 bgr_11_0.V_TOP.n29 bgr_11_0.V_TOP.n28 301.933
R16936 bgr_11_0.V_TOP.n27 bgr_11_0.V_TOP.n26 301.933
R16937 bgr_11_0.V_TOP.n24 bgr_11_0.V_TOP.n20 297.433
R16938 bgr_11_0.V_TOP.n19 bgr_11_0.V_TOP.t13 108.424
R16939 bgr_11_0.V_TOP.n32 bgr_11_0.V_TOP.t8 99.5675
R16940 bgr_11_0.V_TOP.n22 bgr_11_0.V_TOP.t10 39.4005
R16941 bgr_11_0.V_TOP.n22 bgr_11_0.V_TOP.t5 39.4005
R16942 bgr_11_0.V_TOP.n21 bgr_11_0.V_TOP.t7 39.4005
R16943 bgr_11_0.V_TOP.n21 bgr_11_0.V_TOP.t12 39.4005
R16944 bgr_11_0.V_TOP.n20 bgr_11_0.V_TOP.t11 39.4005
R16945 bgr_11_0.V_TOP.n20 bgr_11_0.V_TOP.t1 39.4005
R16946 bgr_11_0.V_TOP.n30 bgr_11_0.V_TOP.t6 39.4005
R16947 bgr_11_0.V_TOP.n30 bgr_11_0.V_TOP.t9 39.4005
R16948 bgr_11_0.V_TOP.n28 bgr_11_0.V_TOP.t3 39.4005
R16949 bgr_11_0.V_TOP.n28 bgr_11_0.V_TOP.t2 39.4005
R16950 bgr_11_0.V_TOP.n26 bgr_11_0.V_TOP.t4 39.4005
R16951 bgr_11_0.V_TOP.n26 bgr_11_0.V_TOP.t0 39.4005
R16952 bgr_11_0.V_TOP.n19 bgr_11_0.V_TOP.n18 29.1779
R16953 bgr_11_0.V_TOP.n25 bgr_11_0.V_TOP.n19 16.5063
R16954 bgr_11_0.V_TOP.n32 bgr_11_0.V_TOP.n31 4.90675
R16955 bgr_11_0.V_TOP.n8 bgr_11_0.V_TOP.t24 4.8295
R16956 bgr_11_0.V_TOP.n9 bgr_11_0.V_TOP.t46 4.8295
R16957 bgr_11_0.V_TOP.n10 bgr_11_0.V_TOP.t34 4.8295
R16958 bgr_11_0.V_TOP.n11 bgr_11_0.V_TOP.t18 4.8295
R16959 bgr_11_0.V_TOP.n12 bgr_11_0.V_TOP.t22 4.8295
R16960 bgr_11_0.V_TOP.n13 bgr_11_0.V_TOP.t44 4.8295
R16961 bgr_11_0.V_TOP.n14 bgr_11_0.V_TOP.t47 4.8295
R16962 bgr_11_0.V_TOP.n15 bgr_11_0.V_TOP.t35 4.8295
R16963 bgr_11_0.V_TOP.n16 bgr_11_0.V_TOP.t41 4.8295
R16964 bgr_11_0.V_TOP.n8 bgr_11_0.V_TOP.t32 4.5005
R16965 bgr_11_0.V_TOP.n9 bgr_11_0.V_TOP.t19 4.5005
R16966 bgr_11_0.V_TOP.n10 bgr_11_0.V_TOP.t40 4.5005
R16967 bgr_11_0.V_TOP.n11 bgr_11_0.V_TOP.t31 4.5005
R16968 bgr_11_0.V_TOP.n12 bgr_11_0.V_TOP.t30 4.5005
R16969 bgr_11_0.V_TOP.n13 bgr_11_0.V_TOP.t17 4.5005
R16970 bgr_11_0.V_TOP.n14 bgr_11_0.V_TOP.t16 4.5005
R16971 bgr_11_0.V_TOP.n15 bgr_11_0.V_TOP.t43 4.5005
R16972 bgr_11_0.V_TOP.n18 bgr_11_0.V_TOP.t20 4.5005
R16973 bgr_11_0.V_TOP.n17 bgr_11_0.V_TOP.t28 4.5005
R16974 bgr_11_0.V_TOP.n16 bgr_11_0.V_TOP.t15 4.5005
R16975 bgr_11_0.V_TOP.n7 bgr_11_0.V_TOP.n6 4.5005
R16976 bgr_11_0.V_TOP.n33 bgr_11_0.V_TOP.n0 4.5005
R16977 bgr_11_0.V_TOP.n35 bgr_11_0.V_TOP.n34 4.5005
R16978 bgr_11_0.V_TOP.n25 bgr_11_0.V_TOP.n24 4.5005
R16979 bgr_11_0.V_TOP.n24 bgr_11_0.V_TOP.n23 1.59425
R16980 bgr_11_0.V_TOP.n33 bgr_11_0.V_TOP.n32 1.21925
R16981 bgr_11_0.V_TOP.n27 bgr_11_0.V_TOP.n25 1.1255
R16982 bgr_11_0.V_TOP.n29 bgr_11_0.V_TOP.n27 1.1255
R16983 bgr_11_0.V_TOP.n31 bgr_11_0.V_TOP.n29 1.1255
R16984 bgr_11_0.V_TOP.n9 bgr_11_0.V_TOP.n8 0.3295
R16985 bgr_11_0.V_TOP.n11 bgr_11_0.V_TOP.n10 0.3295
R16986 bgr_11_0.V_TOP.n13 bgr_11_0.V_TOP.n12 0.3295
R16987 bgr_11_0.V_TOP.n15 bgr_11_0.V_TOP.n14 0.3295
R16988 bgr_11_0.V_TOP.n18 bgr_11_0.V_TOP.n17 0.3295
R16989 bgr_11_0.V_TOP.n17 bgr_11_0.V_TOP.n16 0.3295
R16990 bgr_11_0.V_TOP.n11 bgr_11_0.V_TOP.n9 0.2825
R16991 bgr_11_0.V_TOP.n13 bgr_11_0.V_TOP.n11 0.2825
R16992 bgr_11_0.V_TOP.n15 bgr_11_0.V_TOP.n13 0.2825
R16993 bgr_11_0.V_TOP.n16 bgr_11_0.V_TOP.n15 0.2825
R16994 bgr_11_0.V_TOP.n2 bgr_11_0.V_TOP.n1 0.28175
R16995 bgr_11_0.V_TOP.n3 bgr_11_0.V_TOP.n2 0.28175
R16996 bgr_11_0.V_TOP.n4 bgr_11_0.V_TOP.n3 0.28175
R16997 bgr_11_0.V_TOP.n5 bgr_11_0.V_TOP.n4 0.28175
R16998 bgr_11_0.V_TOP.n6 bgr_11_0.V_TOP.n5 0.28175
R16999 bgr_11_0.V_TOP.n36 bgr_11_0.V_TOP.n35 0.28175
R17000 bgr_11_0.V_TOP.n37 bgr_11_0.V_TOP.n36 0.28175
R17001 bgr_11_0.V_TOP.n38 bgr_11_0.V_TOP.n37 0.28175
R17002 bgr_11_0.V_TOP.n39 bgr_11_0.V_TOP.n38 0.28175
R17003 bgr_11_0.V_TOP.n40 bgr_11_0.V_TOP.n39 0.28175
R17004 bgr_11_0.V_TOP.n41 bgr_11_0.V_TOP.n40 0.28175
R17005 bgr_11_0.V_TOP.n42 bgr_11_0.V_TOP.n41 0.28175
R17006 bgr_11_0.V_TOP.n6 bgr_11_0.V_TOP.n0 0.141125
R17007 bgr_11_0.V_TOP.n35 bgr_11_0.V_TOP.n0 0.141125
R17008 bgr_11_0.V_TOP bgr_11_0.V_TOP.n42 0.141125
R17009 bgr_11_0.V_TOP.n33 bgr_11_0.V_TOP.n7 0.141125
R17010 bgr_11_0.V_TOP.n34 bgr_11_0.V_TOP.n33 0.141125
R17011 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref.n7 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref.t7 651.343
R17012 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref.n7 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref.t8 647.968
R17013 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref.n0 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref.t9 537.922
R17014 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref.n0 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref.t4 117.243
R17015 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref.n3 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref.n1 107.266
R17016 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref.n5 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref.n4 105.016
R17017 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref.n3 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref.n2 105.016
R17018 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref.n4 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref.t2 13.1338
R17019 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref.n4 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref.t6 13.1338
R17020 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref.n2 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref.t3 13.1338
R17021 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref.n2 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref.t0 13.1338
R17022 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref.n1 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref.t5 13.1338
R17023 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref.n1 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref.t1 13.1338
R17024 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref.n6 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref.n5 7.32862
R17025 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref two_stage_opamp_dummy_magic_29_0.V_err_amp_ref.n6 3.98488
R17026 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref.n5 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref.n3 2.2505
R17027 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref.n6 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref.n0 1.73488
R17028 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref two_stage_opamp_dummy_magic_29_0.V_err_amp_ref.n7 1.53175
R17029 two_stage_opamp_dummy_magic_29_0.cap_res_X two_stage_opamp_dummy_magic_29_0.cap_res_X.t143 49.8942
R17030 two_stage_opamp_dummy_magic_29_0.cap_res_X two_stage_opamp_dummy_magic_29_0.cap_res_X.t30 0.9405
R17031 two_stage_opamp_dummy_magic_29_0.cap_res_X.t25 two_stage_opamp_dummy_magic_29_0.cap_res_X.t131 0.1603
R17032 two_stage_opamp_dummy_magic_29_0.cap_res_X.t50 two_stage_opamp_dummy_magic_29_0.cap_res_X.t18 0.1603
R17033 two_stage_opamp_dummy_magic_29_0.cap_res_X.t31 two_stage_opamp_dummy_magic_29_0.cap_res_X.t137 0.1603
R17034 two_stage_opamp_dummy_magic_29_0.cap_res_X.t132 two_stage_opamp_dummy_magic_29_0.cap_res_X.t99 0.1603
R17035 two_stage_opamp_dummy_magic_29_0.cap_res_X.t19 two_stage_opamp_dummy_magic_29_0.cap_res_X.t123 0.1603
R17036 two_stage_opamp_dummy_magic_29_0.cap_res_X.t119 two_stage_opamp_dummy_magic_29_0.cap_res_X.t82 0.1603
R17037 two_stage_opamp_dummy_magic_29_0.cap_res_X.t80 two_stage_opamp_dummy_magic_29_0.cap_res_X.t44 0.1603
R17038 two_stage_opamp_dummy_magic_29_0.cap_res_X.t75 two_stage_opamp_dummy_magic_29_0.cap_res_X.t97 0.1603
R17039 two_stage_opamp_dummy_magic_29_0.cap_res_X.t117 two_stage_opamp_dummy_magic_29_0.cap_res_X.t92 0.1603
R17040 two_stage_opamp_dummy_magic_29_0.cap_res_X.t37 two_stage_opamp_dummy_magic_29_0.cap_res_X.t63 0.1603
R17041 two_stage_opamp_dummy_magic_29_0.cap_res_X.t141 two_stage_opamp_dummy_magic_29_0.cap_res_X.t52 0.1603
R17042 two_stage_opamp_dummy_magic_29_0.cap_res_X.t72 two_stage_opamp_dummy_magic_29_0.cap_res_X.t20 0.1603
R17043 two_stage_opamp_dummy_magic_29_0.cap_res_X.t38 two_stage_opamp_dummy_magic_29_0.cap_res_X.t89 0.1603
R17044 two_stage_opamp_dummy_magic_29_0.cap_res_X.t110 two_stage_opamp_dummy_magic_29_0.cap_res_X.t60 0.1603
R17045 two_stage_opamp_dummy_magic_29_0.cap_res_X.t2 two_stage_opamp_dummy_magic_29_0.cap_res_X.t58 0.1603
R17046 two_stage_opamp_dummy_magic_29_0.cap_res_X.t77 two_stage_opamp_dummy_magic_29_0.cap_res_X.t23 0.1603
R17047 two_stage_opamp_dummy_magic_29_0.cap_res_X.t43 two_stage_opamp_dummy_magic_29_0.cap_res_X.t96 0.1603
R17048 two_stage_opamp_dummy_magic_29_0.cap_res_X.t116 two_stage_opamp_dummy_magic_29_0.cap_res_X.t65 0.1603
R17049 two_stage_opamp_dummy_magic_29_0.cap_res_X.t84 two_stage_opamp_dummy_magic_29_0.cap_res_X.t135 0.1603
R17050 two_stage_opamp_dummy_magic_29_0.cap_res_X.t16 two_stage_opamp_dummy_magic_29_0.cap_res_X.t105 0.1603
R17051 two_stage_opamp_dummy_magic_29_0.cap_res_X.t51 two_stage_opamp_dummy_magic_29_0.cap_res_X.t103 0.1603
R17052 two_stage_opamp_dummy_magic_29_0.cap_res_X.t121 two_stage_opamp_dummy_magic_29_0.cap_res_X.t71 0.1603
R17053 two_stage_opamp_dummy_magic_29_0.cap_res_X.t88 two_stage_opamp_dummy_magic_29_0.cap_res_X.t142 0.1603
R17054 two_stage_opamp_dummy_magic_29_0.cap_res_X.t21 two_stage_opamp_dummy_magic_29_0.cap_res_X.t108 0.1603
R17055 two_stage_opamp_dummy_magic_29_0.cap_res_X.t127 two_stage_opamp_dummy_magic_29_0.cap_res_X.t40 0.1603
R17056 two_stage_opamp_dummy_magic_29_0.cap_res_X.t61 two_stage_opamp_dummy_magic_29_0.cap_res_X.t7 0.1603
R17057 two_stage_opamp_dummy_magic_29_0.cap_res_X.t27 two_stage_opamp_dummy_magic_29_0.cap_res_X.t81 0.1603
R17058 two_stage_opamp_dummy_magic_29_0.cap_res_X.t100 two_stage_opamp_dummy_magic_29_0.cap_res_X.t48 0.1603
R17059 two_stage_opamp_dummy_magic_29_0.cap_res_X.t134 two_stage_opamp_dummy_magic_29_0.cap_res_X.t45 0.1603
R17060 two_stage_opamp_dummy_magic_29_0.cap_res_X.t68 two_stage_opamp_dummy_magic_29_0.cap_res_X.t13 0.1603
R17061 two_stage_opamp_dummy_magic_29_0.cap_res_X.t34 two_stage_opamp_dummy_magic_29_0.cap_res_X.t85 0.1603
R17062 two_stage_opamp_dummy_magic_29_0.cap_res_X.t106 two_stage_opamp_dummy_magic_29_0.cap_res_X.t54 0.1603
R17063 two_stage_opamp_dummy_magic_29_0.cap_res_X.t76 two_stage_opamp_dummy_magic_29_0.cap_res_X.t125 0.1603
R17064 two_stage_opamp_dummy_magic_29_0.cap_res_X.t0 two_stage_opamp_dummy_magic_29_0.cap_res_X.t93 0.1603
R17065 two_stage_opamp_dummy_magic_29_0.cap_res_X.t39 two_stage_opamp_dummy_magic_29_0.cap_res_X.t90 0.1603
R17066 two_stage_opamp_dummy_magic_29_0.cap_res_X.t111 two_stage_opamp_dummy_magic_29_0.cap_res_X.t59 0.1603
R17067 two_stage_opamp_dummy_magic_29_0.cap_res_X.t12 two_stage_opamp_dummy_magic_29_0.cap_res_X.t57 0.1603
R17068 two_stage_opamp_dummy_magic_29_0.cap_res_X.t115 two_stage_opamp_dummy_magic_29_0.cap_res_X.t74 0.1603
R17069 two_stage_opamp_dummy_magic_29_0.cap_res_X.t70 two_stage_opamp_dummy_magic_29_0.cap_res_X.t120 0.1603
R17070 two_stage_opamp_dummy_magic_29_0.cap_res_X.t138 two_stage_opamp_dummy_magic_29_0.cap_res_X.t87 0.1603
R17071 two_stage_opamp_dummy_magic_29_0.cap_res_X.t104 two_stage_opamp_dummy_magic_29_0.cap_res_X.t14 0.1603
R17072 two_stage_opamp_dummy_magic_29_0.cap_res_X.t32 two_stage_opamp_dummy_magic_29_0.cap_res_X.t124 0.1603
R17073 two_stage_opamp_dummy_magic_29_0.cap_res_X.t47 two_stage_opamp_dummy_magic_29_0.cap_res_X.t6 0.1603
R17074 two_stage_opamp_dummy_magic_29_0.cap_res_X.t73 two_stage_opamp_dummy_magic_29_0.cap_res_X.t28 0.1603
R17075 two_stage_opamp_dummy_magic_29_0.cap_res_X.t53 two_stage_opamp_dummy_magic_29_0.cap_res_X.t11 0.1603
R17076 two_stage_opamp_dummy_magic_29_0.cap_res_X.t15 two_stage_opamp_dummy_magic_29_0.cap_res_X.t114 0.1603
R17077 two_stage_opamp_dummy_magic_29_0.cap_res_X.t35 two_stage_opamp_dummy_magic_29_0.cap_res_X.t136 0.1603
R17078 two_stage_opamp_dummy_magic_29_0.cap_res_X.t139 two_stage_opamp_dummy_magic_29_0.cap_res_X.t98 0.1603
R17079 two_stage_opamp_dummy_magic_29_0.cap_res_X.t102 two_stage_opamp_dummy_magic_29_0.cap_res_X.t62 0.1603
R17080 two_stage_opamp_dummy_magic_29_0.cap_res_X.t64 two_stage_opamp_dummy_magic_29_0.cap_res_X.t22 0.1603
R17081 two_stage_opamp_dummy_magic_29_0.cap_res_X.t83 two_stage_opamp_dummy_magic_29_0.cap_res_X.t42 0.1603
R17082 two_stage_opamp_dummy_magic_29_0.cap_res_X.t46 two_stage_opamp_dummy_magic_29_0.cap_res_X.t4 0.1603
R17083 two_stage_opamp_dummy_magic_29_0.cap_res_X.t8 two_stage_opamp_dummy_magic_29_0.cap_res_X.t109 0.1603
R17084 two_stage_opamp_dummy_magic_29_0.cap_res_X.t29 two_stage_opamp_dummy_magic_29_0.cap_res_X.t128 0.1603
R17085 two_stage_opamp_dummy_magic_29_0.cap_res_X.t95 two_stage_opamp_dummy_magic_29_0.cap_res_X.t118 0.1603
R17086 two_stage_opamp_dummy_magic_29_0.cap_res_X.t56 two_stage_opamp_dummy_magic_29_0.cap_res_X.t78 0.1603
R17087 two_stage_opamp_dummy_magic_29_0.cap_res_X.t126 two_stage_opamp_dummy_magic_29_0.cap_res_X.t10 0.1603
R17088 two_stage_opamp_dummy_magic_29_0.cap_res_X.t129 two_stage_opamp_dummy_magic_29_0.cap_res_X.t86 0.1603
R17089 two_stage_opamp_dummy_magic_29_0.cap_res_X.t24 two_stage_opamp_dummy_magic_29_0.cap_res_X.t129 0.1603
R17090 two_stage_opamp_dummy_magic_29_0.cap_res_X.t26 two_stage_opamp_dummy_magic_29_0.cap_res_X.t122 0.1603
R17091 two_stage_opamp_dummy_magic_29_0.cap_res_X.t67 two_stage_opamp_dummy_magic_29_0.cap_res_X.t26 0.1603
R17092 two_stage_opamp_dummy_magic_29_0.cap_res_X.t5 two_stage_opamp_dummy_magic_29_0.cap_res_X.t41 0.1603
R17093 two_stage_opamp_dummy_magic_29_0.cap_res_X.t30 two_stage_opamp_dummy_magic_29_0.cap_res_X.t5 0.1603
R17094 two_stage_opamp_dummy_magic_29_0.cap_res_X.t130 two_stage_opamp_dummy_magic_29_0.cap_res_X.n11 0.159278
R17095 two_stage_opamp_dummy_magic_29_0.cap_res_X.t69 two_stage_opamp_dummy_magic_29_0.cap_res_X.n12 0.159278
R17096 two_stage_opamp_dummy_magic_29_0.cap_res_X.t33 two_stage_opamp_dummy_magic_29_0.cap_res_X.n13 0.159278
R17097 two_stage_opamp_dummy_magic_29_0.cap_res_X.t66 two_stage_opamp_dummy_magic_29_0.cap_res_X.n14 0.159278
R17098 two_stage_opamp_dummy_magic_29_0.cap_res_X.t3 two_stage_opamp_dummy_magic_29_0.cap_res_X.n15 0.159278
R17099 two_stage_opamp_dummy_magic_29_0.cap_res_X.t36 two_stage_opamp_dummy_magic_29_0.cap_res_X.n16 0.159278
R17100 two_stage_opamp_dummy_magic_29_0.cap_res_X.t140 two_stage_opamp_dummy_magic_29_0.cap_res_X.n17 0.159278
R17101 two_stage_opamp_dummy_magic_29_0.cap_res_X.t101 two_stage_opamp_dummy_magic_29_0.cap_res_X.n18 0.159278
R17102 two_stage_opamp_dummy_magic_29_0.cap_res_X.t133 two_stage_opamp_dummy_magic_29_0.cap_res_X.n19 0.159278
R17103 two_stage_opamp_dummy_magic_29_0.cap_res_X.t94 two_stage_opamp_dummy_magic_29_0.cap_res_X.n20 0.159278
R17104 two_stage_opamp_dummy_magic_29_0.cap_res_X.t55 two_stage_opamp_dummy_magic_29_0.cap_res_X.n21 0.159278
R17105 two_stage_opamp_dummy_magic_29_0.cap_res_X.t17 two_stage_opamp_dummy_magic_29_0.cap_res_X.n22 0.159278
R17106 two_stage_opamp_dummy_magic_29_0.cap_res_X.t49 two_stage_opamp_dummy_magic_29_0.cap_res_X.n23 0.159278
R17107 two_stage_opamp_dummy_magic_29_0.cap_res_X.t9 two_stage_opamp_dummy_magic_29_0.cap_res_X.n24 0.159278
R17108 two_stage_opamp_dummy_magic_29_0.cap_res_X.t112 two_stage_opamp_dummy_magic_29_0.cap_res_X.n25 0.159278
R17109 two_stage_opamp_dummy_magic_29_0.cap_res_X.t1 two_stage_opamp_dummy_magic_29_0.cap_res_X.n26 0.159278
R17110 two_stage_opamp_dummy_magic_29_0.cap_res_X.t107 two_stage_opamp_dummy_magic_29_0.cap_res_X.n27 0.159278
R17111 two_stage_opamp_dummy_magic_29_0.cap_res_X.t79 two_stage_opamp_dummy_magic_29_0.cap_res_X.n28 0.159278
R17112 two_stage_opamp_dummy_magic_29_0.cap_res_X.t113 two_stage_opamp_dummy_magic_29_0.cap_res_X.n29 0.159278
R17113 two_stage_opamp_dummy_magic_29_0.cap_res_X.n30 two_stage_opamp_dummy_magic_29_0.cap_res_X.t75 0.1368
R17114 two_stage_opamp_dummy_magic_29_0.cap_res_X.n29 two_stage_opamp_dummy_magic_29_0.cap_res_X.t117 0.1368
R17115 two_stage_opamp_dummy_magic_29_0.cap_res_X.n29 two_stage_opamp_dummy_magic_29_0.cap_res_X.t37 0.1368
R17116 two_stage_opamp_dummy_magic_29_0.cap_res_X.n28 two_stage_opamp_dummy_magic_29_0.cap_res_X.t141 0.1368
R17117 two_stage_opamp_dummy_magic_29_0.cap_res_X.n28 two_stage_opamp_dummy_magic_29_0.cap_res_X.t72 0.1368
R17118 two_stage_opamp_dummy_magic_29_0.cap_res_X.n27 two_stage_opamp_dummy_magic_29_0.cap_res_X.t38 0.1368
R17119 two_stage_opamp_dummy_magic_29_0.cap_res_X.n27 two_stage_opamp_dummy_magic_29_0.cap_res_X.t110 0.1368
R17120 two_stage_opamp_dummy_magic_29_0.cap_res_X.n26 two_stage_opamp_dummy_magic_29_0.cap_res_X.t2 0.1368
R17121 two_stage_opamp_dummy_magic_29_0.cap_res_X.n26 two_stage_opamp_dummy_magic_29_0.cap_res_X.t77 0.1368
R17122 two_stage_opamp_dummy_magic_29_0.cap_res_X.n25 two_stage_opamp_dummy_magic_29_0.cap_res_X.t43 0.1368
R17123 two_stage_opamp_dummy_magic_29_0.cap_res_X.n25 two_stage_opamp_dummy_magic_29_0.cap_res_X.t116 0.1368
R17124 two_stage_opamp_dummy_magic_29_0.cap_res_X.n24 two_stage_opamp_dummy_magic_29_0.cap_res_X.t84 0.1368
R17125 two_stage_opamp_dummy_magic_29_0.cap_res_X.n24 two_stage_opamp_dummy_magic_29_0.cap_res_X.t16 0.1368
R17126 two_stage_opamp_dummy_magic_29_0.cap_res_X.n23 two_stage_opamp_dummy_magic_29_0.cap_res_X.t51 0.1368
R17127 two_stage_opamp_dummy_magic_29_0.cap_res_X.n23 two_stage_opamp_dummy_magic_29_0.cap_res_X.t121 0.1368
R17128 two_stage_opamp_dummy_magic_29_0.cap_res_X.n22 two_stage_opamp_dummy_magic_29_0.cap_res_X.t88 0.1368
R17129 two_stage_opamp_dummy_magic_29_0.cap_res_X.n22 two_stage_opamp_dummy_magic_29_0.cap_res_X.t21 0.1368
R17130 two_stage_opamp_dummy_magic_29_0.cap_res_X.n21 two_stage_opamp_dummy_magic_29_0.cap_res_X.t127 0.1368
R17131 two_stage_opamp_dummy_magic_29_0.cap_res_X.n21 two_stage_opamp_dummy_magic_29_0.cap_res_X.t61 0.1368
R17132 two_stage_opamp_dummy_magic_29_0.cap_res_X.n20 two_stage_opamp_dummy_magic_29_0.cap_res_X.t27 0.1368
R17133 two_stage_opamp_dummy_magic_29_0.cap_res_X.n20 two_stage_opamp_dummy_magic_29_0.cap_res_X.t100 0.1368
R17134 two_stage_opamp_dummy_magic_29_0.cap_res_X.n19 two_stage_opamp_dummy_magic_29_0.cap_res_X.t134 0.1368
R17135 two_stage_opamp_dummy_magic_29_0.cap_res_X.n19 two_stage_opamp_dummy_magic_29_0.cap_res_X.t68 0.1368
R17136 two_stage_opamp_dummy_magic_29_0.cap_res_X.n18 two_stage_opamp_dummy_magic_29_0.cap_res_X.t34 0.1368
R17137 two_stage_opamp_dummy_magic_29_0.cap_res_X.n18 two_stage_opamp_dummy_magic_29_0.cap_res_X.t106 0.1368
R17138 two_stage_opamp_dummy_magic_29_0.cap_res_X.n17 two_stage_opamp_dummy_magic_29_0.cap_res_X.t76 0.1368
R17139 two_stage_opamp_dummy_magic_29_0.cap_res_X.n17 two_stage_opamp_dummy_magic_29_0.cap_res_X.t0 0.1368
R17140 two_stage_opamp_dummy_magic_29_0.cap_res_X.n16 two_stage_opamp_dummy_magic_29_0.cap_res_X.t39 0.1368
R17141 two_stage_opamp_dummy_magic_29_0.cap_res_X.n16 two_stage_opamp_dummy_magic_29_0.cap_res_X.t111 0.1368
R17142 two_stage_opamp_dummy_magic_29_0.cap_res_X.n15 two_stage_opamp_dummy_magic_29_0.cap_res_X.t12 0.1368
R17143 two_stage_opamp_dummy_magic_29_0.cap_res_X.n15 two_stage_opamp_dummy_magic_29_0.cap_res_X.t115 0.1368
R17144 two_stage_opamp_dummy_magic_29_0.cap_res_X.n14 two_stage_opamp_dummy_magic_29_0.cap_res_X.t70 0.1368
R17145 two_stage_opamp_dummy_magic_29_0.cap_res_X.n14 two_stage_opamp_dummy_magic_29_0.cap_res_X.t138 0.1368
R17146 two_stage_opamp_dummy_magic_29_0.cap_res_X.n13 two_stage_opamp_dummy_magic_29_0.cap_res_X.t104 0.1368
R17147 two_stage_opamp_dummy_magic_29_0.cap_res_X.n13 two_stage_opamp_dummy_magic_29_0.cap_res_X.t32 0.1368
R17148 two_stage_opamp_dummy_magic_29_0.cap_res_X.n12 two_stage_opamp_dummy_magic_29_0.cap_res_X.t95 0.1368
R17149 two_stage_opamp_dummy_magic_29_0.cap_res_X.n11 two_stage_opamp_dummy_magic_29_0.cap_res_X.t56 0.1368
R17150 two_stage_opamp_dummy_magic_29_0.cap_res_X.t10 two_stage_opamp_dummy_magic_29_0.cap_res_X.n30 0.1368
R17151 two_stage_opamp_dummy_magic_29_0.cap_res_X.n31 two_stage_opamp_dummy_magic_29_0.cap_res_X.t126 0.1368
R17152 two_stage_opamp_dummy_magic_29_0.cap_res_X.n33 two_stage_opamp_dummy_magic_29_0.cap_res_X.t25 0.114322
R17153 two_stage_opamp_dummy_magic_29_0.cap_res_X.n0 two_stage_opamp_dummy_magic_29_0.cap_res_X.t47 0.114322
R17154 two_stage_opamp_dummy_magic_29_0.cap_res_X.n34 two_stage_opamp_dummy_magic_29_0.cap_res_X.n33 0.1133
R17155 two_stage_opamp_dummy_magic_29_0.cap_res_X.n35 two_stage_opamp_dummy_magic_29_0.cap_res_X.n34 0.1133
R17156 two_stage_opamp_dummy_magic_29_0.cap_res_X.n36 two_stage_opamp_dummy_magic_29_0.cap_res_X.n35 0.1133
R17157 two_stage_opamp_dummy_magic_29_0.cap_res_X.n37 two_stage_opamp_dummy_magic_29_0.cap_res_X.n36 0.1133
R17158 two_stage_opamp_dummy_magic_29_0.cap_res_X.n38 two_stage_opamp_dummy_magic_29_0.cap_res_X.n37 0.1133
R17159 two_stage_opamp_dummy_magic_29_0.cap_res_X.n1 two_stage_opamp_dummy_magic_29_0.cap_res_X.n0 0.1133
R17160 two_stage_opamp_dummy_magic_29_0.cap_res_X.n2 two_stage_opamp_dummy_magic_29_0.cap_res_X.n1 0.1133
R17161 two_stage_opamp_dummy_magic_29_0.cap_res_X.n3 two_stage_opamp_dummy_magic_29_0.cap_res_X.n2 0.1133
R17162 two_stage_opamp_dummy_magic_29_0.cap_res_X.n4 two_stage_opamp_dummy_magic_29_0.cap_res_X.n3 0.1133
R17163 two_stage_opamp_dummy_magic_29_0.cap_res_X.n5 two_stage_opamp_dummy_magic_29_0.cap_res_X.n4 0.1133
R17164 two_stage_opamp_dummy_magic_29_0.cap_res_X.n6 two_stage_opamp_dummy_magic_29_0.cap_res_X.n5 0.1133
R17165 two_stage_opamp_dummy_magic_29_0.cap_res_X.n7 two_stage_opamp_dummy_magic_29_0.cap_res_X.n6 0.1133
R17166 two_stage_opamp_dummy_magic_29_0.cap_res_X.n8 two_stage_opamp_dummy_magic_29_0.cap_res_X.n7 0.1133
R17167 two_stage_opamp_dummy_magic_29_0.cap_res_X.n9 two_stage_opamp_dummy_magic_29_0.cap_res_X.n8 0.1133
R17168 two_stage_opamp_dummy_magic_29_0.cap_res_X.n10 two_stage_opamp_dummy_magic_29_0.cap_res_X.n9 0.1133
R17169 two_stage_opamp_dummy_magic_29_0.cap_res_X.n12 two_stage_opamp_dummy_magic_29_0.cap_res_X.n10 0.1133
R17170 two_stage_opamp_dummy_magic_29_0.cap_res_X.n32 two_stage_opamp_dummy_magic_29_0.cap_res_X.n31 0.1133
R17171 two_stage_opamp_dummy_magic_29_0.cap_res_X.n39 two_stage_opamp_dummy_magic_29_0.cap_res_X.n32 0.1133
R17172 two_stage_opamp_dummy_magic_29_0.cap_res_X.n39 two_stage_opamp_dummy_magic_29_0.cap_res_X.n38 0.1133
R17173 two_stage_opamp_dummy_magic_29_0.cap_res_X.n33 two_stage_opamp_dummy_magic_29_0.cap_res_X.t50 0.00152174
R17174 two_stage_opamp_dummy_magic_29_0.cap_res_X.n34 two_stage_opamp_dummy_magic_29_0.cap_res_X.t31 0.00152174
R17175 two_stage_opamp_dummy_magic_29_0.cap_res_X.n35 two_stage_opamp_dummy_magic_29_0.cap_res_X.t132 0.00152174
R17176 two_stage_opamp_dummy_magic_29_0.cap_res_X.n36 two_stage_opamp_dummy_magic_29_0.cap_res_X.t19 0.00152174
R17177 two_stage_opamp_dummy_magic_29_0.cap_res_X.n37 two_stage_opamp_dummy_magic_29_0.cap_res_X.t119 0.00152174
R17178 two_stage_opamp_dummy_magic_29_0.cap_res_X.n38 two_stage_opamp_dummy_magic_29_0.cap_res_X.t80 0.00152174
R17179 two_stage_opamp_dummy_magic_29_0.cap_res_X.n0 two_stage_opamp_dummy_magic_29_0.cap_res_X.t73 0.00152174
R17180 two_stage_opamp_dummy_magic_29_0.cap_res_X.n1 two_stage_opamp_dummy_magic_29_0.cap_res_X.t53 0.00152174
R17181 two_stage_opamp_dummy_magic_29_0.cap_res_X.n2 two_stage_opamp_dummy_magic_29_0.cap_res_X.t15 0.00152174
R17182 two_stage_opamp_dummy_magic_29_0.cap_res_X.n3 two_stage_opamp_dummy_magic_29_0.cap_res_X.t35 0.00152174
R17183 two_stage_opamp_dummy_magic_29_0.cap_res_X.n4 two_stage_opamp_dummy_magic_29_0.cap_res_X.t139 0.00152174
R17184 two_stage_opamp_dummy_magic_29_0.cap_res_X.n5 two_stage_opamp_dummy_magic_29_0.cap_res_X.t102 0.00152174
R17185 two_stage_opamp_dummy_magic_29_0.cap_res_X.n6 two_stage_opamp_dummy_magic_29_0.cap_res_X.t64 0.00152174
R17186 two_stage_opamp_dummy_magic_29_0.cap_res_X.n7 two_stage_opamp_dummy_magic_29_0.cap_res_X.t83 0.00152174
R17187 two_stage_opamp_dummy_magic_29_0.cap_res_X.n8 two_stage_opamp_dummy_magic_29_0.cap_res_X.t46 0.00152174
R17188 two_stage_opamp_dummy_magic_29_0.cap_res_X.n9 two_stage_opamp_dummy_magic_29_0.cap_res_X.t8 0.00152174
R17189 two_stage_opamp_dummy_magic_29_0.cap_res_X.n10 two_stage_opamp_dummy_magic_29_0.cap_res_X.t29 0.00152174
R17190 two_stage_opamp_dummy_magic_29_0.cap_res_X.n11 two_stage_opamp_dummy_magic_29_0.cap_res_X.t91 0.00152174
R17191 two_stage_opamp_dummy_magic_29_0.cap_res_X.n12 two_stage_opamp_dummy_magic_29_0.cap_res_X.t130 0.00152174
R17192 two_stage_opamp_dummy_magic_29_0.cap_res_X.n13 two_stage_opamp_dummy_magic_29_0.cap_res_X.t69 0.00152174
R17193 two_stage_opamp_dummy_magic_29_0.cap_res_X.n14 two_stage_opamp_dummy_magic_29_0.cap_res_X.t33 0.00152174
R17194 two_stage_opamp_dummy_magic_29_0.cap_res_X.n15 two_stage_opamp_dummy_magic_29_0.cap_res_X.t66 0.00152174
R17195 two_stage_opamp_dummy_magic_29_0.cap_res_X.n16 two_stage_opamp_dummy_magic_29_0.cap_res_X.t3 0.00152174
R17196 two_stage_opamp_dummy_magic_29_0.cap_res_X.n17 two_stage_opamp_dummy_magic_29_0.cap_res_X.t36 0.00152174
R17197 two_stage_opamp_dummy_magic_29_0.cap_res_X.n18 two_stage_opamp_dummy_magic_29_0.cap_res_X.t140 0.00152174
R17198 two_stage_opamp_dummy_magic_29_0.cap_res_X.n19 two_stage_opamp_dummy_magic_29_0.cap_res_X.t101 0.00152174
R17199 two_stage_opamp_dummy_magic_29_0.cap_res_X.n20 two_stage_opamp_dummy_magic_29_0.cap_res_X.t133 0.00152174
R17200 two_stage_opamp_dummy_magic_29_0.cap_res_X.n21 two_stage_opamp_dummy_magic_29_0.cap_res_X.t94 0.00152174
R17201 two_stage_opamp_dummy_magic_29_0.cap_res_X.n22 two_stage_opamp_dummy_magic_29_0.cap_res_X.t55 0.00152174
R17202 two_stage_opamp_dummy_magic_29_0.cap_res_X.n23 two_stage_opamp_dummy_magic_29_0.cap_res_X.t17 0.00152174
R17203 two_stage_opamp_dummy_magic_29_0.cap_res_X.n24 two_stage_opamp_dummy_magic_29_0.cap_res_X.t49 0.00152174
R17204 two_stage_opamp_dummy_magic_29_0.cap_res_X.n25 two_stage_opamp_dummy_magic_29_0.cap_res_X.t9 0.00152174
R17205 two_stage_opamp_dummy_magic_29_0.cap_res_X.n26 two_stage_opamp_dummy_magic_29_0.cap_res_X.t112 0.00152174
R17206 two_stage_opamp_dummy_magic_29_0.cap_res_X.n27 two_stage_opamp_dummy_magic_29_0.cap_res_X.t1 0.00152174
R17207 two_stage_opamp_dummy_magic_29_0.cap_res_X.n28 two_stage_opamp_dummy_magic_29_0.cap_res_X.t107 0.00152174
R17208 two_stage_opamp_dummy_magic_29_0.cap_res_X.n29 two_stage_opamp_dummy_magic_29_0.cap_res_X.t79 0.00152174
R17209 two_stage_opamp_dummy_magic_29_0.cap_res_X.n30 two_stage_opamp_dummy_magic_29_0.cap_res_X.t113 0.00152174
R17210 two_stage_opamp_dummy_magic_29_0.cap_res_X.n31 two_stage_opamp_dummy_magic_29_0.cap_res_X.t24 0.00152174
R17211 two_stage_opamp_dummy_magic_29_0.cap_res_X.n32 two_stage_opamp_dummy_magic_29_0.cap_res_X.t67 0.00152174
R17212 two_stage_opamp_dummy_magic_29_0.cap_res_X.t41 two_stage_opamp_dummy_magic_29_0.cap_res_X.n39 0.00152174
R17213 two_stage_opamp_dummy_magic_29_0.X.n70 two_stage_opamp_dummy_magic_29_0.X.t37 1172.87
R17214 two_stage_opamp_dummy_magic_29_0.X.n66 two_stage_opamp_dummy_magic_29_0.X.t32 1172.87
R17215 two_stage_opamp_dummy_magic_29_0.X.n70 two_stage_opamp_dummy_magic_29_0.X.t54 996.134
R17216 two_stage_opamp_dummy_magic_29_0.X.n71 two_stage_opamp_dummy_magic_29_0.X.t42 996.134
R17217 two_stage_opamp_dummy_magic_29_0.X.n72 two_stage_opamp_dummy_magic_29_0.X.t53 996.134
R17218 two_stage_opamp_dummy_magic_29_0.X.n73 two_stage_opamp_dummy_magic_29_0.X.t41 996.134
R17219 two_stage_opamp_dummy_magic_29_0.X.n69 two_stage_opamp_dummy_magic_29_0.X.t27 996.134
R17220 two_stage_opamp_dummy_magic_29_0.X.n68 two_stage_opamp_dummy_magic_29_0.X.t45 996.134
R17221 two_stage_opamp_dummy_magic_29_0.X.n67 two_stage_opamp_dummy_magic_29_0.X.t30 996.134
R17222 two_stage_opamp_dummy_magic_29_0.X.n66 two_stage_opamp_dummy_magic_29_0.X.t47 996.134
R17223 two_stage_opamp_dummy_magic_29_0.X.n37 two_stage_opamp_dummy_magic_29_0.X.t33 690.867
R17224 two_stage_opamp_dummy_magic_29_0.X.n36 two_stage_opamp_dummy_magic_29_0.X.t29 690.867
R17225 two_stage_opamp_dummy_magic_29_0.X.n46 two_stage_opamp_dummy_magic_29_0.X.t34 530.201
R17226 two_stage_opamp_dummy_magic_29_0.X.n45 two_stage_opamp_dummy_magic_29_0.X.t31 530.201
R17227 two_stage_opamp_dummy_magic_29_0.X.n43 two_stage_opamp_dummy_magic_29_0.X.t26 514.134
R17228 two_stage_opamp_dummy_magic_29_0.X.n42 two_stage_opamp_dummy_magic_29_0.X.t40 514.134
R17229 two_stage_opamp_dummy_magic_29_0.X.n41 two_stage_opamp_dummy_magic_29_0.X.t52 514.134
R17230 two_stage_opamp_dummy_magic_29_0.X.n40 two_stage_opamp_dummy_magic_29_0.X.t35 514.134
R17231 two_stage_opamp_dummy_magic_29_0.X.n39 two_stage_opamp_dummy_magic_29_0.X.t48 514.134
R17232 two_stage_opamp_dummy_magic_29_0.X.n38 two_stage_opamp_dummy_magic_29_0.X.t36 514.134
R17233 two_stage_opamp_dummy_magic_29_0.X.n37 two_stage_opamp_dummy_magic_29_0.X.t49 514.134
R17234 two_stage_opamp_dummy_magic_29_0.X.n36 two_stage_opamp_dummy_magic_29_0.X.t44 514.134
R17235 two_stage_opamp_dummy_magic_29_0.X.n46 two_stage_opamp_dummy_magic_29_0.X.t51 353.467
R17236 two_stage_opamp_dummy_magic_29_0.X.n47 two_stage_opamp_dummy_magic_29_0.X.t39 353.467
R17237 two_stage_opamp_dummy_magic_29_0.X.n48 two_stage_opamp_dummy_magic_29_0.X.t50 353.467
R17238 two_stage_opamp_dummy_magic_29_0.X.n49 two_stage_opamp_dummy_magic_29_0.X.t38 353.467
R17239 two_stage_opamp_dummy_magic_29_0.X.n50 two_stage_opamp_dummy_magic_29_0.X.t25 353.467
R17240 two_stage_opamp_dummy_magic_29_0.X.n51 two_stage_opamp_dummy_magic_29_0.X.t43 353.467
R17241 two_stage_opamp_dummy_magic_29_0.X.n52 two_stage_opamp_dummy_magic_29_0.X.t28 353.467
R17242 two_stage_opamp_dummy_magic_29_0.X.n45 two_stage_opamp_dummy_magic_29_0.X.t46 353.467
R17243 two_stage_opamp_dummy_magic_29_0.X.n69 two_stage_opamp_dummy_magic_29_0.X.n68 176.733
R17244 two_stage_opamp_dummy_magic_29_0.X.n68 two_stage_opamp_dummy_magic_29_0.X.n67 176.733
R17245 two_stage_opamp_dummy_magic_29_0.X.n67 two_stage_opamp_dummy_magic_29_0.X.n66 176.733
R17246 two_stage_opamp_dummy_magic_29_0.X.n71 two_stage_opamp_dummy_magic_29_0.X.n70 176.733
R17247 two_stage_opamp_dummy_magic_29_0.X.n72 two_stage_opamp_dummy_magic_29_0.X.n71 176.733
R17248 two_stage_opamp_dummy_magic_29_0.X.n73 two_stage_opamp_dummy_magic_29_0.X.n72 176.733
R17249 two_stage_opamp_dummy_magic_29_0.X.n47 two_stage_opamp_dummy_magic_29_0.X.n46 176.733
R17250 two_stage_opamp_dummy_magic_29_0.X.n48 two_stage_opamp_dummy_magic_29_0.X.n47 176.733
R17251 two_stage_opamp_dummy_magic_29_0.X.n49 two_stage_opamp_dummy_magic_29_0.X.n48 176.733
R17252 two_stage_opamp_dummy_magic_29_0.X.n50 two_stage_opamp_dummy_magic_29_0.X.n49 176.733
R17253 two_stage_opamp_dummy_magic_29_0.X.n51 two_stage_opamp_dummy_magic_29_0.X.n50 176.733
R17254 two_stage_opamp_dummy_magic_29_0.X.n52 two_stage_opamp_dummy_magic_29_0.X.n51 176.733
R17255 two_stage_opamp_dummy_magic_29_0.X.n38 two_stage_opamp_dummy_magic_29_0.X.n37 176.733
R17256 two_stage_opamp_dummy_magic_29_0.X.n39 two_stage_opamp_dummy_magic_29_0.X.n38 176.733
R17257 two_stage_opamp_dummy_magic_29_0.X.n40 two_stage_opamp_dummy_magic_29_0.X.n39 176.733
R17258 two_stage_opamp_dummy_magic_29_0.X.n41 two_stage_opamp_dummy_magic_29_0.X.n40 176.733
R17259 two_stage_opamp_dummy_magic_29_0.X.n42 two_stage_opamp_dummy_magic_29_0.X.n41 176.733
R17260 two_stage_opamp_dummy_magic_29_0.X.n43 two_stage_opamp_dummy_magic_29_0.X.n42 176.733
R17261 two_stage_opamp_dummy_magic_29_0.X.n54 two_stage_opamp_dummy_magic_29_0.X.n53 165.472
R17262 two_stage_opamp_dummy_magic_29_0.X.n54 two_stage_opamp_dummy_magic_29_0.X.n44 165.472
R17263 two_stage_opamp_dummy_magic_29_0.X.n76 two_stage_opamp_dummy_magic_29_0.X.n75 152
R17264 two_stage_opamp_dummy_magic_29_0.X.n77 two_stage_opamp_dummy_magic_29_0.X.n76 131.571
R17265 two_stage_opamp_dummy_magic_29_0.X.n76 two_stage_opamp_dummy_magic_29_0.X.n74 124.517
R17266 two_stage_opamp_dummy_magic_29_0.X.n81 two_stage_opamp_dummy_magic_29_0.X.n54 74.5362
R17267 two_stage_opamp_dummy_magic_29_0.X.n13 two_stage_opamp_dummy_magic_29_0.X.n12 66.0338
R17268 two_stage_opamp_dummy_magic_29_0.X.n29 two_stage_opamp_dummy_magic_29_0.X.n28 66.0338
R17269 two_stage_opamp_dummy_magic_29_0.X.n26 two_stage_opamp_dummy_magic_29_0.X.n25 66.0338
R17270 two_stage_opamp_dummy_magic_29_0.X.n23 two_stage_opamp_dummy_magic_29_0.X.n22 66.0338
R17271 two_stage_opamp_dummy_magic_29_0.X.n19 two_stage_opamp_dummy_magic_29_0.X.n18 66.0338
R17272 two_stage_opamp_dummy_magic_29_0.X.n16 two_stage_opamp_dummy_magic_29_0.X.n15 66.0338
R17273 two_stage_opamp_dummy_magic_29_0.X.n110 two_stage_opamp_dummy_magic_29_0.X.n108 54.7984
R17274 two_stage_opamp_dummy_magic_29_0.X.n118 two_stage_opamp_dummy_magic_29_0.X.n117 54.4547
R17275 two_stage_opamp_dummy_magic_29_0.X.n116 two_stage_opamp_dummy_magic_29_0.X.n115 54.4547
R17276 two_stage_opamp_dummy_magic_29_0.X.n114 two_stage_opamp_dummy_magic_29_0.X.n113 54.4547
R17277 two_stage_opamp_dummy_magic_29_0.X.n112 two_stage_opamp_dummy_magic_29_0.X.n111 54.4547
R17278 two_stage_opamp_dummy_magic_29_0.X.n110 two_stage_opamp_dummy_magic_29_0.X.n109 54.4547
R17279 two_stage_opamp_dummy_magic_29_0.X.n60 two_stage_opamp_dummy_magic_29_0.X.t8 41.0384
R17280 two_stage_opamp_dummy_magic_29_0.X.n74 two_stage_opamp_dummy_magic_29_0.X.n69 40.1672
R17281 two_stage_opamp_dummy_magic_29_0.X.n74 two_stage_opamp_dummy_magic_29_0.X.n73 40.1672
R17282 two_stage_opamp_dummy_magic_29_0.X.n53 two_stage_opamp_dummy_magic_29_0.X.n45 40.1672
R17283 two_stage_opamp_dummy_magic_29_0.X.n53 two_stage_opamp_dummy_magic_29_0.X.n52 40.1672
R17284 two_stage_opamp_dummy_magic_29_0.X.n44 two_stage_opamp_dummy_magic_29_0.X.n36 40.1672
R17285 two_stage_opamp_dummy_magic_29_0.X.n44 two_stage_opamp_dummy_magic_29_0.X.n43 40.1672
R17286 two_stage_opamp_dummy_magic_29_0.X.n78 two_stage_opamp_dummy_magic_29_0.X.n77 16.3217
R17287 two_stage_opamp_dummy_magic_29_0.X.n117 two_stage_opamp_dummy_magic_29_0.X.t0 16.0005
R17288 two_stage_opamp_dummy_magic_29_0.X.n117 two_stage_opamp_dummy_magic_29_0.X.t6 16.0005
R17289 two_stage_opamp_dummy_magic_29_0.X.n115 two_stage_opamp_dummy_magic_29_0.X.t1 16.0005
R17290 two_stage_opamp_dummy_magic_29_0.X.n115 two_stage_opamp_dummy_magic_29_0.X.t22 16.0005
R17291 two_stage_opamp_dummy_magic_29_0.X.n113 two_stage_opamp_dummy_magic_29_0.X.t4 16.0005
R17292 two_stage_opamp_dummy_magic_29_0.X.n113 two_stage_opamp_dummy_magic_29_0.X.t5 16.0005
R17293 two_stage_opamp_dummy_magic_29_0.X.n111 two_stage_opamp_dummy_magic_29_0.X.t24 16.0005
R17294 two_stage_opamp_dummy_magic_29_0.X.n111 two_stage_opamp_dummy_magic_29_0.X.t3 16.0005
R17295 two_stage_opamp_dummy_magic_29_0.X.n109 two_stage_opamp_dummy_magic_29_0.X.t11 16.0005
R17296 two_stage_opamp_dummy_magic_29_0.X.n109 two_stage_opamp_dummy_magic_29_0.X.t9 16.0005
R17297 two_stage_opamp_dummy_magic_29_0.X.n108 two_stage_opamp_dummy_magic_29_0.X.t7 16.0005
R17298 two_stage_opamp_dummy_magic_29_0.X.n108 two_stage_opamp_dummy_magic_29_0.X.t10 16.0005
R17299 two_stage_opamp_dummy_magic_29_0.X.n75 two_stage_opamp_dummy_magic_29_0.X.n65 12.8005
R17300 two_stage_opamp_dummy_magic_29_0.X.n12 two_stage_opamp_dummy_magic_29_0.X.t2 11.2576
R17301 two_stage_opamp_dummy_magic_29_0.X.n12 two_stage_opamp_dummy_magic_29_0.X.t20 11.2576
R17302 two_stage_opamp_dummy_magic_29_0.X.n28 two_stage_opamp_dummy_magic_29_0.X.t12 11.2576
R17303 two_stage_opamp_dummy_magic_29_0.X.n28 two_stage_opamp_dummy_magic_29_0.X.t23 11.2576
R17304 two_stage_opamp_dummy_magic_29_0.X.n25 two_stage_opamp_dummy_magic_29_0.X.t17 11.2576
R17305 two_stage_opamp_dummy_magic_29_0.X.n25 two_stage_opamp_dummy_magic_29_0.X.t14 11.2576
R17306 two_stage_opamp_dummy_magic_29_0.X.n22 two_stage_opamp_dummy_magic_29_0.X.t13 11.2576
R17307 two_stage_opamp_dummy_magic_29_0.X.n22 two_stage_opamp_dummy_magic_29_0.X.t16 11.2576
R17308 two_stage_opamp_dummy_magic_29_0.X.n18 two_stage_opamp_dummy_magic_29_0.X.t19 11.2576
R17309 two_stage_opamp_dummy_magic_29_0.X.n18 two_stage_opamp_dummy_magic_29_0.X.t18 11.2576
R17310 two_stage_opamp_dummy_magic_29_0.X.n15 two_stage_opamp_dummy_magic_29_0.X.t15 11.2576
R17311 two_stage_opamp_dummy_magic_29_0.X.n15 two_stage_opamp_dummy_magic_29_0.X.t21 11.2576
R17312 two_stage_opamp_dummy_magic_29_0.X.n119 two_stage_opamp_dummy_magic_29_0.X.n118 11.1099
R17313 two_stage_opamp_dummy_magic_29_0.X.n75 two_stage_opamp_dummy_magic_29_0.X.n63 9.36264
R17314 two_stage_opamp_dummy_magic_29_0.X.n65 two_stage_opamp_dummy_magic_29_0.X.n64 9.3005
R17315 two_stage_opamp_dummy_magic_29_0.X.n103 two_stage_opamp_dummy_magic_29_0.X.n3 5.78175
R17316 two_stage_opamp_dummy_magic_29_0.X.n29 two_stage_opamp_dummy_magic_29_0.X.n27 5.66717
R17317 two_stage_opamp_dummy_magic_29_0.X.n14 two_stage_opamp_dummy_magic_29_0.X.n13 5.66717
R17318 two_stage_opamp_dummy_magic_29_0.X.n17 two_stage_opamp_dummy_magic_29_0.X.n13 5.66717
R17319 two_stage_opamp_dummy_magic_29_0.X.n120 two_stage_opamp_dummy_magic_29_0.X.n119 5.46373
R17320 two_stage_opamp_dummy_magic_29_0.X.n103 two_stage_opamp_dummy_magic_29_0.X.n102 5.438
R17321 two_stage_opamp_dummy_magic_29_0.X.n104 two_stage_opamp_dummy_magic_29_0.X.n2 5.438
R17322 two_stage_opamp_dummy_magic_29_0.X.n123 two_stage_opamp_dummy_magic_29_0.X.n105 5.438
R17323 two_stage_opamp_dummy_magic_29_0.X.n107 two_stage_opamp_dummy_magic_29_0.X.n106 5.438
R17324 two_stage_opamp_dummy_magic_29_0.X.n77 two_stage_opamp_dummy_magic_29_0.X.n65 5.33141
R17325 two_stage_opamp_dummy_magic_29_0.X.n30 two_stage_opamp_dummy_magic_29_0.X.n29 5.29217
R17326 two_stage_opamp_dummy_magic_29_0.X.n26 two_stage_opamp_dummy_magic_29_0.X.n10 5.29217
R17327 two_stage_opamp_dummy_magic_29_0.X.n27 two_stage_opamp_dummy_magic_29_0.X.n26 5.29217
R17328 two_stage_opamp_dummy_magic_29_0.X.n23 two_stage_opamp_dummy_magic_29_0.X.n21 5.29217
R17329 two_stage_opamp_dummy_magic_29_0.X.n24 two_stage_opamp_dummy_magic_29_0.X.n23 5.29217
R17330 two_stage_opamp_dummy_magic_29_0.X.n20 two_stage_opamp_dummy_magic_29_0.X.n19 5.29217
R17331 two_stage_opamp_dummy_magic_29_0.X.n19 two_stage_opamp_dummy_magic_29_0.X.n11 5.29217
R17332 two_stage_opamp_dummy_magic_29_0.X.n17 two_stage_opamp_dummy_magic_29_0.X.n16 5.29217
R17333 two_stage_opamp_dummy_magic_29_0.X.n16 two_stage_opamp_dummy_magic_29_0.X.n14 5.29217
R17334 two_stage_opamp_dummy_magic_29_0.X.n93 two_stage_opamp_dummy_magic_29_0.X.n9 4.5005
R17335 two_stage_opamp_dummy_magic_29_0.X.n93 two_stage_opamp_dummy_magic_29_0.X.n90 4.5005
R17336 two_stage_opamp_dummy_magic_29_0.X.n93 two_stage_opamp_dummy_magic_29_0.X.n88 4.5005
R17337 two_stage_opamp_dummy_magic_29_0.X.n93 two_stage_opamp_dummy_magic_29_0.X.n92 4.5005
R17338 two_stage_opamp_dummy_magic_29_0.X.n86 two_stage_opamp_dummy_magic_29_0.X.n31 4.5005
R17339 two_stage_opamp_dummy_magic_29_0.X.n80 two_stage_opamp_dummy_magic_29_0.X.n33 4.5005
R17340 two_stage_opamp_dummy_magic_29_0.X.n82 two_stage_opamp_dummy_magic_29_0.X.n81 4.5005
R17341 two_stage_opamp_dummy_magic_29_0.X.n81 two_stage_opamp_dummy_magic_29_0.X.n80 4.5005
R17342 two_stage_opamp_dummy_magic_29_0.X.n79 two_stage_opamp_dummy_magic_29_0.X.n78 4.5005
R17343 two_stage_opamp_dummy_magic_29_0.X.n57 two_stage_opamp_dummy_magic_29_0.X.n56 4.5005
R17344 two_stage_opamp_dummy_magic_29_0.X.n95 two_stage_opamp_dummy_magic_29_0.X.n30 2.35465
R17345 two_stage_opamp_dummy_magic_29_0.X.n59 two_stage_opamp_dummy_magic_29_0.X.n58 2.26187
R17346 two_stage_opamp_dummy_magic_29_0.X.n58 two_stage_opamp_dummy_magic_29_0.X.n55 2.26187
R17347 two_stage_opamp_dummy_magic_29_0.X.n95 two_stage_opamp_dummy_magic_29_0.X.n94 2.24654
R17348 two_stage_opamp_dummy_magic_29_0.X.n85 two_stage_opamp_dummy_magic_29_0.X.n6 2.24654
R17349 two_stage_opamp_dummy_magic_29_0.X.n89 two_stage_opamp_dummy_magic_29_0.X.n31 2.24063
R17350 two_stage_opamp_dummy_magic_29_0.X.n91 two_stage_opamp_dummy_magic_29_0.X.n31 2.24063
R17351 two_stage_opamp_dummy_magic_29_0.X.n93 two_stage_opamp_dummy_magic_29_0.X.n87 2.24063
R17352 two_stage_opamp_dummy_magic_29_0.X.n83 two_stage_opamp_dummy_magic_29_0.X.n82 2.24063
R17353 two_stage_opamp_dummy_magic_29_0.X.n35 two_stage_opamp_dummy_magic_29_0.X.n34 2.24063
R17354 two_stage_opamp_dummy_magic_29_0.X.n97 two_stage_opamp_dummy_magic_29_0.X.n96 2.24063
R17355 two_stage_opamp_dummy_magic_29_0.X.n97 two_stage_opamp_dummy_magic_29_0.X.n8 2.24063
R17356 two_stage_opamp_dummy_magic_29_0.X.n97 two_stage_opamp_dummy_magic_29_0.X.n7 2.24063
R17357 two_stage_opamp_dummy_magic_29_0.X.n84 two_stage_opamp_dummy_magic_29_0.X.n32 2.24063
R17358 two_stage_opamp_dummy_magic_29_0.X.n60 two_stage_opamp_dummy_magic_29_0.X.n59 2.24063
R17359 two_stage_opamp_dummy_magic_29_0.X.n62 two_stage_opamp_dummy_magic_29_0.X.n61 2.24063
R17360 two_stage_opamp_dummy_magic_29_0.X.n79 two_stage_opamp_dummy_magic_29_0.X.n63 2.22018
R17361 two_stage_opamp_dummy_magic_29_0.X.n79 two_stage_opamp_dummy_magic_29_0.X.n62 0.682792
R17362 two_stage_opamp_dummy_magic_29_0.X.n122 two_stage_opamp_dummy_magic_29_0.X.n121 0.643357
R17363 two_stage_opamp_dummy_magic_29_0.X.n123 two_stage_opamp_dummy_magic_29_0.X.n1 0.643357
R17364 two_stage_opamp_dummy_magic_29_0.X.n125 two_stage_opamp_dummy_magic_29_0.X.n124 0.643357
R17365 two_stage_opamp_dummy_magic_29_0.X.n2 two_stage_opamp_dummy_magic_29_0.X.n0 0.643357
R17366 two_stage_opamp_dummy_magic_29_0.X.n100 two_stage_opamp_dummy_magic_29_0.X.n5 0.643357
R17367 two_stage_opamp_dummy_magic_29_0.X.n102 two_stage_opamp_dummy_magic_29_0.X.n101 0.643357
R17368 two_stage_opamp_dummy_magic_29_0.X.n99 two_stage_opamp_dummy_magic_29_0.X.n4 0.643357
R17369 two_stage_opamp_dummy_magic_29_0.X.n98 two_stage_opamp_dummy_magic_29_0.X.n3 0.643357
R17370 two_stage_opamp_dummy_magic_29_0.X.n85 two_stage_opamp_dummy_magic_29_0.X.n84 0.479667
R17371 two_stage_opamp_dummy_magic_29_0.X.n80 two_stage_opamp_dummy_magic_29_0.X.n79 0.46925
R17372 two_stage_opamp_dummy_magic_29_0.X.n14 two_stage_opamp_dummy_magic_29_0.X.n11 0.3755
R17373 two_stage_opamp_dummy_magic_29_0.X.n24 two_stage_opamp_dummy_magic_29_0.X.n11 0.3755
R17374 two_stage_opamp_dummy_magic_29_0.X.n27 two_stage_opamp_dummy_magic_29_0.X.n24 0.3755
R17375 two_stage_opamp_dummy_magic_29_0.X.n20 two_stage_opamp_dummy_magic_29_0.X.n17 0.3755
R17376 two_stage_opamp_dummy_magic_29_0.X.n21 two_stage_opamp_dummy_magic_29_0.X.n20 0.3755
R17377 two_stage_opamp_dummy_magic_29_0.X.n21 two_stage_opamp_dummy_magic_29_0.X.n10 0.3755
R17378 two_stage_opamp_dummy_magic_29_0.X.n30 two_stage_opamp_dummy_magic_29_0.X.n10 0.3755
R17379 two_stage_opamp_dummy_magic_29_0.X.n112 two_stage_opamp_dummy_magic_29_0.X.n110 0.34425
R17380 two_stage_opamp_dummy_magic_29_0.X.n114 two_stage_opamp_dummy_magic_29_0.X.n112 0.34425
R17381 two_stage_opamp_dummy_magic_29_0.X.n116 two_stage_opamp_dummy_magic_29_0.X.n114 0.34425
R17382 two_stage_opamp_dummy_magic_29_0.X.n118 two_stage_opamp_dummy_magic_29_0.X.n116 0.34425
R17383 two_stage_opamp_dummy_magic_29_0.X.n104 two_stage_opamp_dummy_magic_29_0.X.n103 0.34425
R17384 two_stage_opamp_dummy_magic_29_0.X.n105 two_stage_opamp_dummy_magic_29_0.X.n104 0.34425
R17385 two_stage_opamp_dummy_magic_29_0.X.n107 two_stage_opamp_dummy_magic_29_0.X.n105 0.34425
R17386 two_stage_opamp_dummy_magic_29_0.X.n119 two_stage_opamp_dummy_magic_29_0.X.n107 0.34425
R17387 two_stage_opamp_dummy_magic_29_0.X.n98 two_stage_opamp_dummy_magic_29_0.X.n97 0.270589
R17388 two_stage_opamp_dummy_magic_29_0.X.n121 two_stage_opamp_dummy_magic_29_0.X.n120 0.242602
R17389 two_stage_opamp_dummy_magic_29_0.X.n78 two_stage_opamp_dummy_magic_29_0.X.n64 0.1255
R17390 two_stage_opamp_dummy_magic_29_0.X.n64 two_stage_opamp_dummy_magic_29_0.X.n63 0.0626438
R17391 two_stage_opamp_dummy_magic_29_0.X.n82 two_stage_opamp_dummy_magic_29_0.X.n34 0.0421667
R17392 two_stage_opamp_dummy_magic_29_0.X.n4 two_stage_opamp_dummy_magic_29_0.X.n3 0.0250536
R17393 two_stage_opamp_dummy_magic_29_0.X.n102 two_stage_opamp_dummy_magic_29_0.X.n4 0.0250536
R17394 two_stage_opamp_dummy_magic_29_0.X.n102 two_stage_opamp_dummy_magic_29_0.X.n5 0.0250536
R17395 two_stage_opamp_dummy_magic_29_0.X.n5 two_stage_opamp_dummy_magic_29_0.X.n2 0.0250536
R17396 two_stage_opamp_dummy_magic_29_0.X.n124 two_stage_opamp_dummy_magic_29_0.X.n2 0.0250536
R17397 two_stage_opamp_dummy_magic_29_0.X.n124 two_stage_opamp_dummy_magic_29_0.X.n123 0.0250536
R17398 two_stage_opamp_dummy_magic_29_0.X.n123 two_stage_opamp_dummy_magic_29_0.X.n122 0.0250536
R17399 two_stage_opamp_dummy_magic_29_0.X.n122 two_stage_opamp_dummy_magic_29_0.X.n106 0.0250536
R17400 two_stage_opamp_dummy_magic_29_0.X.n99 two_stage_opamp_dummy_magic_29_0.X.n98 0.0250536
R17401 two_stage_opamp_dummy_magic_29_0.X.n101 two_stage_opamp_dummy_magic_29_0.X.n99 0.0250536
R17402 two_stage_opamp_dummy_magic_29_0.X.n101 two_stage_opamp_dummy_magic_29_0.X.n100 0.0250536
R17403 two_stage_opamp_dummy_magic_29_0.X.n100 two_stage_opamp_dummy_magic_29_0.X.n0 0.0250536
R17404 two_stage_opamp_dummy_magic_29_0.X.n125 two_stage_opamp_dummy_magic_29_0.X.n1 0.0250536
R17405 two_stage_opamp_dummy_magic_29_0.X.n121 two_stage_opamp_dummy_magic_29_0.X.n1 0.0250536
R17406 two_stage_opamp_dummy_magic_29_0.X.n120 two_stage_opamp_dummy_magic_29_0.X.n106 0.0241021
R17407 two_stage_opamp_dummy_magic_29_0.X.n90 two_stage_opamp_dummy_magic_29_0.X.n89 0.0217373
R17408 two_stage_opamp_dummy_magic_29_0.X.n92 two_stage_opamp_dummy_magic_29_0.X.n91 0.0217373
R17409 two_stage_opamp_dummy_magic_29_0.X.n87 two_stage_opamp_dummy_magic_29_0.X.n86 0.0217373
R17410 two_stage_opamp_dummy_magic_29_0.X.n84 two_stage_opamp_dummy_magic_29_0.X.n83 0.0217373
R17411 two_stage_opamp_dummy_magic_29_0.X.n81 two_stage_opamp_dummy_magic_29_0.X.n35 0.0217373
R17412 two_stage_opamp_dummy_magic_29_0.X.n89 two_stage_opamp_dummy_magic_29_0.X.n9 0.0217373
R17413 two_stage_opamp_dummy_magic_29_0.X.n91 two_stage_opamp_dummy_magic_29_0.X.n88 0.0217373
R17414 two_stage_opamp_dummy_magic_29_0.X.n87 two_stage_opamp_dummy_magic_29_0.X.n85 0.0217373
R17415 two_stage_opamp_dummy_magic_29_0.X.n62 two_stage_opamp_dummy_magic_29_0.X.n55 0.0217373
R17416 two_stage_opamp_dummy_magic_29_0.X.n83 two_stage_opamp_dummy_magic_29_0.X.n33 0.0217373
R17417 two_stage_opamp_dummy_magic_29_0.X.n35 two_stage_opamp_dummy_magic_29_0.X.n33 0.0217373
R17418 two_stage_opamp_dummy_magic_29_0.X.n58 two_stage_opamp_dummy_magic_29_0.X.n56 0.0217373
R17419 two_stage_opamp_dummy_magic_29_0.X.n57 two_stage_opamp_dummy_magic_29_0.X.n55 0.0217373
R17420 two_stage_opamp_dummy_magic_29_0.X.n96 two_stage_opamp_dummy_magic_29_0.X.n9 0.0217373
R17421 two_stage_opamp_dummy_magic_29_0.X.n88 two_stage_opamp_dummy_magic_29_0.X.n8 0.0217373
R17422 two_stage_opamp_dummy_magic_29_0.X.n86 two_stage_opamp_dummy_magic_29_0.X.n7 0.0217373
R17423 two_stage_opamp_dummy_magic_29_0.X.n96 two_stage_opamp_dummy_magic_29_0.X.n95 0.0217373
R17424 two_stage_opamp_dummy_magic_29_0.X.n90 two_stage_opamp_dummy_magic_29_0.X.n8 0.0217373
R17425 two_stage_opamp_dummy_magic_29_0.X.n92 two_stage_opamp_dummy_magic_29_0.X.n7 0.0217373
R17426 two_stage_opamp_dummy_magic_29_0.X.n59 two_stage_opamp_dummy_magic_29_0.X.n57 0.0217373
R17427 two_stage_opamp_dummy_magic_29_0.X.n80 two_stage_opamp_dummy_magic_29_0.X.n32 0.0217373
R17428 two_stage_opamp_dummy_magic_29_0.X.n34 two_stage_opamp_dummy_magic_29_0.X.n32 0.0217373
R17429 two_stage_opamp_dummy_magic_29_0.X.n61 two_stage_opamp_dummy_magic_29_0.X.n56 0.0217373
R17430 two_stage_opamp_dummy_magic_29_0.X.n61 two_stage_opamp_dummy_magic_29_0.X.n60 0.0217373
R17431 two_stage_opamp_dummy_magic_29_0.X two_stage_opamp_dummy_magic_29_0.X.n125 0.016125
R17432 two_stage_opamp_dummy_magic_29_0.X.n94 two_stage_opamp_dummy_magic_29_0.X.n31 0.00991089
R17433 two_stage_opamp_dummy_magic_29_0.X.n97 two_stage_opamp_dummy_magic_29_0.X.n6 0.00991089
R17434 two_stage_opamp_dummy_magic_29_0.X.n94 two_stage_opamp_dummy_magic_29_0.X.n93 0.00991089
R17435 two_stage_opamp_dummy_magic_29_0.X.n31 two_stage_opamp_dummy_magic_29_0.X.n6 0.00991089
R17436 two_stage_opamp_dummy_magic_29_0.X two_stage_opamp_dummy_magic_29_0.X.n0 0.00942857
R17437 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n8 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n7 301.983
R17438 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n10 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n9 297.151
R17439 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n6 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n5 297.151
R17440 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n27 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n26 118.861
R17441 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n29 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n28 118.861
R17442 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n33 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n32 118.861
R17443 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n36 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n35 118.861
R17444 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n39 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n38 118.861
R17445 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n41 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.t0 115.672
R17446 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n9 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.t15 39.4005
R17447 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n9 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.t12 39.4005
R17448 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n7 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.t14 39.4005
R17449 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n7 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.t13 39.4005
R17450 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n5 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.t11 39.4005
R17451 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n5 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.t16 39.4005
R17452 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n26 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.t3 19.7005
R17453 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n26 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.t8 19.7005
R17454 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n28 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.t4 19.7005
R17455 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n28 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.t9 19.7005
R17456 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n32 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.t6 19.7005
R17457 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n32 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.t10 19.7005
R17458 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n35 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.t5 19.7005
R17459 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n35 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.t2 19.7005
R17460 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n38 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.t7 19.7005
R17461 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n38 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.t1 19.7005
R17462 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n12 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n11 13.2304
R17463 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n11 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n6 12.339
R17464 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n11 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n10 11.6515
R17465 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n30 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n27 5.60467
R17466 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n39 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n37 5.54217
R17467 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n27 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n25 5.54217
R17468 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n8 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n6 5.39633
R17469 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n10 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n8 5.39633
R17470 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n30 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n29 5.04217
R17471 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n33 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n31 5.04217
R17472 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n36 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n24 5.04217
R17473 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n40 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n39 5.04217
R17474 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n29 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n25 4.97967
R17475 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n34 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n33 4.97967
R17476 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n37 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n36 4.97967
R17477 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n14 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n4 4.5005
R17478 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n16 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n15 4.5005
R17479 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n15 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n14 4.5005
R17480 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n21 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n20 4.5005
R17481 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n41 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n40 2.99085
R17482 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n18 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n0 2.26187
R17483 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n19 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n18 2.26187
R17484 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n16 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n2 2.24063
R17485 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n3 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n1 2.24063
R17486 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n22 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n17 2.24063
R17487 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n23 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n0 2.24063
R17488 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n13 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n12 2.24063
R17489 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n37 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n34 0.563
R17490 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n34 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n25 0.563
R17491 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n23 0.443208
R17492 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n40 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n24 0.34425
R17493 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n31 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n24 0.34425
R17494 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n31 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n30 0.34425
R17495 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n17 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n16 0.078625
R17496 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n16 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n1 0.0421667
R17497 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n12 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n2 0.0217373
R17498 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n15 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n3 0.0217373
R17499 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n4 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n2 0.0217373
R17500 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n4 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n3 0.0217373
R17501 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n22 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n21 0.0217373
R17502 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n20 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n0 0.0217373
R17503 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n23 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n22 0.0217373
R17504 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n14 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n13 0.0217373
R17505 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n20 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n19 0.0217373
R17506 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n13 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n1 0.0217373
R17507 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n21 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n18 0.0217373
R17508 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n19 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n17 0.0217373
R17509 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n41 0.0213333
R17510 bgr_11_0.1st_Vout_1.n12 bgr_11_0.1st_Vout_1.t29 363.909
R17511 bgr_11_0.1st_Vout_1 bgr_11_0.1st_Vout_1.t13 351.88
R17512 bgr_11_0.1st_Vout_1.n0 bgr_11_0.1st_Vout_1.n22 299.25
R17513 bgr_11_0.1st_Vout_1.n14 bgr_11_0.1st_Vout_1.n13 299.25
R17514 bgr_11_0.1st_Vout_1.n18 bgr_11_0.1st_Vout_1.n17 297.807
R17515 bgr_11_0.1st_Vout_1.n20 bgr_11_0.1st_Vout_1.t30 194.809
R17516 bgr_11_0.1st_Vout_1.n20 bgr_11_0.1st_Vout_1.t10 194.809
R17517 bgr_11_0.1st_Vout_1.n15 bgr_11_0.1st_Vout_1.t28 194.809
R17518 bgr_11_0.1st_Vout_1.n15 bgr_11_0.1st_Vout_1.t19 194.809
R17519 bgr_11_0.1st_Vout_1.n21 bgr_11_0.1st_Vout_1.n20 163.097
R17520 bgr_11_0.1st_Vout_1.n16 bgr_11_0.1st_Vout_1.n15 163.097
R17521 bgr_11_0.1st_Vout_1.n18 bgr_11_0.1st_Vout_1.t3 49.4474
R17522 bgr_11_0.1st_Vout_1.n22 bgr_11_0.1st_Vout_1.t2 39.4005
R17523 bgr_11_0.1st_Vout_1.n22 bgr_11_0.1st_Vout_1.t4 39.4005
R17524 bgr_11_0.1st_Vout_1.n13 bgr_11_0.1st_Vout_1.t6 39.4005
R17525 bgr_11_0.1st_Vout_1.n13 bgr_11_0.1st_Vout_1.t5 39.4005
R17526 bgr_11_0.1st_Vout_1.n17 bgr_11_0.1st_Vout_1.t1 39.4005
R17527 bgr_11_0.1st_Vout_1.n17 bgr_11_0.1st_Vout_1.t0 39.4005
R17528 bgr_11_0.1st_Vout_1.n2 bgr_11_0.1st_Vout_1.t27 4.8295
R17529 bgr_11_0.1st_Vout_1.n1 bgr_11_0.1st_Vout_1.t14 4.8295
R17530 bgr_11_0.1st_Vout_1.n4 bgr_11_0.1st_Vout_1.t32 4.8295
R17531 bgr_11_0.1st_Vout_1.n3 bgr_11_0.1st_Vout_1.t22 4.8295
R17532 bgr_11_0.1st_Vout_1.n6 bgr_11_0.1st_Vout_1.t25 4.8295
R17533 bgr_11_0.1st_Vout_1.n5 bgr_11_0.1st_Vout_1.t12 4.8295
R17534 bgr_11_0.1st_Vout_1.n8 bgr_11_0.1st_Vout_1.t16 4.8295
R17535 bgr_11_0.1st_Vout_1.n7 bgr_11_0.1st_Vout_1.t7 4.8295
R17536 bgr_11_0.1st_Vout_1.n9 bgr_11_0.1st_Vout_1.t24 4.8295
R17537 bgr_11_0.1st_Vout_1.n2 bgr_11_0.1st_Vout_1.t18 4.5005
R17538 bgr_11_0.1st_Vout_1.n1 bgr_11_0.1st_Vout_1.t23 4.5005
R17539 bgr_11_0.1st_Vout_1.n4 bgr_11_0.1st_Vout_1.t26 4.5005
R17540 bgr_11_0.1st_Vout_1.n3 bgr_11_0.1st_Vout_1.t31 4.5005
R17541 bgr_11_0.1st_Vout_1.n6 bgr_11_0.1st_Vout_1.t17 4.5005
R17542 bgr_11_0.1st_Vout_1.n5 bgr_11_0.1st_Vout_1.t21 4.5005
R17543 bgr_11_0.1st_Vout_1.n8 bgr_11_0.1st_Vout_1.t8 4.5005
R17544 bgr_11_0.1st_Vout_1.n7 bgr_11_0.1st_Vout_1.t11 4.5005
R17545 bgr_11_0.1st_Vout_1.n9 bgr_11_0.1st_Vout_1.t15 4.5005
R17546 bgr_11_0.1st_Vout_1.n10 bgr_11_0.1st_Vout_1.t20 4.5005
R17547 bgr_11_0.1st_Vout_1.n11 bgr_11_0.1st_Vout_1.t9 4.5005
R17548 bgr_11_0.1st_Vout_1.n19 bgr_11_0.1st_Vout_1.n18 1.44719
R17549 bgr_11_0.1st_Vout_1.n2 bgr_11_0.1st_Vout_1.n1 0.3295
R17550 bgr_11_0.1st_Vout_1.n4 bgr_11_0.1st_Vout_1.n3 0.3295
R17551 bgr_11_0.1st_Vout_1.n6 bgr_11_0.1st_Vout_1.n5 0.3295
R17552 bgr_11_0.1st_Vout_1.n8 bgr_11_0.1st_Vout_1.n7 0.3295
R17553 bgr_11_0.1st_Vout_1.n10 bgr_11_0.1st_Vout_1.n9 0.3295
R17554 bgr_11_0.1st_Vout_1.n11 bgr_11_0.1st_Vout_1.n10 0.3295
R17555 bgr_11_0.1st_Vout_1.n4 bgr_11_0.1st_Vout_1.n2 0.2825
R17556 bgr_11_0.1st_Vout_1.n6 bgr_11_0.1st_Vout_1.n4 0.2825
R17557 bgr_11_0.1st_Vout_1.n8 bgr_11_0.1st_Vout_1.n6 0.2825
R17558 bgr_11_0.1st_Vout_1.n9 bgr_11_0.1st_Vout_1.n8 0.2825
R17559 bgr_11_0.1st_Vout_1.n19 bgr_11_0.1st_Vout_1.n16 0.2505
R17560 bgr_11_0.1st_Vout_1.n0 bgr_11_0.1st_Vout_1.n21 0.2505
R17561 bgr_11_0.1st_Vout_1.n14 bgr_11_0.1st_Vout_1.n12 0.21925
R17562 bgr_11_0.1st_Vout_1.n16 bgr_11_0.1st_Vout_1.n14 0.1255
R17563 bgr_11_0.1st_Vout_1.n21 bgr_11_0.1st_Vout_1.n19 0.1255
R17564 bgr_11_0.1st_Vout_1 bgr_11_0.1st_Vout_1.n0 0.09425
R17565 bgr_11_0.1st_Vout_1.n12 bgr_11_0.1st_Vout_1.n11 10.102
R17566 bgr_11_0.cap_res1.t20 bgr_11_0.cap_res1.t13 121.983
R17567 bgr_11_0.cap_res1.t9 bgr_11_0.cap_res1.t17 0.1603
R17568 bgr_11_0.cap_res1.t16 bgr_11_0.cap_res1.t19 0.1603
R17569 bgr_11_0.cap_res1.t8 bgr_11_0.cap_res1.t15 0.1603
R17570 bgr_11_0.cap_res1.t1 bgr_11_0.cap_res1.t7 0.1603
R17571 bgr_11_0.cap_res1.t6 bgr_11_0.cap_res1.t14 0.1603
R17572 bgr_11_0.cap_res1.n1 bgr_11_0.cap_res1.t10 0.159278
R17573 bgr_11_0.cap_res1.n2 bgr_11_0.cap_res1.t3 0.159278
R17574 bgr_11_0.cap_res1.n3 bgr_11_0.cap_res1.t11 0.159278
R17575 bgr_11_0.cap_res1.n4 bgr_11_0.cap_res1.t18 0.159278
R17576 bgr_11_0.cap_res1.n4 bgr_11_0.cap_res1.t9 0.1368
R17577 bgr_11_0.cap_res1.n4 bgr_11_0.cap_res1.t5 0.1368
R17578 bgr_11_0.cap_res1.n3 bgr_11_0.cap_res1.t16 0.1368
R17579 bgr_11_0.cap_res1.n3 bgr_11_0.cap_res1.t12 0.1368
R17580 bgr_11_0.cap_res1.n2 bgr_11_0.cap_res1.t8 0.1368
R17581 bgr_11_0.cap_res1.n2 bgr_11_0.cap_res1.t4 0.1368
R17582 bgr_11_0.cap_res1.n1 bgr_11_0.cap_res1.t1 0.1368
R17583 bgr_11_0.cap_res1.n1 bgr_11_0.cap_res1.t0 0.1368
R17584 bgr_11_0.cap_res1.n0 bgr_11_0.cap_res1.t6 0.1368
R17585 bgr_11_0.cap_res1.n0 bgr_11_0.cap_res1.t2 0.1368
R17586 bgr_11_0.cap_res1.t10 bgr_11_0.cap_res1.n0 0.00152174
R17587 bgr_11_0.cap_res1.t3 bgr_11_0.cap_res1.n1 0.00152174
R17588 bgr_11_0.cap_res1.t11 bgr_11_0.cap_res1.n2 0.00152174
R17589 bgr_11_0.cap_res1.t18 bgr_11_0.cap_res1.n3 0.00152174
R17590 bgr_11_0.cap_res1.t13 bgr_11_0.cap_res1.n4 0.00152174
R17591 bgr_11_0.NFET_GATE_10uA.n3 bgr_11_0.NFET_GATE_10uA.t6 369.534
R17592 bgr_11_0.NFET_GATE_10uA.n2 bgr_11_0.NFET_GATE_10uA.t9 369.534
R17593 bgr_11_0.NFET_GATE_10uA.n8 bgr_11_0.NFET_GATE_10uA.t22 369.534
R17594 bgr_11_0.NFET_GATE_10uA.n7 bgr_11_0.NFET_GATE_10uA.t20 369.534
R17595 bgr_11_0.NFET_GATE_10uA.n15 bgr_11_0.NFET_GATE_10uA.t13 369.534
R17596 bgr_11_0.NFET_GATE_10uA.n12 bgr_11_0.NFET_GATE_10uA.t11 369.534
R17597 bgr_11_0.NFET_GATE_10uA.n18 bgr_11_0.NFET_GATE_10uA.t1 369.534
R17598 bgr_11_0.NFET_GATE_10uA.n0 bgr_11_0.NFET_GATE_10uA.n1 360.288
R17599 bgr_11_0.NFET_GATE_10uA.n19 bgr_11_0.NFET_GATE_10uA.t7 249.034
R17600 bgr_11_0.NFET_GATE_10uA.n5 bgr_11_0.NFET_GATE_10uA.t5 192.8
R17601 bgr_11_0.NFET_GATE_10uA.n4 bgr_11_0.NFET_GATE_10uA.t12 192.8
R17602 bgr_11_0.NFET_GATE_10uA.n3 bgr_11_0.NFET_GATE_10uA.t19 192.8
R17603 bgr_11_0.NFET_GATE_10uA.n2 bgr_11_0.NFET_GATE_10uA.t18 192.8
R17604 bgr_11_0.NFET_GATE_10uA.n9 bgr_11_0.NFET_GATE_10uA.t15 192.8
R17605 bgr_11_0.NFET_GATE_10uA.n8 bgr_11_0.NFET_GATE_10uA.t23 192.8
R17606 bgr_11_0.NFET_GATE_10uA.n7 bgr_11_0.NFET_GATE_10uA.t8 192.8
R17607 bgr_11_0.NFET_GATE_10uA.n15 bgr_11_0.NFET_GATE_10uA.t10 192.8
R17608 bgr_11_0.NFET_GATE_10uA.n12 bgr_11_0.NFET_GATE_10uA.t17 192.8
R17609 bgr_11_0.NFET_GATE_10uA.n13 bgr_11_0.NFET_GATE_10uA.t16 192.8
R17610 bgr_11_0.NFET_GATE_10uA.n14 bgr_11_0.NFET_GATE_10uA.t21 192.8
R17611 bgr_11_0.NFET_GATE_10uA.n18 bgr_11_0.NFET_GATE_10uA.t14 192.8
R17612 bgr_11_0.NFET_GATE_10uA.n5 bgr_11_0.NFET_GATE_10uA.n4 176.733
R17613 bgr_11_0.NFET_GATE_10uA.n4 bgr_11_0.NFET_GATE_10uA.n3 176.733
R17614 bgr_11_0.NFET_GATE_10uA.n9 bgr_11_0.NFET_GATE_10uA.n8 176.733
R17615 bgr_11_0.NFET_GATE_10uA.n13 bgr_11_0.NFET_GATE_10uA.n12 176.733
R17616 bgr_11_0.NFET_GATE_10uA.n14 bgr_11_0.NFET_GATE_10uA.n13 176.733
R17617 bgr_11_0.NFET_GATE_10uA.n11 bgr_11_0.NFET_GATE_10uA.n6 168.014
R17618 bgr_11_0.NFET_GATE_10uA.n11 bgr_11_0.NFET_GATE_10uA.n10 166.343
R17619 bgr_11_0.NFET_GATE_10uA.n17 bgr_11_0.NFET_GATE_10uA.n16 166.343
R17620 bgr_11_0.NFET_GATE_10uA.n0 bgr_11_0.NFET_GATE_10uA.n19 166.343
R17621 bgr_11_0.NFET_GATE_10uA.n20 bgr_11_0.NFET_GATE_10uA.n0 141.752
R17622 bgr_11_0.NFET_GATE_10uA.n6 bgr_11_0.NFET_GATE_10uA.n5 56.2338
R17623 bgr_11_0.NFET_GATE_10uA.n6 bgr_11_0.NFET_GATE_10uA.n2 56.2338
R17624 bgr_11_0.NFET_GATE_10uA.n10 bgr_11_0.NFET_GATE_10uA.n9 56.2338
R17625 bgr_11_0.NFET_GATE_10uA.n10 bgr_11_0.NFET_GATE_10uA.n7 56.2338
R17626 bgr_11_0.NFET_GATE_10uA.n16 bgr_11_0.NFET_GATE_10uA.n15 56.2338
R17627 bgr_11_0.NFET_GATE_10uA.n16 bgr_11_0.NFET_GATE_10uA.n14 56.2338
R17628 bgr_11_0.NFET_GATE_10uA.n19 bgr_11_0.NFET_GATE_10uA.n18 56.2338
R17629 bgr_11_0.NFET_GATE_10uA.n1 bgr_11_0.NFET_GATE_10uA.t4 39.4005
R17630 bgr_11_0.NFET_GATE_10uA.n1 bgr_11_0.NFET_GATE_10uA.t3 39.4005
R17631 bgr_11_0.NFET_GATE_10uA.t0 bgr_11_0.NFET_GATE_10uA.n20 24.0005
R17632 bgr_11_0.NFET_GATE_10uA.n20 bgr_11_0.NFET_GATE_10uA.t2 24.0005
R17633 bgr_11_0.NFET_GATE_10uA.n0 bgr_11_0.NFET_GATE_10uA.n17 2.01612
R17634 bgr_11_0.NFET_GATE_10uA.n17 bgr_11_0.NFET_GATE_10uA.n11 1.5005
R17635 two_stage_opamp_dummy_magic_29_0.VD4.n17 two_stage_opamp_dummy_magic_29_0.VD4.t32 671.418
R17636 two_stage_opamp_dummy_magic_29_0.VD4.n14 two_stage_opamp_dummy_magic_29_0.VD4.t35 671.418
R17637 two_stage_opamp_dummy_magic_29_0.VD4.t36 two_stage_opamp_dummy_magic_29_0.VD4.n15 213.131
R17638 two_stage_opamp_dummy_magic_29_0.VD4.n16 two_stage_opamp_dummy_magic_29_0.VD4.t33 213.131
R17639 two_stage_opamp_dummy_magic_29_0.VD4.t30 two_stage_opamp_dummy_magic_29_0.VD4.t36 146.155
R17640 two_stage_opamp_dummy_magic_29_0.VD4.t16 two_stage_opamp_dummy_magic_29_0.VD4.t30 146.155
R17641 two_stage_opamp_dummy_magic_29_0.VD4.t24 two_stage_opamp_dummy_magic_29_0.VD4.t16 146.155
R17642 two_stage_opamp_dummy_magic_29_0.VD4.t20 two_stage_opamp_dummy_magic_29_0.VD4.t24 146.155
R17643 two_stage_opamp_dummy_magic_29_0.VD4.t26 two_stage_opamp_dummy_magic_29_0.VD4.t20 146.155
R17644 two_stage_opamp_dummy_magic_29_0.VD4.t28 two_stage_opamp_dummy_magic_29_0.VD4.t26 146.155
R17645 two_stage_opamp_dummy_magic_29_0.VD4.t12 two_stage_opamp_dummy_magic_29_0.VD4.t28 146.155
R17646 two_stage_opamp_dummy_magic_29_0.VD4.t18 two_stage_opamp_dummy_magic_29_0.VD4.t12 146.155
R17647 two_stage_opamp_dummy_magic_29_0.VD4.t14 two_stage_opamp_dummy_magic_29_0.VD4.t18 146.155
R17648 two_stage_opamp_dummy_magic_29_0.VD4.t22 two_stage_opamp_dummy_magic_29_0.VD4.t14 146.155
R17649 two_stage_opamp_dummy_magic_29_0.VD4.t33 two_stage_opamp_dummy_magic_29_0.VD4.t22 146.155
R17650 two_stage_opamp_dummy_magic_29_0.VD4.n15 two_stage_opamp_dummy_magic_29_0.VD4.t37 76.2576
R17651 two_stage_opamp_dummy_magic_29_0.VD4.n16 two_stage_opamp_dummy_magic_29_0.VD4.t34 76.2576
R17652 two_stage_opamp_dummy_magic_29_0.VD4.n31 two_stage_opamp_dummy_magic_29_0.VD4.n6 67.013
R17653 two_stage_opamp_dummy_magic_29_0.VD4.n30 two_stage_opamp_dummy_magic_29_0.VD4.n9 67.013
R17654 two_stage_opamp_dummy_magic_29_0.VD4.n13 two_stage_opamp_dummy_magic_29_0.VD4.n12 67.013
R17655 two_stage_opamp_dummy_magic_29_0.VD4.n0 two_stage_opamp_dummy_magic_29_0.VD4.n18 67.013
R17656 two_stage_opamp_dummy_magic_29_0.VD4.n33 two_stage_opamp_dummy_magic_29_0.VD4.n32 67.013
R17657 two_stage_opamp_dummy_magic_29_0.VD4.n28 two_stage_opamp_dummy_magic_29_0.VD4.n27 66.0338
R17658 two_stage_opamp_dummy_magic_29_0.VD4.n25 two_stage_opamp_dummy_magic_29_0.VD4.n24 66.0338
R17659 two_stage_opamp_dummy_magic_29_0.VD4.n11 two_stage_opamp_dummy_magic_29_0.VD4.n10 66.0338
R17660 two_stage_opamp_dummy_magic_29_0.VD4.n8 two_stage_opamp_dummy_magic_29_0.VD4.n7 66.0338
R17661 two_stage_opamp_dummy_magic_29_0.VD4.n5 two_stage_opamp_dummy_magic_29_0.VD4.n4 66.0338
R17662 two_stage_opamp_dummy_magic_29_0.VD4.n20 two_stage_opamp_dummy_magic_29_0.VD4.n19 66.0338
R17663 two_stage_opamp_dummy_magic_29_0.VD4.n6 two_stage_opamp_dummy_magic_29_0.VD4.t25 11.2576
R17664 two_stage_opamp_dummy_magic_29_0.VD4.n6 two_stage_opamp_dummy_magic_29_0.VD4.t21 11.2576
R17665 two_stage_opamp_dummy_magic_29_0.VD4.n9 two_stage_opamp_dummy_magic_29_0.VD4.t27 11.2576
R17666 two_stage_opamp_dummy_magic_29_0.VD4.n9 two_stage_opamp_dummy_magic_29_0.VD4.t29 11.2576
R17667 two_stage_opamp_dummy_magic_29_0.VD4.n12 two_stage_opamp_dummy_magic_29_0.VD4.t13 11.2576
R17668 two_stage_opamp_dummy_magic_29_0.VD4.n12 two_stage_opamp_dummy_magic_29_0.VD4.t19 11.2576
R17669 two_stage_opamp_dummy_magic_29_0.VD4.n27 two_stage_opamp_dummy_magic_29_0.VD4.t4 11.2576
R17670 two_stage_opamp_dummy_magic_29_0.VD4.n27 two_stage_opamp_dummy_magic_29_0.VD4.t10 11.2576
R17671 two_stage_opamp_dummy_magic_29_0.VD4.n24 two_stage_opamp_dummy_magic_29_0.VD4.t8 11.2576
R17672 two_stage_opamp_dummy_magic_29_0.VD4.n24 two_stage_opamp_dummy_magic_29_0.VD4.t3 11.2576
R17673 two_stage_opamp_dummy_magic_29_0.VD4.n10 two_stage_opamp_dummy_magic_29_0.VD4.t7 11.2576
R17674 two_stage_opamp_dummy_magic_29_0.VD4.n10 two_stage_opamp_dummy_magic_29_0.VD4.t1 11.2576
R17675 two_stage_opamp_dummy_magic_29_0.VD4.n7 two_stage_opamp_dummy_magic_29_0.VD4.t2 11.2576
R17676 two_stage_opamp_dummy_magic_29_0.VD4.n7 two_stage_opamp_dummy_magic_29_0.VD4.t0 11.2576
R17677 two_stage_opamp_dummy_magic_29_0.VD4.n4 two_stage_opamp_dummy_magic_29_0.VD4.t6 11.2576
R17678 two_stage_opamp_dummy_magic_29_0.VD4.n4 two_stage_opamp_dummy_magic_29_0.VD4.t9 11.2576
R17679 two_stage_opamp_dummy_magic_29_0.VD4.n19 two_stage_opamp_dummy_magic_29_0.VD4.t11 11.2576
R17680 two_stage_opamp_dummy_magic_29_0.VD4.n19 two_stage_opamp_dummy_magic_29_0.VD4.t5 11.2576
R17681 two_stage_opamp_dummy_magic_29_0.VD4.n18 two_stage_opamp_dummy_magic_29_0.VD4.t15 11.2576
R17682 two_stage_opamp_dummy_magic_29_0.VD4.n18 two_stage_opamp_dummy_magic_29_0.VD4.t23 11.2576
R17683 two_stage_opamp_dummy_magic_29_0.VD4.n32 two_stage_opamp_dummy_magic_29_0.VD4.t31 11.2576
R17684 two_stage_opamp_dummy_magic_29_0.VD4.n32 two_stage_opamp_dummy_magic_29_0.VD4.t17 11.2576
R17685 two_stage_opamp_dummy_magic_29_0.VD4.n21 two_stage_opamp_dummy_magic_29_0.VD4.n20 5.66717
R17686 two_stage_opamp_dummy_magic_29_0.VD4.n28 two_stage_opamp_dummy_magic_29_0.VD4.n26 5.66717
R17687 two_stage_opamp_dummy_magic_29_0.VD4.n26 two_stage_opamp_dummy_magic_29_0.VD4.n25 5.29217
R17688 two_stage_opamp_dummy_magic_29_0.VD4.n23 two_stage_opamp_dummy_magic_29_0.VD4.n11 5.29217
R17689 two_stage_opamp_dummy_magic_29_0.VD4.n22 two_stage_opamp_dummy_magic_29_0.VD4.n8 5.29217
R17690 two_stage_opamp_dummy_magic_29_0.VD4.n21 two_stage_opamp_dummy_magic_29_0.VD4.n5 5.29217
R17691 two_stage_opamp_dummy_magic_29_0.VD4.n15 two_stage_opamp_dummy_magic_29_0.VD4.n14 1.90883
R17692 two_stage_opamp_dummy_magic_29_0.VD4.n17 two_stage_opamp_dummy_magic_29_0.VD4.n16 1.90883
R17693 two_stage_opamp_dummy_magic_29_0.VD4.n25 two_stage_opamp_dummy_magic_29_0.VD4.n13 1.02133
R17694 two_stage_opamp_dummy_magic_29_0.VD4.n30 two_stage_opamp_dummy_magic_29_0.VD4.n11 1.02133
R17695 two_stage_opamp_dummy_magic_29_0.VD4.n31 two_stage_opamp_dummy_magic_29_0.VD4.n8 1.02133
R17696 two_stage_opamp_dummy_magic_29_0.VD4.n33 two_stage_opamp_dummy_magic_29_0.VD4.n5 1.02133
R17697 two_stage_opamp_dummy_magic_29_0.VD4.n20 two_stage_opamp_dummy_magic_29_0.VD4.n2 1.02133
R17698 two_stage_opamp_dummy_magic_29_0.VD4.n0 two_stage_opamp_dummy_magic_29_0.VD4.n28 1.02133
R17699 two_stage_opamp_dummy_magic_29_0.VD4 two_stage_opamp_dummy_magic_29_0.VD4.n2 0.65675
R17700 two_stage_opamp_dummy_magic_29_0.VD4.n30 two_stage_opamp_dummy_magic_29_0.VD4.n29 0.643357
R17701 two_stage_opamp_dummy_magic_29_0.VD4.n31 two_stage_opamp_dummy_magic_29_0.VD4.n3 0.643357
R17702 two_stage_opamp_dummy_magic_29_0.VD4.n34 two_stage_opamp_dummy_magic_29_0.VD4.n33 0.643357
R17703 two_stage_opamp_dummy_magic_29_0.VD4.n1 two_stage_opamp_dummy_magic_29_0.VD4.n0 0.0280497
R17704 two_stage_opamp_dummy_magic_29_0.VD4.n22 two_stage_opamp_dummy_magic_29_0.VD4.n21 0.3755
R17705 two_stage_opamp_dummy_magic_29_0.VD4.n23 two_stage_opamp_dummy_magic_29_0.VD4.n22 0.3755
R17706 two_stage_opamp_dummy_magic_29_0.VD4.n26 two_stage_opamp_dummy_magic_29_0.VD4.n23 0.3755
R17707 two_stage_opamp_dummy_magic_29_0.VD4.n0 two_stage_opamp_dummy_magic_29_0.VD4.n17 0.132669
R17708 two_stage_opamp_dummy_magic_29_0.VD4.n14 two_stage_opamp_dummy_magic_29_0.VD4.n2 0.104667
R17709 two_stage_opamp_dummy_magic_29_0.VD4.n1 two_stage_opamp_dummy_magic_29_0.VD4.n13 0.0473045
R17710 two_stage_opamp_dummy_magic_29_0.VD4.n34 two_stage_opamp_dummy_magic_29_0.VD4.n3 0.0540714
R17711 two_stage_opamp_dummy_magic_29_0.VD4.n29 two_stage_opamp_dummy_magic_29_0.VD4.n3 0.0540714
R17712 two_stage_opamp_dummy_magic_29_0.VD4.n29 two_stage_opamp_dummy_magic_29_0.VD4.n1 0.274553
R17713 two_stage_opamp_dummy_magic_29_0.VD4.n33 two_stage_opamp_dummy_magic_29_0.VD4.n2 0.0540714
R17714 two_stage_opamp_dummy_magic_29_0.VD4.n33 two_stage_opamp_dummy_magic_29_0.VD4.n31 0.0540714
R17715 two_stage_opamp_dummy_magic_29_0.VD4.n31 two_stage_opamp_dummy_magic_29_0.VD4.n30 0.0540714
R17716 two_stage_opamp_dummy_magic_29_0.VD4.n30 two_stage_opamp_dummy_magic_29_0.VD4.n13 0.0540714
R17717 two_stage_opamp_dummy_magic_29_0.VD4 two_stage_opamp_dummy_magic_29_0.VD4.n34 0.0406786
R17718 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n20 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.t14 115.6
R17719 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n2 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n0 107.121
R17720 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n2 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n1 97.4332
R17721 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n2 24.5317
R17722 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n18 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n17 24.288
R17723 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n15 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n14 24.288
R17724 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n12 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n11 24.288
R17725 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n8 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n7 24.288
R17726 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n6 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n5 24.288
R17727 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n0 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.t3 24.0005
R17728 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n0 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.t0 24.0005
R17729 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n1 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.t1 24.0005
R17730 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n1 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.t2 24.0005
R17731 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n17 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.t11 8.0005
R17732 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n17 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.t5 8.0005
R17733 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n14 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.t9 8.0005
R17734 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n14 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.t6 8.0005
R17735 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n11 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.t10 8.0005
R17736 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n11 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.t4 8.0005
R17737 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n7 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.t8 8.0005
R17738 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n7 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.t13 8.0005
R17739 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n5 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.t7 8.0005
R17740 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n5 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.t12 8.0005
R17741 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n6 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n4 5.7505
R17742 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n18 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n16 5.7505
R17743 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n9 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n6 5.53175
R17744 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n15 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n3 5.188
R17745 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n16 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n15 5.188
R17746 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n12 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n10 5.188
R17747 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n13 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n12 5.188
R17748 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n9 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n8 5.188
R17749 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n8 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n4 5.188
R17750 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n19 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n18 5.188
R17751 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n20 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n19 2.38147
R17752 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n13 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n4 0.563
R17753 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n16 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n13 0.563
R17754 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n19 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n3 0.34425
R17755 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n10 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n3 0.34425
R17756 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n10 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n9 0.34425
R17757 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n20 0.0213333
R17758 bgr_11_0.START_UP_NFET1 bgr_11_0.START_UP_NFET1.t0 141.653
R17759 bgr_11_0.V_mir1.n11 bgr_11_0.V_mir1.t18 310.488
R17760 bgr_11_0.V_mir1.n5 bgr_11_0.V_mir1.t13 310.488
R17761 bgr_11_0.V_mir1.n0 bgr_11_0.V_mir1.t17 310.488
R17762 bgr_11_0.V_mir1.n9 bgr_11_0.V_mir1.n8 297.433
R17763 bgr_11_0.V_mir1.n4 bgr_11_0.V_mir1.n3 297.433
R17764 bgr_11_0.V_mir1.n15 bgr_11_0.V_mir1.n14 297.433
R17765 bgr_11_0.V_mir1.n13 bgr_11_0.V_mir1.t11 184.097
R17766 bgr_11_0.V_mir1.n7 bgr_11_0.V_mir1.t9 184.097
R17767 bgr_11_0.V_mir1.n2 bgr_11_0.V_mir1.t7 184.097
R17768 bgr_11_0.V_mir1.n12 bgr_11_0.V_mir1.n11 167.094
R17769 bgr_11_0.V_mir1.n6 bgr_11_0.V_mir1.n5 167.094
R17770 bgr_11_0.V_mir1.n1 bgr_11_0.V_mir1.n0 167.094
R17771 bgr_11_0.V_mir1.n14 bgr_11_0.V_mir1.n13 161.3
R17772 bgr_11_0.V_mir1.n9 bgr_11_0.V_mir1.n7 161.3
R17773 bgr_11_0.V_mir1.n4 bgr_11_0.V_mir1.n2 161.3
R17774 bgr_11_0.V_mir1.n11 bgr_11_0.V_mir1.t14 120.501
R17775 bgr_11_0.V_mir1.n12 bgr_11_0.V_mir1.t5 120.501
R17776 bgr_11_0.V_mir1.n5 bgr_11_0.V_mir1.t15 120.501
R17777 bgr_11_0.V_mir1.n6 bgr_11_0.V_mir1.t3 120.501
R17778 bgr_11_0.V_mir1.n0 bgr_11_0.V_mir1.t16 120.501
R17779 bgr_11_0.V_mir1.n1 bgr_11_0.V_mir1.t1 120.501
R17780 bgr_11_0.V_mir1.n9 bgr_11_0.V_mir1.t0 50.2004
R17781 bgr_11_0.V_mir1.n13 bgr_11_0.V_mir1.n12 40.7027
R17782 bgr_11_0.V_mir1.n7 bgr_11_0.V_mir1.n6 40.7027
R17783 bgr_11_0.V_mir1.n2 bgr_11_0.V_mir1.n1 40.7027
R17784 bgr_11_0.V_mir1.n8 bgr_11_0.V_mir1.t10 39.4005
R17785 bgr_11_0.V_mir1.n8 bgr_11_0.V_mir1.t4 39.4005
R17786 bgr_11_0.V_mir1.n3 bgr_11_0.V_mir1.t8 39.4005
R17787 bgr_11_0.V_mir1.n3 bgr_11_0.V_mir1.t2 39.4005
R17788 bgr_11_0.V_mir1.t12 bgr_11_0.V_mir1.n15 39.4005
R17789 bgr_11_0.V_mir1.n15 bgr_11_0.V_mir1.t6 39.4005
R17790 bgr_11_0.V_mir1.n10 bgr_11_0.V_mir1.n4 6.6255
R17791 bgr_11_0.V_mir1.n14 bgr_11_0.V_mir1.n10 6.6255
R17792 bgr_11_0.V_mir1.n10 bgr_11_0.V_mir1.n9 4.5005
R17793 two_stage_opamp_dummy_magic_29_0.Vb1.n2 two_stage_opamp_dummy_magic_29_0.Vb1.t15 484.212
R17794 two_stage_opamp_dummy_magic_29_0.Vb1.n2 two_stage_opamp_dummy_magic_29_0.Vb1.t26 484.212
R17795 two_stage_opamp_dummy_magic_29_0.Vb1.n2 two_stage_opamp_dummy_magic_29_0.Vb1.t13 484.212
R17796 two_stage_opamp_dummy_magic_29_0.Vb1.n2 two_stage_opamp_dummy_magic_29_0.Vb1.t25 484.212
R17797 two_stage_opamp_dummy_magic_29_0.Vb1.n3 two_stage_opamp_dummy_magic_29_0.Vb1.t12 484.212
R17798 two_stage_opamp_dummy_magic_29_0.Vb1.n3 two_stage_opamp_dummy_magic_29_0.Vb1.t23 484.212
R17799 two_stage_opamp_dummy_magic_29_0.Vb1.n3 two_stage_opamp_dummy_magic_29_0.Vb1.t18 484.212
R17800 two_stage_opamp_dummy_magic_29_0.Vb1.n3 two_stage_opamp_dummy_magic_29_0.Vb1.t24 484.212
R17801 two_stage_opamp_dummy_magic_29_0.Vb1.n7 two_stage_opamp_dummy_magic_29_0.Vb1.t32 484.212
R17802 two_stage_opamp_dummy_magic_29_0.Vb1.n7 two_stage_opamp_dummy_magic_29_0.Vb1.t22 484.212
R17803 two_stage_opamp_dummy_magic_29_0.Vb1.n4 two_stage_opamp_dummy_magic_29_0.Vb1.t20 484.212
R17804 two_stage_opamp_dummy_magic_29_0.Vb1.n4 two_stage_opamp_dummy_magic_29_0.Vb1.t30 484.212
R17805 two_stage_opamp_dummy_magic_29_0.Vb1.n4 two_stage_opamp_dummy_magic_29_0.Vb1.t19 484.212
R17806 two_stage_opamp_dummy_magic_29_0.Vb1.n4 two_stage_opamp_dummy_magic_29_0.Vb1.t28 484.212
R17807 two_stage_opamp_dummy_magic_29_0.Vb1.n5 two_stage_opamp_dummy_magic_29_0.Vb1.t16 484.212
R17808 two_stage_opamp_dummy_magic_29_0.Vb1.n5 two_stage_opamp_dummy_magic_29_0.Vb1.t29 484.212
R17809 two_stage_opamp_dummy_magic_29_0.Vb1.n5 two_stage_opamp_dummy_magic_29_0.Vb1.t17 484.212
R17810 two_stage_opamp_dummy_magic_29_0.Vb1.n5 two_stage_opamp_dummy_magic_29_0.Vb1.t27 484.212
R17811 two_stage_opamp_dummy_magic_29_0.Vb1.n6 two_stage_opamp_dummy_magic_29_0.Vb1.t14 484.212
R17812 two_stage_opamp_dummy_magic_29_0.Vb1.n6 two_stage_opamp_dummy_magic_29_0.Vb1.t21 484.212
R17813 two_stage_opamp_dummy_magic_29_0.Vb1.n9 two_stage_opamp_dummy_magic_29_0.Vb1.t9 449.868
R17814 two_stage_opamp_dummy_magic_29_0.Vb1.n8 two_stage_opamp_dummy_magic_29_0.Vb1.t3 449.868
R17815 two_stage_opamp_dummy_magic_29_0.Vb1.n9 two_stage_opamp_dummy_magic_29_0.Vb1.t7 273.134
R17816 two_stage_opamp_dummy_magic_29_0.Vb1.n8 two_stage_opamp_dummy_magic_29_0.Vb1.t5 273.134
R17817 two_stage_opamp_dummy_magic_29_0.Vb1.n12 two_stage_opamp_dummy_magic_29_0.Vb1.t31 161.363
R17818 two_stage_opamp_dummy_magic_29_0.Vb1.n1 two_stage_opamp_dummy_magic_29_0.Vb1.n10 161.3
R17819 two_stage_opamp_dummy_magic_29_0.Vb1 two_stage_opamp_dummy_magic_29_0.Vb1.n19 151.863
R17820 two_stage_opamp_dummy_magic_29_0.Vb1.n15 two_stage_opamp_dummy_magic_29_0.Vb1.n14 49.3505
R17821 two_stage_opamp_dummy_magic_29_0.Vb1.n1 two_stage_opamp_dummy_magic_29_0.Vb1.n11 49.3505
R17822 two_stage_opamp_dummy_magic_29_0.Vb1.n18 two_stage_opamp_dummy_magic_29_0.Vb1.n17 49.3505
R17823 two_stage_opamp_dummy_magic_29_0.Vb1.n10 two_stage_opamp_dummy_magic_29_0.Vb1.n9 45.5227
R17824 two_stage_opamp_dummy_magic_29_0.Vb1.n10 two_stage_opamp_dummy_magic_29_0.Vb1.n8 45.5227
R17825 two_stage_opamp_dummy_magic_29_0.Vb1.n2 two_stage_opamp_dummy_magic_29_0.Vb1.n0 21.4927
R17826 two_stage_opamp_dummy_magic_29_0.Vb1.n13 two_stage_opamp_dummy_magic_29_0.Vb1.n6 21.4927
R17827 two_stage_opamp_dummy_magic_29_0.Vb1.n19 two_stage_opamp_dummy_magic_29_0.Vb1.t2 19.7005
R17828 two_stage_opamp_dummy_magic_29_0.Vb1.n19 two_stage_opamp_dummy_magic_29_0.Vb1.t11 19.7005
R17829 two_stage_opamp_dummy_magic_29_0.Vb1.n14 two_stage_opamp_dummy_magic_29_0.Vb1.t0 16.0005
R17830 two_stage_opamp_dummy_magic_29_0.Vb1.n14 two_stage_opamp_dummy_magic_29_0.Vb1.t4 16.0005
R17831 two_stage_opamp_dummy_magic_29_0.Vb1.n11 two_stage_opamp_dummy_magic_29_0.Vb1.t6 16.0005
R17832 two_stage_opamp_dummy_magic_29_0.Vb1.n11 two_stage_opamp_dummy_magic_29_0.Vb1.t8 16.0005
R17833 two_stage_opamp_dummy_magic_29_0.Vb1.n17 two_stage_opamp_dummy_magic_29_0.Vb1.t10 16.0005
R17834 two_stage_opamp_dummy_magic_29_0.Vb1.n17 two_stage_opamp_dummy_magic_29_0.Vb1.t1 16.0005
R17835 two_stage_opamp_dummy_magic_29_0.Vb1.n16 two_stage_opamp_dummy_magic_29_0.Vb1.n15 5.28175
R17836 two_stage_opamp_dummy_magic_29_0.Vb1.n18 two_stage_opamp_dummy_magic_29_0.Vb1.n16 5.28175
R17837 two_stage_opamp_dummy_magic_29_0.Vb1.n0 two_stage_opamp_dummy_magic_29_0.Vb1.n18 4.938
R17838 two_stage_opamp_dummy_magic_29_0.Vb1.n15 two_stage_opamp_dummy_magic_29_0.Vb1.n13 4.938
R17839 two_stage_opamp_dummy_magic_29_0.Vb1.n1 two_stage_opamp_dummy_magic_29_0.Vb1.n0 4.5005
R17840 two_stage_opamp_dummy_magic_29_0.Vb1.n16 two_stage_opamp_dummy_magic_29_0.Vb1.n12 2.23569
R17841 two_stage_opamp_dummy_magic_29_0.Vb1.n5 two_stage_opamp_dummy_magic_29_0.Vb1.n4 1.03175
R17842 two_stage_opamp_dummy_magic_29_0.Vb1.n3 two_stage_opamp_dummy_magic_29_0.Vb1.n2 1.03175
R17843 two_stage_opamp_dummy_magic_29_0.Vb1.n12 two_stage_opamp_dummy_magic_29_0.Vb1.n1 0.937224
R17844 two_stage_opamp_dummy_magic_29_0.Vb1 two_stage_opamp_dummy_magic_29_0.Vb1.n4 0.852062
R17845 two_stage_opamp_dummy_magic_29_0.Vb1 two_stage_opamp_dummy_magic_29_0.Vb1.n7 0.852062
R17846 two_stage_opamp_dummy_magic_29_0.Vb1.n13 two_stage_opamp_dummy_magic_29_0.Vb1.n0 0.688
R17847 two_stage_opamp_dummy_magic_29_0.Vb1.n7 two_stage_opamp_dummy_magic_29_0.Vb1.n3 0.516125
R17848 two_stage_opamp_dummy_magic_29_0.Vb1.n6 two_stage_opamp_dummy_magic_29_0.Vb1.n5 0.516125
R17849 two_stage_opamp_dummy_magic_29_0.Vb1_2 two_stage_opamp_dummy_magic_29_0.Vb1_2.t4 74.8571
R17850 two_stage_opamp_dummy_magic_29_0.Vb1_2 two_stage_opamp_dummy_magic_29_0.Vb1_2.n1 54.689
R17851 two_stage_opamp_dummy_magic_29_0.Vb1_2 two_stage_opamp_dummy_magic_29_0.Vb1_2.n0 54.689
R17852 two_stage_opamp_dummy_magic_29_0.Vb1_2.n0 two_stage_opamp_dummy_magic_29_0.Vb1_2.t2 16.0005
R17853 two_stage_opamp_dummy_magic_29_0.Vb1_2.n0 two_stage_opamp_dummy_magic_29_0.Vb1_2.t0 16.0005
R17854 two_stage_opamp_dummy_magic_29_0.Vb1_2.n1 two_stage_opamp_dummy_magic_29_0.Vb1_2.t1 16.0005
R17855 two_stage_opamp_dummy_magic_29_0.Vb1_2.n1 two_stage_opamp_dummy_magic_29_0.Vb1_2.t3 16.0005
R17856 two_stage_opamp_dummy_magic_29_0.VD2.n27 two_stage_opamp_dummy_magic_29_0.VD2.n9 49.7255
R17857 two_stage_opamp_dummy_magic_29_0.VD2.n21 two_stage_opamp_dummy_magic_29_0.VD2.n12 49.7255
R17858 two_stage_opamp_dummy_magic_29_0.VD2.n11 two_stage_opamp_dummy_magic_29_0.VD2.n10 49.7255
R17859 two_stage_opamp_dummy_magic_29_0.VD2.n25 two_stage_opamp_dummy_magic_29_0.VD2.n24 49.7255
R17860 two_stage_opamp_dummy_magic_29_0.VD2.n1 two_stage_opamp_dummy_magic_29_0.VD2.n0 49.7255
R17861 two_stage_opamp_dummy_magic_29_0.VD2.n15 two_stage_opamp_dummy_magic_29_0.VD2.n14 49.3505
R17862 two_stage_opamp_dummy_magic_29_0.VD2.n18 two_stage_opamp_dummy_magic_29_0.VD2.n17 49.3505
R17863 two_stage_opamp_dummy_magic_29_0.VD2.n5 two_stage_opamp_dummy_magic_29_0.VD2.n4 49.3505
R17864 two_stage_opamp_dummy_magic_29_0.VD2.n8 two_stage_opamp_dummy_magic_29_0.VD2.n7 49.3505
R17865 two_stage_opamp_dummy_magic_29_0.VD2.n31 two_stage_opamp_dummy_magic_29_0.VD2.n30 49.3505
R17866 two_stage_opamp_dummy_magic_29_0.VD2.n35 two_stage_opamp_dummy_magic_29_0.VD2.n34 49.3505
R17867 two_stage_opamp_dummy_magic_29_0.VD2.n14 two_stage_opamp_dummy_magic_29_0.VD2.t2 16.0005
R17868 two_stage_opamp_dummy_magic_29_0.VD2.n14 two_stage_opamp_dummy_magic_29_0.VD2.t17 16.0005
R17869 two_stage_opamp_dummy_magic_29_0.VD2.n17 two_stage_opamp_dummy_magic_29_0.VD2.t18 16.0005
R17870 two_stage_opamp_dummy_magic_29_0.VD2.n17 two_stage_opamp_dummy_magic_29_0.VD2.t16 16.0005
R17871 two_stage_opamp_dummy_magic_29_0.VD2.n4 two_stage_opamp_dummy_magic_29_0.VD2.t19 16.0005
R17872 two_stage_opamp_dummy_magic_29_0.VD2.n4 two_stage_opamp_dummy_magic_29_0.VD2.t4 16.0005
R17873 two_stage_opamp_dummy_magic_29_0.VD2.n7 two_stage_opamp_dummy_magic_29_0.VD2.t1 16.0005
R17874 two_stage_opamp_dummy_magic_29_0.VD2.n7 two_stage_opamp_dummy_magic_29_0.VD2.t3 16.0005
R17875 two_stage_opamp_dummy_magic_29_0.VD2.n30 two_stage_opamp_dummy_magic_29_0.VD2.t20 16.0005
R17876 two_stage_opamp_dummy_magic_29_0.VD2.n30 two_stage_opamp_dummy_magic_29_0.VD2.t5 16.0005
R17877 two_stage_opamp_dummy_magic_29_0.VD2.n9 two_stage_opamp_dummy_magic_29_0.VD2.t7 16.0005
R17878 two_stage_opamp_dummy_magic_29_0.VD2.n9 two_stage_opamp_dummy_magic_29_0.VD2.t13 16.0005
R17879 two_stage_opamp_dummy_magic_29_0.VD2.n12 two_stage_opamp_dummy_magic_29_0.VD2.t9 16.0005
R17880 two_stage_opamp_dummy_magic_29_0.VD2.n12 two_stage_opamp_dummy_magic_29_0.VD2.t12 16.0005
R17881 two_stage_opamp_dummy_magic_29_0.VD2.n10 two_stage_opamp_dummy_magic_29_0.VD2.t11 16.0005
R17882 two_stage_opamp_dummy_magic_29_0.VD2.n10 two_stage_opamp_dummy_magic_29_0.VD2.t6 16.0005
R17883 two_stage_opamp_dummy_magic_29_0.VD2.n24 two_stage_opamp_dummy_magic_29_0.VD2.t8 16.0005
R17884 two_stage_opamp_dummy_magic_29_0.VD2.n24 two_stage_opamp_dummy_magic_29_0.VD2.t14 16.0005
R17885 two_stage_opamp_dummy_magic_29_0.VD2.n34 two_stage_opamp_dummy_magic_29_0.VD2.t21 16.0005
R17886 two_stage_opamp_dummy_magic_29_0.VD2.n34 two_stage_opamp_dummy_magic_29_0.VD2.t0 16.0005
R17887 two_stage_opamp_dummy_magic_29_0.VD2.n0 two_stage_opamp_dummy_magic_29_0.VD2.t10 16.0005
R17888 two_stage_opamp_dummy_magic_29_0.VD2.n0 two_stage_opamp_dummy_magic_29_0.VD2.t15 16.0005
R17889 two_stage_opamp_dummy_magic_29_0.VD2.n28 two_stage_opamp_dummy_magic_29_0.VD2.n27 8.89633
R17890 two_stage_opamp_dummy_magic_29_0.VD2.n21 two_stage_opamp_dummy_magic_29_0.VD2.n20 8.89633
R17891 two_stage_opamp_dummy_magic_29_0.VD2.n13 two_stage_opamp_dummy_magic_29_0.VD2.n11 8.89633
R17892 two_stage_opamp_dummy_magic_29_0.VD2.n25 two_stage_opamp_dummy_magic_29_0.VD2.n3 8.89633
R17893 two_stage_opamp_dummy_magic_29_0.VD2.n32 two_stage_opamp_dummy_magic_29_0.VD2.n8 5.438
R17894 two_stage_opamp_dummy_magic_29_0.VD2.n16 two_stage_opamp_dummy_magic_29_0.VD2.n15 5.438
R17895 two_stage_opamp_dummy_magic_29_0.VD2.n28 two_stage_opamp_dummy_magic_29_0.VD2.n8 5.31821
R17896 two_stage_opamp_dummy_magic_29_0.VD2.n15 two_stage_opamp_dummy_magic_29_0.VD2.n13 5.31821
R17897 two_stage_opamp_dummy_magic_29_0.VD2.n19 two_stage_opamp_dummy_magic_29_0.VD2.n18 5.08383
R17898 two_stage_opamp_dummy_magic_29_0.VD2.n5 two_stage_opamp_dummy_magic_29_0.VD2.n2 5.08383
R17899 two_stage_opamp_dummy_magic_29_0.VD2.n31 two_stage_opamp_dummy_magic_29_0.VD2.n29 5.08383
R17900 two_stage_opamp_dummy_magic_29_0.VD2.n36 two_stage_opamp_dummy_magic_29_0.VD2.n35 5.08383
R17901 two_stage_opamp_dummy_magic_29_0.VD2.n27 two_stage_opamp_dummy_magic_29_0.VD2.n26 5.063
R17902 two_stage_opamp_dummy_magic_29_0.VD2.n22 two_stage_opamp_dummy_magic_29_0.VD2.n11 5.063
R17903 two_stage_opamp_dummy_magic_29_0.VD2.n18 two_stage_opamp_dummy_magic_29_0.VD2.n16 4.8755
R17904 two_stage_opamp_dummy_magic_29_0.VD2.n6 two_stage_opamp_dummy_magic_29_0.VD2.n5 4.8755
R17905 two_stage_opamp_dummy_magic_29_0.VD2.n32 two_stage_opamp_dummy_magic_29_0.VD2.n31 4.8755
R17906 two_stage_opamp_dummy_magic_29_0.VD2.n35 two_stage_opamp_dummy_magic_29_0.VD2.n33 4.8755
R17907 two_stage_opamp_dummy_magic_29_0.VD2 two_stage_opamp_dummy_magic_29_0.VD2.n37 4.60467
R17908 two_stage_opamp_dummy_magic_29_0.VD2.n22 two_stage_opamp_dummy_magic_29_0.VD2.n21 4.5005
R17909 two_stage_opamp_dummy_magic_29_0.VD2.n26 two_stage_opamp_dummy_magic_29_0.VD2.n25 4.5005
R17910 two_stage_opamp_dummy_magic_29_0.VD2.n23 two_stage_opamp_dummy_magic_29_0.VD2.n1 4.5005
R17911 two_stage_opamp_dummy_magic_29_0.VD2 two_stage_opamp_dummy_magic_29_0.VD2.n1 4.29217
R17912 two_stage_opamp_dummy_magic_29_0.VD2.n23 two_stage_opamp_dummy_magic_29_0.VD2.n22 0.563
R17913 two_stage_opamp_dummy_magic_29_0.VD2.n26 two_stage_opamp_dummy_magic_29_0.VD2.n23 0.563
R17914 two_stage_opamp_dummy_magic_29_0.VD2.n33 two_stage_opamp_dummy_magic_29_0.VD2.n32 0.563
R17915 two_stage_opamp_dummy_magic_29_0.VD2.n33 two_stage_opamp_dummy_magic_29_0.VD2.n6 0.563
R17916 two_stage_opamp_dummy_magic_29_0.VD2.n16 two_stage_opamp_dummy_magic_29_0.VD2.n6 0.563
R17917 two_stage_opamp_dummy_magic_29_0.VD2.n37 two_stage_opamp_dummy_magic_29_0.VD2.n36 0.234875
R17918 two_stage_opamp_dummy_magic_29_0.VD2.n36 two_stage_opamp_dummy_magic_29_0.VD2.n3 0.234875
R17919 two_stage_opamp_dummy_magic_29_0.VD2.n29 two_stage_opamp_dummy_magic_29_0.VD2.n3 0.234875
R17920 two_stage_opamp_dummy_magic_29_0.VD2.n29 two_stage_opamp_dummy_magic_29_0.VD2.n28 0.234875
R17921 two_stage_opamp_dummy_magic_29_0.VD2.n19 two_stage_opamp_dummy_magic_29_0.VD2.n13 0.234875
R17922 two_stage_opamp_dummy_magic_29_0.VD2.n20 two_stage_opamp_dummy_magic_29_0.VD2.n19 0.234875
R17923 two_stage_opamp_dummy_magic_29_0.VD2.n20 two_stage_opamp_dummy_magic_29_0.VD2.n2 0.234875
R17924 two_stage_opamp_dummy_magic_29_0.VD2.n37 two_stage_opamp_dummy_magic_29_0.VD2.n2 0.234875
R17925 two_stage_opamp_dummy_magic_29_0.VD3.n3 two_stage_opamp_dummy_magic_29_0.VD3.t3 671.418
R17926 two_stage_opamp_dummy_magic_29_0.VD3.n15 two_stage_opamp_dummy_magic_29_0.VD3.t6 671.418
R17927 two_stage_opamp_dummy_magic_29_0.VD3.n14 two_stage_opamp_dummy_magic_29_0.VD3.t7 213.131
R17928 two_stage_opamp_dummy_magic_29_0.VD3.t4 two_stage_opamp_dummy_magic_29_0.VD3.n13 213.131
R17929 two_stage_opamp_dummy_magic_29_0.VD3.t7 two_stage_opamp_dummy_magic_29_0.VD3.t29 146.155
R17930 two_stage_opamp_dummy_magic_29_0.VD3.t29 two_stage_opamp_dummy_magic_29_0.VD3.t33 146.155
R17931 two_stage_opamp_dummy_magic_29_0.VD3.t33 two_stage_opamp_dummy_magic_29_0.VD3.t19 146.155
R17932 two_stage_opamp_dummy_magic_29_0.VD3.t19 two_stage_opamp_dummy_magic_29_0.VD3.t23 146.155
R17933 two_stage_opamp_dummy_magic_29_0.VD3.t23 two_stage_opamp_dummy_magic_29_0.VD3.t25 146.155
R17934 two_stage_opamp_dummy_magic_29_0.VD3.t25 two_stage_opamp_dummy_magic_29_0.VD3.t27 146.155
R17935 two_stage_opamp_dummy_magic_29_0.VD3.t27 two_stage_opamp_dummy_magic_29_0.VD3.t31 146.155
R17936 two_stage_opamp_dummy_magic_29_0.VD3.t31 two_stage_opamp_dummy_magic_29_0.VD3.t35 146.155
R17937 two_stage_opamp_dummy_magic_29_0.VD3.t35 two_stage_opamp_dummy_magic_29_0.VD3.t21 146.155
R17938 two_stage_opamp_dummy_magic_29_0.VD3.t21 two_stage_opamp_dummy_magic_29_0.VD3.t17 146.155
R17939 two_stage_opamp_dummy_magic_29_0.VD3.t17 two_stage_opamp_dummy_magic_29_0.VD3.t4 146.155
R17940 two_stage_opamp_dummy_magic_29_0.VD3.n14 two_stage_opamp_dummy_magic_29_0.VD3.t8 76.2576
R17941 two_stage_opamp_dummy_magic_29_0.VD3.n13 two_stage_opamp_dummy_magic_29_0.VD3.t5 76.2576
R17942 two_stage_opamp_dummy_magic_29_0.VD3.n0 two_stage_opamp_dummy_magic_29_0.VD3.n19 67.013
R17943 two_stage_opamp_dummy_magic_29_0.VD3.n28 two_stage_opamp_dummy_magic_29_0.VD3.n16 67.013
R17944 two_stage_opamp_dummy_magic_29_0.VD3.n12 two_stage_opamp_dummy_magic_29_0.VD3.n11 67.013
R17945 two_stage_opamp_dummy_magic_29_0.VD3.n33 two_stage_opamp_dummy_magic_29_0.VD3.n6 67.013
R17946 two_stage_opamp_dummy_magic_29_0.VD3.n32 two_stage_opamp_dummy_magic_29_0.VD3.n31 67.013
R17947 two_stage_opamp_dummy_magic_29_0.VD3.n5 two_stage_opamp_dummy_magic_29_0.VD3.n4 66.0338
R17948 two_stage_opamp_dummy_magic_29_0.VD3.n8 two_stage_opamp_dummy_magic_29_0.VD3.n7 66.0338
R17949 two_stage_opamp_dummy_magic_29_0.VD3.n10 two_stage_opamp_dummy_magic_29_0.VD3.n9 66.0338
R17950 two_stage_opamp_dummy_magic_29_0.VD3.n23 two_stage_opamp_dummy_magic_29_0.VD3.n22 66.0338
R17951 two_stage_opamp_dummy_magic_29_0.VD3.n18 two_stage_opamp_dummy_magic_29_0.VD3.n17 66.0338
R17952 two_stage_opamp_dummy_magic_29_0.VD3.n27 two_stage_opamp_dummy_magic_29_0.VD3.n26 66.0338
R17953 two_stage_opamp_dummy_magic_29_0.VD3.n19 two_stage_opamp_dummy_magic_29_0.VD3.t30 11.2576
R17954 two_stage_opamp_dummy_magic_29_0.VD3.n19 two_stage_opamp_dummy_magic_29_0.VD3.t34 11.2576
R17955 two_stage_opamp_dummy_magic_29_0.VD3.n16 two_stage_opamp_dummy_magic_29_0.VD3.t20 11.2576
R17956 two_stage_opamp_dummy_magic_29_0.VD3.n16 two_stage_opamp_dummy_magic_29_0.VD3.t24 11.2576
R17957 two_stage_opamp_dummy_magic_29_0.VD3.n11 two_stage_opamp_dummy_magic_29_0.VD3.t26 11.2576
R17958 two_stage_opamp_dummy_magic_29_0.VD3.n11 two_stage_opamp_dummy_magic_29_0.VD3.t28 11.2576
R17959 two_stage_opamp_dummy_magic_29_0.VD3.n6 two_stage_opamp_dummy_magic_29_0.VD3.t22 11.2576
R17960 two_stage_opamp_dummy_magic_29_0.VD3.n6 two_stage_opamp_dummy_magic_29_0.VD3.t18 11.2576
R17961 two_stage_opamp_dummy_magic_29_0.VD3.n4 two_stage_opamp_dummy_magic_29_0.VD3.t12 11.2576
R17962 two_stage_opamp_dummy_magic_29_0.VD3.n4 two_stage_opamp_dummy_magic_29_0.VD3.t15 11.2576
R17963 two_stage_opamp_dummy_magic_29_0.VD3.n7 two_stage_opamp_dummy_magic_29_0.VD3.t14 11.2576
R17964 two_stage_opamp_dummy_magic_29_0.VD3.n7 two_stage_opamp_dummy_magic_29_0.VD3.t2 11.2576
R17965 two_stage_opamp_dummy_magic_29_0.VD3.n9 two_stage_opamp_dummy_magic_29_0.VD3.t1 11.2576
R17966 two_stage_opamp_dummy_magic_29_0.VD3.n9 two_stage_opamp_dummy_magic_29_0.VD3.t10 11.2576
R17967 two_stage_opamp_dummy_magic_29_0.VD3.n22 two_stage_opamp_dummy_magic_29_0.VD3.t13 11.2576
R17968 two_stage_opamp_dummy_magic_29_0.VD3.n22 two_stage_opamp_dummy_magic_29_0.VD3.t9 11.2576
R17969 two_stage_opamp_dummy_magic_29_0.VD3.n17 two_stage_opamp_dummy_magic_29_0.VD3.t37 11.2576
R17970 two_stage_opamp_dummy_magic_29_0.VD3.n17 two_stage_opamp_dummy_magic_29_0.VD3.t11 11.2576
R17971 two_stage_opamp_dummy_magic_29_0.VD3.n26 two_stage_opamp_dummy_magic_29_0.VD3.t16 11.2576
R17972 two_stage_opamp_dummy_magic_29_0.VD3.n26 two_stage_opamp_dummy_magic_29_0.VD3.t0 11.2576
R17973 two_stage_opamp_dummy_magic_29_0.VD3.n31 two_stage_opamp_dummy_magic_29_0.VD3.t32 11.2576
R17974 two_stage_opamp_dummy_magic_29_0.VD3.n31 two_stage_opamp_dummy_magic_29_0.VD3.t36 11.2576
R17975 two_stage_opamp_dummy_magic_29_0.VD3.n27 two_stage_opamp_dummy_magic_29_0.VD3.n25 5.66717
R17976 two_stage_opamp_dummy_magic_29_0.VD3.n20 two_stage_opamp_dummy_magic_29_0.VD3.n5 5.66717
R17977 two_stage_opamp_dummy_magic_29_0.VD3.n20 two_stage_opamp_dummy_magic_29_0.VD3.n8 5.29217
R17978 two_stage_opamp_dummy_magic_29_0.VD3.n21 two_stage_opamp_dummy_magic_29_0.VD3.n10 5.29217
R17979 two_stage_opamp_dummy_magic_29_0.VD3.n24 two_stage_opamp_dummy_magic_29_0.VD3.n23 5.29217
R17980 two_stage_opamp_dummy_magic_29_0.VD3.n25 two_stage_opamp_dummy_magic_29_0.VD3.n18 5.29217
R17981 two_stage_opamp_dummy_magic_29_0.VD3.n15 two_stage_opamp_dummy_magic_29_0.VD3.n14 1.90883
R17982 two_stage_opamp_dummy_magic_29_0.VD3.n13 two_stage_opamp_dummy_magic_29_0.VD3.n3 1.90883
R17983 two_stage_opamp_dummy_magic_29_0.VD3.n33 two_stage_opamp_dummy_magic_29_0.VD3.n8 1.02133
R17984 two_stage_opamp_dummy_magic_29_0.VD3.n32 two_stage_opamp_dummy_magic_29_0.VD3.n10 1.02133
R17985 two_stage_opamp_dummy_magic_29_0.VD3.n23 two_stage_opamp_dummy_magic_29_0.VD3.n12 1.02133
R17986 two_stage_opamp_dummy_magic_29_0.VD3.n28 two_stage_opamp_dummy_magic_29_0.VD3.n18 1.02133
R17987 two_stage_opamp_dummy_magic_29_0.VD3.n0 two_stage_opamp_dummy_magic_29_0.VD3.n27 1.02133
R17988 two_stage_opamp_dummy_magic_29_0.VD3.n34 two_stage_opamp_dummy_magic_29_0.VD3.n5 1.02133
R17989 two_stage_opamp_dummy_magic_29_0.VD3 two_stage_opamp_dummy_magic_29_0.VD3.n34 0.65675
R17990 two_stage_opamp_dummy_magic_29_0.VD3.n33 two_stage_opamp_dummy_magic_29_0.VD3.n2 0.643357
R17991 two_stage_opamp_dummy_magic_29_0.VD3.n32 two_stage_opamp_dummy_magic_29_0.VD3.n30 0.643357
R17992 two_stage_opamp_dummy_magic_29_0.VD3.n29 two_stage_opamp_dummy_magic_29_0.VD3.n12 0.643357
R17993 two_stage_opamp_dummy_magic_29_0.VD3.n1 two_stage_opamp_dummy_magic_29_0.VD3.n0 0.0279681
R17994 two_stage_opamp_dummy_magic_29_0.VD3.n25 two_stage_opamp_dummy_magic_29_0.VD3.n24 0.3755
R17995 two_stage_opamp_dummy_magic_29_0.VD3.n24 two_stage_opamp_dummy_magic_29_0.VD3.n21 0.3755
R17996 two_stage_opamp_dummy_magic_29_0.VD3.n21 two_stage_opamp_dummy_magic_29_0.VD3.n20 0.3755
R17997 two_stage_opamp_dummy_magic_29_0.VD3.n0 two_stage_opamp_dummy_magic_29_0.VD3.n15 0.131952
R17998 two_stage_opamp_dummy_magic_29_0.VD3.n34 two_stage_opamp_dummy_magic_29_0.VD3.n3 0.104667
R17999 two_stage_opamp_dummy_magic_29_0.VD3.n28 two_stage_opamp_dummy_magic_29_0.VD3.n1 0.0471695
R18000 two_stage_opamp_dummy_magic_29_0.VD3.n29 two_stage_opamp_dummy_magic_29_0.VD3.n1 0.274589
R18001 two_stage_opamp_dummy_magic_29_0.VD3.n30 two_stage_opamp_dummy_magic_29_0.VD3.n29 0.0540714
R18002 two_stage_opamp_dummy_magic_29_0.VD3.n30 two_stage_opamp_dummy_magic_29_0.VD3.n2 0.0540714
R18003 two_stage_opamp_dummy_magic_29_0.VD3.n28 two_stage_opamp_dummy_magic_29_0.VD3.n12 0.0540714
R18004 two_stage_opamp_dummy_magic_29_0.VD3.n32 two_stage_opamp_dummy_magic_29_0.VD3.n12 0.0540714
R18005 two_stage_opamp_dummy_magic_29_0.VD3.n33 two_stage_opamp_dummy_magic_29_0.VD3.n32 0.0540714
R18006 two_stage_opamp_dummy_magic_29_0.VD3.n34 two_stage_opamp_dummy_magic_29_0.VD3.n33 0.0540714
R18007 two_stage_opamp_dummy_magic_29_0.VD3 two_stage_opamp_dummy_magic_29_0.VD3.n2 0.0406786
R18008 two_stage_opamp_dummy_magic_29_0.Vb3.n16 two_stage_opamp_dummy_magic_29_0.Vb3.t19 793.28
R18009 two_stage_opamp_dummy_magic_29_0.Vb3.n9 two_stage_opamp_dummy_magic_29_0.Vb3.t22 752.422
R18010 two_stage_opamp_dummy_magic_29_0.Vb3.n0 two_stage_opamp_dummy_magic_29_0.Vb3.t28 752.422
R18011 two_stage_opamp_dummy_magic_29_0.Vb3.n9 two_stage_opamp_dummy_magic_29_0.Vb3.t18 752.234
R18012 two_stage_opamp_dummy_magic_29_0.Vb3.n9 two_stage_opamp_dummy_magic_29_0.Vb3.t25 752.234
R18013 two_stage_opamp_dummy_magic_29_0.Vb3.n8 two_stage_opamp_dummy_magic_29_0.Vb3.t11 752.234
R18014 two_stage_opamp_dummy_magic_29_0.Vb3.n6 two_stage_opamp_dummy_magic_29_0.Vb3.t14 752.234
R18015 two_stage_opamp_dummy_magic_29_0.Vb3.n7 two_stage_opamp_dummy_magic_29_0.Vb3.t20 752.234
R18016 two_stage_opamp_dummy_magic_29_0.Vb3.n7 two_stage_opamp_dummy_magic_29_0.Vb3.t26 752.234
R18017 two_stage_opamp_dummy_magic_29_0.Vb3.n20 two_stage_opamp_dummy_magic_29_0.Vb3.t8 752.234
R18018 two_stage_opamp_dummy_magic_29_0.Vb3.n5 two_stage_opamp_dummy_magic_29_0.Vb3.t17 752.234
R18019 two_stage_opamp_dummy_magic_29_0.Vb3.n5 two_stage_opamp_dummy_magic_29_0.Vb3.t24 752.234
R18020 two_stage_opamp_dummy_magic_29_0.Vb3.n4 two_stage_opamp_dummy_magic_29_0.Vb3.t21 752.234
R18021 two_stage_opamp_dummy_magic_29_0.Vb3.n4 two_stage_opamp_dummy_magic_29_0.Vb3.t27 752.234
R18022 two_stage_opamp_dummy_magic_29_0.Vb3.n1 two_stage_opamp_dummy_magic_29_0.Vb3.t12 752.234
R18023 two_stage_opamp_dummy_magic_29_0.Vb3.n1 two_stage_opamp_dummy_magic_29_0.Vb3.t15 752.234
R18024 two_stage_opamp_dummy_magic_29_0.Vb3.n0 two_stage_opamp_dummy_magic_29_0.Vb3.t23 752.234
R18025 two_stage_opamp_dummy_magic_29_0.Vb3.n18 two_stage_opamp_dummy_magic_29_0.Vb3.t13 747.734
R18026 two_stage_opamp_dummy_magic_29_0.Vb3.n19 two_stage_opamp_dummy_magic_29_0.Vb3.t16 747.734
R18027 two_stage_opamp_dummy_magic_29_0.Vb3.n3 two_stage_opamp_dummy_magic_29_0.Vb3.t10 747.827
R18028 two_stage_opamp_dummy_magic_29_0.Vb3.n12 two_stage_opamp_dummy_magic_29_0.Vb3.n10 139.639
R18029 two_stage_opamp_dummy_magic_29_0.Vb3.n12 two_stage_opamp_dummy_magic_29_0.Vb3.n11 139.638
R18030 two_stage_opamp_dummy_magic_29_0.Vb3.n14 two_stage_opamp_dummy_magic_29_0.Vb3.n13 134.577
R18031 two_stage_opamp_dummy_magic_29_0.Vb3.n16 two_stage_opamp_dummy_magic_29_0.Vb3.n15 72.612
R18032 bgr_11_0.VB3_CUR_BIAS two_stage_opamp_dummy_magic_29_0.Vb3.n21 44.688
R18033 bgr_11_0.VB3_CUR_BIAS two_stage_opamp_dummy_magic_29_0.Vb3.n14 43.0317
R18034 two_stage_opamp_dummy_magic_29_0.Vb3.n11 two_stage_opamp_dummy_magic_29_0.Vb3.t1 24.0005
R18035 two_stage_opamp_dummy_magic_29_0.Vb3.n11 two_stage_opamp_dummy_magic_29_0.Vb3.t2 24.0005
R18036 two_stage_opamp_dummy_magic_29_0.Vb3.n10 two_stage_opamp_dummy_magic_29_0.Vb3.t0 24.0005
R18037 two_stage_opamp_dummy_magic_29_0.Vb3.n10 two_stage_opamp_dummy_magic_29_0.Vb3.t3 24.0005
R18038 two_stage_opamp_dummy_magic_29_0.Vb3.n13 two_stage_opamp_dummy_magic_29_0.Vb3.t5 24.0005
R18039 two_stage_opamp_dummy_magic_29_0.Vb3.n13 two_stage_opamp_dummy_magic_29_0.Vb3.t4 24.0005
R18040 two_stage_opamp_dummy_magic_29_0.Vb3.n15 two_stage_opamp_dummy_magic_29_0.Vb3.t6 11.2576
R18041 two_stage_opamp_dummy_magic_29_0.Vb3.n15 two_stage_opamp_dummy_magic_29_0.Vb3.t7 11.2576
R18042 two_stage_opamp_dummy_magic_29_0.Vb3.n17 two_stage_opamp_dummy_magic_29_0.Vb3.n16 11.2036
R18043 two_stage_opamp_dummy_magic_29_0.Vb3.n21 two_stage_opamp_dummy_magic_29_0.Vb3.n17 6.14112
R18044 two_stage_opamp_dummy_magic_29_0.Vb3.n2 two_stage_opamp_dummy_magic_29_0.Vb3.n3 2.20508
R18045 two_stage_opamp_dummy_magic_29_0.Vb3.n6 two_stage_opamp_dummy_magic_29_0.Vb3.n19 4.5005
R18046 two_stage_opamp_dummy_magic_29_0.Vb3.n18 two_stage_opamp_dummy_magic_29_0.Vb3.n8 4.5005
R18047 two_stage_opamp_dummy_magic_29_0.Vb3.n14 two_stage_opamp_dummy_magic_29_0.Vb3.n12 4.5005
R18048 two_stage_opamp_dummy_magic_29_0.Vb3.n17 two_stage_opamp_dummy_magic_29_0.Vb3.n5 3.21925
R18049 two_stage_opamp_dummy_magic_29_0.Vb3.n21 two_stage_opamp_dummy_magic_29_0.Vb3.n20 0.641125
R18050 two_stage_opamp_dummy_magic_29_0.Vb3.n8 two_stage_opamp_dummy_magic_29_0.Vb3.n9 0.3755
R18051 two_stage_opamp_dummy_magic_29_0.Vb3.n6 two_stage_opamp_dummy_magic_29_0.Vb3.n8 0.3755
R18052 two_stage_opamp_dummy_magic_29_0.Vb3.n7 two_stage_opamp_dummy_magic_29_0.Vb3.n6 0.3755
R18053 two_stage_opamp_dummy_magic_29_0.Vb3.n20 two_stage_opamp_dummy_magic_29_0.Vb3.n7 0.3755
R18054 two_stage_opamp_dummy_magic_29_0.Vb3.n5 two_stage_opamp_dummy_magic_29_0.Vb3.n4 0.3755
R18055 two_stage_opamp_dummy_magic_29_0.Vb3.n4 two_stage_opamp_dummy_magic_29_0.Vb3.n2 0.3755
R18056 two_stage_opamp_dummy_magic_29_0.Vb3.n2 two_stage_opamp_dummy_magic_29_0.Vb3.n1 0.3755
R18057 two_stage_opamp_dummy_magic_29_0.Vb3.n19 two_stage_opamp_dummy_magic_29_0.Vb3.n18 0.188
R18058 two_stage_opamp_dummy_magic_29_0.Vb3.t9 two_stage_opamp_dummy_magic_29_0.Vb3.n3 747.827
R18059 two_stage_opamp_dummy_magic_29_0.Vb3.n1 two_stage_opamp_dummy_magic_29_0.Vb3.n0 0.3755
R18060 a_6350_30238.t0 a_6350_30238.t1 178.133
R18061 bgr_11_0.Vin+ bgr_11_0.Vin+.t6 529.879
R18062 bgr_11_0.Vin+.n0 bgr_11_0.Vin+.t5 148.653
R18063 bgr_11_0.Vin+.n0 bgr_11_0.Vin+.t4 125.418
R18064 bgr_11_0.Vin+.n3 bgr_11_0.Vin+.n1 106.609
R18065 bgr_11_0.Vin+.n3 bgr_11_0.Vin+.n2 104.484
R18066 bgr_11_0.Vin+.n4 bgr_11_0.Vin+.n0 25.0809
R18067 bgr_11_0.Vin+.n4 bgr_11_0.Vin+.n3 18.7817
R18068 bgr_11_0.Vin+.n2 bgr_11_0.Vin+.t2 13.1338
R18069 bgr_11_0.Vin+.n2 bgr_11_0.Vin+.t1 13.1338
R18070 bgr_11_0.Vin+.n1 bgr_11_0.Vin+.t0 13.1338
R18071 bgr_11_0.Vin+.n1 bgr_11_0.Vin+.t3 13.1338
R18072 bgr_11_0.Vin+ bgr_11_0.Vin+.n4 6.53175
R18073 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n3 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n2 301.983
R18074 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n5 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n4 297.151
R18075 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n1 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n0 297.151
R18076 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n16 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n15 118.861
R18077 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n18 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n17 118.861
R18078 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n22 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n21 118.861
R18079 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n25 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n24 118.861
R18080 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n28 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n27 118.861
R18081 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n30 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.t0 115.672
R18082 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n4 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.t5 39.4005
R18083 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n4 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.t4 39.4005
R18084 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n2 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.t2 39.4005
R18085 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n2 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.t1 39.4005
R18086 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n0 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.t3 39.4005
R18087 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n0 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.t6 39.4005
R18088 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n15 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.t14 19.7005
R18089 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n15 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.t7 19.7005
R18090 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n17 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.t11 19.7005
R18091 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n17 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.t16 19.7005
R18092 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n21 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.t10 19.7005
R18093 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n21 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.t15 19.7005
R18094 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n24 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.t13 19.7005
R18095 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n24 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.t9 19.7005
R18096 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n27 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.t12 19.7005
R18097 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n27 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.t8 19.7005
R18098 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n41 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n40 13.2453
R18099 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n41 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n5 11.912
R18100 bgr_11_0.V_CMFB_S3 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n41 9.8755
R18101 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n28 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n26 5.54217
R18102 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n16 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n14 5.54217
R18103 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n3 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n1 5.39633
R18104 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n5 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n3 5.39633
R18105 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n19 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n16 5.38592
R18106 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n19 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n18 5.04217
R18107 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n22 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n20 5.04217
R18108 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n25 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n13 5.04217
R18109 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n29 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n28 5.04217
R18110 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n18 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n14 4.97967
R18111 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n23 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n22 4.97967
R18112 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n26 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n25 4.97967
R18113 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n36 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n7 4.5005
R18114 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n38 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n37 4.5005
R18115 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n37 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n36 4.5005
R18116 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n12 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n11 4.5005
R18117 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n30 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n29 2.99007
R18118 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n33 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n32 2.26187
R18119 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n34 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n33 2.26187
R18120 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n39 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n38 2.24063
R18121 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n9 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n8 2.24063
R18122 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n31 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n10 2.24063
R18123 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n40 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n6 2.24063
R18124 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n35 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n34 2.24063
R18125 bgr_11_0.V_CMFB_S3 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n1 1.34946
R18126 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n26 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n23 0.563
R18127 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n23 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n14 0.563
R18128 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n31 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n30 0.464042
R18129 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n20 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n19 0.34425
R18130 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n20 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n13 0.34425
R18131 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n29 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n13 0.34425
R18132 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n36 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n35 0.078625
R18133 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n38 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n8 0.0421667
R18134 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n40 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n39 0.0217373
R18135 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n37 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n9 0.0217373
R18136 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n35 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n10 0.0217373
R18137 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n39 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n7 0.0217373
R18138 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n9 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n7 0.0217373
R18139 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n32 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n11 0.0217373
R18140 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n12 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n10 0.0217373
R18141 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n32 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n31 0.0217373
R18142 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n33 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n12 0.0217373
R18143 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n36 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n6 0.0217373
R18144 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n8 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n6 0.0217373
R18145 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n34 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n11 0.0217373
R18146 two_stage_opamp_dummy_magic_29_0.V_err_gate.n2 two_stage_opamp_dummy_magic_29_0.V_err_gate.t7 479.322
R18147 two_stage_opamp_dummy_magic_29_0.V_err_gate.n2 two_stage_opamp_dummy_magic_29_0.V_err_gate.t9 479.322
R18148 two_stage_opamp_dummy_magic_29_0.V_err_gate.n6 two_stage_opamp_dummy_magic_29_0.V_err_gate.t6 479.322
R18149 two_stage_opamp_dummy_magic_29_0.V_err_gate.n6 two_stage_opamp_dummy_magic_29_0.V_err_gate.t8 479.322
R18150 two_stage_opamp_dummy_magic_29_0.V_err_gate.n3 two_stage_opamp_dummy_magic_29_0.V_err_gate.n1 178.075
R18151 two_stage_opamp_dummy_magic_29_0.V_err_gate.n5 two_stage_opamp_dummy_magic_29_0.V_err_gate.n4 177.434
R18152 two_stage_opamp_dummy_magic_29_0.V_err_gate two_stage_opamp_dummy_magic_29_0.V_err_gate.n0 170.357
R18153 two_stage_opamp_dummy_magic_29_0.V_err_gate.n3 two_stage_opamp_dummy_magic_29_0.V_err_gate.n2 165.8
R18154 two_stage_opamp_dummy_magic_29_0.V_err_gate two_stage_opamp_dummy_magic_29_0.V_err_gate.n6 165.8
R18155 two_stage_opamp_dummy_magic_29_0.V_err_gate.n0 two_stage_opamp_dummy_magic_29_0.V_err_gate.t1 24.0005
R18156 two_stage_opamp_dummy_magic_29_0.V_err_gate.n0 two_stage_opamp_dummy_magic_29_0.V_err_gate.t2 24.0005
R18157 two_stage_opamp_dummy_magic_29_0.V_err_gate.n4 two_stage_opamp_dummy_magic_29_0.V_err_gate.t3 15.7605
R18158 two_stage_opamp_dummy_magic_29_0.V_err_gate.n4 two_stage_opamp_dummy_magic_29_0.V_err_gate.t5 15.7605
R18159 two_stage_opamp_dummy_magic_29_0.V_err_gate.n1 two_stage_opamp_dummy_magic_29_0.V_err_gate.t0 15.7605
R18160 two_stage_opamp_dummy_magic_29_0.V_err_gate.n1 two_stage_opamp_dummy_magic_29_0.V_err_gate.t4 15.7605
R18161 two_stage_opamp_dummy_magic_29_0.V_err_gate two_stage_opamp_dummy_magic_29_0.V_err_gate.n5 1.76612
R18162 two_stage_opamp_dummy_magic_29_0.V_err_gate.n5 two_stage_opamp_dummy_magic_29_0.V_err_gate.n3 0.641125
R18163 a_6540_22450.n11 a_6540_22450.t18 310.488
R18164 a_6540_22450.n5 a_6540_22450.t13 310.488
R18165 a_6540_22450.n0 a_6540_22450.t14 310.488
R18166 a_6540_22450.n9 a_6540_22450.n8 297.433
R18167 a_6540_22450.n4 a_6540_22450.n3 297.433
R18168 a_6540_22450.n15 a_6540_22450.n14 297.433
R18169 a_6540_22450.n13 a_6540_22450.t7 184.097
R18170 a_6540_22450.n7 a_6540_22450.t5 184.097
R18171 a_6540_22450.n2 a_6540_22450.t3 184.097
R18172 a_6540_22450.n12 a_6540_22450.n11 167.094
R18173 a_6540_22450.n6 a_6540_22450.n5 167.094
R18174 a_6540_22450.n1 a_6540_22450.n0 167.094
R18175 a_6540_22450.n14 a_6540_22450.n13 161.3
R18176 a_6540_22450.n9 a_6540_22450.n7 161.3
R18177 a_6540_22450.n4 a_6540_22450.n2 161.3
R18178 a_6540_22450.n11 a_6540_22450.t15 120.501
R18179 a_6540_22450.n12 a_6540_22450.t11 120.501
R18180 a_6540_22450.n5 a_6540_22450.t17 120.501
R18181 a_6540_22450.n6 a_6540_22450.t1 120.501
R18182 a_6540_22450.n0 a_6540_22450.t16 120.501
R18183 a_6540_22450.n1 a_6540_22450.t9 120.501
R18184 a_6540_22450.n9 a_6540_22450.t0 50.2004
R18185 a_6540_22450.n13 a_6540_22450.n12 40.7027
R18186 a_6540_22450.n7 a_6540_22450.n6 40.7027
R18187 a_6540_22450.n2 a_6540_22450.n1 40.7027
R18188 a_6540_22450.n8 a_6540_22450.t2 39.4005
R18189 a_6540_22450.n8 a_6540_22450.t6 39.4005
R18190 a_6540_22450.n3 a_6540_22450.t10 39.4005
R18191 a_6540_22450.n3 a_6540_22450.t4 39.4005
R18192 a_6540_22450.t12 a_6540_22450.n15 39.4005
R18193 a_6540_22450.n15 a_6540_22450.t8 39.4005
R18194 a_6540_22450.n10 a_6540_22450.n4 6.6255
R18195 a_6540_22450.n14 a_6540_22450.n10 6.6255
R18196 a_6540_22450.n10 a_6540_22450.n9 4.5005
R18197 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n20 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.t1 115.6
R18198 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n2 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n0 107.121
R18199 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n2 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n1 97.4332
R18200 bgr_11_0.V_CMFB_S4 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n2 28.6724
R18201 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n6 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n5 24.288
R18202 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n8 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n7 24.288
R18203 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n12 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n11 24.288
R18204 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n15 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n14 24.288
R18205 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n18 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n17 24.288
R18206 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n0 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.t0 24.0005
R18207 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n0 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.t4 24.0005
R18208 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n1 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.t3 24.0005
R18209 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n1 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.t2 24.0005
R18210 bgr_11_0.V_CMFB_S4 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n20 19.0422
R18211 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n5 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.t13 8.0005
R18212 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n5 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.t6 8.0005
R18213 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n7 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.t10 8.0005
R18214 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n7 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.t5 8.0005
R18215 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n11 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.t9 8.0005
R18216 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n11 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.t14 8.0005
R18217 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n14 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.t12 8.0005
R18218 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n14 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.t8 8.0005
R18219 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n17 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.t11 8.0005
R18220 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n17 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.t7 8.0005
R18221 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n18 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n16 5.7505
R18222 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n6 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n4 5.7505
R18223 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n9 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n6 5.53175
R18224 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n9 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n8 5.188
R18225 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n8 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n4 5.188
R18226 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n12 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n10 5.188
R18227 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n13 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n12 5.188
R18228 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n15 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n3 5.188
R18229 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n16 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n15 5.188
R18230 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n19 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n18 5.188
R18231 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n20 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n19 2.38069
R18232 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n16 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n13 0.563
R18233 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n13 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n4 0.563
R18234 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n10 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n9 0.34425
R18235 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n10 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n3 0.34425
R18236 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n19 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n3 0.34425
R18237 VIN+.n0 VIN+.t10 1097.62
R18238 VIN+ VIN+.n9 433.019
R18239 VIN+.n9 VIN+.t5 273.134
R18240 VIN+.n0 VIN+.t7 273.134
R18241 VIN+.n8 VIN+.t1 273.134
R18242 VIN+.n7 VIN+.t4 273.134
R18243 VIN+.n6 VIN+.t0 273.134
R18244 VIN+.n5 VIN+.t3 273.134
R18245 VIN+.n4 VIN+.t8 273.134
R18246 VIN+.n3 VIN+.t6 273.134
R18247 VIN+.n2 VIN+.t9 273.134
R18248 VIN+.n1 VIN+.t2 273.134
R18249 VIN+.n1 VIN+.n0 176.733
R18250 VIN+.n2 VIN+.n1 176.733
R18251 VIN+.n3 VIN+.n2 176.733
R18252 VIN+.n4 VIN+.n3 176.733
R18253 VIN+.n5 VIN+.n4 176.733
R18254 VIN+.n6 VIN+.n5 176.733
R18255 VIN+.n7 VIN+.n6 176.733
R18256 VIN+.n8 VIN+.n7 176.733
R18257 VIN+.n9 VIN+.n8 176.733
R18258 two_stage_opamp_dummy_magic_29_0.V_source.n56 two_stage_opamp_dummy_magic_29_0.V_source.t23 67.545
R18259 two_stage_opamp_dummy_magic_29_0.V_source.n15 two_stage_opamp_dummy_magic_29_0.V_source.n14 49.3505
R18260 two_stage_opamp_dummy_magic_29_0.V_source.n17 two_stage_opamp_dummy_magic_29_0.V_source.n16 49.3505
R18261 two_stage_opamp_dummy_magic_29_0.V_source.n21 two_stage_opamp_dummy_magic_29_0.V_source.n20 49.3505
R18262 two_stage_opamp_dummy_magic_29_0.V_source.n33 two_stage_opamp_dummy_magic_29_0.V_source.n32 49.3505
R18263 two_stage_opamp_dummy_magic_29_0.V_source.n30 two_stage_opamp_dummy_magic_29_0.V_source.n29 49.3505
R18264 two_stage_opamp_dummy_magic_29_0.V_source.n27 two_stage_opamp_dummy_magic_29_0.V_source.n26 49.3505
R18265 two_stage_opamp_dummy_magic_29_0.V_source.n25 two_stage_opamp_dummy_magic_29_0.V_source.n24 49.3505
R18266 two_stage_opamp_dummy_magic_29_0.V_source.n42 two_stage_opamp_dummy_magic_29_0.V_source.n41 49.3505
R18267 two_stage_opamp_dummy_magic_29_0.V_source.n36 two_stage_opamp_dummy_magic_29_0.V_source.n35 49.3505
R18268 two_stage_opamp_dummy_magic_29_0.V_source.n38 two_stage_opamp_dummy_magic_29_0.V_source.n37 49.3505
R18269 two_stage_opamp_dummy_magic_29_0.V_source.n60 two_stage_opamp_dummy_magic_29_0.V_source.n59 32.3838
R18270 two_stage_opamp_dummy_magic_29_0.V_source.n48 two_stage_opamp_dummy_magic_29_0.V_source.n47 32.3838
R18271 two_stage_opamp_dummy_magic_29_0.V_source.n46 two_stage_opamp_dummy_magic_29_0.V_source.n45 32.3838
R18272 two_stage_opamp_dummy_magic_29_0.V_source.n5 two_stage_opamp_dummy_magic_29_0.V_source.n4 32.3838
R18273 two_stage_opamp_dummy_magic_29_0.V_source.n50 two_stage_opamp_dummy_magic_29_0.V_source.n49 32.3838
R18274 two_stage_opamp_dummy_magic_29_0.V_source.n53 two_stage_opamp_dummy_magic_29_0.V_source.n52 32.3838
R18275 two_stage_opamp_dummy_magic_29_0.V_source.n8 two_stage_opamp_dummy_magic_29_0.V_source.n7 32.3838
R18276 two_stage_opamp_dummy_magic_29_0.V_source.n63 two_stage_opamp_dummy_magic_29_0.V_source.n62 32.3838
R18277 two_stage_opamp_dummy_magic_29_0.V_source.n66 two_stage_opamp_dummy_magic_29_0.V_source.n65 32.3838
R18278 two_stage_opamp_dummy_magic_29_0.V_source.n70 two_stage_opamp_dummy_magic_29_0.V_source.n69 32.3838
R18279 two_stage_opamp_dummy_magic_29_0.V_source.n14 two_stage_opamp_dummy_magic_29_0.V_source.t15 16.0005
R18280 two_stage_opamp_dummy_magic_29_0.V_source.n14 two_stage_opamp_dummy_magic_29_0.V_source.t24 16.0005
R18281 two_stage_opamp_dummy_magic_29_0.V_source.n16 two_stage_opamp_dummy_magic_29_0.V_source.t3 16.0005
R18282 two_stage_opamp_dummy_magic_29_0.V_source.n16 two_stage_opamp_dummy_magic_29_0.V_source.t14 16.0005
R18283 two_stage_opamp_dummy_magic_29_0.V_source.n20 two_stage_opamp_dummy_magic_29_0.V_source.t10 16.0005
R18284 two_stage_opamp_dummy_magic_29_0.V_source.n20 two_stage_opamp_dummy_magic_29_0.V_source.t19 16.0005
R18285 two_stage_opamp_dummy_magic_29_0.V_source.n32 two_stage_opamp_dummy_magic_29_0.V_source.t28 16.0005
R18286 two_stage_opamp_dummy_magic_29_0.V_source.n32 two_stage_opamp_dummy_magic_29_0.V_source.t31 16.0005
R18287 two_stage_opamp_dummy_magic_29_0.V_source.n29 two_stage_opamp_dummy_magic_29_0.V_source.t30 16.0005
R18288 two_stage_opamp_dummy_magic_29_0.V_source.n29 two_stage_opamp_dummy_magic_29_0.V_source.t35 16.0005
R18289 two_stage_opamp_dummy_magic_29_0.V_source.n26 two_stage_opamp_dummy_magic_29_0.V_source.t39 16.0005
R18290 two_stage_opamp_dummy_magic_29_0.V_source.n26 two_stage_opamp_dummy_magic_29_0.V_source.t9 16.0005
R18291 two_stage_opamp_dummy_magic_29_0.V_source.n24 two_stage_opamp_dummy_magic_29_0.V_source.t4 16.0005
R18292 two_stage_opamp_dummy_magic_29_0.V_source.n24 two_stage_opamp_dummy_magic_29_0.V_source.t6 16.0005
R18293 two_stage_opamp_dummy_magic_29_0.V_source.n41 two_stage_opamp_dummy_magic_29_0.V_source.t29 16.0005
R18294 two_stage_opamp_dummy_magic_29_0.V_source.n41 two_stage_opamp_dummy_magic_29_0.V_source.t34 16.0005
R18295 two_stage_opamp_dummy_magic_29_0.V_source.n35 two_stage_opamp_dummy_magic_29_0.V_source.t36 16.0005
R18296 two_stage_opamp_dummy_magic_29_0.V_source.n35 two_stage_opamp_dummy_magic_29_0.V_source.t32 16.0005
R18297 two_stage_opamp_dummy_magic_29_0.V_source.n37 two_stage_opamp_dummy_magic_29_0.V_source.t37 16.0005
R18298 two_stage_opamp_dummy_magic_29_0.V_source.n37 two_stage_opamp_dummy_magic_29_0.V_source.t33 16.0005
R18299 two_stage_opamp_dummy_magic_29_0.V_source.n59 two_stage_opamp_dummy_magic_29_0.V_source.t17 9.6005
R18300 two_stage_opamp_dummy_magic_29_0.V_source.n59 two_stage_opamp_dummy_magic_29_0.V_source.t12 9.6005
R18301 two_stage_opamp_dummy_magic_29_0.V_source.n47 two_stage_opamp_dummy_magic_29_0.V_source.t8 9.6005
R18302 two_stage_opamp_dummy_magic_29_0.V_source.n47 two_stage_opamp_dummy_magic_29_0.V_source.t38 9.6005
R18303 two_stage_opamp_dummy_magic_29_0.V_source.n45 two_stage_opamp_dummy_magic_29_0.V_source.t16 9.6005
R18304 two_stage_opamp_dummy_magic_29_0.V_source.n45 two_stage_opamp_dummy_magic_29_0.V_source.t25 9.6005
R18305 two_stage_opamp_dummy_magic_29_0.V_source.n4 two_stage_opamp_dummy_magic_29_0.V_source.t40 9.6005
R18306 two_stage_opamp_dummy_magic_29_0.V_source.n4 two_stage_opamp_dummy_magic_29_0.V_source.t22 9.6005
R18307 two_stage_opamp_dummy_magic_29_0.V_source.n49 two_stage_opamp_dummy_magic_29_0.V_source.t11 9.6005
R18308 two_stage_opamp_dummy_magic_29_0.V_source.n49 two_stage_opamp_dummy_magic_29_0.V_source.t20 9.6005
R18309 two_stage_opamp_dummy_magic_29_0.V_source.n52 two_stage_opamp_dummy_magic_29_0.V_source.t18 9.6005
R18310 two_stage_opamp_dummy_magic_29_0.V_source.n52 two_stage_opamp_dummy_magic_29_0.V_source.t2 9.6005
R18311 two_stage_opamp_dummy_magic_29_0.V_source.n7 two_stage_opamp_dummy_magic_29_0.V_source.t21 9.6005
R18312 two_stage_opamp_dummy_magic_29_0.V_source.n7 two_stage_opamp_dummy_magic_29_0.V_source.t27 9.6005
R18313 two_stage_opamp_dummy_magic_29_0.V_source.n62 two_stage_opamp_dummy_magic_29_0.V_source.t13 9.6005
R18314 two_stage_opamp_dummy_magic_29_0.V_source.n62 two_stage_opamp_dummy_magic_29_0.V_source.t1 9.6005
R18315 two_stage_opamp_dummy_magic_29_0.V_source.n65 two_stage_opamp_dummy_magic_29_0.V_source.t7 9.6005
R18316 two_stage_opamp_dummy_magic_29_0.V_source.n65 two_stage_opamp_dummy_magic_29_0.V_source.t26 9.6005
R18317 two_stage_opamp_dummy_magic_29_0.V_source.n69 two_stage_opamp_dummy_magic_29_0.V_source.t5 9.6005
R18318 two_stage_opamp_dummy_magic_29_0.V_source.n69 two_stage_opamp_dummy_magic_29_0.V_source.t0 9.6005
R18319 two_stage_opamp_dummy_magic_29_0.V_source.n72 two_stage_opamp_dummy_magic_29_0.V_source.n5 5.85227
R18320 two_stage_opamp_dummy_magic_29_0.V_source.n36 two_stage_opamp_dummy_magic_29_0.V_source.n12 5.51092
R18321 two_stage_opamp_dummy_magic_29_0.V_source.n18 two_stage_opamp_dummy_magic_29_0.V_source.n15 5.51092
R18322 two_stage_opamp_dummy_magic_29_0.V_source.n39 two_stage_opamp_dummy_magic_29_0.V_source.n36 5.45883
R18323 two_stage_opamp_dummy_magic_29_0.V_source.n15 two_stage_opamp_dummy_magic_29_0.V_source.n13 5.45883
R18324 two_stage_opamp_dummy_magic_29_0.V_source.n63 two_stage_opamp_dummy_magic_29_0.V_source.n61 5.188
R18325 two_stage_opamp_dummy_magic_29_0.V_source.n66 two_stage_opamp_dummy_magic_29_0.V_source.n6 5.188
R18326 two_stage_opamp_dummy_magic_29_0.V_source.n71 two_stage_opamp_dummy_magic_29_0.V_source.n70 5.188
R18327 two_stage_opamp_dummy_magic_29_0.V_source.n18 two_stage_opamp_dummy_magic_29_0.V_source.n17 5.16717
R18328 two_stage_opamp_dummy_magic_29_0.V_source.n21 two_stage_opamp_dummy_magic_29_0.V_source.n19 5.16717
R18329 two_stage_opamp_dummy_magic_29_0.V_source.n43 two_stage_opamp_dummy_magic_29_0.V_source.n42 5.16717
R18330 two_stage_opamp_dummy_magic_29_0.V_source.n38 two_stage_opamp_dummy_magic_29_0.V_source.n12 5.16717
R18331 two_stage_opamp_dummy_magic_29_0.V_source.n17 two_stage_opamp_dummy_magic_29_0.V_source.n13 4.89633
R18332 two_stage_opamp_dummy_magic_29_0.V_source.n22 two_stage_opamp_dummy_magic_29_0.V_source.n21 4.89633
R18333 two_stage_opamp_dummy_magic_29_0.V_source.n31 two_stage_opamp_dummy_magic_29_0.V_source.n30 4.89633
R18334 two_stage_opamp_dummy_magic_29_0.V_source.n28 two_stage_opamp_dummy_magic_29_0.V_source.n27 4.89633
R18335 two_stage_opamp_dummy_magic_29_0.V_source.n25 two_stage_opamp_dummy_magic_29_0.V_source.n23 4.89633
R18336 two_stage_opamp_dummy_magic_29_0.V_source.n34 two_stage_opamp_dummy_magic_29_0.V_source.n33 4.89633
R18337 two_stage_opamp_dummy_magic_29_0.V_source.n42 two_stage_opamp_dummy_magic_29_0.V_source.n40 4.89633
R18338 two_stage_opamp_dummy_magic_29_0.V_source.n39 two_stage_opamp_dummy_magic_29_0.V_source.n38 4.89633
R18339 two_stage_opamp_dummy_magic_29_0.V_source.n31 two_stage_opamp_dummy_magic_29_0.V_source.n28 3.6255
R18340 two_stage_opamp_dummy_magic_29_0.V_source.n48 two_stage_opamp_dummy_magic_29_0.V_source.n10 2.98664
R18341 two_stage_opamp_dummy_magic_29_0.V_source.n60 two_stage_opamp_dummy_magic_29_0.V_source.n58 2.98664
R18342 two_stage_opamp_dummy_magic_29_0.V_source.n51 two_stage_opamp_dummy_magic_29_0.V_source.n50 2.98664
R18343 two_stage_opamp_dummy_magic_29_0.V_source.n54 two_stage_opamp_dummy_magic_29_0.V_source.n53 2.98664
R18344 two_stage_opamp_dummy_magic_29_0.V_source.n9 two_stage_opamp_dummy_magic_29_0.V_source.n8 2.98664
R18345 two_stage_opamp_dummy_magic_29_0.V_source.n64 two_stage_opamp_dummy_magic_29_0.V_source.n63 2.98664
R18346 two_stage_opamp_dummy_magic_29_0.V_source.n67 two_stage_opamp_dummy_magic_29_0.V_source.n66 2.98664
R18347 two_stage_opamp_dummy_magic_29_0.V_source.n70 two_stage_opamp_dummy_magic_29_0.V_source.n68 2.98664
R18348 two_stage_opamp_dummy_magic_29_0.V_source.n55 two_stage_opamp_dummy_magic_29_0.V_source.n5 2.98664
R18349 two_stage_opamp_dummy_magic_29_0.V_source.n57 two_stage_opamp_dummy_magic_29_0.V_source.n46 2.98628
R18350 two_stage_opamp_dummy_magic_29_0.V_source.n44 two_stage_opamp_dummy_magic_29_0.V_source.n11 2.2076
R18351 two_stage_opamp_dummy_magic_29_0.V_source.n11 two_stage_opamp_dummy_magic_29_0.V_source.n0 2.16822
R18352 two_stage_opamp_dummy_magic_29_0.V_source.n2 two_stage_opamp_dummy_magic_29_0.V_source.n44 2.16822
R18353 two_stage_opamp_dummy_magic_29_0.V_source.n61 two_stage_opamp_dummy_magic_29_0.V_source.n3 2.02255
R18354 two_stage_opamp_dummy_magic_29_0.V_source.n1 two_stage_opamp_dummy_magic_29_0.V_source.n72 1.36007
R18355 two_stage_opamp_dummy_magic_29_0.V_source.n57 two_stage_opamp_dummy_magic_29_0.V_source.n56 2.96976
R18356 two_stage_opamp_dummy_magic_29_0.V_source.n56 two_stage_opamp_dummy_magic_29_0.V_source.n55 2.52416
R18357 two_stage_opamp_dummy_magic_29_0.V_source.n72 two_stage_opamp_dummy_magic_29_0.V_source.n71 0.664374
R18358 two_stage_opamp_dummy_magic_29_0.V_source.n8 two_stage_opamp_dummy_magic_29_0.V_source.n1 0.6255
R18359 two_stage_opamp_dummy_magic_29_0.V_source.n53 two_stage_opamp_dummy_magic_29_0.V_source.n1 0.6255
R18360 two_stage_opamp_dummy_magic_29_0.V_source.n50 two_stage_opamp_dummy_magic_29_0.V_source.n1 0.6255
R18361 two_stage_opamp_dummy_magic_29_0.V_source.n3 two_stage_opamp_dummy_magic_29_0.V_source.n46 0.6255
R18362 two_stage_opamp_dummy_magic_29_0.V_source.n3 two_stage_opamp_dummy_magic_29_0.V_source.n48 0.6255
R18363 two_stage_opamp_dummy_magic_29_0.V_source.n3 two_stage_opamp_dummy_magic_29_0.V_source.n60 0.6255
R18364 two_stage_opamp_dummy_magic_29_0.V_source.n30 two_stage_opamp_dummy_magic_29_0.V_source.n2 0.604667
R18365 two_stage_opamp_dummy_magic_29_0.V_source.n0 two_stage_opamp_dummy_magic_29_0.V_source.n25 0.604667
R18366 two_stage_opamp_dummy_magic_29_0.V_source.n27 two_stage_opamp_dummy_magic_29_0.V_source.n0 0.604667
R18367 two_stage_opamp_dummy_magic_29_0.V_source.n33 two_stage_opamp_dummy_magic_29_0.V_source.n2 0.604667
R18368 two_stage_opamp_dummy_magic_29_0.V_source.n40 two_stage_opamp_dummy_magic_29_0.V_source.n39 0.563
R18369 two_stage_opamp_dummy_magic_29_0.V_source.n40 two_stage_opamp_dummy_magic_29_0.V_source.n34 0.563
R18370 two_stage_opamp_dummy_magic_29_0.V_source.n34 two_stage_opamp_dummy_magic_29_0.V_source.n31 0.563
R18371 two_stage_opamp_dummy_magic_29_0.V_source.n28 two_stage_opamp_dummy_magic_29_0.V_source.n23 0.563
R18372 two_stage_opamp_dummy_magic_29_0.V_source.n23 two_stage_opamp_dummy_magic_29_0.V_source.n22 0.563
R18373 two_stage_opamp_dummy_magic_29_0.V_source.n22 two_stage_opamp_dummy_magic_29_0.V_source.n13 0.563
R18374 two_stage_opamp_dummy_magic_29_0.V_source.n19 two_stage_opamp_dummy_magic_29_0.V_source.n11 0.510302
R18375 two_stage_opamp_dummy_magic_29_0.V_source.n44 two_stage_opamp_dummy_magic_29_0.V_source.n43 0.510302
R18376 two_stage_opamp_dummy_magic_29_0.V_source.n71 two_stage_opamp_dummy_magic_29_0.V_source.n6 0.34425
R18377 two_stage_opamp_dummy_magic_29_0.V_source.n61 two_stage_opamp_dummy_magic_29_0.V_source.n6 0.34425
R18378 two_stage_opamp_dummy_magic_29_0.V_source.n19 two_stage_opamp_dummy_magic_29_0.V_source.n18 0.34425
R18379 two_stage_opamp_dummy_magic_29_0.V_source.n43 two_stage_opamp_dummy_magic_29_0.V_source.n12 0.34425
R18380 two_stage_opamp_dummy_magic_29_0.V_source.n3 two_stage_opamp_dummy_magic_29_0.V_source.n2 0.216846
R18381 two_stage_opamp_dummy_magic_29_0.V_source two_stage_opamp_dummy_magic_29_0.V_source.n0 0.120692
R18382 two_stage_opamp_dummy_magic_29_0.V_source.n55 two_stage_opamp_dummy_magic_29_0.V_source.n54 0.115083
R18383 two_stage_opamp_dummy_magic_29_0.V_source.n54 two_stage_opamp_dummy_magic_29_0.V_source.n51 0.115083
R18384 two_stage_opamp_dummy_magic_29_0.V_source.n51 two_stage_opamp_dummy_magic_29_0.V_source.n9 0.115083
R18385 two_stage_opamp_dummy_magic_29_0.V_source.n68 two_stage_opamp_dummy_magic_29_0.V_source.n9 0.115083
R18386 two_stage_opamp_dummy_magic_29_0.V_source.n68 two_stage_opamp_dummy_magic_29_0.V_source.n67 0.115083
R18387 two_stage_opamp_dummy_magic_29_0.V_source.n67 two_stage_opamp_dummy_magic_29_0.V_source.n64 0.115083
R18388 two_stage_opamp_dummy_magic_29_0.V_source.n64 two_stage_opamp_dummy_magic_29_0.V_source.n10 0.115083
R18389 two_stage_opamp_dummy_magic_29_0.V_source.n58 two_stage_opamp_dummy_magic_29_0.V_source.n10 0.115083
R18390 two_stage_opamp_dummy_magic_29_0.V_source.n58 two_stage_opamp_dummy_magic_29_0.V_source.n57 0.115083
R18391 two_stage_opamp_dummy_magic_29_0.V_source two_stage_opamp_dummy_magic_29_0.V_source.n1 0.0966538
R18392 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n27 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t29 610.534
R18393 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n6 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t27 610.534
R18394 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n27 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t18 433.8
R18395 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n28 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t15 433.8
R18396 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n29 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t24 433.8
R18397 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n30 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t12 433.8
R18398 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n31 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t21 433.8
R18399 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n32 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t31 433.8
R18400 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n33 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t20 433.8
R18401 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n34 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t30 433.8
R18402 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n35 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t13 433.8
R18403 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n12 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t28 433.8
R18404 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n11 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t17 433.8
R18405 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n10 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t26 433.8
R18406 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n9 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t16 433.8
R18407 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n8 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t25 433.8
R18408 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n7 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t14 433.8
R18409 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n6 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t23 433.8
R18410 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n26 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t22 433.8
R18411 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n25 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t19 433.8
R18412 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n2 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n14 287.264
R18413 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n19 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n18 287.264
R18414 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n16 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n15 287.264
R18415 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n22 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n21 287.264
R18416 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n35 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n34 176.733
R18417 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n34 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n33 176.733
R18418 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n33 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n32 176.733
R18419 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n32 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n31 176.733
R18420 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n31 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n30 176.733
R18421 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n30 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n29 176.733
R18422 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n29 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n28 176.733
R18423 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n28 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n27 176.733
R18424 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n7 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n6 176.733
R18425 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n8 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n7 176.733
R18426 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n9 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n8 176.733
R18427 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n10 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n9 176.733
R18428 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n11 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n10 176.733
R18429 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n12 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n11 176.733
R18430 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n26 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n25 176.733
R18431 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n37 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n36 161.986
R18432 two_stage_opamp_dummy_magic_29_0.V_tail_gate two_stage_opamp_dummy_magic_29_0.V_tail_gate.n13 161.986
R18433 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n0 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n22 63.1753
R18434 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n19 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n0 63.1745
R18435 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n3 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n2 63.1745
R18436 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n17 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n2 52.5725
R18437 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n22 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n20 52.5725
R18438 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n20 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n19 52.01
R18439 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n17 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n16 52.01
R18440 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n24 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n23 49.7255
R18441 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n5 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n4 49.7255
R18442 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n16 two_stage_opamp_dummy_magic_29_0.V_tail_gate 46.7517
R18443 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n36 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n35 45.5227
R18444 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n13 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n12 45.5227
R18445 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n25 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n13 45.5227
R18446 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n36 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n26 45.5227
R18447 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n21 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t8 39.4005
R18448 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n21 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t4 39.4005
R18449 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n18 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t10 39.4005
R18450 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n18 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t7 39.4005
R18451 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n15 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t9 39.4005
R18452 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n15 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t5 39.4005
R18453 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n14 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t6 39.4005
R18454 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n14 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t11 39.4005
R18455 two_stage_opamp_dummy_magic_29_0.V_tail_gate two_stage_opamp_dummy_magic_29_0.V_tail_gate.n3 16.4233
R18456 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n23 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t3 16.0005
R18457 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n23 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t1 16.0005
R18458 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n4 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t2 16.0005
R18459 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n4 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t0 16.0005
R18460 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n24 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n5 9.563
R18461 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n1 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n0 6.53418
R18462 two_stage_opamp_dummy_magic_29_0.V_tail_gate two_stage_opamp_dummy_magic_29_0.V_tail_gate.n1 1.56177
R18463 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n1 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n37 1.44719
R18464 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n37 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n24 0.842037
R18465 two_stage_opamp_dummy_magic_29_0.V_tail_gate two_stage_opamp_dummy_magic_29_0.V_tail_gate.n5 0.842037
R18466 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n20 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n17 0.563
R18467 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n3 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n0 0.340844
R18468 a_14420_3878.t0 a_14420_3878.t1 294.339
R18469 two_stage_opamp_dummy_magic_29_0.V_tot.n2 two_stage_opamp_dummy_magic_29_0.V_tot.t4 648.343
R18470 two_stage_opamp_dummy_magic_29_0.V_tot.n3 two_stage_opamp_dummy_magic_29_0.V_tot.t5 648.343
R18471 two_stage_opamp_dummy_magic_29_0.V_tot.n1 two_stage_opamp_dummy_magic_29_0.V_tot.t2 117.591
R18472 two_stage_opamp_dummy_magic_29_0.V_tot.n0 two_stage_opamp_dummy_magic_29_0.V_tot.t1 117.591
R18473 two_stage_opamp_dummy_magic_29_0.V_tot.n0 two_stage_opamp_dummy_magic_29_0.V_tot.t3 108.424
R18474 two_stage_opamp_dummy_magic_29_0.V_tot.n1 two_stage_opamp_dummy_magic_29_0.V_tot.t0 108.424
R18475 two_stage_opamp_dummy_magic_29_0.V_tot.n2 two_stage_opamp_dummy_magic_29_0.V_tot.n1 31.2036
R18476 two_stage_opamp_dummy_magic_29_0.V_tot two_stage_opamp_dummy_magic_29_0.V_tot.n0 29.5027
R18477 two_stage_opamp_dummy_magic_29_0.V_tot two_stage_opamp_dummy_magic_29_0.V_tot.n3 1.70362
R18478 two_stage_opamp_dummy_magic_29_0.V_tot.n3 two_stage_opamp_dummy_magic_29_0.V_tot.n2 0.84425
R18479 bgr_11_0.cap_res2.t0 bgr_11_0.cap_res2.t15 121.931
R18480 bgr_11_0.cap_res2.t10 bgr_11_0.cap_res2.t4 0.1603
R18481 bgr_11_0.cap_res2.t14 bgr_11_0.cap_res2.t9 0.1603
R18482 bgr_11_0.cap_res2.t8 bgr_11_0.cap_res2.t3 0.1603
R18483 bgr_11_0.cap_res2.t2 bgr_11_0.cap_res2.t16 0.1603
R18484 bgr_11_0.cap_res2.t6 bgr_11_0.cap_res2.t1 0.1603
R18485 bgr_11_0.cap_res2.n1 bgr_11_0.cap_res2.t11 0.159278
R18486 bgr_11_0.cap_res2.n2 bgr_11_0.cap_res2.t7 0.159278
R18487 bgr_11_0.cap_res2.n3 bgr_11_0.cap_res2.t13 0.159278
R18488 bgr_11_0.cap_res2.n4 bgr_11_0.cap_res2.t19 0.159278
R18489 bgr_11_0.cap_res2.n4 bgr_11_0.cap_res2.t20 0.1368
R18490 bgr_11_0.cap_res2.n4 bgr_11_0.cap_res2.t10 0.1368
R18491 bgr_11_0.cap_res2.n3 bgr_11_0.cap_res2.t5 0.1368
R18492 bgr_11_0.cap_res2.n3 bgr_11_0.cap_res2.t14 0.1368
R18493 bgr_11_0.cap_res2.n2 bgr_11_0.cap_res2.t18 0.1368
R18494 bgr_11_0.cap_res2.n2 bgr_11_0.cap_res2.t8 0.1368
R18495 bgr_11_0.cap_res2.n1 bgr_11_0.cap_res2.t12 0.1368
R18496 bgr_11_0.cap_res2.n1 bgr_11_0.cap_res2.t2 0.1368
R18497 bgr_11_0.cap_res2.n0 bgr_11_0.cap_res2.t17 0.1368
R18498 bgr_11_0.cap_res2.n0 bgr_11_0.cap_res2.t6 0.1368
R18499 bgr_11_0.cap_res2.t11 bgr_11_0.cap_res2.n0 0.00152174
R18500 bgr_11_0.cap_res2.t7 bgr_11_0.cap_res2.n1 0.00152174
R18501 bgr_11_0.cap_res2.t13 bgr_11_0.cap_res2.n2 0.00152174
R18502 bgr_11_0.cap_res2.t19 bgr_11_0.cap_res2.n3 0.00152174
R18503 bgr_11_0.cap_res2.t15 bgr_11_0.cap_res2.n4 0.00152174
R18504 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n141 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n140 807.99
R18505 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n33 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t8 172.969
R18506 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n142 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n141 84.0884
R18507 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n71 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n70 83.5719
R18508 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n69 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n44 83.5719
R18509 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n68 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n67 83.5719
R18510 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n59 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 83.5719
R18511 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n52 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n48 83.5719
R18512 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n54 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n53 83.5719
R18513 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n41 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n40 83.5719
R18514 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n39 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n38 83.5719
R18515 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n37 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n36 83.5719
R18516 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n89 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n88 83.5719
R18517 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n87 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n86 83.5719
R18518 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n23 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n22 83.5719
R18519 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n97 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n96 83.5719
R18520 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n18 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n16 83.5719
R18521 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n102 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n15 83.5719
R18522 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n110 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n109 83.5719
R18523 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n13 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n12 83.5719
R18524 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n125 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n124 83.5719
R18525 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n123 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n122 83.5719
R18526 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n121 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n120 83.5719
R18527 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n139 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n1 83.5719
R18528 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n138 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n0 83.5719
R18529 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n137 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n136 83.5719
R18530 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n70 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n43 73.8495
R18531 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n83 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n22 73.8495
R18532 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n61 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 73.3165
R18533 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n40 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n32 73.3165
R18534 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n96 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n95 73.3165
R18535 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n109 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n108 73.3165
R18536 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n126 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n125 73.3165
R18537 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n68 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n45 73.19
R18538 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n53 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n51 73.19
R18539 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n37 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n35 73.19
R18540 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n88 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n19 73.19
R18541 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n104 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n15 73.19
R18542 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n121 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n9 73.19
R18543 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t6 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n10 65.0299
R18544 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n134 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t7 65.0299
R18545 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n70 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n69 26.074
R18546 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n52 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 26.074
R18547 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n40 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n39 26.074
R18548 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n87 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n22 26.074
R18549 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n96 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n18 26.074
R18550 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n109 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n13 26.074
R18551 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n125 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n123 26.074
R18552 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n138 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n137 26.074
R18553 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n139 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n138 26.074
R18554 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n141 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n139 26.074
R18555 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t5 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n68 25.7843
R18556 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n53 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t1 25.7843
R18557 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t2 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n37 25.7843
R18558 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n88 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t3 25.7843
R18559 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t0 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n15 25.7843
R18560 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t4 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n121 25.7843
R18561 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n127 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n115 9.3005
R18562 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n115 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n7 9.3005
R18563 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n115 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n8 9.3005
R18564 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n131 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n115 9.3005
R18565 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n117 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n7 9.3005
R18566 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n117 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n8 9.3005
R18567 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n117 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n5 9.3005
R18568 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n131 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n117 9.3005
R18569 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n132 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n7 9.3005
R18570 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n132 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n6 9.3005
R18571 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n132 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n8 9.3005
R18572 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n132 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n5 9.3005
R18573 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n132 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n131 9.3005
R18574 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n131 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n119 9.3005
R18575 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n119 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n5 9.3005
R18576 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n119 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n8 9.3005
R18577 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n119 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n6 9.3005
R18578 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n131 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 9.3005
R18579 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n5 9.3005
R18580 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n8 9.3005
R18581 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n6 9.3005
R18582 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n127 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 9.3005
R18583 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n130 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n7 9.3005
R18584 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n130 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n6 9.3005
R18585 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n130 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n8 9.3005
R18586 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n131 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n130 9.3005
R18587 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n80 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n79 9.3005
R18588 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n79 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n78 9.3005
R18589 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n79 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n28 9.3005
R18590 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n79 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n25 9.3005
R18591 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n79 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n26 9.3005
R18592 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n78 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n76 9.3005
R18593 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n76 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n28 9.3005
R18594 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n76 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n25 9.3005
R18595 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n76 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n26 9.3005
R18596 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n78 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n75 9.3005
R18597 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n75 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n28 9.3005
R18598 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n75 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n25 9.3005
R18599 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n75 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n27 9.3005
R18600 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n75 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n26 9.3005
R18601 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n29 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n26 9.3005
R18602 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n29 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n27 9.3005
R18603 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n29 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n25 9.3005
R18604 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n29 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n28 9.3005
R18605 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n81 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n26 9.3005
R18606 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n81 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n27 9.3005
R18607 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n81 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n25 9.3005
R18608 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n81 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n28 9.3005
R18609 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n81 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n80 9.3005
R18610 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n78 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n77 9.3005
R18611 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n77 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n28 9.3005
R18612 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n77 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n25 9.3005
R18613 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n77 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n27 9.3005
R18614 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n77 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n26 9.3005
R18615 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n129 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n5 4.64654
R18616 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n116 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n6 4.64654
R18617 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n127 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n4 4.64654
R18618 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n118 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n7 4.64654
R18619 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n128 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n127 4.64654
R18620 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n34 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n27 4.64654
R18621 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n80 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n31 4.64654
R18622 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n78 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n24 4.64654
R18623 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n80 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n30 4.64654
R18624 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n63 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n45 2.36206
R18625 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n51 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n3 2.36206
R18626 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n92 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n19 2.36206
R18627 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n105 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n104 2.36206
R18628 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n62 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n61 2.19742
R18629 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n95 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n93 2.19742
R18630 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n108 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n106 2.19742
R18631 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n12 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n10 1.56363
R18632 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n136 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n134 1.56363
R18633 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n107 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n11 1.5505
R18634 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n112 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n111 1.5505
R18635 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n94 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 1.5505
R18636 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n99 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n98 1.5505
R18637 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n101 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n100 1.5505
R18638 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n103 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n14 1.5505
R18639 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n85 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n84 1.5505
R18640 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n91 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n90 1.5505
R18641 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n21 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n20 1.5505
R18642 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n60 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n46 1.5505
R18643 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n58 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n57 1.5505
R18644 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n56 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n55 1.5505
R18645 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n50 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n49 1.5505
R18646 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n73 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n72 1.5505
R18647 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n66 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n42 1.5505
R18648 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n65 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n64 1.5505
R18649 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n143 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n142 1.5505
R18650 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n145 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n144 1.5505
R18651 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n135 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n2 1.5505
R18652 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n67 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n65 1.25468
R18653 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n54 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n50 1.25468
R18654 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n36 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n27 1.25468
R18655 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n90 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n89 1.25468
R18656 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n103 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n102 1.25468
R18657 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n120 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n5 1.25468
R18658 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n61 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n60 1.19225
R18659 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n78 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n32 1.19225
R18660 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n95 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n94 1.19225
R18661 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n108 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n107 1.19225
R18662 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n126 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n7 1.19225
R18663 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n142 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n1 1.14402
R18664 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n66 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n44 1.07024
R18665 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n55 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n48 1.07024
R18666 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n38 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n25 1.07024
R18667 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n86 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n21 1.07024
R18668 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n101 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n16 1.07024
R18669 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n122 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n8 1.07024
R18670 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n65 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n45 1.0237
R18671 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n51 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n50 1.0237
R18672 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n35 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n27 1.0237
R18673 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n90 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n19 1.0237
R18674 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n104 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n103 1.0237
R18675 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n9 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n5 1.0237
R18676 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n72 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n71 0.885803
R18677 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n59 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n58 0.885803
R18678 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n41 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n28 0.885803
R18679 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n85 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n23 0.885803
R18680 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n98 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n97 0.885803
R18681 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n111 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n110 0.885803
R18682 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n124 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n6 0.885803
R18683 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n135 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n0 0.885803
R18684 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n35 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n26 0.812055
R18685 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n131 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n9 0.812055
R18686 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n72 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n44 0.77514
R18687 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n58 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n48 0.77514
R18688 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n38 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n28 0.77514
R18689 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n86 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n85 0.77514
R18690 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n98 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n16 0.77514
R18691 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n111 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n12 0.77514
R18692 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n122 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n6 0.77514
R18693 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n136 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n135 0.77514
R18694 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n71 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.756696
R18695 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n59 0.756696
R18696 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n41 0.756696
R18697 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n23 0.756696
R18698 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n97 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.756696
R18699 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n110 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.756696
R18700 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n124 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.756696
R18701 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n0 0.756696
R18702 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n84 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n83 0.711459
R18703 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n73 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n43 0.711459
R18704 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n145 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n1 0.701365
R18705 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n80 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n32 0.647417
R18706 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n127 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n126 0.647417
R18707 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n67 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n66 0.590702
R18708 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n55 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n54 0.590702
R18709 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n36 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n25 0.590702
R18710 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n89 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n21 0.590702
R18711 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n102 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n101 0.590702
R18712 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n120 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n8 0.590702
R18713 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n43 0.576566
R18714 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n83 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.576566
R18715 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n113 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n10 0.530034
R18716 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n134 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n133 0.530034
R18717 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n69 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t5 0.290206
R18718 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t1 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n52 0.290206
R18719 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n39 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t2 0.290206
R18720 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t3 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n87 0.290206
R18721 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n18 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t0 0.290206
R18722 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n13 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t6 0.290206
R18723 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n123 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t4 0.290206
R18724 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n137 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t7 0.290206
R18725 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n60 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.203382
R18726 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n78 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.203382
R18727 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n94 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.203382
R18728 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n107 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.203382
R18729 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n7 0.203382
R18730 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n145 0.203382
R18731 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n106 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n105 0.154071
R18732 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n93 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n92 0.154071
R18733 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n143 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n3 0.154071
R18734 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n63 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n62 0.154071
R18735 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n133 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n132 0.137464
R18736 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n75 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n74 0.137464
R18737 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n113 0.134964
R18738 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n82 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n81 0.134964
R18739 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n112 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n11 0.0183571
R18740 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n106 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n11 0.0183571
R18741 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n105 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n14 0.0183571
R18742 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n100 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n14 0.0183571
R18743 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n100 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n99 0.0183571
R18744 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n99 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 0.0183571
R18745 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n93 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 0.0183571
R18746 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n92 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n91 0.0183571
R18747 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n91 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n20 0.0183571
R18748 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n144 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n2 0.0183571
R18749 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n144 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n143 0.0183571
R18750 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n49 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n3 0.0183571
R18751 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n56 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n49 0.0183571
R18752 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n57 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n56 0.0183571
R18753 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n57 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n46 0.0183571
R18754 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n62 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n46 0.0183571
R18755 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n64 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n63 0.0183571
R18756 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n64 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n42 0.0183571
R18757 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n82 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n20 0.0106786
R18758 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n77 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n33 0.0106786
R18759 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n74 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n42 0.0106786
R18760 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n119 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n118 0.00992001
R18761 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n130 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n128 0.00992001
R18762 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n129 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n115 0.00992001
R18763 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n117 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n116 0.00992001
R18764 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n132 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n4 0.00992001
R18765 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n116 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n115 0.00992001
R18766 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n117 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n4 0.00992001
R18767 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n128 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n119 0.00992001
R18768 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n118 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 0.00992001
R18769 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n130 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n129 0.00992001
R18770 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n29 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n24 0.00992001
R18771 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n77 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n30 0.00992001
R18772 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n76 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n34 0.00992001
R18773 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n75 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n31 0.00992001
R18774 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n79 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n34 0.00992001
R18775 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n76 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n31 0.00992001
R18776 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n30 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n29 0.00992001
R18777 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n81 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n24 0.00992001
R18778 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n113 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n112 0.00817857
R18779 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n84 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n82 0.00817857
R18780 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n79 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n33 0.00817857
R18781 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n133 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n2 0.00817857
R18782 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n74 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n73 0.00817857
R18783 a_3230_3878.t0 a_3230_3878.t1 169.905
R18784 two_stage_opamp_dummy_magic_29_0.err_amp_mir.n1 two_stage_opamp_dummy_magic_29_0.err_amp_mir.t5 573.044
R18785 two_stage_opamp_dummy_magic_29_0.err_amp_mir.n1 two_stage_opamp_dummy_magic_29_0.err_amp_mir.t2 433.8
R18786 two_stage_opamp_dummy_magic_29_0.err_amp_mir.n2 two_stage_opamp_dummy_magic_29_0.err_amp_mir.n0 184.09
R18787 two_stage_opamp_dummy_magic_29_0.err_amp_mir.n2 two_stage_opamp_dummy_magic_29_0.err_amp_mir.n1 163.978
R18788 two_stage_opamp_dummy_magic_29_0.err_amp_mir.n3 two_stage_opamp_dummy_magic_29_0.err_amp_mir.n2 33.0088
R18789 two_stage_opamp_dummy_magic_29_0.err_amp_mir.n0 two_stage_opamp_dummy_magic_29_0.err_amp_mir.t4 15.7605
R18790 two_stage_opamp_dummy_magic_29_0.err_amp_mir.n0 two_stage_opamp_dummy_magic_29_0.err_amp_mir.t1 15.7605
R18791 two_stage_opamp_dummy_magic_29_0.err_amp_mir.n3 two_stage_opamp_dummy_magic_29_0.err_amp_mir.t3 9.6005
R18792 two_stage_opamp_dummy_magic_29_0.err_amp_mir.t0 two_stage_opamp_dummy_magic_29_0.err_amp_mir.n3 9.6005
R18793 two_stage_opamp_dummy_magic_29_0.err_amp_out.n0 two_stage_opamp_dummy_magic_29_0.err_amp_out.t4 610.534
R18794 two_stage_opamp_dummy_magic_29_0.err_amp_out.n0 two_stage_opamp_dummy_magic_29_0.err_amp_out.t5 433.8
R18795 two_stage_opamp_dummy_magic_29_0.err_amp_out two_stage_opamp_dummy_magic_29_0.err_amp_out.n0 267.139
R18796 two_stage_opamp_dummy_magic_29_0.err_amp_out.n3 two_stage_opamp_dummy_magic_29_0.err_amp_out.n2 178.829
R18797 two_stage_opamp_dummy_magic_29_0.err_amp_out.n3 two_stage_opamp_dummy_magic_29_0.err_amp_out.n1 38.5609
R18798 two_stage_opamp_dummy_magic_29_0.err_amp_out.n2 two_stage_opamp_dummy_magic_29_0.err_amp_out.t2 15.7605
R18799 two_stage_opamp_dummy_magic_29_0.err_amp_out.n2 two_stage_opamp_dummy_magic_29_0.err_amp_out.t0 15.7605
R18800 two_stage_opamp_dummy_magic_29_0.err_amp_out.n1 two_stage_opamp_dummy_magic_29_0.err_amp_out.t1 9.6005
R18801 two_stage_opamp_dummy_magic_29_0.err_amp_out.n1 two_stage_opamp_dummy_magic_29_0.err_amp_out.t3 9.6005
R18802 two_stage_opamp_dummy_magic_29_0.err_amp_out two_stage_opamp_dummy_magic_29_0.err_amp_out.n3 0.922375
R18803 two_stage_opamp_dummy_magic_29_0.VD1.n1 two_stage_opamp_dummy_magic_29_0.VD1.n0 49.7255
R18804 two_stage_opamp_dummy_magic_29_0.VD1.n25 two_stage_opamp_dummy_magic_29_0.VD1.n24 49.7255
R18805 two_stage_opamp_dummy_magic_29_0.VD1.n27 two_stage_opamp_dummy_magic_29_0.VD1.n9 49.7255
R18806 two_stage_opamp_dummy_magic_29_0.VD1.n21 two_stage_opamp_dummy_magic_29_0.VD1.n12 49.7255
R18807 two_stage_opamp_dummy_magic_29_0.VD1.n11 two_stage_opamp_dummy_magic_29_0.VD1.n10 49.7255
R18808 two_stage_opamp_dummy_magic_29_0.VD1.n15 two_stage_opamp_dummy_magic_29_0.VD1.n14 49.3505
R18809 two_stage_opamp_dummy_magic_29_0.VD1.n8 two_stage_opamp_dummy_magic_29_0.VD1.n7 49.3505
R18810 two_stage_opamp_dummy_magic_29_0.VD1.n31 two_stage_opamp_dummy_magic_29_0.VD1.n30 49.3505
R18811 two_stage_opamp_dummy_magic_29_0.VD1.n35 two_stage_opamp_dummy_magic_29_0.VD1.n34 49.3505
R18812 two_stage_opamp_dummy_magic_29_0.VD1.n5 two_stage_opamp_dummy_magic_29_0.VD1.n4 49.3505
R18813 two_stage_opamp_dummy_magic_29_0.VD1.n18 two_stage_opamp_dummy_magic_29_0.VD1.n17 49.3505
R18814 two_stage_opamp_dummy_magic_29_0.VD1.n14 two_stage_opamp_dummy_magic_29_0.VD1.t6 16.0005
R18815 two_stage_opamp_dummy_magic_29_0.VD1.n14 two_stage_opamp_dummy_magic_29_0.VD1.t8 16.0005
R18816 two_stage_opamp_dummy_magic_29_0.VD1.n7 two_stage_opamp_dummy_magic_29_0.VD1.t3 16.0005
R18817 two_stage_opamp_dummy_magic_29_0.VD1.n7 two_stage_opamp_dummy_magic_29_0.VD1.t5 16.0005
R18818 two_stage_opamp_dummy_magic_29_0.VD1.n30 two_stage_opamp_dummy_magic_29_0.VD1.t2 16.0005
R18819 two_stage_opamp_dummy_magic_29_0.VD1.n30 two_stage_opamp_dummy_magic_29_0.VD1.t21 16.0005
R18820 two_stage_opamp_dummy_magic_29_0.VD1.n34 two_stage_opamp_dummy_magic_29_0.VD1.t9 16.0005
R18821 two_stage_opamp_dummy_magic_29_0.VD1.n34 two_stage_opamp_dummy_magic_29_0.VD1.t1 16.0005
R18822 two_stage_opamp_dummy_magic_29_0.VD1.n4 two_stage_opamp_dummy_magic_29_0.VD1.t7 16.0005
R18823 two_stage_opamp_dummy_magic_29_0.VD1.n4 two_stage_opamp_dummy_magic_29_0.VD1.t4 16.0005
R18824 two_stage_opamp_dummy_magic_29_0.VD1.n0 two_stage_opamp_dummy_magic_29_0.VD1.t11 16.0005
R18825 two_stage_opamp_dummy_magic_29_0.VD1.n0 two_stage_opamp_dummy_magic_29_0.VD1.t18 16.0005
R18826 two_stage_opamp_dummy_magic_29_0.VD1.n24 two_stage_opamp_dummy_magic_29_0.VD1.t12 16.0005
R18827 two_stage_opamp_dummy_magic_29_0.VD1.n24 two_stage_opamp_dummy_magic_29_0.VD1.t16 16.0005
R18828 two_stage_opamp_dummy_magic_29_0.VD1.n9 two_stage_opamp_dummy_magic_29_0.VD1.t10 16.0005
R18829 two_stage_opamp_dummy_magic_29_0.VD1.n9 two_stage_opamp_dummy_magic_29_0.VD1.t15 16.0005
R18830 two_stage_opamp_dummy_magic_29_0.VD1.n12 two_stage_opamp_dummy_magic_29_0.VD1.t13 16.0005
R18831 two_stage_opamp_dummy_magic_29_0.VD1.n12 two_stage_opamp_dummy_magic_29_0.VD1.t17 16.0005
R18832 two_stage_opamp_dummy_magic_29_0.VD1.n17 two_stage_opamp_dummy_magic_29_0.VD1.t20 16.0005
R18833 two_stage_opamp_dummy_magic_29_0.VD1.n17 two_stage_opamp_dummy_magic_29_0.VD1.t0 16.0005
R18834 two_stage_opamp_dummy_magic_29_0.VD1.n10 two_stage_opamp_dummy_magic_29_0.VD1.t14 16.0005
R18835 two_stage_opamp_dummy_magic_29_0.VD1.n10 two_stage_opamp_dummy_magic_29_0.VD1.t19 16.0005
R18836 two_stage_opamp_dummy_magic_29_0.VD1.n25 two_stage_opamp_dummy_magic_29_0.VD1.n3 8.89633
R18837 two_stage_opamp_dummy_magic_29_0.VD1.n28 two_stage_opamp_dummy_magic_29_0.VD1.n27 8.89633
R18838 two_stage_opamp_dummy_magic_29_0.VD1.n21 two_stage_opamp_dummy_magic_29_0.VD1.n20 8.89633
R18839 two_stage_opamp_dummy_magic_29_0.VD1.n13 two_stage_opamp_dummy_magic_29_0.VD1.n11 8.89633
R18840 two_stage_opamp_dummy_magic_29_0.VD1.n32 two_stage_opamp_dummy_magic_29_0.VD1.n8 5.438
R18841 two_stage_opamp_dummy_magic_29_0.VD1.n16 two_stage_opamp_dummy_magic_29_0.VD1.n15 5.438
R18842 two_stage_opamp_dummy_magic_29_0.VD1.n28 two_stage_opamp_dummy_magic_29_0.VD1.n8 5.31821
R18843 two_stage_opamp_dummy_magic_29_0.VD1.n15 two_stage_opamp_dummy_magic_29_0.VD1.n13 5.31821
R18844 two_stage_opamp_dummy_magic_29_0.VD1.n31 two_stage_opamp_dummy_magic_29_0.VD1.n29 5.08383
R18845 two_stage_opamp_dummy_magic_29_0.VD1.n36 two_stage_opamp_dummy_magic_29_0.VD1.n35 5.08383
R18846 two_stage_opamp_dummy_magic_29_0.VD1.n5 two_stage_opamp_dummy_magic_29_0.VD1.n2 5.08383
R18847 two_stage_opamp_dummy_magic_29_0.VD1.n19 two_stage_opamp_dummy_magic_29_0.VD1.n18 5.08383
R18848 two_stage_opamp_dummy_magic_29_0.VD1.n27 two_stage_opamp_dummy_magic_29_0.VD1.n26 5.063
R18849 two_stage_opamp_dummy_magic_29_0.VD1.n22 two_stage_opamp_dummy_magic_29_0.VD1.n11 5.063
R18850 two_stage_opamp_dummy_magic_29_0.VD1.n32 two_stage_opamp_dummy_magic_29_0.VD1.n31 4.8755
R18851 two_stage_opamp_dummy_magic_29_0.VD1.n35 two_stage_opamp_dummy_magic_29_0.VD1.n33 4.8755
R18852 two_stage_opamp_dummy_magic_29_0.VD1.n6 two_stage_opamp_dummy_magic_29_0.VD1.n5 4.8755
R18853 two_stage_opamp_dummy_magic_29_0.VD1.n18 two_stage_opamp_dummy_magic_29_0.VD1.n16 4.8755
R18854 two_stage_opamp_dummy_magic_29_0.VD1 two_stage_opamp_dummy_magic_29_0.VD1.n37 4.60467
R18855 two_stage_opamp_dummy_magic_29_0.VD1.n26 two_stage_opamp_dummy_magic_29_0.VD1.n25 4.5005
R18856 two_stage_opamp_dummy_magic_29_0.VD1.n23 two_stage_opamp_dummy_magic_29_0.VD1.n1 4.5005
R18857 two_stage_opamp_dummy_magic_29_0.VD1.n22 two_stage_opamp_dummy_magic_29_0.VD1.n21 4.5005
R18858 two_stage_opamp_dummy_magic_29_0.VD1 two_stage_opamp_dummy_magic_29_0.VD1.n1 4.29217
R18859 two_stage_opamp_dummy_magic_29_0.VD1.n26 two_stage_opamp_dummy_magic_29_0.VD1.n23 0.563
R18860 two_stage_opamp_dummy_magic_29_0.VD1.n23 two_stage_opamp_dummy_magic_29_0.VD1.n22 0.563
R18861 two_stage_opamp_dummy_magic_29_0.VD1.n33 two_stage_opamp_dummy_magic_29_0.VD1.n32 0.563
R18862 two_stage_opamp_dummy_magic_29_0.VD1.n33 two_stage_opamp_dummy_magic_29_0.VD1.n6 0.563
R18863 two_stage_opamp_dummy_magic_29_0.VD1.n16 two_stage_opamp_dummy_magic_29_0.VD1.n6 0.563
R18864 two_stage_opamp_dummy_magic_29_0.VD1.n19 two_stage_opamp_dummy_magic_29_0.VD1.n13 0.234875
R18865 two_stage_opamp_dummy_magic_29_0.VD1.n20 two_stage_opamp_dummy_magic_29_0.VD1.n19 0.234875
R18866 two_stage_opamp_dummy_magic_29_0.VD1.n20 two_stage_opamp_dummy_magic_29_0.VD1.n2 0.234875
R18867 two_stage_opamp_dummy_magic_29_0.VD1.n37 two_stage_opamp_dummy_magic_29_0.VD1.n2 0.234875
R18868 two_stage_opamp_dummy_magic_29_0.VD1.n37 two_stage_opamp_dummy_magic_29_0.VD1.n36 0.234875
R18869 two_stage_opamp_dummy_magic_29_0.VD1.n36 two_stage_opamp_dummy_magic_29_0.VD1.n3 0.234875
R18870 two_stage_opamp_dummy_magic_29_0.VD1.n29 two_stage_opamp_dummy_magic_29_0.VD1.n3 0.234875
R18871 two_stage_opamp_dummy_magic_29_0.VD1.n29 two_stage_opamp_dummy_magic_29_0.VD1.n28 0.234875
R18872 bgr_11_0.START_UP.n4 bgr_11_0.START_UP.t7 238.322
R18873 bgr_11_0.START_UP.n4 bgr_11_0.START_UP.t6 238.322
R18874 bgr_11_0.START_UP.n5 bgr_11_0.START_UP.n4 167.332
R18875 bgr_11_0.START_UP.n0 bgr_11_0.START_UP.t5 130.001
R18876 bgr_11_0.START_UP.n3 bgr_11_0.START_UP.n1 111.796
R18877 bgr_11_0.START_UP.n3 bgr_11_0.START_UP.n2 105.171
R18878 bgr_11_0.START_UP.n0 bgr_11_0.START_UP.t4 81.7074
R18879 bgr_11_0.START_UP bgr_11_0.START_UP.n0 36.8552
R18880 bgr_11_0.START_UP bgr_11_0.START_UP.n5 15.3755
R18881 bgr_11_0.START_UP.n1 bgr_11_0.START_UP.t0 13.1338
R18882 bgr_11_0.START_UP.n1 bgr_11_0.START_UP.t2 13.1338
R18883 bgr_11_0.START_UP.n2 bgr_11_0.START_UP.t1 13.1338
R18884 bgr_11_0.START_UP.n2 bgr_11_0.START_UP.t3 13.1338
R18885 bgr_11_0.START_UP.n5 bgr_11_0.START_UP.n3 4.21925
R18886 a_11420_30238.t0 a_11420_30238.t1 178.133
R18887 bgr_11_0.Vin-.n8 bgr_11_0.Vin-.t8 539.797
R18888 bgr_11_0.Vin-.n7 bgr_11_0.Vin-.n6 351.865
R18889 bgr_11_0.Vin-.n18 bgr_11_0.Vin-.n17 141.667
R18890 bgr_11_0.Vin-.n9 bgr_11_0.Vin-.t5 117.817
R18891 bgr_11_0.Vin-.n5 bgr_11_0.Vin-.n3 109.204
R18892 bgr_11_0.Vin-.n5 bgr_11_0.Vin-.n4 104.829
R18893 bgr_11_0.Vin-.n19 bgr_11_0.Vin-.n18 84.0884
R18894 bgr_11_0.Vin-.n14 bgr_11_0.Vin-.n13 83.5719
R18895 bgr_11_0.Vin-.n15 bgr_11_0.Vin-.n0 83.5719
R18896 bgr_11_0.Vin-.n16 bgr_11_0.Vin-.n1 83.5719
R18897 bgr_11_0.Vin-.n11 bgr_11_0.Vin-.t4 65.0299
R18898 bgr_11_0.Vin-.n6 bgr_11_0.Vin-.t7 39.4005
R18899 bgr_11_0.Vin-.n6 bgr_11_0.Vin-.t6 39.4005
R18900 bgr_11_0.Vin-.n15 bgr_11_0.Vin-.n14 26.074
R18901 bgr_11_0.Vin-.n16 bgr_11_0.Vin-.n15 26.074
R18902 bgr_11_0.Vin-.n18 bgr_11_0.Vin-.n16 26.074
R18903 bgr_11_0.Vin-.n10 bgr_11_0.Vin-.n9 24.3755
R18904 bgr_11_0.Vin-.n9 bgr_11_0.Vin-.n8 17.6255
R18905 bgr_11_0.Vin-.n4 bgr_11_0.Vin-.t1 13.1338
R18906 bgr_11_0.Vin-.n4 bgr_11_0.Vin-.t2 13.1338
R18907 bgr_11_0.Vin-.n3 bgr_11_0.Vin-.t3 13.1338
R18908 bgr_11_0.Vin-.n3 bgr_11_0.Vin-.t0 13.1338
R18909 bgr_11_0.Vin-.n8 bgr_11_0.Vin-.n7 11.6567
R18910 bgr_11_0.Vin-.n7 bgr_11_0.Vin-.n5 3.8755
R18911 bgr_11_0.Vin-.n20 bgr_11_0.Vin-.n19 1.56836
R18912 bgr_11_0.Vin-.n13 bgr_11_0.Vin-.n11 1.56363
R18913 bgr_11_0.Vin-.n21 bgr_11_0.Vin-.n20 1.5505
R18914 bgr_11_0.Vin-.n12 bgr_11_0.Vin-.n2 1.5505
R18915 bgr_11_0.Vin-.n19 bgr_11_0.Vin-.n1 1.14402
R18916 bgr_11_0.Vin-.n12 bgr_11_0.Vin-.n0 0.885803
R18917 bgr_11_0.Vin-.n13 bgr_11_0.Vin-.n12 0.77514
R18918 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_23.Emitter bgr_11_0.Vin-.n0 0.756696
R18919 bgr_11_0.Vin-.n21 bgr_11_0.Vin-.n1 0.701365
R18920 bgr_11_0.Vin-.n11 bgr_11_0.Vin-.n10 0.530034
R18921 bgr_11_0.Vin-.n14 bgr_11_0.Vin-.t4 0.290206
R18922 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_23.Emitter bgr_11_0.Vin-.n21 0.203382
R18923 bgr_11_0.Vin-.n20 bgr_11_0.Vin-.n2 0.0183571
R18924 bgr_11_0.Vin-.n10 bgr_11_0.Vin-.n2 0.00817857
R18925 a_11950_28880.t0 a_11950_28880.t1 178.133
R18926 two_stage_opamp_dummy_magic_29_0.V_err_p.n1 two_stage_opamp_dummy_magic_29_0.V_err_p.n0 363.962
R18927 two_stage_opamp_dummy_magic_29_0.V_err_p.n0 two_stage_opamp_dummy_magic_29_0.V_err_p.t3 15.7605
R18928 two_stage_opamp_dummy_magic_29_0.V_err_p.n0 two_stage_opamp_dummy_magic_29_0.V_err_p.t1 15.7605
R18929 two_stage_opamp_dummy_magic_29_0.V_err_p.n1 two_stage_opamp_dummy_magic_29_0.V_err_p.t0 15.7605
R18930 two_stage_opamp_dummy_magic_29_0.V_err_p.t2 two_stage_opamp_dummy_magic_29_0.V_err_p.n1 15.7605
R18931 VIN-.n0 VIN-.t7 1097.62
R18932 VIN- VIN-.n9 433.019
R18933 VIN-.n9 VIN-.t10 273.134
R18934 VIN-.n0 VIN-.t9 273.134
R18935 VIN-.n1 VIN-.t3 273.134
R18936 VIN-.n2 VIN-.t8 273.134
R18937 VIN-.n3 VIN-.t1 273.134
R18938 VIN-.n4 VIN-.t5 273.134
R18939 VIN-.n5 VIN-.t2 273.134
R18940 VIN-.n6 VIN-.t6 273.134
R18941 VIN-.n7 VIN-.t0 273.134
R18942 VIN-.n8 VIN-.t4 273.134
R18943 VIN-.n9 VIN-.n8 176.733
R18944 VIN-.n8 VIN-.n7 176.733
R18945 VIN-.n7 VIN-.n6 176.733
R18946 VIN-.n6 VIN-.n5 176.733
R18947 VIN-.n5 VIN-.n4 176.733
R18948 VIN-.n4 VIN-.n3 176.733
R18949 VIN-.n3 VIN-.n2 176.733
R18950 VIN-.n2 VIN-.n1 176.733
R18951 VIN-.n1 VIN-.n0 176.733
R18952 VDDA_2.n174 VDDA_2.n80 2100
R18953 VDDA_2.n172 VDDA_2.n80 2070
R18954 VDDA_2.n174 VDDA_2.n81 1830
R18955 VDDA_2.n172 VDDA_2.n81 1800
R18956 VDDA_2.n183 VDDA_2.t3 605.143
R18957 VDDA_2.n163 VDDA_2.t0 589.076
R18958 VDDA_2.n168 VDDA_2.t2 461.389
R18959 VDDA_2.t2 VDDA_2.n167 461.389
R18960 VDDA_2.t6 VDDA_2.n180 461.389
R18961 VDDA_2.n181 VDDA_2.t6 461.389
R18962 VDDA_2.t1 VDDA_2.n172 279.298
R18963 VDDA_2.n174 VDDA_2.t4 279.298
R18964 VDDA_2.n175 VDDA_2.n79 195.201
R18965 VDDA_2.n171 VDDA_2.n79 192
R18966 VDDA_2.n176 VDDA_2.n175 163.201
R18967 VDDA_2.n171 VDDA_2.n170 163.201
R18968 VDDA_2.n74 VDDA_2.n73 149.112
R18969 VDDA_2.t4 VDDA_2.t7 117.416
R18970 VDDA_2.n173 VDDA_2.t1 112.079
R18971 VDDA_2.n80 VDDA_2.n78 92.5005
R18972 VDDA_2.n173 VDDA_2.n80 92.5005
R18973 VDDA_2.n175 VDDA_2.n174 92.5005
R18974 VDDA_2.n81 VDDA_2.n79 92.5005
R18975 VDDA_2.n173 VDDA_2.n81 92.5005
R18976 VDDA_2.n172 VDDA_2.n171 92.5005
R18977 VDDA_2.n176 VDDA_2.n78 48.0005
R18978 VDDA_2.n170 VDDA_2.n78 44.8005
R18979 VDDA_2.n169 VDDA_2.n168 21.6365
R18980 VDDA_2.n167 VDDA_2.n164 21.6365
R18981 VDDA_2.n180 VDDA_2.n177 21.6365
R18982 VDDA_2.n182 VDDA_2.n181 21.6365
R18983 VDDA_2.n166 VDDA_2.n83 21.3338
R18984 VDDA_2.n179 VDDA_2.n77 21.3338
R18985 VDDA_2.n73 VDDA_2.t8 19.7005
R18986 VDDA_2.n73 VDDA_2.t5 19.7005
R18987 VDDA_2.n177 VDDA_2.n176 9.8005
R18988 VDDA_2.n170 VDDA_2.n169 9.8005
R18989 VDDA_2.n77 VDDA_2.n76 9.3005
R18990 VDDA_2.n179 VDDA_2.n178 9.3005
R18991 VDDA_2.n166 VDDA_2.n165 9.3005
R18992 VDDA_2.n83 VDDA_2.n82 9.3005
R18993 VDDA_2.n168 VDDA_2.n83 8.68224
R18994 VDDA_2.n167 VDDA_2.n166 8.68224
R18995 VDDA_2.n180 VDDA_2.n179 8.68224
R18996 VDDA_2.n181 VDDA_2.n77 8.68224
R18997 VDDA_2.n162 VDDA_2.n161 7.61355
R18998 VDDA_2.n185 VDDA_2.n74 7.51355
R18999 VDDA_2.n185 VDDA_2.n184 7.51355
R19000 VDDA_2.t7 VDDA_2.n173 5.33758
R19001 VDDA_2.n161 VDDA_2.n160 4.5005
R19002 VDDA_2.n85 VDDA_2.n84 4.5005
R19003 VDDA_2.n107 VDDA_2.n87 4.5005
R19004 VDDA_2.n108 VDDA_2.n88 4.5005
R19005 VDDA_2.n109 VDDA_2.n89 4.5005
R19006 VDDA_2.n110 VDDA_2.n90 4.5005
R19007 VDDA_2.n111 VDDA_2.n91 4.5005
R19008 VDDA_2.n112 VDDA_2.n92 4.5005
R19009 VDDA_2.n113 VDDA_2.n93 4.5005
R19010 VDDA_2.n114 VDDA_2.n94 4.5005
R19011 VDDA_2.n115 VDDA_2.n95 4.5005
R19012 VDDA_2.n116 VDDA_2.n96 4.5005
R19013 VDDA_2.n117 VDDA_2.n97 4.5005
R19014 VDDA_2.n118 VDDA_2.n98 4.5005
R19015 VDDA_2.n119 VDDA_2.n99 4.5005
R19016 VDDA_2.n120 VDDA_2.n100 4.5005
R19017 VDDA_2.n121 VDDA_2.n101 4.5005
R19018 VDDA_2.n122 VDDA_2.n102 4.5005
R19019 VDDA_2.n123 VDDA_2.n103 4.5005
R19020 VDDA_2.n124 VDDA_2.n104 4.5005
R19021 VDDA_2.n125 VDDA_2.n105 4.5005
R19022 VDDA_2.n127 VDDA_2.n126 3.49225
R19023 VDDA_2.n160 VDDA_2.n159 3.44359
R19024 VDDA_2.n128 VDDA_2.n106 3.4105
R19025 VDDA_2.n130 VDDA_2.n105 3.4105
R19026 VDDA_2.n131 VDDA_2.n104 3.4105
R19027 VDDA_2.n133 VDDA_2.n103 3.4105
R19028 VDDA_2.n134 VDDA_2.n102 3.4105
R19029 VDDA_2.n136 VDDA_2.n101 3.4105
R19030 VDDA_2.n137 VDDA_2.n100 3.4105
R19031 VDDA_2.n139 VDDA_2.n99 3.4105
R19032 VDDA_2.n140 VDDA_2.n98 3.4105
R19033 VDDA_2.n142 VDDA_2.n97 3.4105
R19034 VDDA_2.n143 VDDA_2.n96 3.4105
R19035 VDDA_2.n145 VDDA_2.n95 3.4105
R19036 VDDA_2.n146 VDDA_2.n94 3.4105
R19037 VDDA_2.n148 VDDA_2.n93 3.4105
R19038 VDDA_2.n149 VDDA_2.n92 3.4105
R19039 VDDA_2.n151 VDDA_2.n91 3.4105
R19040 VDDA_2.n152 VDDA_2.n90 3.4105
R19041 VDDA_2.n154 VDDA_2.n89 3.4105
R19042 VDDA_2.n155 VDDA_2.n88 3.4105
R19043 VDDA_2.n157 VDDA_2.n87 3.4105
R19044 VDDA_2.n158 VDDA_2.n85 3.4105
R19045 VDDA_2.n127 VDDA_2.n86 3.4105
R19046 VDDA_2.n186 VDDA_2.n33 3.4105
R19047 VDDA_2.n236 VDDA_2.n235 3.4105
R19048 VDDA_2.n333 VDDA_2.n268 3.4105
R19049 VDDA_2.n317 VDDA_2.n268 3.4105
R19050 VDDA_2.n268 VDDA_2.n32 3.4105
R19051 VDDA_2.n336 VDDA_2.n268 3.4105
R19052 VDDA_2.n336 VDDA_2.n286 3.4105
R19053 VDDA_2.n317 VDDA_2.n252 3.4105
R19054 VDDA_2.n252 VDDA_2.n17 3.4105
R19055 VDDA_2.n252 VDDA_2.n15 3.4105
R19056 VDDA_2.n252 VDDA_2.n18 3.4105
R19057 VDDA_2.n252 VDDA_2.n14 3.4105
R19058 VDDA_2.n252 VDDA_2.n19 3.4105
R19059 VDDA_2.n252 VDDA_2.n13 3.4105
R19060 VDDA_2.n252 VDDA_2.n20 3.4105
R19061 VDDA_2.n252 VDDA_2.n12 3.4105
R19062 VDDA_2.n252 VDDA_2.n21 3.4105
R19063 VDDA_2.n252 VDDA_2.n11 3.4105
R19064 VDDA_2.n252 VDDA_2.n22 3.4105
R19065 VDDA_2.n252 VDDA_2.n10 3.4105
R19066 VDDA_2.n252 VDDA_2.n23 3.4105
R19067 VDDA_2.n252 VDDA_2.n9 3.4105
R19068 VDDA_2.n252 VDDA_2.n24 3.4105
R19069 VDDA_2.n252 VDDA_2.n8 3.4105
R19070 VDDA_2.n252 VDDA_2.n25 3.4105
R19071 VDDA_2.n252 VDDA_2.n7 3.4105
R19072 VDDA_2.n252 VDDA_2.n26 3.4105
R19073 VDDA_2.n252 VDDA_2.n6 3.4105
R19074 VDDA_2.n252 VDDA_2.n27 3.4105
R19075 VDDA_2.n252 VDDA_2.n5 3.4105
R19076 VDDA_2.n252 VDDA_2.n28 3.4105
R19077 VDDA_2.n252 VDDA_2.n4 3.4105
R19078 VDDA_2.n252 VDDA_2.n29 3.4105
R19079 VDDA_2.n252 VDDA_2.n3 3.4105
R19080 VDDA_2.n252 VDDA_2.n30 3.4105
R19081 VDDA_2.n252 VDDA_2.n2 3.4105
R19082 VDDA_2.n252 VDDA_2.n31 3.4105
R19083 VDDA_2.n252 VDDA_2.n1 3.4105
R19084 VDDA_2.n252 VDDA_2.n32 3.4105
R19085 VDDA_2.n336 VDDA_2.n252 3.4105
R19086 VDDA_2.n317 VDDA_2.n288 3.4105
R19087 VDDA_2.n288 VDDA_2.n17 3.4105
R19088 VDDA_2.n288 VDDA_2.n15 3.4105
R19089 VDDA_2.n288 VDDA_2.n18 3.4105
R19090 VDDA_2.n288 VDDA_2.n14 3.4105
R19091 VDDA_2.n288 VDDA_2.n19 3.4105
R19092 VDDA_2.n288 VDDA_2.n13 3.4105
R19093 VDDA_2.n288 VDDA_2.n20 3.4105
R19094 VDDA_2.n288 VDDA_2.n12 3.4105
R19095 VDDA_2.n288 VDDA_2.n21 3.4105
R19096 VDDA_2.n288 VDDA_2.n11 3.4105
R19097 VDDA_2.n288 VDDA_2.n22 3.4105
R19098 VDDA_2.n288 VDDA_2.n10 3.4105
R19099 VDDA_2.n288 VDDA_2.n23 3.4105
R19100 VDDA_2.n288 VDDA_2.n9 3.4105
R19101 VDDA_2.n288 VDDA_2.n24 3.4105
R19102 VDDA_2.n288 VDDA_2.n8 3.4105
R19103 VDDA_2.n288 VDDA_2.n25 3.4105
R19104 VDDA_2.n288 VDDA_2.n7 3.4105
R19105 VDDA_2.n288 VDDA_2.n26 3.4105
R19106 VDDA_2.n288 VDDA_2.n6 3.4105
R19107 VDDA_2.n288 VDDA_2.n27 3.4105
R19108 VDDA_2.n288 VDDA_2.n5 3.4105
R19109 VDDA_2.n288 VDDA_2.n28 3.4105
R19110 VDDA_2.n288 VDDA_2.n4 3.4105
R19111 VDDA_2.n288 VDDA_2.n29 3.4105
R19112 VDDA_2.n288 VDDA_2.n3 3.4105
R19113 VDDA_2.n288 VDDA_2.n30 3.4105
R19114 VDDA_2.n288 VDDA_2.n2 3.4105
R19115 VDDA_2.n288 VDDA_2.n31 3.4105
R19116 VDDA_2.n288 VDDA_2.n1 3.4105
R19117 VDDA_2.n288 VDDA_2.n32 3.4105
R19118 VDDA_2.n336 VDDA_2.n288 3.4105
R19119 VDDA_2.n317 VDDA_2.n251 3.4105
R19120 VDDA_2.n251 VDDA_2.n17 3.4105
R19121 VDDA_2.n251 VDDA_2.n15 3.4105
R19122 VDDA_2.n251 VDDA_2.n18 3.4105
R19123 VDDA_2.n251 VDDA_2.n14 3.4105
R19124 VDDA_2.n251 VDDA_2.n19 3.4105
R19125 VDDA_2.n251 VDDA_2.n13 3.4105
R19126 VDDA_2.n251 VDDA_2.n20 3.4105
R19127 VDDA_2.n251 VDDA_2.n12 3.4105
R19128 VDDA_2.n251 VDDA_2.n21 3.4105
R19129 VDDA_2.n251 VDDA_2.n11 3.4105
R19130 VDDA_2.n251 VDDA_2.n22 3.4105
R19131 VDDA_2.n251 VDDA_2.n10 3.4105
R19132 VDDA_2.n251 VDDA_2.n23 3.4105
R19133 VDDA_2.n251 VDDA_2.n9 3.4105
R19134 VDDA_2.n251 VDDA_2.n24 3.4105
R19135 VDDA_2.n251 VDDA_2.n8 3.4105
R19136 VDDA_2.n251 VDDA_2.n25 3.4105
R19137 VDDA_2.n251 VDDA_2.n7 3.4105
R19138 VDDA_2.n251 VDDA_2.n26 3.4105
R19139 VDDA_2.n251 VDDA_2.n6 3.4105
R19140 VDDA_2.n251 VDDA_2.n27 3.4105
R19141 VDDA_2.n251 VDDA_2.n5 3.4105
R19142 VDDA_2.n251 VDDA_2.n28 3.4105
R19143 VDDA_2.n251 VDDA_2.n4 3.4105
R19144 VDDA_2.n251 VDDA_2.n29 3.4105
R19145 VDDA_2.n251 VDDA_2.n3 3.4105
R19146 VDDA_2.n251 VDDA_2.n30 3.4105
R19147 VDDA_2.n251 VDDA_2.n2 3.4105
R19148 VDDA_2.n251 VDDA_2.n31 3.4105
R19149 VDDA_2.n251 VDDA_2.n1 3.4105
R19150 VDDA_2.n251 VDDA_2.n32 3.4105
R19151 VDDA_2.n336 VDDA_2.n251 3.4105
R19152 VDDA_2.n317 VDDA_2.n290 3.4105
R19153 VDDA_2.n290 VDDA_2.n17 3.4105
R19154 VDDA_2.n290 VDDA_2.n15 3.4105
R19155 VDDA_2.n290 VDDA_2.n18 3.4105
R19156 VDDA_2.n290 VDDA_2.n14 3.4105
R19157 VDDA_2.n290 VDDA_2.n19 3.4105
R19158 VDDA_2.n290 VDDA_2.n13 3.4105
R19159 VDDA_2.n290 VDDA_2.n20 3.4105
R19160 VDDA_2.n290 VDDA_2.n12 3.4105
R19161 VDDA_2.n290 VDDA_2.n21 3.4105
R19162 VDDA_2.n290 VDDA_2.n11 3.4105
R19163 VDDA_2.n290 VDDA_2.n22 3.4105
R19164 VDDA_2.n290 VDDA_2.n10 3.4105
R19165 VDDA_2.n290 VDDA_2.n23 3.4105
R19166 VDDA_2.n290 VDDA_2.n9 3.4105
R19167 VDDA_2.n290 VDDA_2.n24 3.4105
R19168 VDDA_2.n290 VDDA_2.n8 3.4105
R19169 VDDA_2.n290 VDDA_2.n25 3.4105
R19170 VDDA_2.n290 VDDA_2.n7 3.4105
R19171 VDDA_2.n290 VDDA_2.n26 3.4105
R19172 VDDA_2.n290 VDDA_2.n6 3.4105
R19173 VDDA_2.n290 VDDA_2.n27 3.4105
R19174 VDDA_2.n290 VDDA_2.n5 3.4105
R19175 VDDA_2.n290 VDDA_2.n28 3.4105
R19176 VDDA_2.n290 VDDA_2.n4 3.4105
R19177 VDDA_2.n290 VDDA_2.n29 3.4105
R19178 VDDA_2.n290 VDDA_2.n3 3.4105
R19179 VDDA_2.n290 VDDA_2.n30 3.4105
R19180 VDDA_2.n290 VDDA_2.n2 3.4105
R19181 VDDA_2.n290 VDDA_2.n31 3.4105
R19182 VDDA_2.n290 VDDA_2.n1 3.4105
R19183 VDDA_2.n290 VDDA_2.n32 3.4105
R19184 VDDA_2.n336 VDDA_2.n290 3.4105
R19185 VDDA_2.n317 VDDA_2.n250 3.4105
R19186 VDDA_2.n250 VDDA_2.n17 3.4105
R19187 VDDA_2.n250 VDDA_2.n15 3.4105
R19188 VDDA_2.n250 VDDA_2.n18 3.4105
R19189 VDDA_2.n250 VDDA_2.n14 3.4105
R19190 VDDA_2.n250 VDDA_2.n19 3.4105
R19191 VDDA_2.n250 VDDA_2.n13 3.4105
R19192 VDDA_2.n250 VDDA_2.n20 3.4105
R19193 VDDA_2.n250 VDDA_2.n12 3.4105
R19194 VDDA_2.n250 VDDA_2.n21 3.4105
R19195 VDDA_2.n250 VDDA_2.n11 3.4105
R19196 VDDA_2.n250 VDDA_2.n22 3.4105
R19197 VDDA_2.n250 VDDA_2.n10 3.4105
R19198 VDDA_2.n250 VDDA_2.n23 3.4105
R19199 VDDA_2.n250 VDDA_2.n9 3.4105
R19200 VDDA_2.n250 VDDA_2.n24 3.4105
R19201 VDDA_2.n250 VDDA_2.n8 3.4105
R19202 VDDA_2.n250 VDDA_2.n25 3.4105
R19203 VDDA_2.n250 VDDA_2.n7 3.4105
R19204 VDDA_2.n250 VDDA_2.n26 3.4105
R19205 VDDA_2.n250 VDDA_2.n6 3.4105
R19206 VDDA_2.n250 VDDA_2.n27 3.4105
R19207 VDDA_2.n250 VDDA_2.n5 3.4105
R19208 VDDA_2.n250 VDDA_2.n28 3.4105
R19209 VDDA_2.n250 VDDA_2.n4 3.4105
R19210 VDDA_2.n250 VDDA_2.n29 3.4105
R19211 VDDA_2.n250 VDDA_2.n3 3.4105
R19212 VDDA_2.n250 VDDA_2.n30 3.4105
R19213 VDDA_2.n250 VDDA_2.n2 3.4105
R19214 VDDA_2.n250 VDDA_2.n31 3.4105
R19215 VDDA_2.n250 VDDA_2.n1 3.4105
R19216 VDDA_2.n250 VDDA_2.n32 3.4105
R19217 VDDA_2.n336 VDDA_2.n250 3.4105
R19218 VDDA_2.n317 VDDA_2.n292 3.4105
R19219 VDDA_2.n292 VDDA_2.n17 3.4105
R19220 VDDA_2.n292 VDDA_2.n15 3.4105
R19221 VDDA_2.n292 VDDA_2.n18 3.4105
R19222 VDDA_2.n292 VDDA_2.n14 3.4105
R19223 VDDA_2.n292 VDDA_2.n19 3.4105
R19224 VDDA_2.n292 VDDA_2.n13 3.4105
R19225 VDDA_2.n292 VDDA_2.n20 3.4105
R19226 VDDA_2.n292 VDDA_2.n12 3.4105
R19227 VDDA_2.n292 VDDA_2.n21 3.4105
R19228 VDDA_2.n292 VDDA_2.n11 3.4105
R19229 VDDA_2.n292 VDDA_2.n22 3.4105
R19230 VDDA_2.n292 VDDA_2.n10 3.4105
R19231 VDDA_2.n292 VDDA_2.n23 3.4105
R19232 VDDA_2.n292 VDDA_2.n9 3.4105
R19233 VDDA_2.n292 VDDA_2.n24 3.4105
R19234 VDDA_2.n292 VDDA_2.n8 3.4105
R19235 VDDA_2.n292 VDDA_2.n25 3.4105
R19236 VDDA_2.n292 VDDA_2.n7 3.4105
R19237 VDDA_2.n292 VDDA_2.n26 3.4105
R19238 VDDA_2.n292 VDDA_2.n6 3.4105
R19239 VDDA_2.n292 VDDA_2.n27 3.4105
R19240 VDDA_2.n292 VDDA_2.n5 3.4105
R19241 VDDA_2.n292 VDDA_2.n28 3.4105
R19242 VDDA_2.n292 VDDA_2.n4 3.4105
R19243 VDDA_2.n292 VDDA_2.n29 3.4105
R19244 VDDA_2.n292 VDDA_2.n3 3.4105
R19245 VDDA_2.n292 VDDA_2.n30 3.4105
R19246 VDDA_2.n292 VDDA_2.n2 3.4105
R19247 VDDA_2.n292 VDDA_2.n31 3.4105
R19248 VDDA_2.n292 VDDA_2.n1 3.4105
R19249 VDDA_2.n292 VDDA_2.n32 3.4105
R19250 VDDA_2.n336 VDDA_2.n292 3.4105
R19251 VDDA_2.n317 VDDA_2.n249 3.4105
R19252 VDDA_2.n249 VDDA_2.n17 3.4105
R19253 VDDA_2.n249 VDDA_2.n15 3.4105
R19254 VDDA_2.n249 VDDA_2.n18 3.4105
R19255 VDDA_2.n249 VDDA_2.n14 3.4105
R19256 VDDA_2.n249 VDDA_2.n19 3.4105
R19257 VDDA_2.n249 VDDA_2.n13 3.4105
R19258 VDDA_2.n249 VDDA_2.n20 3.4105
R19259 VDDA_2.n249 VDDA_2.n12 3.4105
R19260 VDDA_2.n249 VDDA_2.n21 3.4105
R19261 VDDA_2.n249 VDDA_2.n11 3.4105
R19262 VDDA_2.n249 VDDA_2.n22 3.4105
R19263 VDDA_2.n249 VDDA_2.n10 3.4105
R19264 VDDA_2.n249 VDDA_2.n23 3.4105
R19265 VDDA_2.n249 VDDA_2.n9 3.4105
R19266 VDDA_2.n249 VDDA_2.n24 3.4105
R19267 VDDA_2.n249 VDDA_2.n8 3.4105
R19268 VDDA_2.n249 VDDA_2.n25 3.4105
R19269 VDDA_2.n249 VDDA_2.n7 3.4105
R19270 VDDA_2.n249 VDDA_2.n26 3.4105
R19271 VDDA_2.n249 VDDA_2.n6 3.4105
R19272 VDDA_2.n249 VDDA_2.n27 3.4105
R19273 VDDA_2.n249 VDDA_2.n5 3.4105
R19274 VDDA_2.n249 VDDA_2.n28 3.4105
R19275 VDDA_2.n249 VDDA_2.n4 3.4105
R19276 VDDA_2.n249 VDDA_2.n29 3.4105
R19277 VDDA_2.n249 VDDA_2.n3 3.4105
R19278 VDDA_2.n249 VDDA_2.n30 3.4105
R19279 VDDA_2.n249 VDDA_2.n2 3.4105
R19280 VDDA_2.n249 VDDA_2.n31 3.4105
R19281 VDDA_2.n249 VDDA_2.n1 3.4105
R19282 VDDA_2.n249 VDDA_2.n32 3.4105
R19283 VDDA_2.n336 VDDA_2.n249 3.4105
R19284 VDDA_2.n317 VDDA_2.n294 3.4105
R19285 VDDA_2.n294 VDDA_2.n17 3.4105
R19286 VDDA_2.n294 VDDA_2.n15 3.4105
R19287 VDDA_2.n294 VDDA_2.n18 3.4105
R19288 VDDA_2.n294 VDDA_2.n14 3.4105
R19289 VDDA_2.n294 VDDA_2.n19 3.4105
R19290 VDDA_2.n294 VDDA_2.n13 3.4105
R19291 VDDA_2.n294 VDDA_2.n20 3.4105
R19292 VDDA_2.n294 VDDA_2.n12 3.4105
R19293 VDDA_2.n294 VDDA_2.n21 3.4105
R19294 VDDA_2.n294 VDDA_2.n11 3.4105
R19295 VDDA_2.n294 VDDA_2.n22 3.4105
R19296 VDDA_2.n294 VDDA_2.n10 3.4105
R19297 VDDA_2.n294 VDDA_2.n23 3.4105
R19298 VDDA_2.n294 VDDA_2.n9 3.4105
R19299 VDDA_2.n294 VDDA_2.n24 3.4105
R19300 VDDA_2.n294 VDDA_2.n8 3.4105
R19301 VDDA_2.n294 VDDA_2.n25 3.4105
R19302 VDDA_2.n294 VDDA_2.n7 3.4105
R19303 VDDA_2.n294 VDDA_2.n26 3.4105
R19304 VDDA_2.n294 VDDA_2.n6 3.4105
R19305 VDDA_2.n294 VDDA_2.n27 3.4105
R19306 VDDA_2.n294 VDDA_2.n5 3.4105
R19307 VDDA_2.n294 VDDA_2.n28 3.4105
R19308 VDDA_2.n294 VDDA_2.n4 3.4105
R19309 VDDA_2.n294 VDDA_2.n29 3.4105
R19310 VDDA_2.n294 VDDA_2.n3 3.4105
R19311 VDDA_2.n294 VDDA_2.n30 3.4105
R19312 VDDA_2.n294 VDDA_2.n2 3.4105
R19313 VDDA_2.n294 VDDA_2.n31 3.4105
R19314 VDDA_2.n294 VDDA_2.n1 3.4105
R19315 VDDA_2.n294 VDDA_2.n32 3.4105
R19316 VDDA_2.n336 VDDA_2.n294 3.4105
R19317 VDDA_2.n317 VDDA_2.n248 3.4105
R19318 VDDA_2.n248 VDDA_2.n17 3.4105
R19319 VDDA_2.n248 VDDA_2.n15 3.4105
R19320 VDDA_2.n248 VDDA_2.n18 3.4105
R19321 VDDA_2.n248 VDDA_2.n14 3.4105
R19322 VDDA_2.n248 VDDA_2.n19 3.4105
R19323 VDDA_2.n248 VDDA_2.n13 3.4105
R19324 VDDA_2.n248 VDDA_2.n20 3.4105
R19325 VDDA_2.n248 VDDA_2.n12 3.4105
R19326 VDDA_2.n248 VDDA_2.n21 3.4105
R19327 VDDA_2.n248 VDDA_2.n11 3.4105
R19328 VDDA_2.n248 VDDA_2.n22 3.4105
R19329 VDDA_2.n248 VDDA_2.n10 3.4105
R19330 VDDA_2.n248 VDDA_2.n23 3.4105
R19331 VDDA_2.n248 VDDA_2.n9 3.4105
R19332 VDDA_2.n248 VDDA_2.n24 3.4105
R19333 VDDA_2.n248 VDDA_2.n8 3.4105
R19334 VDDA_2.n248 VDDA_2.n25 3.4105
R19335 VDDA_2.n248 VDDA_2.n7 3.4105
R19336 VDDA_2.n248 VDDA_2.n26 3.4105
R19337 VDDA_2.n248 VDDA_2.n6 3.4105
R19338 VDDA_2.n248 VDDA_2.n27 3.4105
R19339 VDDA_2.n248 VDDA_2.n5 3.4105
R19340 VDDA_2.n248 VDDA_2.n28 3.4105
R19341 VDDA_2.n248 VDDA_2.n4 3.4105
R19342 VDDA_2.n248 VDDA_2.n29 3.4105
R19343 VDDA_2.n248 VDDA_2.n3 3.4105
R19344 VDDA_2.n248 VDDA_2.n30 3.4105
R19345 VDDA_2.n248 VDDA_2.n2 3.4105
R19346 VDDA_2.n248 VDDA_2.n31 3.4105
R19347 VDDA_2.n248 VDDA_2.n1 3.4105
R19348 VDDA_2.n248 VDDA_2.n32 3.4105
R19349 VDDA_2.n336 VDDA_2.n248 3.4105
R19350 VDDA_2.n317 VDDA_2.n296 3.4105
R19351 VDDA_2.n296 VDDA_2.n17 3.4105
R19352 VDDA_2.n296 VDDA_2.n15 3.4105
R19353 VDDA_2.n296 VDDA_2.n18 3.4105
R19354 VDDA_2.n296 VDDA_2.n14 3.4105
R19355 VDDA_2.n296 VDDA_2.n19 3.4105
R19356 VDDA_2.n296 VDDA_2.n13 3.4105
R19357 VDDA_2.n296 VDDA_2.n20 3.4105
R19358 VDDA_2.n296 VDDA_2.n12 3.4105
R19359 VDDA_2.n296 VDDA_2.n21 3.4105
R19360 VDDA_2.n296 VDDA_2.n11 3.4105
R19361 VDDA_2.n296 VDDA_2.n22 3.4105
R19362 VDDA_2.n296 VDDA_2.n10 3.4105
R19363 VDDA_2.n296 VDDA_2.n23 3.4105
R19364 VDDA_2.n296 VDDA_2.n9 3.4105
R19365 VDDA_2.n296 VDDA_2.n24 3.4105
R19366 VDDA_2.n296 VDDA_2.n8 3.4105
R19367 VDDA_2.n296 VDDA_2.n25 3.4105
R19368 VDDA_2.n296 VDDA_2.n7 3.4105
R19369 VDDA_2.n296 VDDA_2.n26 3.4105
R19370 VDDA_2.n296 VDDA_2.n6 3.4105
R19371 VDDA_2.n296 VDDA_2.n27 3.4105
R19372 VDDA_2.n296 VDDA_2.n5 3.4105
R19373 VDDA_2.n296 VDDA_2.n28 3.4105
R19374 VDDA_2.n296 VDDA_2.n4 3.4105
R19375 VDDA_2.n296 VDDA_2.n29 3.4105
R19376 VDDA_2.n296 VDDA_2.n3 3.4105
R19377 VDDA_2.n296 VDDA_2.n30 3.4105
R19378 VDDA_2.n296 VDDA_2.n2 3.4105
R19379 VDDA_2.n296 VDDA_2.n31 3.4105
R19380 VDDA_2.n296 VDDA_2.n1 3.4105
R19381 VDDA_2.n296 VDDA_2.n32 3.4105
R19382 VDDA_2.n336 VDDA_2.n296 3.4105
R19383 VDDA_2.n317 VDDA_2.n247 3.4105
R19384 VDDA_2.n247 VDDA_2.n17 3.4105
R19385 VDDA_2.n247 VDDA_2.n15 3.4105
R19386 VDDA_2.n247 VDDA_2.n18 3.4105
R19387 VDDA_2.n247 VDDA_2.n14 3.4105
R19388 VDDA_2.n247 VDDA_2.n19 3.4105
R19389 VDDA_2.n247 VDDA_2.n13 3.4105
R19390 VDDA_2.n247 VDDA_2.n20 3.4105
R19391 VDDA_2.n247 VDDA_2.n12 3.4105
R19392 VDDA_2.n247 VDDA_2.n21 3.4105
R19393 VDDA_2.n247 VDDA_2.n11 3.4105
R19394 VDDA_2.n247 VDDA_2.n22 3.4105
R19395 VDDA_2.n247 VDDA_2.n10 3.4105
R19396 VDDA_2.n247 VDDA_2.n23 3.4105
R19397 VDDA_2.n247 VDDA_2.n9 3.4105
R19398 VDDA_2.n247 VDDA_2.n24 3.4105
R19399 VDDA_2.n247 VDDA_2.n8 3.4105
R19400 VDDA_2.n247 VDDA_2.n25 3.4105
R19401 VDDA_2.n247 VDDA_2.n7 3.4105
R19402 VDDA_2.n247 VDDA_2.n26 3.4105
R19403 VDDA_2.n247 VDDA_2.n6 3.4105
R19404 VDDA_2.n247 VDDA_2.n27 3.4105
R19405 VDDA_2.n247 VDDA_2.n5 3.4105
R19406 VDDA_2.n247 VDDA_2.n28 3.4105
R19407 VDDA_2.n247 VDDA_2.n4 3.4105
R19408 VDDA_2.n247 VDDA_2.n29 3.4105
R19409 VDDA_2.n247 VDDA_2.n3 3.4105
R19410 VDDA_2.n247 VDDA_2.n30 3.4105
R19411 VDDA_2.n247 VDDA_2.n2 3.4105
R19412 VDDA_2.n247 VDDA_2.n31 3.4105
R19413 VDDA_2.n247 VDDA_2.n1 3.4105
R19414 VDDA_2.n247 VDDA_2.n32 3.4105
R19415 VDDA_2.n336 VDDA_2.n247 3.4105
R19416 VDDA_2.n317 VDDA_2.n298 3.4105
R19417 VDDA_2.n298 VDDA_2.n17 3.4105
R19418 VDDA_2.n298 VDDA_2.n15 3.4105
R19419 VDDA_2.n298 VDDA_2.n18 3.4105
R19420 VDDA_2.n298 VDDA_2.n14 3.4105
R19421 VDDA_2.n298 VDDA_2.n19 3.4105
R19422 VDDA_2.n298 VDDA_2.n13 3.4105
R19423 VDDA_2.n298 VDDA_2.n20 3.4105
R19424 VDDA_2.n298 VDDA_2.n12 3.4105
R19425 VDDA_2.n298 VDDA_2.n21 3.4105
R19426 VDDA_2.n298 VDDA_2.n11 3.4105
R19427 VDDA_2.n298 VDDA_2.n22 3.4105
R19428 VDDA_2.n298 VDDA_2.n10 3.4105
R19429 VDDA_2.n298 VDDA_2.n23 3.4105
R19430 VDDA_2.n298 VDDA_2.n9 3.4105
R19431 VDDA_2.n298 VDDA_2.n24 3.4105
R19432 VDDA_2.n298 VDDA_2.n8 3.4105
R19433 VDDA_2.n298 VDDA_2.n25 3.4105
R19434 VDDA_2.n298 VDDA_2.n7 3.4105
R19435 VDDA_2.n298 VDDA_2.n26 3.4105
R19436 VDDA_2.n298 VDDA_2.n6 3.4105
R19437 VDDA_2.n298 VDDA_2.n27 3.4105
R19438 VDDA_2.n298 VDDA_2.n5 3.4105
R19439 VDDA_2.n298 VDDA_2.n28 3.4105
R19440 VDDA_2.n298 VDDA_2.n4 3.4105
R19441 VDDA_2.n298 VDDA_2.n29 3.4105
R19442 VDDA_2.n298 VDDA_2.n3 3.4105
R19443 VDDA_2.n298 VDDA_2.n30 3.4105
R19444 VDDA_2.n298 VDDA_2.n2 3.4105
R19445 VDDA_2.n298 VDDA_2.n31 3.4105
R19446 VDDA_2.n298 VDDA_2.n1 3.4105
R19447 VDDA_2.n298 VDDA_2.n32 3.4105
R19448 VDDA_2.n336 VDDA_2.n298 3.4105
R19449 VDDA_2.n317 VDDA_2.n246 3.4105
R19450 VDDA_2.n246 VDDA_2.n17 3.4105
R19451 VDDA_2.n246 VDDA_2.n15 3.4105
R19452 VDDA_2.n246 VDDA_2.n18 3.4105
R19453 VDDA_2.n246 VDDA_2.n14 3.4105
R19454 VDDA_2.n246 VDDA_2.n19 3.4105
R19455 VDDA_2.n246 VDDA_2.n13 3.4105
R19456 VDDA_2.n246 VDDA_2.n20 3.4105
R19457 VDDA_2.n246 VDDA_2.n12 3.4105
R19458 VDDA_2.n246 VDDA_2.n21 3.4105
R19459 VDDA_2.n246 VDDA_2.n11 3.4105
R19460 VDDA_2.n246 VDDA_2.n22 3.4105
R19461 VDDA_2.n246 VDDA_2.n10 3.4105
R19462 VDDA_2.n246 VDDA_2.n23 3.4105
R19463 VDDA_2.n246 VDDA_2.n9 3.4105
R19464 VDDA_2.n246 VDDA_2.n24 3.4105
R19465 VDDA_2.n246 VDDA_2.n8 3.4105
R19466 VDDA_2.n246 VDDA_2.n25 3.4105
R19467 VDDA_2.n246 VDDA_2.n7 3.4105
R19468 VDDA_2.n246 VDDA_2.n26 3.4105
R19469 VDDA_2.n246 VDDA_2.n6 3.4105
R19470 VDDA_2.n246 VDDA_2.n27 3.4105
R19471 VDDA_2.n246 VDDA_2.n5 3.4105
R19472 VDDA_2.n246 VDDA_2.n28 3.4105
R19473 VDDA_2.n246 VDDA_2.n4 3.4105
R19474 VDDA_2.n246 VDDA_2.n29 3.4105
R19475 VDDA_2.n246 VDDA_2.n3 3.4105
R19476 VDDA_2.n246 VDDA_2.n30 3.4105
R19477 VDDA_2.n246 VDDA_2.n2 3.4105
R19478 VDDA_2.n246 VDDA_2.n31 3.4105
R19479 VDDA_2.n246 VDDA_2.n1 3.4105
R19480 VDDA_2.n246 VDDA_2.n32 3.4105
R19481 VDDA_2.n336 VDDA_2.n246 3.4105
R19482 VDDA_2.n317 VDDA_2.n300 3.4105
R19483 VDDA_2.n300 VDDA_2.n17 3.4105
R19484 VDDA_2.n300 VDDA_2.n15 3.4105
R19485 VDDA_2.n300 VDDA_2.n18 3.4105
R19486 VDDA_2.n300 VDDA_2.n14 3.4105
R19487 VDDA_2.n300 VDDA_2.n19 3.4105
R19488 VDDA_2.n300 VDDA_2.n13 3.4105
R19489 VDDA_2.n300 VDDA_2.n20 3.4105
R19490 VDDA_2.n300 VDDA_2.n12 3.4105
R19491 VDDA_2.n300 VDDA_2.n21 3.4105
R19492 VDDA_2.n300 VDDA_2.n11 3.4105
R19493 VDDA_2.n300 VDDA_2.n22 3.4105
R19494 VDDA_2.n300 VDDA_2.n10 3.4105
R19495 VDDA_2.n300 VDDA_2.n23 3.4105
R19496 VDDA_2.n300 VDDA_2.n9 3.4105
R19497 VDDA_2.n300 VDDA_2.n24 3.4105
R19498 VDDA_2.n300 VDDA_2.n8 3.4105
R19499 VDDA_2.n300 VDDA_2.n25 3.4105
R19500 VDDA_2.n300 VDDA_2.n7 3.4105
R19501 VDDA_2.n300 VDDA_2.n26 3.4105
R19502 VDDA_2.n300 VDDA_2.n6 3.4105
R19503 VDDA_2.n300 VDDA_2.n27 3.4105
R19504 VDDA_2.n300 VDDA_2.n5 3.4105
R19505 VDDA_2.n300 VDDA_2.n28 3.4105
R19506 VDDA_2.n300 VDDA_2.n4 3.4105
R19507 VDDA_2.n300 VDDA_2.n29 3.4105
R19508 VDDA_2.n300 VDDA_2.n3 3.4105
R19509 VDDA_2.n300 VDDA_2.n30 3.4105
R19510 VDDA_2.n300 VDDA_2.n2 3.4105
R19511 VDDA_2.n300 VDDA_2.n31 3.4105
R19512 VDDA_2.n300 VDDA_2.n1 3.4105
R19513 VDDA_2.n300 VDDA_2.n32 3.4105
R19514 VDDA_2.n336 VDDA_2.n300 3.4105
R19515 VDDA_2.n317 VDDA_2.n245 3.4105
R19516 VDDA_2.n245 VDDA_2.n17 3.4105
R19517 VDDA_2.n245 VDDA_2.n15 3.4105
R19518 VDDA_2.n245 VDDA_2.n18 3.4105
R19519 VDDA_2.n245 VDDA_2.n14 3.4105
R19520 VDDA_2.n245 VDDA_2.n19 3.4105
R19521 VDDA_2.n245 VDDA_2.n13 3.4105
R19522 VDDA_2.n245 VDDA_2.n20 3.4105
R19523 VDDA_2.n245 VDDA_2.n12 3.4105
R19524 VDDA_2.n245 VDDA_2.n21 3.4105
R19525 VDDA_2.n245 VDDA_2.n11 3.4105
R19526 VDDA_2.n245 VDDA_2.n22 3.4105
R19527 VDDA_2.n245 VDDA_2.n10 3.4105
R19528 VDDA_2.n245 VDDA_2.n23 3.4105
R19529 VDDA_2.n245 VDDA_2.n9 3.4105
R19530 VDDA_2.n245 VDDA_2.n24 3.4105
R19531 VDDA_2.n245 VDDA_2.n8 3.4105
R19532 VDDA_2.n245 VDDA_2.n25 3.4105
R19533 VDDA_2.n245 VDDA_2.n7 3.4105
R19534 VDDA_2.n245 VDDA_2.n26 3.4105
R19535 VDDA_2.n245 VDDA_2.n6 3.4105
R19536 VDDA_2.n245 VDDA_2.n27 3.4105
R19537 VDDA_2.n245 VDDA_2.n5 3.4105
R19538 VDDA_2.n245 VDDA_2.n28 3.4105
R19539 VDDA_2.n245 VDDA_2.n4 3.4105
R19540 VDDA_2.n245 VDDA_2.n29 3.4105
R19541 VDDA_2.n245 VDDA_2.n3 3.4105
R19542 VDDA_2.n245 VDDA_2.n30 3.4105
R19543 VDDA_2.n245 VDDA_2.n2 3.4105
R19544 VDDA_2.n245 VDDA_2.n31 3.4105
R19545 VDDA_2.n245 VDDA_2.n1 3.4105
R19546 VDDA_2.n245 VDDA_2.n32 3.4105
R19547 VDDA_2.n336 VDDA_2.n245 3.4105
R19548 VDDA_2.n317 VDDA_2.n302 3.4105
R19549 VDDA_2.n302 VDDA_2.n17 3.4105
R19550 VDDA_2.n302 VDDA_2.n15 3.4105
R19551 VDDA_2.n302 VDDA_2.n18 3.4105
R19552 VDDA_2.n302 VDDA_2.n14 3.4105
R19553 VDDA_2.n302 VDDA_2.n19 3.4105
R19554 VDDA_2.n302 VDDA_2.n13 3.4105
R19555 VDDA_2.n302 VDDA_2.n20 3.4105
R19556 VDDA_2.n302 VDDA_2.n12 3.4105
R19557 VDDA_2.n302 VDDA_2.n21 3.4105
R19558 VDDA_2.n302 VDDA_2.n11 3.4105
R19559 VDDA_2.n302 VDDA_2.n22 3.4105
R19560 VDDA_2.n302 VDDA_2.n10 3.4105
R19561 VDDA_2.n302 VDDA_2.n23 3.4105
R19562 VDDA_2.n302 VDDA_2.n9 3.4105
R19563 VDDA_2.n302 VDDA_2.n24 3.4105
R19564 VDDA_2.n302 VDDA_2.n8 3.4105
R19565 VDDA_2.n302 VDDA_2.n25 3.4105
R19566 VDDA_2.n302 VDDA_2.n7 3.4105
R19567 VDDA_2.n302 VDDA_2.n26 3.4105
R19568 VDDA_2.n302 VDDA_2.n6 3.4105
R19569 VDDA_2.n302 VDDA_2.n27 3.4105
R19570 VDDA_2.n302 VDDA_2.n5 3.4105
R19571 VDDA_2.n302 VDDA_2.n28 3.4105
R19572 VDDA_2.n302 VDDA_2.n4 3.4105
R19573 VDDA_2.n302 VDDA_2.n29 3.4105
R19574 VDDA_2.n302 VDDA_2.n3 3.4105
R19575 VDDA_2.n302 VDDA_2.n30 3.4105
R19576 VDDA_2.n302 VDDA_2.n2 3.4105
R19577 VDDA_2.n302 VDDA_2.n31 3.4105
R19578 VDDA_2.n302 VDDA_2.n1 3.4105
R19579 VDDA_2.n302 VDDA_2.n32 3.4105
R19580 VDDA_2.n336 VDDA_2.n302 3.4105
R19581 VDDA_2.n317 VDDA_2.n244 3.4105
R19582 VDDA_2.n244 VDDA_2.n17 3.4105
R19583 VDDA_2.n244 VDDA_2.n15 3.4105
R19584 VDDA_2.n244 VDDA_2.n18 3.4105
R19585 VDDA_2.n244 VDDA_2.n14 3.4105
R19586 VDDA_2.n244 VDDA_2.n19 3.4105
R19587 VDDA_2.n244 VDDA_2.n13 3.4105
R19588 VDDA_2.n244 VDDA_2.n20 3.4105
R19589 VDDA_2.n244 VDDA_2.n12 3.4105
R19590 VDDA_2.n244 VDDA_2.n21 3.4105
R19591 VDDA_2.n244 VDDA_2.n11 3.4105
R19592 VDDA_2.n244 VDDA_2.n22 3.4105
R19593 VDDA_2.n244 VDDA_2.n10 3.4105
R19594 VDDA_2.n244 VDDA_2.n23 3.4105
R19595 VDDA_2.n244 VDDA_2.n9 3.4105
R19596 VDDA_2.n244 VDDA_2.n24 3.4105
R19597 VDDA_2.n244 VDDA_2.n8 3.4105
R19598 VDDA_2.n244 VDDA_2.n25 3.4105
R19599 VDDA_2.n244 VDDA_2.n7 3.4105
R19600 VDDA_2.n244 VDDA_2.n26 3.4105
R19601 VDDA_2.n244 VDDA_2.n6 3.4105
R19602 VDDA_2.n244 VDDA_2.n27 3.4105
R19603 VDDA_2.n244 VDDA_2.n5 3.4105
R19604 VDDA_2.n244 VDDA_2.n28 3.4105
R19605 VDDA_2.n244 VDDA_2.n4 3.4105
R19606 VDDA_2.n244 VDDA_2.n29 3.4105
R19607 VDDA_2.n244 VDDA_2.n3 3.4105
R19608 VDDA_2.n244 VDDA_2.n30 3.4105
R19609 VDDA_2.n244 VDDA_2.n2 3.4105
R19610 VDDA_2.n244 VDDA_2.n31 3.4105
R19611 VDDA_2.n244 VDDA_2.n1 3.4105
R19612 VDDA_2.n244 VDDA_2.n32 3.4105
R19613 VDDA_2.n336 VDDA_2.n244 3.4105
R19614 VDDA_2.n317 VDDA_2.n304 3.4105
R19615 VDDA_2.n304 VDDA_2.n17 3.4105
R19616 VDDA_2.n304 VDDA_2.n15 3.4105
R19617 VDDA_2.n304 VDDA_2.n18 3.4105
R19618 VDDA_2.n304 VDDA_2.n14 3.4105
R19619 VDDA_2.n304 VDDA_2.n19 3.4105
R19620 VDDA_2.n304 VDDA_2.n13 3.4105
R19621 VDDA_2.n304 VDDA_2.n20 3.4105
R19622 VDDA_2.n304 VDDA_2.n12 3.4105
R19623 VDDA_2.n304 VDDA_2.n21 3.4105
R19624 VDDA_2.n304 VDDA_2.n11 3.4105
R19625 VDDA_2.n304 VDDA_2.n22 3.4105
R19626 VDDA_2.n304 VDDA_2.n10 3.4105
R19627 VDDA_2.n304 VDDA_2.n23 3.4105
R19628 VDDA_2.n304 VDDA_2.n9 3.4105
R19629 VDDA_2.n304 VDDA_2.n24 3.4105
R19630 VDDA_2.n304 VDDA_2.n8 3.4105
R19631 VDDA_2.n304 VDDA_2.n25 3.4105
R19632 VDDA_2.n304 VDDA_2.n7 3.4105
R19633 VDDA_2.n304 VDDA_2.n26 3.4105
R19634 VDDA_2.n304 VDDA_2.n6 3.4105
R19635 VDDA_2.n304 VDDA_2.n27 3.4105
R19636 VDDA_2.n304 VDDA_2.n5 3.4105
R19637 VDDA_2.n304 VDDA_2.n28 3.4105
R19638 VDDA_2.n304 VDDA_2.n4 3.4105
R19639 VDDA_2.n304 VDDA_2.n29 3.4105
R19640 VDDA_2.n304 VDDA_2.n3 3.4105
R19641 VDDA_2.n304 VDDA_2.n30 3.4105
R19642 VDDA_2.n304 VDDA_2.n2 3.4105
R19643 VDDA_2.n304 VDDA_2.n31 3.4105
R19644 VDDA_2.n304 VDDA_2.n1 3.4105
R19645 VDDA_2.n304 VDDA_2.n32 3.4105
R19646 VDDA_2.n336 VDDA_2.n304 3.4105
R19647 VDDA_2.n317 VDDA_2.n243 3.4105
R19648 VDDA_2.n243 VDDA_2.n17 3.4105
R19649 VDDA_2.n243 VDDA_2.n15 3.4105
R19650 VDDA_2.n243 VDDA_2.n18 3.4105
R19651 VDDA_2.n243 VDDA_2.n14 3.4105
R19652 VDDA_2.n243 VDDA_2.n19 3.4105
R19653 VDDA_2.n243 VDDA_2.n13 3.4105
R19654 VDDA_2.n243 VDDA_2.n20 3.4105
R19655 VDDA_2.n243 VDDA_2.n12 3.4105
R19656 VDDA_2.n243 VDDA_2.n21 3.4105
R19657 VDDA_2.n243 VDDA_2.n11 3.4105
R19658 VDDA_2.n243 VDDA_2.n22 3.4105
R19659 VDDA_2.n243 VDDA_2.n10 3.4105
R19660 VDDA_2.n243 VDDA_2.n23 3.4105
R19661 VDDA_2.n243 VDDA_2.n9 3.4105
R19662 VDDA_2.n243 VDDA_2.n24 3.4105
R19663 VDDA_2.n243 VDDA_2.n8 3.4105
R19664 VDDA_2.n243 VDDA_2.n25 3.4105
R19665 VDDA_2.n243 VDDA_2.n7 3.4105
R19666 VDDA_2.n243 VDDA_2.n26 3.4105
R19667 VDDA_2.n243 VDDA_2.n6 3.4105
R19668 VDDA_2.n243 VDDA_2.n27 3.4105
R19669 VDDA_2.n243 VDDA_2.n5 3.4105
R19670 VDDA_2.n243 VDDA_2.n28 3.4105
R19671 VDDA_2.n243 VDDA_2.n4 3.4105
R19672 VDDA_2.n243 VDDA_2.n29 3.4105
R19673 VDDA_2.n243 VDDA_2.n3 3.4105
R19674 VDDA_2.n243 VDDA_2.n30 3.4105
R19675 VDDA_2.n243 VDDA_2.n2 3.4105
R19676 VDDA_2.n243 VDDA_2.n31 3.4105
R19677 VDDA_2.n243 VDDA_2.n1 3.4105
R19678 VDDA_2.n243 VDDA_2.n32 3.4105
R19679 VDDA_2.n336 VDDA_2.n243 3.4105
R19680 VDDA_2.n317 VDDA_2.n306 3.4105
R19681 VDDA_2.n306 VDDA_2.n17 3.4105
R19682 VDDA_2.n306 VDDA_2.n15 3.4105
R19683 VDDA_2.n306 VDDA_2.n18 3.4105
R19684 VDDA_2.n306 VDDA_2.n14 3.4105
R19685 VDDA_2.n306 VDDA_2.n19 3.4105
R19686 VDDA_2.n306 VDDA_2.n13 3.4105
R19687 VDDA_2.n306 VDDA_2.n20 3.4105
R19688 VDDA_2.n306 VDDA_2.n12 3.4105
R19689 VDDA_2.n306 VDDA_2.n21 3.4105
R19690 VDDA_2.n306 VDDA_2.n11 3.4105
R19691 VDDA_2.n306 VDDA_2.n22 3.4105
R19692 VDDA_2.n306 VDDA_2.n10 3.4105
R19693 VDDA_2.n306 VDDA_2.n23 3.4105
R19694 VDDA_2.n306 VDDA_2.n9 3.4105
R19695 VDDA_2.n306 VDDA_2.n24 3.4105
R19696 VDDA_2.n306 VDDA_2.n8 3.4105
R19697 VDDA_2.n306 VDDA_2.n25 3.4105
R19698 VDDA_2.n306 VDDA_2.n7 3.4105
R19699 VDDA_2.n306 VDDA_2.n26 3.4105
R19700 VDDA_2.n306 VDDA_2.n6 3.4105
R19701 VDDA_2.n306 VDDA_2.n27 3.4105
R19702 VDDA_2.n306 VDDA_2.n5 3.4105
R19703 VDDA_2.n306 VDDA_2.n28 3.4105
R19704 VDDA_2.n306 VDDA_2.n4 3.4105
R19705 VDDA_2.n306 VDDA_2.n29 3.4105
R19706 VDDA_2.n306 VDDA_2.n3 3.4105
R19707 VDDA_2.n306 VDDA_2.n30 3.4105
R19708 VDDA_2.n306 VDDA_2.n2 3.4105
R19709 VDDA_2.n306 VDDA_2.n31 3.4105
R19710 VDDA_2.n306 VDDA_2.n1 3.4105
R19711 VDDA_2.n306 VDDA_2.n32 3.4105
R19712 VDDA_2.n336 VDDA_2.n306 3.4105
R19713 VDDA_2.n317 VDDA_2.n242 3.4105
R19714 VDDA_2.n242 VDDA_2.n17 3.4105
R19715 VDDA_2.n242 VDDA_2.n15 3.4105
R19716 VDDA_2.n242 VDDA_2.n18 3.4105
R19717 VDDA_2.n242 VDDA_2.n14 3.4105
R19718 VDDA_2.n242 VDDA_2.n19 3.4105
R19719 VDDA_2.n242 VDDA_2.n13 3.4105
R19720 VDDA_2.n242 VDDA_2.n20 3.4105
R19721 VDDA_2.n242 VDDA_2.n12 3.4105
R19722 VDDA_2.n242 VDDA_2.n21 3.4105
R19723 VDDA_2.n242 VDDA_2.n11 3.4105
R19724 VDDA_2.n242 VDDA_2.n22 3.4105
R19725 VDDA_2.n242 VDDA_2.n10 3.4105
R19726 VDDA_2.n242 VDDA_2.n23 3.4105
R19727 VDDA_2.n242 VDDA_2.n9 3.4105
R19728 VDDA_2.n242 VDDA_2.n24 3.4105
R19729 VDDA_2.n242 VDDA_2.n8 3.4105
R19730 VDDA_2.n242 VDDA_2.n25 3.4105
R19731 VDDA_2.n242 VDDA_2.n7 3.4105
R19732 VDDA_2.n242 VDDA_2.n26 3.4105
R19733 VDDA_2.n242 VDDA_2.n6 3.4105
R19734 VDDA_2.n242 VDDA_2.n27 3.4105
R19735 VDDA_2.n242 VDDA_2.n5 3.4105
R19736 VDDA_2.n242 VDDA_2.n28 3.4105
R19737 VDDA_2.n242 VDDA_2.n4 3.4105
R19738 VDDA_2.n242 VDDA_2.n29 3.4105
R19739 VDDA_2.n242 VDDA_2.n3 3.4105
R19740 VDDA_2.n242 VDDA_2.n30 3.4105
R19741 VDDA_2.n242 VDDA_2.n2 3.4105
R19742 VDDA_2.n242 VDDA_2.n31 3.4105
R19743 VDDA_2.n242 VDDA_2.n1 3.4105
R19744 VDDA_2.n242 VDDA_2.n32 3.4105
R19745 VDDA_2.n336 VDDA_2.n242 3.4105
R19746 VDDA_2.n317 VDDA_2.n308 3.4105
R19747 VDDA_2.n308 VDDA_2.n17 3.4105
R19748 VDDA_2.n308 VDDA_2.n15 3.4105
R19749 VDDA_2.n308 VDDA_2.n18 3.4105
R19750 VDDA_2.n308 VDDA_2.n14 3.4105
R19751 VDDA_2.n308 VDDA_2.n19 3.4105
R19752 VDDA_2.n308 VDDA_2.n13 3.4105
R19753 VDDA_2.n308 VDDA_2.n20 3.4105
R19754 VDDA_2.n308 VDDA_2.n12 3.4105
R19755 VDDA_2.n308 VDDA_2.n21 3.4105
R19756 VDDA_2.n308 VDDA_2.n11 3.4105
R19757 VDDA_2.n308 VDDA_2.n22 3.4105
R19758 VDDA_2.n308 VDDA_2.n10 3.4105
R19759 VDDA_2.n308 VDDA_2.n23 3.4105
R19760 VDDA_2.n308 VDDA_2.n9 3.4105
R19761 VDDA_2.n308 VDDA_2.n24 3.4105
R19762 VDDA_2.n308 VDDA_2.n8 3.4105
R19763 VDDA_2.n308 VDDA_2.n25 3.4105
R19764 VDDA_2.n308 VDDA_2.n7 3.4105
R19765 VDDA_2.n308 VDDA_2.n26 3.4105
R19766 VDDA_2.n308 VDDA_2.n6 3.4105
R19767 VDDA_2.n308 VDDA_2.n27 3.4105
R19768 VDDA_2.n308 VDDA_2.n5 3.4105
R19769 VDDA_2.n308 VDDA_2.n28 3.4105
R19770 VDDA_2.n308 VDDA_2.n4 3.4105
R19771 VDDA_2.n308 VDDA_2.n29 3.4105
R19772 VDDA_2.n308 VDDA_2.n3 3.4105
R19773 VDDA_2.n308 VDDA_2.n30 3.4105
R19774 VDDA_2.n308 VDDA_2.n2 3.4105
R19775 VDDA_2.n308 VDDA_2.n31 3.4105
R19776 VDDA_2.n308 VDDA_2.n1 3.4105
R19777 VDDA_2.n308 VDDA_2.n32 3.4105
R19778 VDDA_2.n336 VDDA_2.n308 3.4105
R19779 VDDA_2.n317 VDDA_2.n241 3.4105
R19780 VDDA_2.n241 VDDA_2.n17 3.4105
R19781 VDDA_2.n241 VDDA_2.n15 3.4105
R19782 VDDA_2.n241 VDDA_2.n18 3.4105
R19783 VDDA_2.n241 VDDA_2.n14 3.4105
R19784 VDDA_2.n241 VDDA_2.n19 3.4105
R19785 VDDA_2.n241 VDDA_2.n13 3.4105
R19786 VDDA_2.n241 VDDA_2.n20 3.4105
R19787 VDDA_2.n241 VDDA_2.n12 3.4105
R19788 VDDA_2.n241 VDDA_2.n21 3.4105
R19789 VDDA_2.n241 VDDA_2.n11 3.4105
R19790 VDDA_2.n241 VDDA_2.n22 3.4105
R19791 VDDA_2.n241 VDDA_2.n10 3.4105
R19792 VDDA_2.n241 VDDA_2.n23 3.4105
R19793 VDDA_2.n241 VDDA_2.n9 3.4105
R19794 VDDA_2.n241 VDDA_2.n24 3.4105
R19795 VDDA_2.n241 VDDA_2.n8 3.4105
R19796 VDDA_2.n241 VDDA_2.n25 3.4105
R19797 VDDA_2.n241 VDDA_2.n7 3.4105
R19798 VDDA_2.n241 VDDA_2.n26 3.4105
R19799 VDDA_2.n241 VDDA_2.n6 3.4105
R19800 VDDA_2.n241 VDDA_2.n27 3.4105
R19801 VDDA_2.n241 VDDA_2.n5 3.4105
R19802 VDDA_2.n241 VDDA_2.n28 3.4105
R19803 VDDA_2.n241 VDDA_2.n4 3.4105
R19804 VDDA_2.n241 VDDA_2.n29 3.4105
R19805 VDDA_2.n241 VDDA_2.n3 3.4105
R19806 VDDA_2.n241 VDDA_2.n30 3.4105
R19807 VDDA_2.n241 VDDA_2.n2 3.4105
R19808 VDDA_2.n241 VDDA_2.n31 3.4105
R19809 VDDA_2.n241 VDDA_2.n1 3.4105
R19810 VDDA_2.n241 VDDA_2.n32 3.4105
R19811 VDDA_2.n336 VDDA_2.n241 3.4105
R19812 VDDA_2.n317 VDDA_2.n310 3.4105
R19813 VDDA_2.n310 VDDA_2.n17 3.4105
R19814 VDDA_2.n310 VDDA_2.n15 3.4105
R19815 VDDA_2.n310 VDDA_2.n18 3.4105
R19816 VDDA_2.n310 VDDA_2.n14 3.4105
R19817 VDDA_2.n310 VDDA_2.n19 3.4105
R19818 VDDA_2.n310 VDDA_2.n13 3.4105
R19819 VDDA_2.n310 VDDA_2.n20 3.4105
R19820 VDDA_2.n310 VDDA_2.n12 3.4105
R19821 VDDA_2.n310 VDDA_2.n21 3.4105
R19822 VDDA_2.n310 VDDA_2.n11 3.4105
R19823 VDDA_2.n310 VDDA_2.n22 3.4105
R19824 VDDA_2.n310 VDDA_2.n10 3.4105
R19825 VDDA_2.n310 VDDA_2.n23 3.4105
R19826 VDDA_2.n310 VDDA_2.n9 3.4105
R19827 VDDA_2.n310 VDDA_2.n24 3.4105
R19828 VDDA_2.n310 VDDA_2.n8 3.4105
R19829 VDDA_2.n310 VDDA_2.n25 3.4105
R19830 VDDA_2.n310 VDDA_2.n7 3.4105
R19831 VDDA_2.n310 VDDA_2.n26 3.4105
R19832 VDDA_2.n310 VDDA_2.n6 3.4105
R19833 VDDA_2.n310 VDDA_2.n27 3.4105
R19834 VDDA_2.n310 VDDA_2.n5 3.4105
R19835 VDDA_2.n310 VDDA_2.n28 3.4105
R19836 VDDA_2.n310 VDDA_2.n4 3.4105
R19837 VDDA_2.n310 VDDA_2.n29 3.4105
R19838 VDDA_2.n310 VDDA_2.n3 3.4105
R19839 VDDA_2.n310 VDDA_2.n30 3.4105
R19840 VDDA_2.n310 VDDA_2.n2 3.4105
R19841 VDDA_2.n310 VDDA_2.n31 3.4105
R19842 VDDA_2.n310 VDDA_2.n1 3.4105
R19843 VDDA_2.n310 VDDA_2.n32 3.4105
R19844 VDDA_2.n336 VDDA_2.n310 3.4105
R19845 VDDA_2.n317 VDDA_2.n240 3.4105
R19846 VDDA_2.n240 VDDA_2.n17 3.4105
R19847 VDDA_2.n240 VDDA_2.n15 3.4105
R19848 VDDA_2.n240 VDDA_2.n18 3.4105
R19849 VDDA_2.n240 VDDA_2.n14 3.4105
R19850 VDDA_2.n240 VDDA_2.n19 3.4105
R19851 VDDA_2.n240 VDDA_2.n13 3.4105
R19852 VDDA_2.n240 VDDA_2.n20 3.4105
R19853 VDDA_2.n240 VDDA_2.n12 3.4105
R19854 VDDA_2.n240 VDDA_2.n21 3.4105
R19855 VDDA_2.n240 VDDA_2.n11 3.4105
R19856 VDDA_2.n240 VDDA_2.n22 3.4105
R19857 VDDA_2.n240 VDDA_2.n10 3.4105
R19858 VDDA_2.n240 VDDA_2.n23 3.4105
R19859 VDDA_2.n240 VDDA_2.n9 3.4105
R19860 VDDA_2.n240 VDDA_2.n24 3.4105
R19861 VDDA_2.n240 VDDA_2.n8 3.4105
R19862 VDDA_2.n240 VDDA_2.n25 3.4105
R19863 VDDA_2.n240 VDDA_2.n7 3.4105
R19864 VDDA_2.n240 VDDA_2.n26 3.4105
R19865 VDDA_2.n240 VDDA_2.n6 3.4105
R19866 VDDA_2.n240 VDDA_2.n27 3.4105
R19867 VDDA_2.n240 VDDA_2.n5 3.4105
R19868 VDDA_2.n240 VDDA_2.n28 3.4105
R19869 VDDA_2.n240 VDDA_2.n4 3.4105
R19870 VDDA_2.n240 VDDA_2.n29 3.4105
R19871 VDDA_2.n240 VDDA_2.n3 3.4105
R19872 VDDA_2.n240 VDDA_2.n30 3.4105
R19873 VDDA_2.n240 VDDA_2.n2 3.4105
R19874 VDDA_2.n240 VDDA_2.n31 3.4105
R19875 VDDA_2.n240 VDDA_2.n1 3.4105
R19876 VDDA_2.n240 VDDA_2.n32 3.4105
R19877 VDDA_2.n336 VDDA_2.n240 3.4105
R19878 VDDA_2.n317 VDDA_2.n312 3.4105
R19879 VDDA_2.n312 VDDA_2.n17 3.4105
R19880 VDDA_2.n312 VDDA_2.n15 3.4105
R19881 VDDA_2.n312 VDDA_2.n18 3.4105
R19882 VDDA_2.n312 VDDA_2.n14 3.4105
R19883 VDDA_2.n312 VDDA_2.n19 3.4105
R19884 VDDA_2.n312 VDDA_2.n13 3.4105
R19885 VDDA_2.n312 VDDA_2.n20 3.4105
R19886 VDDA_2.n312 VDDA_2.n12 3.4105
R19887 VDDA_2.n312 VDDA_2.n21 3.4105
R19888 VDDA_2.n312 VDDA_2.n11 3.4105
R19889 VDDA_2.n312 VDDA_2.n22 3.4105
R19890 VDDA_2.n312 VDDA_2.n10 3.4105
R19891 VDDA_2.n312 VDDA_2.n23 3.4105
R19892 VDDA_2.n312 VDDA_2.n9 3.4105
R19893 VDDA_2.n312 VDDA_2.n24 3.4105
R19894 VDDA_2.n312 VDDA_2.n8 3.4105
R19895 VDDA_2.n312 VDDA_2.n25 3.4105
R19896 VDDA_2.n312 VDDA_2.n7 3.4105
R19897 VDDA_2.n312 VDDA_2.n26 3.4105
R19898 VDDA_2.n312 VDDA_2.n6 3.4105
R19899 VDDA_2.n312 VDDA_2.n27 3.4105
R19900 VDDA_2.n312 VDDA_2.n5 3.4105
R19901 VDDA_2.n312 VDDA_2.n28 3.4105
R19902 VDDA_2.n312 VDDA_2.n4 3.4105
R19903 VDDA_2.n312 VDDA_2.n29 3.4105
R19904 VDDA_2.n312 VDDA_2.n3 3.4105
R19905 VDDA_2.n312 VDDA_2.n30 3.4105
R19906 VDDA_2.n312 VDDA_2.n2 3.4105
R19907 VDDA_2.n312 VDDA_2.n31 3.4105
R19908 VDDA_2.n312 VDDA_2.n1 3.4105
R19909 VDDA_2.n312 VDDA_2.n32 3.4105
R19910 VDDA_2.n336 VDDA_2.n312 3.4105
R19911 VDDA_2.n317 VDDA_2.n239 3.4105
R19912 VDDA_2.n239 VDDA_2.n17 3.4105
R19913 VDDA_2.n239 VDDA_2.n15 3.4105
R19914 VDDA_2.n239 VDDA_2.n18 3.4105
R19915 VDDA_2.n239 VDDA_2.n14 3.4105
R19916 VDDA_2.n239 VDDA_2.n19 3.4105
R19917 VDDA_2.n239 VDDA_2.n13 3.4105
R19918 VDDA_2.n239 VDDA_2.n20 3.4105
R19919 VDDA_2.n239 VDDA_2.n12 3.4105
R19920 VDDA_2.n239 VDDA_2.n21 3.4105
R19921 VDDA_2.n239 VDDA_2.n11 3.4105
R19922 VDDA_2.n239 VDDA_2.n22 3.4105
R19923 VDDA_2.n239 VDDA_2.n10 3.4105
R19924 VDDA_2.n239 VDDA_2.n23 3.4105
R19925 VDDA_2.n239 VDDA_2.n9 3.4105
R19926 VDDA_2.n239 VDDA_2.n24 3.4105
R19927 VDDA_2.n239 VDDA_2.n8 3.4105
R19928 VDDA_2.n239 VDDA_2.n25 3.4105
R19929 VDDA_2.n239 VDDA_2.n7 3.4105
R19930 VDDA_2.n239 VDDA_2.n26 3.4105
R19931 VDDA_2.n239 VDDA_2.n6 3.4105
R19932 VDDA_2.n239 VDDA_2.n27 3.4105
R19933 VDDA_2.n239 VDDA_2.n5 3.4105
R19934 VDDA_2.n239 VDDA_2.n28 3.4105
R19935 VDDA_2.n239 VDDA_2.n4 3.4105
R19936 VDDA_2.n239 VDDA_2.n29 3.4105
R19937 VDDA_2.n239 VDDA_2.n3 3.4105
R19938 VDDA_2.n239 VDDA_2.n30 3.4105
R19939 VDDA_2.n239 VDDA_2.n2 3.4105
R19940 VDDA_2.n239 VDDA_2.n31 3.4105
R19941 VDDA_2.n239 VDDA_2.n1 3.4105
R19942 VDDA_2.n239 VDDA_2.n32 3.4105
R19943 VDDA_2.n336 VDDA_2.n239 3.4105
R19944 VDDA_2.n317 VDDA_2.n314 3.4105
R19945 VDDA_2.n314 VDDA_2.n17 3.4105
R19946 VDDA_2.n314 VDDA_2.n15 3.4105
R19947 VDDA_2.n314 VDDA_2.n18 3.4105
R19948 VDDA_2.n314 VDDA_2.n14 3.4105
R19949 VDDA_2.n314 VDDA_2.n19 3.4105
R19950 VDDA_2.n314 VDDA_2.n13 3.4105
R19951 VDDA_2.n314 VDDA_2.n20 3.4105
R19952 VDDA_2.n314 VDDA_2.n12 3.4105
R19953 VDDA_2.n314 VDDA_2.n21 3.4105
R19954 VDDA_2.n314 VDDA_2.n11 3.4105
R19955 VDDA_2.n314 VDDA_2.n22 3.4105
R19956 VDDA_2.n314 VDDA_2.n10 3.4105
R19957 VDDA_2.n314 VDDA_2.n23 3.4105
R19958 VDDA_2.n314 VDDA_2.n9 3.4105
R19959 VDDA_2.n314 VDDA_2.n24 3.4105
R19960 VDDA_2.n314 VDDA_2.n8 3.4105
R19961 VDDA_2.n314 VDDA_2.n25 3.4105
R19962 VDDA_2.n314 VDDA_2.n7 3.4105
R19963 VDDA_2.n314 VDDA_2.n26 3.4105
R19964 VDDA_2.n314 VDDA_2.n6 3.4105
R19965 VDDA_2.n314 VDDA_2.n27 3.4105
R19966 VDDA_2.n314 VDDA_2.n5 3.4105
R19967 VDDA_2.n314 VDDA_2.n28 3.4105
R19968 VDDA_2.n314 VDDA_2.n4 3.4105
R19969 VDDA_2.n314 VDDA_2.n29 3.4105
R19970 VDDA_2.n314 VDDA_2.n3 3.4105
R19971 VDDA_2.n314 VDDA_2.n30 3.4105
R19972 VDDA_2.n314 VDDA_2.n2 3.4105
R19973 VDDA_2.n314 VDDA_2.n31 3.4105
R19974 VDDA_2.n314 VDDA_2.n1 3.4105
R19975 VDDA_2.n314 VDDA_2.n32 3.4105
R19976 VDDA_2.n336 VDDA_2.n314 3.4105
R19977 VDDA_2.n317 VDDA_2.n238 3.4105
R19978 VDDA_2.n238 VDDA_2.n17 3.4105
R19979 VDDA_2.n238 VDDA_2.n15 3.4105
R19980 VDDA_2.n238 VDDA_2.n18 3.4105
R19981 VDDA_2.n238 VDDA_2.n14 3.4105
R19982 VDDA_2.n238 VDDA_2.n19 3.4105
R19983 VDDA_2.n238 VDDA_2.n13 3.4105
R19984 VDDA_2.n238 VDDA_2.n20 3.4105
R19985 VDDA_2.n238 VDDA_2.n12 3.4105
R19986 VDDA_2.n238 VDDA_2.n21 3.4105
R19987 VDDA_2.n238 VDDA_2.n11 3.4105
R19988 VDDA_2.n238 VDDA_2.n22 3.4105
R19989 VDDA_2.n238 VDDA_2.n10 3.4105
R19990 VDDA_2.n238 VDDA_2.n23 3.4105
R19991 VDDA_2.n238 VDDA_2.n9 3.4105
R19992 VDDA_2.n238 VDDA_2.n24 3.4105
R19993 VDDA_2.n238 VDDA_2.n8 3.4105
R19994 VDDA_2.n238 VDDA_2.n25 3.4105
R19995 VDDA_2.n238 VDDA_2.n7 3.4105
R19996 VDDA_2.n238 VDDA_2.n26 3.4105
R19997 VDDA_2.n238 VDDA_2.n6 3.4105
R19998 VDDA_2.n238 VDDA_2.n27 3.4105
R19999 VDDA_2.n238 VDDA_2.n5 3.4105
R20000 VDDA_2.n238 VDDA_2.n28 3.4105
R20001 VDDA_2.n238 VDDA_2.n4 3.4105
R20002 VDDA_2.n238 VDDA_2.n29 3.4105
R20003 VDDA_2.n238 VDDA_2.n3 3.4105
R20004 VDDA_2.n238 VDDA_2.n30 3.4105
R20005 VDDA_2.n238 VDDA_2.n2 3.4105
R20006 VDDA_2.n238 VDDA_2.n31 3.4105
R20007 VDDA_2.n238 VDDA_2.n1 3.4105
R20008 VDDA_2.n238 VDDA_2.n32 3.4105
R20009 VDDA_2.n336 VDDA_2.n238 3.4105
R20010 VDDA_2.n335 VDDA_2.n317 3.4105
R20011 VDDA_2.n335 VDDA_2.n17 3.4105
R20012 VDDA_2.n335 VDDA_2.n15 3.4105
R20013 VDDA_2.n335 VDDA_2.n18 3.4105
R20014 VDDA_2.n335 VDDA_2.n14 3.4105
R20015 VDDA_2.n335 VDDA_2.n19 3.4105
R20016 VDDA_2.n335 VDDA_2.n13 3.4105
R20017 VDDA_2.n335 VDDA_2.n20 3.4105
R20018 VDDA_2.n335 VDDA_2.n12 3.4105
R20019 VDDA_2.n335 VDDA_2.n21 3.4105
R20020 VDDA_2.n335 VDDA_2.n11 3.4105
R20021 VDDA_2.n335 VDDA_2.n22 3.4105
R20022 VDDA_2.n335 VDDA_2.n10 3.4105
R20023 VDDA_2.n335 VDDA_2.n23 3.4105
R20024 VDDA_2.n335 VDDA_2.n9 3.4105
R20025 VDDA_2.n335 VDDA_2.n24 3.4105
R20026 VDDA_2.n335 VDDA_2.n8 3.4105
R20027 VDDA_2.n335 VDDA_2.n25 3.4105
R20028 VDDA_2.n335 VDDA_2.n7 3.4105
R20029 VDDA_2.n335 VDDA_2.n26 3.4105
R20030 VDDA_2.n335 VDDA_2.n6 3.4105
R20031 VDDA_2.n335 VDDA_2.n27 3.4105
R20032 VDDA_2.n335 VDDA_2.n5 3.4105
R20033 VDDA_2.n335 VDDA_2.n28 3.4105
R20034 VDDA_2.n335 VDDA_2.n4 3.4105
R20035 VDDA_2.n335 VDDA_2.n29 3.4105
R20036 VDDA_2.n335 VDDA_2.n3 3.4105
R20037 VDDA_2.n335 VDDA_2.n30 3.4105
R20038 VDDA_2.n335 VDDA_2.n2 3.4105
R20039 VDDA_2.n335 VDDA_2.n31 3.4105
R20040 VDDA_2.n335 VDDA_2.n1 3.4105
R20041 VDDA_2.n335 VDDA_2.n32 3.4105
R20042 VDDA_2.n336 VDDA_2.n335 3.4105
R20043 VDDA_2.n317 VDDA_2.n237 3.4105
R20044 VDDA_2.n237 VDDA_2.n17 3.4105
R20045 VDDA_2.n237 VDDA_2.n15 3.4105
R20046 VDDA_2.n237 VDDA_2.n18 3.4105
R20047 VDDA_2.n237 VDDA_2.n14 3.4105
R20048 VDDA_2.n237 VDDA_2.n19 3.4105
R20049 VDDA_2.n237 VDDA_2.n13 3.4105
R20050 VDDA_2.n237 VDDA_2.n20 3.4105
R20051 VDDA_2.n237 VDDA_2.n12 3.4105
R20052 VDDA_2.n237 VDDA_2.n21 3.4105
R20053 VDDA_2.n237 VDDA_2.n11 3.4105
R20054 VDDA_2.n237 VDDA_2.n22 3.4105
R20055 VDDA_2.n237 VDDA_2.n10 3.4105
R20056 VDDA_2.n237 VDDA_2.n23 3.4105
R20057 VDDA_2.n237 VDDA_2.n9 3.4105
R20058 VDDA_2.n237 VDDA_2.n24 3.4105
R20059 VDDA_2.n237 VDDA_2.n8 3.4105
R20060 VDDA_2.n237 VDDA_2.n25 3.4105
R20061 VDDA_2.n237 VDDA_2.n7 3.4105
R20062 VDDA_2.n237 VDDA_2.n26 3.4105
R20063 VDDA_2.n237 VDDA_2.n6 3.4105
R20064 VDDA_2.n237 VDDA_2.n27 3.4105
R20065 VDDA_2.n237 VDDA_2.n5 3.4105
R20066 VDDA_2.n237 VDDA_2.n28 3.4105
R20067 VDDA_2.n237 VDDA_2.n4 3.4105
R20068 VDDA_2.n237 VDDA_2.n29 3.4105
R20069 VDDA_2.n237 VDDA_2.n3 3.4105
R20070 VDDA_2.n237 VDDA_2.n30 3.4105
R20071 VDDA_2.n237 VDDA_2.n2 3.4105
R20072 VDDA_2.n237 VDDA_2.n31 3.4105
R20073 VDDA_2.n237 VDDA_2.n1 3.4105
R20074 VDDA_2.n237 VDDA_2.n32 3.4105
R20075 VDDA_2.n336 VDDA_2.n237 3.4105
R20076 VDDA_2.n337 VDDA_2.n17 3.4105
R20077 VDDA_2.n337 VDDA_2.n15 3.4105
R20078 VDDA_2.n337 VDDA_2.n18 3.4105
R20079 VDDA_2.n337 VDDA_2.n14 3.4105
R20080 VDDA_2.n337 VDDA_2.n19 3.4105
R20081 VDDA_2.n337 VDDA_2.n13 3.4105
R20082 VDDA_2.n337 VDDA_2.n20 3.4105
R20083 VDDA_2.n337 VDDA_2.n12 3.4105
R20084 VDDA_2.n337 VDDA_2.n21 3.4105
R20085 VDDA_2.n337 VDDA_2.n11 3.4105
R20086 VDDA_2.n337 VDDA_2.n22 3.4105
R20087 VDDA_2.n337 VDDA_2.n10 3.4105
R20088 VDDA_2.n337 VDDA_2.n23 3.4105
R20089 VDDA_2.n337 VDDA_2.n9 3.4105
R20090 VDDA_2.n337 VDDA_2.n24 3.4105
R20091 VDDA_2.n337 VDDA_2.n8 3.4105
R20092 VDDA_2.n337 VDDA_2.n25 3.4105
R20093 VDDA_2.n337 VDDA_2.n7 3.4105
R20094 VDDA_2.n337 VDDA_2.n26 3.4105
R20095 VDDA_2.n337 VDDA_2.n6 3.4105
R20096 VDDA_2.n337 VDDA_2.n27 3.4105
R20097 VDDA_2.n337 VDDA_2.n5 3.4105
R20098 VDDA_2.n337 VDDA_2.n28 3.4105
R20099 VDDA_2.n337 VDDA_2.n4 3.4105
R20100 VDDA_2.n337 VDDA_2.n29 3.4105
R20101 VDDA_2.n337 VDDA_2.n3 3.4105
R20102 VDDA_2.n337 VDDA_2.n30 3.4105
R20103 VDDA_2.n337 VDDA_2.n2 3.4105
R20104 VDDA_2.n337 VDDA_2.n31 3.4105
R20105 VDDA_2.n337 VDDA_2.n1 3.4105
R20106 VDDA_2.n337 VDDA_2.n32 3.4105
R20107 VDDA_2.n337 VDDA_2.n336 3.4105
R20108 VDDA_2.n126 VDDA_2.n125 2.426
R20109 VDDA_2.n188 VDDA_2.n187 2.2505
R20110 VDDA_2.n189 VDDA_2.n69 2.2505
R20111 VDDA_2.n191 VDDA_2.n190 2.2505
R20112 VDDA_2.n192 VDDA_2.n68 2.2505
R20113 VDDA_2.n197 VDDA_2.n196 2.2505
R20114 VDDA_2.n198 VDDA_2.n64 2.2505
R20115 VDDA_2.n200 VDDA_2.n199 2.2505
R20116 VDDA_2.n201 VDDA_2.n63 2.2505
R20117 VDDA_2.n206 VDDA_2.n205 2.2505
R20118 VDDA_2.n207 VDDA_2.n59 2.2505
R20119 VDDA_2.n209 VDDA_2.n208 2.2505
R20120 VDDA_2.n210 VDDA_2.n58 2.2505
R20121 VDDA_2.n215 VDDA_2.n214 2.2505
R20122 VDDA_2.n216 VDDA_2.n54 2.2505
R20123 VDDA_2.n218 VDDA_2.n217 2.2505
R20124 VDDA_2.n219 VDDA_2.n53 2.2505
R20125 VDDA_2.n224 VDDA_2.n223 2.2505
R20126 VDDA_2.n225 VDDA_2.n49 2.2505
R20127 VDDA_2.n227 VDDA_2.n226 2.2505
R20128 VDDA_2.n228 VDDA_2.n48 2.2505
R20129 VDDA_2.n233 VDDA_2.n232 2.2505
R20130 VDDA_2.n235 VDDA_2.n234 1.74133
R20131 VDDA_2.n270 VDDA_2.n269 1.70567
R20132 VDDA_2.n333 VDDA_2.n332 1.70567
R20133 VDDA_2.n287 VDDA_2.n269 1.70567
R20134 VDDA_2.n333 VDDA_2.n331 1.70567
R20135 VDDA_2.n289 VDDA_2.n269 1.70567
R20136 VDDA_2.n333 VDDA_2.n330 1.70567
R20137 VDDA_2.n291 VDDA_2.n269 1.70567
R20138 VDDA_2.n333 VDDA_2.n329 1.70567
R20139 VDDA_2.n293 VDDA_2.n269 1.70567
R20140 VDDA_2.n333 VDDA_2.n328 1.70567
R20141 VDDA_2.n295 VDDA_2.n269 1.70567
R20142 VDDA_2.n333 VDDA_2.n327 1.70567
R20143 VDDA_2.n297 VDDA_2.n269 1.70567
R20144 VDDA_2.n333 VDDA_2.n326 1.70567
R20145 VDDA_2.n299 VDDA_2.n269 1.70567
R20146 VDDA_2.n333 VDDA_2.n325 1.70567
R20147 VDDA_2.n301 VDDA_2.n269 1.70567
R20148 VDDA_2.n333 VDDA_2.n324 1.70567
R20149 VDDA_2.n303 VDDA_2.n269 1.70567
R20150 VDDA_2.n333 VDDA_2.n323 1.70567
R20151 VDDA_2.n305 VDDA_2.n269 1.70567
R20152 VDDA_2.n333 VDDA_2.n322 1.70567
R20153 VDDA_2.n307 VDDA_2.n269 1.70567
R20154 VDDA_2.n333 VDDA_2.n321 1.70567
R20155 VDDA_2.n309 VDDA_2.n269 1.70567
R20156 VDDA_2.n333 VDDA_2.n320 1.70567
R20157 VDDA_2.n311 VDDA_2.n269 1.70567
R20158 VDDA_2.n333 VDDA_2.n319 1.70567
R20159 VDDA_2.n313 VDDA_2.n269 1.70567
R20160 VDDA_2.n333 VDDA_2.n318 1.70567
R20161 VDDA_2.n315 VDDA_2.n269 1.70567
R20162 VDDA_2.n334 VDDA_2.n333 1.70567
R20163 VDDA_2.n269 VDDA_2.n0 1.70567
R20164 VDDA_2.n268 VDDA_2.n267 1.70566
R20165 VDDA_2.n268 VDDA_2.n266 1.70566
R20166 VDDA_2.n268 VDDA_2.n265 1.70566
R20167 VDDA_2.n268 VDDA_2.n264 1.70566
R20168 VDDA_2.n268 VDDA_2.n263 1.70566
R20169 VDDA_2.n268 VDDA_2.n262 1.70566
R20170 VDDA_2.n268 VDDA_2.n261 1.70566
R20171 VDDA_2.n268 VDDA_2.n260 1.70566
R20172 VDDA_2.n268 VDDA_2.n259 1.70566
R20173 VDDA_2.n268 VDDA_2.n258 1.70566
R20174 VDDA_2.n268 VDDA_2.n257 1.70566
R20175 VDDA_2.n268 VDDA_2.n256 1.70566
R20176 VDDA_2.n268 VDDA_2.n255 1.70566
R20177 VDDA_2.n268 VDDA_2.n254 1.70566
R20178 VDDA_2.n268 VDDA_2.n253 1.70566
R20179 VDDA_2.n316 VDDA_2.n286 1.70566
R20180 VDDA_2.n286 VDDA_2.n285 1.70566
R20181 VDDA_2.n286 VDDA_2.n284 1.70566
R20182 VDDA_2.n286 VDDA_2.n283 1.70566
R20183 VDDA_2.n286 VDDA_2.n282 1.70566
R20184 VDDA_2.n286 VDDA_2.n281 1.70566
R20185 VDDA_2.n286 VDDA_2.n280 1.70566
R20186 VDDA_2.n286 VDDA_2.n279 1.70566
R20187 VDDA_2.n286 VDDA_2.n278 1.70566
R20188 VDDA_2.n286 VDDA_2.n277 1.70566
R20189 VDDA_2.n286 VDDA_2.n276 1.70566
R20190 VDDA_2.n286 VDDA_2.n275 1.70566
R20191 VDDA_2.n286 VDDA_2.n274 1.70566
R20192 VDDA_2.n286 VDDA_2.n273 1.70566
R20193 VDDA_2.n286 VDDA_2.n272 1.70566
R20194 VDDA_2.n286 VDDA_2.n271 1.70566
R20195 VDDA_2.n337 VDDA_2.n16 1.70566
R20196 VDDA_2.n47 VDDA_2.n46 1.7055
R20197 VDDA_2.n232 VDDA_2.n231 1.7055
R20198 VDDA_2.n229 VDDA_2.n228 1.7055
R20199 VDDA_2.n227 VDDA_2.n52 1.7055
R20200 VDDA_2.n50 VDDA_2.n49 1.7055
R20201 VDDA_2.n223 VDDA_2.n222 1.7055
R20202 VDDA_2.n220 VDDA_2.n219 1.7055
R20203 VDDA_2.n218 VDDA_2.n57 1.7055
R20204 VDDA_2.n55 VDDA_2.n54 1.7055
R20205 VDDA_2.n214 VDDA_2.n213 1.7055
R20206 VDDA_2.n211 VDDA_2.n210 1.7055
R20207 VDDA_2.n209 VDDA_2.n62 1.7055
R20208 VDDA_2.n60 VDDA_2.n59 1.7055
R20209 VDDA_2.n205 VDDA_2.n204 1.7055
R20210 VDDA_2.n202 VDDA_2.n201 1.7055
R20211 VDDA_2.n200 VDDA_2.n67 1.7055
R20212 VDDA_2.n65 VDDA_2.n64 1.7055
R20213 VDDA_2.n196 VDDA_2.n195 1.7055
R20214 VDDA_2.n193 VDDA_2.n192 1.7055
R20215 VDDA_2.n191 VDDA_2.n72 1.7055
R20216 VDDA_2.n70 VDDA_2.n69 1.7055
R20217 VDDA_2.n187 VDDA_2.n186 1.7055
R20218 VDDA_2.n236 VDDA_2.n36 1.69989
R20219 VDDA_2.n236 VDDA_2.n39 1.69989
R20220 VDDA_2.n236 VDDA_2.n42 1.69989
R20221 VDDA_2.n51 VDDA_2.n33 1.69938
R20222 VDDA_2.n221 VDDA_2.n33 1.69938
R20223 VDDA_2.n212 VDDA_2.n33 1.69938
R20224 VDDA_2.n61 VDDA_2.n33 1.69938
R20225 VDDA_2.n66 VDDA_2.n33 1.69938
R20226 VDDA_2.n194 VDDA_2.n33 1.69938
R20227 VDDA_2.n45 VDDA_2.n33 1.69938
R20228 VDDA_2.n236 VDDA_2.n34 1.69888
R20229 VDDA_2.n230 VDDA_2.n33 1.69888
R20230 VDDA_2.n236 VDDA_2.n35 1.69888
R20231 VDDA_2.n236 VDDA_2.n37 1.69888
R20232 VDDA_2.n56 VDDA_2.n33 1.69888
R20233 VDDA_2.n236 VDDA_2.n38 1.69888
R20234 VDDA_2.n236 VDDA_2.n40 1.69888
R20235 VDDA_2.n203 VDDA_2.n33 1.69888
R20236 VDDA_2.n236 VDDA_2.n41 1.69888
R20237 VDDA_2.n236 VDDA_2.n43 1.69888
R20238 VDDA_2.n71 VDDA_2.n33 1.69888
R20239 VDDA_2.n236 VDDA_2.n44 1.69888
R20240 VDDA_2.n135 VDDA_2.n86 1.69202
R20241 VDDA_2.n144 VDDA_2.n86 1.69202
R20242 VDDA_2.n153 VDDA_2.n86 1.69202
R20243 VDDA_2.n129 VDDA_2.n86 1.68971
R20244 VDDA_2.n132 VDDA_2.n86 1.68971
R20245 VDDA_2.n138 VDDA_2.n86 1.68971
R20246 VDDA_2.n141 VDDA_2.n86 1.68971
R20247 VDDA_2.n147 VDDA_2.n86 1.68971
R20248 VDDA_2.n150 VDDA_2.n86 1.68971
R20249 VDDA_2.n156 VDDA_2.n86 1.68971
R20250 VDDA_2.n159 VDDA_2.n86 1.68971
R20251 VDDA_2.n162 VDDA_2.n75 1.56177
R20252 VDDA_2.n184 VDDA_2.n75 1.50969
R20253 VDDA_2.n75 VDDA_2.n74 1.44719
R20254 VDDA_2.n336 VDDA_2.n236 1.22957
R20255 VDDA_2.n234 VDDA_2.n233 1.20209
R20256 VDDA_2.n183 VDDA_2.n182 0.229667
R20257 VDDA_2.n164 VDDA_2.n163 0.229667
R20258 VDDA_2.n178 VDDA_2.n177 0.208833
R20259 VDDA_2.n178 VDDA_2.n76 0.208833
R20260 VDDA_2.n182 VDDA_2.n76 0.208833
R20261 VDDA_2.n169 VDDA_2.n82 0.208833
R20262 VDDA_2.n165 VDDA_2.n82 0.208833
R20263 VDDA_2.n165 VDDA_2.n164 0.208833
R20264 VDDA_2.n161 VDDA_2.n84 0.1755
R20265 VDDA_2.n107 VDDA_2.n84 0.1755
R20266 VDDA_2.n108 VDDA_2.n107 0.1755
R20267 VDDA_2.n112 VDDA_2.n111 0.1755
R20268 VDDA_2.n113 VDDA_2.n112 0.1755
R20269 VDDA_2.n114 VDDA_2.n113 0.1755
R20270 VDDA_2.n118 VDDA_2.n117 0.1755
R20271 VDDA_2.n119 VDDA_2.n118 0.1755
R20272 VDDA_2.n120 VDDA_2.n119 0.1755
R20273 VDDA_2.n124 VDDA_2.n123 0.1755
R20274 VDDA_2.n125 VDDA_2.n124 0.1755
R20275 VDDA_2.n160 VDDA_2.n85 0.1755
R20276 VDDA_2.n87 VDDA_2.n85 0.1755
R20277 VDDA_2.n88 VDDA_2.n87 0.1755
R20278 VDDA_2.n92 VDDA_2.n91 0.1755
R20279 VDDA_2.n93 VDDA_2.n92 0.1755
R20280 VDDA_2.n94 VDDA_2.n93 0.1755
R20281 VDDA_2.n98 VDDA_2.n97 0.1755
R20282 VDDA_2.n99 VDDA_2.n98 0.1755
R20283 VDDA_2.n100 VDDA_2.n99 0.1755
R20284 VDDA_2.n104 VDDA_2.n103 0.1755
R20285 VDDA_2.n105 VDDA_2.n104 0.1755
R20286 VDDA_2.n106 VDDA_2.n105 0.1755
R20287 VDDA_2.n109 VDDA_2.n108 0.163
R20288 VDDA_2.n111 VDDA_2.n110 0.163
R20289 VDDA_2.n115 VDDA_2.n114 0.163
R20290 VDDA_2.n117 VDDA_2.n116 0.163
R20291 VDDA_2.n121 VDDA_2.n120 0.163
R20292 VDDA_2.n123 VDDA_2.n122 0.163
R20293 VDDA_2.n89 VDDA_2.n88 0.163
R20294 VDDA_2.n91 VDDA_2.n90 0.163
R20295 VDDA_2.n95 VDDA_2.n94 0.163
R20296 VDDA_2.n97 VDDA_2.n96 0.163
R20297 VDDA_2.n101 VDDA_2.n100 0.163
R20298 VDDA_2.n103 VDDA_2.n102 0.163
R20299 VDDA_2.n110 VDDA_2.n109 0.1505
R20300 VDDA_2.n116 VDDA_2.n115 0.1505
R20301 VDDA_2.n122 VDDA_2.n121 0.1505
R20302 VDDA_2.n90 VDDA_2.n89 0.1505
R20303 VDDA_2.n96 VDDA_2.n95 0.1505
R20304 VDDA_2.n102 VDDA_2.n101 0.1505
R20305 VDDA_2.n184 VDDA_2.n183 0.123287
R20306 VDDA_2.n163 VDDA_2.n162 0.123287
R20307 VDDA_2.n126 VDDA_2.n106 0.0794182
R20308 VDDA_2.n187 VDDA_2.n69 0.076587
R20309 VDDA_2.n191 VDDA_2.n69 0.076587
R20310 VDDA_2.n192 VDDA_2.n191 0.076587
R20311 VDDA_2.n201 VDDA_2.n200 0.076587
R20312 VDDA_2.n205 VDDA_2.n201 0.076587
R20313 VDDA_2.n205 VDDA_2.n59 0.076587
R20314 VDDA_2.n214 VDDA_2.n54 0.076587
R20315 VDDA_2.n218 VDDA_2.n54 0.076587
R20316 VDDA_2.n219 VDDA_2.n218 0.076587
R20317 VDDA_2.n228 VDDA_2.n227 0.076587
R20318 VDDA_2.n232 VDDA_2.n228 0.076587
R20319 VDDA_2.n232 VDDA_2.n47 0.076587
R20320 VDDA_2.n189 VDDA_2.n188 0.076587
R20321 VDDA_2.n190 VDDA_2.n189 0.076587
R20322 VDDA_2.n190 VDDA_2.n68 0.076587
R20323 VDDA_2.n199 VDDA_2.n63 0.076587
R20324 VDDA_2.n206 VDDA_2.n63 0.076587
R20325 VDDA_2.n207 VDDA_2.n206 0.076587
R20326 VDDA_2.n216 VDDA_2.n215 0.076587
R20327 VDDA_2.n217 VDDA_2.n216 0.076587
R20328 VDDA_2.n217 VDDA_2.n53 0.076587
R20329 VDDA_2.n226 VDDA_2.n48 0.076587
R20330 VDDA_2.n233 VDDA_2.n48 0.076587
R20331 VDDA_2.n196 VDDA_2.n192 0.0711522
R20332 VDDA_2.n200 VDDA_2.n64 0.0711522
R20333 VDDA_2.n209 VDDA_2.n59 0.0711522
R20334 VDDA_2.n214 VDDA_2.n210 0.0711522
R20335 VDDA_2.n223 VDDA_2.n219 0.0711522
R20336 VDDA_2.n227 VDDA_2.n49 0.0711522
R20337 VDDA_2.n197 VDDA_2.n68 0.0711522
R20338 VDDA_2.n199 VDDA_2.n198 0.0711522
R20339 VDDA_2.n208 VDDA_2.n207 0.0711522
R20340 VDDA_2.n215 VDDA_2.n58 0.0711522
R20341 VDDA_2.n224 VDDA_2.n53 0.0711522
R20342 VDDA_2.n226 VDDA_2.n225 0.0711522
R20343 VDDA_2.n158 VDDA_2.n157 0.0663
R20344 VDDA_2.n149 VDDA_2.n148 0.0663
R20345 VDDA_2.n140 VDDA_2.n139 0.0663
R20346 VDDA_2.n131 VDDA_2.n130 0.0663
R20347 VDDA_2.n196 VDDA_2.n64 0.0657174
R20348 VDDA_2.n210 VDDA_2.n209 0.0657174
R20349 VDDA_2.n223 VDDA_2.n49 0.0657174
R20350 VDDA_2.n198 VDDA_2.n197 0.0657174
R20351 VDDA_2.n208 VDDA_2.n58 0.0657174
R20352 VDDA_2.n225 VDDA_2.n224 0.0657174
R20353 VDDA_2.n155 VDDA_2.n154 0.0616
R20354 VDDA_2.n152 VDDA_2.n151 0.0616
R20355 VDDA_2.n146 VDDA_2.n145 0.0616
R20356 VDDA_2.n143 VDDA_2.n142 0.0616
R20357 VDDA_2.n137 VDDA_2.n136 0.0616
R20358 VDDA_2.n134 VDDA_2.n133 0.0616
R20359 VDDA_2.n128 VDDA_2.n127 0.0616
R20360 VDDA_2.n188 VDDA_2.n185 0.0439783
R20361 VDDA_2.n234 VDDA_2.n47 0.0352506
R20362 VDDA_2.n159 VDDA_2.n158 0.0335856
R20363 VDDA_2.n156 VDDA_2.n155 0.0335856
R20364 VDDA_2.n150 VDDA_2.n149 0.0335856
R20365 VDDA_2.n147 VDDA_2.n146 0.0335856
R20366 VDDA_2.n141 VDDA_2.n140 0.0335856
R20367 VDDA_2.n138 VDDA_2.n137 0.0335856
R20368 VDDA_2.n132 VDDA_2.n131 0.0335856
R20369 VDDA_2.n129 VDDA_2.n128 0.0335856
R20370 VDDA_2.n130 VDDA_2.n129 0.0335856
R20371 VDDA_2.n133 VDDA_2.n132 0.0335856
R20372 VDDA_2.n139 VDDA_2.n138 0.0335856
R20373 VDDA_2.n142 VDDA_2.n141 0.0335856
R20374 VDDA_2.n148 VDDA_2.n147 0.0335856
R20375 VDDA_2.n151 VDDA_2.n150 0.0335856
R20376 VDDA_2.n157 VDDA_2.n156 0.0335856
R20377 VDDA_2.n153 VDDA_2.n152 0.0289687
R20378 VDDA_2.n144 VDDA_2.n143 0.0289687
R20379 VDDA_2.n135 VDDA_2.n134 0.0289687
R20380 VDDA_2.n136 VDDA_2.n135 0.0289687
R20381 VDDA_2.n145 VDDA_2.n144 0.0289687
R20382 VDDA_2.n154 VDDA_2.n153 0.0289687
R20383 VDDA_2 VDDA_2.n337 0.0159953
R20384 VDDA_2.n70 VDDA_2.n44 0.0152446
R20385 VDDA_2.n72 VDDA_2.n71 0.0152446
R20386 VDDA_2.n193 VDDA_2.n43 0.0152446
R20387 VDDA_2.n202 VDDA_2.n41 0.0152446
R20388 VDDA_2.n204 VDDA_2.n203 0.0152446
R20389 VDDA_2.n60 VDDA_2.n40 0.0152446
R20390 VDDA_2.n55 VDDA_2.n38 0.0152446
R20391 VDDA_2.n57 VDDA_2.n56 0.0152446
R20392 VDDA_2.n220 VDDA_2.n37 0.0152446
R20393 VDDA_2.n229 VDDA_2.n35 0.0152446
R20394 VDDA_2.n231 VDDA_2.n230 0.0152446
R20395 VDDA_2.n46 VDDA_2.n34 0.0152446
R20396 VDDA_2.n231 VDDA_2.n34 0.0152446
R20397 VDDA_2.n230 VDDA_2.n229 0.0152446
R20398 VDDA_2.n52 VDDA_2.n35 0.0152446
R20399 VDDA_2.n57 VDDA_2.n37 0.0152446
R20400 VDDA_2.n56 VDDA_2.n55 0.0152446
R20401 VDDA_2.n213 VDDA_2.n38 0.0152446
R20402 VDDA_2.n204 VDDA_2.n40 0.0152446
R20403 VDDA_2.n203 VDDA_2.n202 0.0152446
R20404 VDDA_2.n67 VDDA_2.n41 0.0152446
R20405 VDDA_2.n72 VDDA_2.n43 0.0152446
R20406 VDDA_2.n71 VDDA_2.n70 0.0152446
R20407 VDDA_2.n186 VDDA_2.n44 0.0152446
R20408 VDDA_2.n195 VDDA_2.n194 0.0142311
R20409 VDDA_2.n67 VDDA_2.n66 0.0142311
R20410 VDDA_2.n62 VDDA_2.n61 0.0142311
R20411 VDDA_2.n213 VDDA_2.n212 0.0142311
R20412 VDDA_2.n222 VDDA_2.n221 0.0142311
R20413 VDDA_2.n52 VDDA_2.n51 0.0142311
R20414 VDDA_2.n235 VDDA_2.n45 0.0142311
R20415 VDDA_2.n46 VDDA_2.n45 0.0142311
R20416 VDDA_2.n51 VDDA_2.n50 0.0142311
R20417 VDDA_2.n221 VDDA_2.n220 0.0142311
R20418 VDDA_2.n212 VDDA_2.n211 0.0142311
R20419 VDDA_2.n61 VDDA_2.n60 0.0142311
R20420 VDDA_2.n66 VDDA_2.n65 0.0142311
R20421 VDDA_2.n194 VDDA_2.n193 0.0142311
R20422 VDDA_2.n65 VDDA_2.n42 0.0132169
R20423 VDDA_2.n211 VDDA_2.n39 0.0132169
R20424 VDDA_2.n50 VDDA_2.n36 0.0132169
R20425 VDDA_2.n222 VDDA_2.n36 0.0132169
R20426 VDDA_2.n62 VDDA_2.n39 0.0132169
R20427 VDDA_2.n195 VDDA_2.n42 0.0132169
R20428 VDDA_2.n86 VDDA_2.n33 0.00384628
R20429 VDDA_2.n236 VDDA_2.n33 0.00232524
R20430 VDDA_2.n336 VDDA_2.n269 0.00186893
R20431 VDDA_2.n269 VDDA_2.n32 0.00186893
R20432 VDDA_2.n271 VDDA_2.n1 0.00168433
R20433 VDDA_2.n253 VDDA_2.n1 0.00168433
R20434 VDDA_2.n272 VDDA_2.n2 0.00168433
R20435 VDDA_2.n254 VDDA_2.n2 0.00168433
R20436 VDDA_2.n273 VDDA_2.n3 0.00168433
R20437 VDDA_2.n255 VDDA_2.n3 0.00168433
R20438 VDDA_2.n274 VDDA_2.n4 0.00168433
R20439 VDDA_2.n256 VDDA_2.n4 0.00168433
R20440 VDDA_2.n275 VDDA_2.n5 0.00168433
R20441 VDDA_2.n257 VDDA_2.n5 0.00168433
R20442 VDDA_2.n276 VDDA_2.n6 0.00168433
R20443 VDDA_2.n258 VDDA_2.n6 0.00168433
R20444 VDDA_2.n277 VDDA_2.n7 0.00168433
R20445 VDDA_2.n259 VDDA_2.n7 0.00168433
R20446 VDDA_2.n278 VDDA_2.n8 0.00168433
R20447 VDDA_2.n260 VDDA_2.n8 0.00168433
R20448 VDDA_2.n279 VDDA_2.n9 0.00168433
R20449 VDDA_2.n261 VDDA_2.n9 0.00168433
R20450 VDDA_2.n280 VDDA_2.n10 0.00168433
R20451 VDDA_2.n262 VDDA_2.n10 0.00168433
R20452 VDDA_2.n281 VDDA_2.n11 0.00168433
R20453 VDDA_2.n263 VDDA_2.n11 0.00168433
R20454 VDDA_2.n282 VDDA_2.n12 0.00168433
R20455 VDDA_2.n264 VDDA_2.n12 0.00168433
R20456 VDDA_2.n283 VDDA_2.n13 0.00168433
R20457 VDDA_2.n265 VDDA_2.n13 0.00168433
R20458 VDDA_2.n284 VDDA_2.n14 0.00168433
R20459 VDDA_2.n266 VDDA_2.n14 0.00168433
R20460 VDDA_2.n285 VDDA_2.n15 0.00168433
R20461 VDDA_2.n267 VDDA_2.n15 0.00168433
R20462 VDDA_2.n317 VDDA_2.n316 0.00168433
R20463 VDDA_2.n333 VDDA_2.n16 0.00168433
R20464 VDDA_2.n267 VDDA_2.n17 0.00168433
R20465 VDDA_2.n266 VDDA_2.n18 0.00168433
R20466 VDDA_2.n265 VDDA_2.n19 0.00168433
R20467 VDDA_2.n264 VDDA_2.n20 0.00168433
R20468 VDDA_2.n263 VDDA_2.n21 0.00168433
R20469 VDDA_2.n262 VDDA_2.n22 0.00168433
R20470 VDDA_2.n261 VDDA_2.n23 0.00168433
R20471 VDDA_2.n260 VDDA_2.n24 0.00168433
R20472 VDDA_2.n259 VDDA_2.n25 0.00168433
R20473 VDDA_2.n258 VDDA_2.n26 0.00168433
R20474 VDDA_2.n257 VDDA_2.n27 0.00168433
R20475 VDDA_2.n256 VDDA_2.n28 0.00168433
R20476 VDDA_2.n255 VDDA_2.n29 0.00168433
R20477 VDDA_2.n254 VDDA_2.n30 0.00168433
R20478 VDDA_2.n253 VDDA_2.n31 0.00168433
R20479 VDDA_2.n316 VDDA_2.n17 0.00168433
R20480 VDDA_2.n285 VDDA_2.n18 0.00168433
R20481 VDDA_2.n284 VDDA_2.n19 0.00168433
R20482 VDDA_2.n283 VDDA_2.n20 0.00168433
R20483 VDDA_2.n282 VDDA_2.n21 0.00168433
R20484 VDDA_2.n281 VDDA_2.n22 0.00168433
R20485 VDDA_2.n280 VDDA_2.n23 0.00168433
R20486 VDDA_2.n279 VDDA_2.n24 0.00168433
R20487 VDDA_2.n278 VDDA_2.n25 0.00168433
R20488 VDDA_2.n277 VDDA_2.n26 0.00168433
R20489 VDDA_2.n276 VDDA_2.n27 0.00168433
R20490 VDDA_2.n275 VDDA_2.n28 0.00168433
R20491 VDDA_2.n274 VDDA_2.n29 0.00168433
R20492 VDDA_2.n273 VDDA_2.n30 0.00168433
R20493 VDDA_2.n272 VDDA_2.n31 0.00168433
R20494 VDDA_2.n271 VDDA_2.n32 0.00168433
R20495 VDDA_2.n317 VDDA_2.n16 0.00168433
R20496 VDDA_2.n286 VDDA_2.n270 0.00166081
R20497 VDDA_2.n332 VDDA_2.n252 0.00166081
R20498 VDDA_2.n288 VDDA_2.n287 0.00166081
R20499 VDDA_2.n331 VDDA_2.n251 0.00166081
R20500 VDDA_2.n290 VDDA_2.n289 0.00166081
R20501 VDDA_2.n330 VDDA_2.n250 0.00166081
R20502 VDDA_2.n292 VDDA_2.n291 0.00166081
R20503 VDDA_2.n329 VDDA_2.n249 0.00166081
R20504 VDDA_2.n294 VDDA_2.n293 0.00166081
R20505 VDDA_2.n328 VDDA_2.n248 0.00166081
R20506 VDDA_2.n296 VDDA_2.n295 0.00166081
R20507 VDDA_2.n327 VDDA_2.n247 0.00166081
R20508 VDDA_2.n298 VDDA_2.n297 0.00166081
R20509 VDDA_2.n326 VDDA_2.n246 0.00166081
R20510 VDDA_2.n300 VDDA_2.n299 0.00166081
R20511 VDDA_2.n325 VDDA_2.n245 0.00166081
R20512 VDDA_2.n302 VDDA_2.n301 0.00166081
R20513 VDDA_2.n324 VDDA_2.n244 0.00166081
R20514 VDDA_2.n304 VDDA_2.n303 0.00166081
R20515 VDDA_2.n323 VDDA_2.n243 0.00166081
R20516 VDDA_2.n306 VDDA_2.n305 0.00166081
R20517 VDDA_2.n322 VDDA_2.n242 0.00166081
R20518 VDDA_2.n308 VDDA_2.n307 0.00166081
R20519 VDDA_2.n321 VDDA_2.n241 0.00166081
R20520 VDDA_2.n310 VDDA_2.n309 0.00166081
R20521 VDDA_2.n320 VDDA_2.n240 0.00166081
R20522 VDDA_2.n312 VDDA_2.n311 0.00166081
R20523 VDDA_2.n319 VDDA_2.n239 0.00166081
R20524 VDDA_2.n314 VDDA_2.n313 0.00166081
R20525 VDDA_2.n318 VDDA_2.n238 0.00166081
R20526 VDDA_2.n335 VDDA_2.n315 0.00166081
R20527 VDDA_2.n334 VDDA_2.n237 0.00166081
R20528 VDDA_2.n337 VDDA_2.n0 0.00166081
R20529 VDDA_2.n270 VDDA_2.n268 0.00166081
R20530 VDDA_2.n332 VDDA_2.n286 0.00166081
R20531 VDDA_2.n287 VDDA_2.n252 0.00166081
R20532 VDDA_2.n331 VDDA_2.n288 0.00166081
R20533 VDDA_2.n289 VDDA_2.n251 0.00166081
R20534 VDDA_2.n330 VDDA_2.n290 0.00166081
R20535 VDDA_2.n291 VDDA_2.n250 0.00166081
R20536 VDDA_2.n329 VDDA_2.n292 0.00166081
R20537 VDDA_2.n293 VDDA_2.n249 0.00166081
R20538 VDDA_2.n328 VDDA_2.n294 0.00166081
R20539 VDDA_2.n295 VDDA_2.n248 0.00166081
R20540 VDDA_2.n327 VDDA_2.n296 0.00166081
R20541 VDDA_2.n297 VDDA_2.n247 0.00166081
R20542 VDDA_2.n326 VDDA_2.n298 0.00166081
R20543 VDDA_2.n299 VDDA_2.n246 0.00166081
R20544 VDDA_2.n325 VDDA_2.n300 0.00166081
R20545 VDDA_2.n301 VDDA_2.n245 0.00166081
R20546 VDDA_2.n324 VDDA_2.n302 0.00166081
R20547 VDDA_2.n303 VDDA_2.n244 0.00166081
R20548 VDDA_2.n323 VDDA_2.n304 0.00166081
R20549 VDDA_2.n305 VDDA_2.n243 0.00166081
R20550 VDDA_2.n322 VDDA_2.n306 0.00166081
R20551 VDDA_2.n307 VDDA_2.n242 0.00166081
R20552 VDDA_2.n321 VDDA_2.n308 0.00166081
R20553 VDDA_2.n309 VDDA_2.n241 0.00166081
R20554 VDDA_2.n320 VDDA_2.n310 0.00166081
R20555 VDDA_2.n311 VDDA_2.n240 0.00166081
R20556 VDDA_2.n319 VDDA_2.n312 0.00166081
R20557 VDDA_2.n313 VDDA_2.n239 0.00166081
R20558 VDDA_2.n318 VDDA_2.n314 0.00166081
R20559 VDDA_2.n315 VDDA_2.n238 0.00166081
R20560 VDDA_2.n335 VDDA_2.n334 0.00166081
R20561 VDDA_2.n237 VDDA_2.n0 0.00166081
R20562 two_stage_opamp_dummy_magic_29_0.V_err_mir_p two_stage_opamp_dummy_magic_29_0.V_err_mir_p.n1 186.762
R20563 two_stage_opamp_dummy_magic_29_0.V_err_mir_p two_stage_opamp_dummy_magic_29_0.V_err_mir_p.n0 177.201
R20564 two_stage_opamp_dummy_magic_29_0.V_err_mir_p.n0 two_stage_opamp_dummy_magic_29_0.V_err_mir_p.t3 15.7605
R20565 two_stage_opamp_dummy_magic_29_0.V_err_mir_p.n0 two_stage_opamp_dummy_magic_29_0.V_err_mir_p.t0 15.7605
R20566 two_stage_opamp_dummy_magic_29_0.V_err_mir_p.n1 two_stage_opamp_dummy_magic_29_0.V_err_mir_p.t1 15.7605
R20567 two_stage_opamp_dummy_magic_29_0.V_err_mir_p.n1 two_stage_opamp_dummy_magic_29_0.V_err_mir_p.t2 15.7605
R20568 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.n3 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.t4 661.375
R20569 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.n0 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.t1 661.375
R20570 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.t2 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.n1 213.131
R20571 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.n2 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.t5 213.131
R20572 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.t9 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.t2 146.155
R20573 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.t5 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.t9 146.155
R20574 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.n1 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.t3 76.2576
R20575 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.n2 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.t7 76.2576
R20576 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.n7 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.n6 66.0338
R20577 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.n9 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.n8 66.0338
R20578 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.n9 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.n7 13.3963
R20579 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.n6 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.t10 11.2576
R20580 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.n6 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.t6 11.2576
R20581 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.n8 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.t0 11.2576
R20582 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.n8 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.t8 11.2576
R20583 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.n9 6.72967
R20584 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.n5 5.57862
R20585 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.n4 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.n0 5.1255
R20586 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.n4 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.n3 4.7505
R20587 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.n5 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.n4 4.5005
R20588 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.n1 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.n0 1.888
R20589 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.n3 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.n2 1.888
R20590 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.n7 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.n5 0.854667
R20591 a_3110_3878.t0 a_3110_3878.t1 294.339
R20592 a_13940_76.t0 a_13940_76.t1 169.905
R20593 a_11300_28630.t0 a_11300_28630.t1 178.133
R20594 two_stage_opamp_dummy_magic_29_0.V_p_mir.n1 two_stage_opamp_dummy_magic_29_0.V_p_mir.n0 95.5151
R20595 two_stage_opamp_dummy_magic_29_0.V_p_mir.n0 two_stage_opamp_dummy_magic_29_0.V_p_mir.t2 16.0005
R20596 two_stage_opamp_dummy_magic_29_0.V_p_mir.n0 two_stage_opamp_dummy_magic_29_0.V_p_mir.t3 16.0005
R20597 two_stage_opamp_dummy_magic_29_0.V_p_mir.t1 two_stage_opamp_dummy_magic_29_0.V_p_mir.n1 9.6005
R20598 two_stage_opamp_dummy_magic_29_0.V_p_mir.n1 two_stage_opamp_dummy_magic_29_0.V_p_mir.t0 9.6005
R20599 bgr_11_0.V_p_1.n0 bgr_11_0.V_p_1.t1 99.8322
R20600 bgr_11_0.V_p_1.t0 bgr_11_0.V_p_1.n0 9.6005
R20601 bgr_11_0.V_p_1.n0 bgr_11_0.V_p_1.t2 9.6005
R20602 a_3830_76.t0 a_3830_76.t1 169.905
R20603 a_5700_30088.t0 a_5700_30088.t1 178.133
R20604 a_5820_28824.t0 a_5820_28824.t1 178.133
R20605 a_6470_28630.t0 a_6470_28630.t1 178.133
R20606 a_12070_30088.t0 a_12070_30088.t1 178.133
R20607 bgr_11_0.V_CUR_REF_REG bgr_11_0.V_CUR_REF_REG.t3 701.501
R20608 bgr_11_0.V_CUR_REF_REG.n1 bgr_11_0.V_CUR_REF_REG.n0 357.647
R20609 bgr_11_0.V_CUR_REF_REG.n1 bgr_11_0.V_CUR_REF_REG.t0 135.239
R20610 bgr_11_0.V_CUR_REF_REG.n0 bgr_11_0.V_CUR_REF_REG.t1 39.4005
R20611 bgr_11_0.V_CUR_REF_REG.n0 bgr_11_0.V_CUR_REF_REG.t2 39.4005
R20612 bgr_11_0.V_CUR_REF_REG bgr_11_0.V_CUR_REF_REG.n1 5.79738
R20613 bgr_11_0.V_p_2.n0 bgr_11_0.V_p_2.t2 142.558
R20614 bgr_11_0.V_p_2.n0 bgr_11_0.V_p_2.t1 9.6005
R20615 bgr_11_0.V_p_2.t0 bgr_11_0.V_p_2.n0 9.6005
R20616 a_14540_3878.t0 a_14540_3878.t1 169.905
R20617 GNDA.n4284 GNDA.n1965 554309
R20618 GNDA.n5388 GNDA.n705 549118
R20619 GNDA.n5390 GNDA.n5389 443417
R20620 GNDA.n4282 GNDA.n4281 438167
R20621 GNDA.n5378 GNDA.n707 396244
R20622 GNDA.n4285 GNDA.n711 235669
R20623 GNDA.n5513 GNDA.n626 215600
R20624 GNDA.n5386 GNDA.n5382 204995
R20625 GNDA.n5386 GNDA.n5385 191583
R20626 GNDA.n4283 GNDA.n4282 182270
R20627 GNDA.n5385 GNDA.n626 151067
R20628 GNDA.n4281 GNDA.n4280 132000
R20629 GNDA.n5389 GNDA.n706 132000
R20630 GNDA.n5379 GNDA.n5378 105027
R20631 GNDA.n5378 GNDA.n5377 71214.8
R20632 GNDA.n4285 GNDA.n4284 70780.9
R20633 GNDA.n1540 GNDA.n707 55733.3
R20634 GNDA.n4280 GNDA.n626 52108.6
R20635 GNDA.n4286 GNDA.n1965 27866.7
R20636 GNDA.n5388 GNDA.n5387 27866.7
R20637 GNDA.n5387 GNDA.n5386 24653.3
R20638 GNDA.n5390 GNDA.n625 24387.2
R20639 GNDA.n709 GNDA.n705 22454.8
R20640 GNDA.n5385 GNDA.n5384 21706.7
R20641 GNDA.n4286 GNDA.n4285 20495.4
R20642 GNDA.n1968 GNDA.n1967 19875.1
R20643 GNDA.n4321 GNDA.n4287 17109.1
R20644 GNDA.n1554 GNDA.n1553 17106.8
R20645 GNDA.n4328 GNDA.n4286 16070.1
R20646 GNDA.n5383 GNDA.n627 14959.6
R20647 GNDA.n709 GNDA.n704 14561.9
R20648 GNDA.n5387 GNDA.n707 13906.7
R20649 GNDA.n5384 GNDA.n710 13566.7
R20650 GNDA.n5382 GNDA.n5381 13527.3
R20651 GNDA.n5381 GNDA.n5380 13460.8
R20652 GNDA.n5382 GNDA.n711 12640.3
R20653 GNDA.n5391 GNDA.n5390 11950.8
R20654 GNDA.n5392 GNDA.n5391 11691.4
R20655 GNDA.n1967 GNDA.n1966 11163
R20656 GNDA.n5395 GNDA.n629 11032
R20657 GNDA.n5510 GNDA.n629 11032
R20658 GNDA.n5511 GNDA.n627 10979
R20659 GNDA.n5394 GNDA.n5392 10979
R20660 GNDA.n5395 GNDA.n628 10933.5
R20661 GNDA.n5510 GNDA.n628 10933.5
R20662 GNDA.n5456 GNDA.n673 10884.2
R20663 GNDA.n5456 GNDA.n674 10884.2
R20664 GNDA.n5464 GNDA.n673 10441
R20665 GNDA.n5464 GNDA.n674 10441
R20666 GNDA.n710 GNDA.n709 10046.7
R20667 GNDA.n5523 GNDA.n39 9850
R20668 GNDA.n5523 GNDA.n38 9751.5
R20669 GNDA.n5377 GNDA.n5376 9511.11
R20670 GNDA.n5376 GNDA.n711 9423.88
R20671 GNDA.n592 GNDA.n39 9406.75
R20672 GNDA.n592 GNDA.n38 9308.25
R20673 GNDA.n3301 GNDA.n706 9121.95
R20674 GNDA.n5393 GNDA.n625 9051.43
R20675 GNDA.n4280 GNDA.n4279 7832.46
R20676 GNDA.n5327 GNDA.n5325 7452.79
R20677 GNDA.n706 GNDA.n625 7266.06
R20678 GNDA.n4284 GNDA.n4283 6794.03
R20679 GNDA.n3301 GNDA.n2115 6760.98
R20680 GNDA.n5513 GNDA.n5512 6495.24
R20681 GNDA.n4283 GNDA.n1966 6475.77
R20682 GNDA.n5512 GNDA.n5511 6285.71
R20683 GNDA.n5394 GNDA.n5393 6285.71
R20684 GNDA.n5384 GNDA.n5383 6010.32
R20685 GNDA.n5516 GNDA.n622 5910
R20686 GNDA.n4279 GNDA.n1968 5805.24
R20687 GNDA.n4282 GNDA.n1967 5681.89
R20688 GNDA.n5520 GNDA.n622 5466.75
R20689 GNDA.n5516 GNDA.n621 5319
R20690 GNDA.n5383 GNDA.n704 5185.26
R20691 GNDA.n5520 GNDA.n621 4875.75
R20692 GNDA.n5379 GNDA.n708 4738.46
R20693 GNDA.n5386 GNDA.n708 4538.62
R20694 GNDA.n5386 GNDA.n710 4538.62
R20695 GNDA.n5027 GNDA.n944 4512.16
R20696 GNDA.n4915 GNDA.n4914 4478.96
R20697 GNDA.n672 GNDA.n671 4375.56
R20698 GNDA.n5376 GNDA.n5375 4106.67
R20699 GNDA.n5380 GNDA.n5377 4106.67
R20700 GNDA.n5473 GNDA.n669 3841.5
R20701 GNDA.n5473 GNDA.n668 3743
R20702 GNDA.n5476 GNDA.n668 3743
R20703 GNDA.n5514 GNDA.n5513 2577.14
R20704 GNDA.n5522 GNDA.n40 2566.67
R20705 GNDA.n5391 GNDA.n705 2306.8
R20706 GNDA.n671 GNDA.n670 2102.22
R20707 GNDA.n5325 GNDA.n753 1874.83
R20708 GNDA.n5389 GNDA.n5388 1860.36
R20709 GNDA.n5465 GNDA.n672 1784.44
R20710 GNDA.n670 GNDA.n40 1417.78
R20711 GNDA.n5515 GNDA.n624 1417.78
R20712 GNDA.n4281 GNDA.n1965 1308.49
R20713 GNDA.n5391 GNDA.n704 1194.29
R20714 GNDA.n5466 GNDA.n5465 1100
R20715 GNDA.n5474 GNDA.n5466 1075.56
R20716 GNDA.n5522 GNDA.n5521 1075.56
R20717 GNDA.n1966 GNDA.n626 1068.57
R20718 GNDA.n5380 GNDA.n5379 1031.25
R20719 GNDA.n5475 GNDA.n669 980.59
R20720 GNDA.n5381 GNDA.n708 854.477
R20721 GNDA.n5521 GNDA.n620 782.222
R20722 GNDA.n2207 GNDA.n2206 749.742
R20723 GNDA.n3619 GNDA.n3618 749.742
R20724 GNDA.n3624 GNDA.n3623 749.742
R20725 GNDA.n2202 GNDA.n2201 747.734
R20726 GNDA.n4846 GNDA.n1171 741.376
R20727 GNDA.n1284 GNDA.n825 741.376
R20728 GNDA.n4846 GNDA.n4845 741.376
R20729 GNDA.n924 GNDA.n825 741.376
R20730 GNDA.n5317 GNDA.n5316 686.717
R20731 GNDA.n5166 GNDA.n5165 686.717
R20732 GNDA.n5156 GNDA.n5043 686.717
R20733 GNDA.n5310 GNDA.n772 686.717
R20734 GNDA.n702 GNDA.n630 678.4
R20735 GNDA.n703 GNDA.n702 678.4
R20736 GNDA.n5458 GNDA.n5457 675.201
R20737 GNDA.n5457 GNDA.n5455 675.201
R20738 GNDA.n5142 GNDA.n5141 669.307
R20739 GNDA.n5058 GNDA.n5057 669.307
R20740 GNDA.n5469 GNDA.n5468 659.367
R20741 GNDA.n5481 GNDA.n5480 659.367
R20742 GNDA.n32 GNDA.n31 659.367
R20743 GNDA.n583 GNDA.n582 659.367
R20744 GNDA.n1116 GNDA.n1115 654.447
R20745 GNDA.n5463 GNDA.n675 646.4
R20746 GNDA.n5463 GNDA.n5462 646.4
R20747 GNDA.n593 GNDA.n591 611.201
R20748 GNDA.n594 GNDA.n593 604.801
R20749 GNDA.n4918 GNDA.n4916 589.494
R20750 GNDA.n5025 GNDA.n5024 585.001
R20751 GNDA.n5017 GNDA.n5016 585.001
R20752 GNDA.n877 GNDA.n876 585.001
R20753 GNDA.n5349 GNDA.n5348 585.001
R20754 GNDA.n821 GNDA.n820 585.001
R20755 GNDA.n5219 GNDA.n5218 585.001
R20756 GNDA.n5339 GNDA.n5338 585.001
R20757 GNDA.n1113 GNDA.n1111 585
R20758 GNDA.n4883 GNDA.n4882 585
R20759 GNDA.n4882 GNDA.n4881 585
R20760 GNDA.n1575 GNDA.n1524 585
R20761 GNDA.n1579 GNDA.n1524 585
R20762 GNDA.n1577 GNDA.n1576 585
R20763 GNDA.n1578 GNDA.n1577 585
R20764 GNDA.n1574 GNDA.n1529 585
R20765 GNDA.n1529 GNDA.n1528 585
R20766 GNDA.n1573 GNDA.n1572 585
R20767 GNDA.n1572 GNDA.n1571 585
R20768 GNDA.n1531 GNDA.n1530 585
R20769 GNDA.n1570 GNDA.n1531 585
R20770 GNDA.n1568 GNDA.n1567 585
R20771 GNDA.n1569 GNDA.n1568 585
R20772 GNDA.n1566 GNDA.n1533 585
R20773 GNDA.n1562 GNDA.n1533 585
R20774 GNDA.n1565 GNDA.n1564 585
R20775 GNDA.n1564 GNDA.n1563 585
R20776 GNDA.n1535 GNDA.n1534 585
R20777 GNDA.n1561 GNDA.n1535 585
R20778 GNDA.n1559 GNDA.n1558 585
R20779 GNDA.n1560 GNDA.n1559 585
R20780 GNDA.n1557 GNDA.n1537 585
R20781 GNDA.n1537 GNDA.n1536 585
R20782 GNDA.n1556 GNDA.n1555 585
R20783 GNDA.n1555 GNDA.n1554 585
R20784 GNDA.n4576 GNDA.n4575 585
R20785 GNDA.n4574 GNDA.n4573 585
R20786 GNDA.n4572 GNDA.n4550 585
R20787 GNDA.n4570 GNDA.n4569 585
R20788 GNDA.n4568 GNDA.n4551 585
R20789 GNDA.n4567 GNDA.n4566 585
R20790 GNDA.n4564 GNDA.n4552 585
R20791 GNDA.n4562 GNDA.n4561 585
R20792 GNDA.n4560 GNDA.n4553 585
R20793 GNDA.n4559 GNDA.n4558 585
R20794 GNDA.n4556 GNDA.n4554 585
R20795 GNDA.n1178 GNDA.n1176 585
R20796 GNDA.n1683 GNDA.n1656 585
R20797 GNDA.n1681 GNDA.n1680 585
R20798 GNDA.n1679 GNDA.n1657 585
R20799 GNDA.n1678 GNDA.n1677 585
R20800 GNDA.n1675 GNDA.n1658 585
R20801 GNDA.n1673 GNDA.n1672 585
R20802 GNDA.n1671 GNDA.n1659 585
R20803 GNDA.n1670 GNDA.n1669 585
R20804 GNDA.n1667 GNDA.n1660 585
R20805 GNDA.n1665 GNDA.n1664 585
R20806 GNDA.n1663 GNDA.n1662 585
R20807 GNDA.n1397 GNDA.n1396 585
R20808 GNDA.n1849 GNDA.n1848 585
R20809 GNDA.n1850 GNDA.n1692 585
R20810 GNDA.n1852 GNDA.n1851 585
R20811 GNDA.n1854 GNDA.n1690 585
R20812 GNDA.n1856 GNDA.n1855 585
R20813 GNDA.n1857 GNDA.n1689 585
R20814 GNDA.n1859 GNDA.n1858 585
R20815 GNDA.n1861 GNDA.n1687 585
R20816 GNDA.n1863 GNDA.n1862 585
R20817 GNDA.n1864 GNDA.n1686 585
R20818 GNDA.n1866 GNDA.n1865 585
R20819 GNDA.n1868 GNDA.n1655 585
R20820 GNDA.n4545 GNDA.n4544 585
R20821 GNDA.n4542 GNDA.n4541 585
R20822 GNDA.n4540 GNDA.n4539 585
R20823 GNDA.n4455 GNDA.n1634 585
R20824 GNDA.n4457 GNDA.n4456 585
R20825 GNDA.n4461 GNDA.n4460 585
R20826 GNDA.n4463 GNDA.n4462 585
R20827 GNDA.n4470 GNDA.n4469 585
R20828 GNDA.n4468 GNDA.n4453 585
R20829 GNDA.n4476 GNDA.n4475 585
R20830 GNDA.n4478 GNDA.n4477 585
R20831 GNDA.n4451 GNDA.n4450 585
R20832 GNDA.n4850 GNDA.n4849 585
R20833 GNDA.n1474 GNDA.n1153 585
R20834 GNDA.n1497 GNDA.n1496 585
R20835 GNDA.n1494 GNDA.n1493 585
R20836 GNDA.n1492 GNDA.n1491 585
R20837 GNDA.n1487 GNDA.n1486 585
R20838 GNDA.n1485 GNDA.n1484 585
R20839 GNDA.n1480 GNDA.n1479 585
R20840 GNDA.n1478 GNDA.n1401 585
R20841 GNDA.n1506 GNDA.n1505 585
R20842 GNDA.n1508 GNDA.n1507 585
R20843 GNDA.n1511 GNDA.n1510 585
R20844 GNDA.n1625 GNDA.n1513 585
R20845 GNDA.n1628 GNDA.n1627 585
R20846 GNDA.n1624 GNDA.n1515 585
R20847 GNDA.n1622 GNDA.n1621 585
R20848 GNDA.n1517 GNDA.n1516 585
R20849 GNDA.n1615 GNDA.n1614 585
R20850 GNDA.n1612 GNDA.n1519 585
R20851 GNDA.n1610 GNDA.n1609 585
R20852 GNDA.n1521 GNDA.n1520 585
R20853 GNDA.n1603 GNDA.n1602 585
R20854 GNDA.n1600 GNDA.n1523 585
R20855 GNDA.n1598 GNDA.n1597 585
R20856 GNDA.n4547 GNDA.n1512 585
R20857 GNDA.n1512 GNDA.n1138 585
R20858 GNDA.n1597 GNDA.n1596 585
R20859 GNDA.n1523 GNDA.n1522 585
R20860 GNDA.n1604 GNDA.n1603 585
R20861 GNDA.n1606 GNDA.n1521 585
R20862 GNDA.n1609 GNDA.n1608 585
R20863 GNDA.n1519 GNDA.n1518 585
R20864 GNDA.n1616 GNDA.n1615 585
R20865 GNDA.n1618 GNDA.n1517 585
R20866 GNDA.n1621 GNDA.n1620 585
R20867 GNDA.n1515 GNDA.n1514 585
R20868 GNDA.n1629 GNDA.n1628 585
R20869 GNDA.n1631 GNDA.n1513 585
R20870 GNDA.n4547 GNDA.n4546 585
R20871 GNDA.n4546 GNDA.n1138 585
R20872 GNDA.n4597 GNDA.n4595 585
R20873 GNDA.n4598 GNDA.n4592 585
R20874 GNDA.n4601 GNDA.n4591 585
R20875 GNDA.n4602 GNDA.n4589 585
R20876 GNDA.n4605 GNDA.n4588 585
R20877 GNDA.n4606 GNDA.n4586 585
R20878 GNDA.n4609 GNDA.n4585 585
R20879 GNDA.n4610 GNDA.n4583 585
R20880 GNDA.n4613 GNDA.n4582 585
R20881 GNDA.n4615 GNDA.n4580 585
R20882 GNDA.n4616 GNDA.n4579 585
R20883 GNDA.n4617 GNDA.n4577 585
R20884 GNDA.n4618 GNDA.n4617 585
R20885 GNDA.n4616 GNDA.n1395 585
R20886 GNDA.n4615 GNDA.n4614 585
R20887 GNDA.n4613 GNDA.n4612 585
R20888 GNDA.n4611 GNDA.n4610 585
R20889 GNDA.n4609 GNDA.n4608 585
R20890 GNDA.n4607 GNDA.n4606 585
R20891 GNDA.n4605 GNDA.n4604 585
R20892 GNDA.n4603 GNDA.n4602 585
R20893 GNDA.n4601 GNDA.n4600 585
R20894 GNDA.n4599 GNDA.n4598 585
R20895 GNDA.n4597 GNDA.n4596 585
R20896 GNDA.n5188 GNDA.n871 585
R20897 GNDA.n5189 GNDA.n869 585
R20898 GNDA.n868 GNDA.n865 585
R20899 GNDA.n5195 GNDA.n864 585
R20900 GNDA.n5196 GNDA.n863 585
R20901 GNDA.n5197 GNDA.n861 585
R20902 GNDA.n860 GNDA.n857 585
R20903 GNDA.n5203 GNDA.n856 585
R20904 GNDA.n5204 GNDA.n855 585
R20905 GNDA.n5205 GNDA.n853 585
R20906 GNDA.n852 GNDA.n848 585
R20907 GNDA.n5210 GNDA.n844 585
R20908 GNDA.n5210 GNDA.n5209 585
R20909 GNDA.n5207 GNDA.n848 585
R20910 GNDA.n5206 GNDA.n5205 585
R20911 GNDA.n5206 GNDA.n712 585
R20912 GNDA.n5204 GNDA.n850 585
R20913 GNDA.n5203 GNDA.n5202 585
R20914 GNDA.n5200 GNDA.n857 585
R20915 GNDA.n5198 GNDA.n5197 585
R20916 GNDA.n5196 GNDA.n858 585
R20917 GNDA.n5195 GNDA.n5194 585
R20918 GNDA.n5192 GNDA.n865 585
R20919 GNDA.n5190 GNDA.n5189 585
R20920 GNDA.n5188 GNDA.n866 585
R20921 GNDA.n866 GNDA.n712 585
R20922 GNDA.n5213 GNDA.n5212 585
R20923 GNDA.n845 GNDA.n843 585
R20924 GNDA.n905 GNDA.n904 585
R20925 GNDA.n907 GNDA.n906 585
R20926 GNDA.n909 GNDA.n908 585
R20927 GNDA.n911 GNDA.n910 585
R20928 GNDA.n913 GNDA.n912 585
R20929 GNDA.n915 GNDA.n914 585
R20930 GNDA.n917 GNDA.n916 585
R20931 GNDA.n919 GNDA.n918 585
R20932 GNDA.n921 GNDA.n920 585
R20933 GNDA.n923 GNDA.n922 585
R20934 GNDA.n1330 GNDA.n1329 585
R20935 GNDA.n1328 GNDA.n1327 585
R20936 GNDA.n1326 GNDA.n1325 585
R20937 GNDA.n1324 GNDA.n1323 585
R20938 GNDA.n1322 GNDA.n1321 585
R20939 GNDA.n1320 GNDA.n1319 585
R20940 GNDA.n1318 GNDA.n1317 585
R20941 GNDA.n1316 GNDA.n1315 585
R20942 GNDA.n1314 GNDA.n1313 585
R20943 GNDA.n1312 GNDA.n1311 585
R20944 GNDA.n1310 GNDA.n1309 585
R20945 GNDA.n849 GNDA.n846 585
R20946 GNDA.n1287 GNDA.n1286 585
R20947 GNDA.n1289 GNDA.n1288 585
R20948 GNDA.n1291 GNDA.n1290 585
R20949 GNDA.n1293 GNDA.n1292 585
R20950 GNDA.n1295 GNDA.n1294 585
R20951 GNDA.n1297 GNDA.n1296 585
R20952 GNDA.n1299 GNDA.n1298 585
R20953 GNDA.n1301 GNDA.n1300 585
R20954 GNDA.n1303 GNDA.n1302 585
R20955 GNDA.n1305 GNDA.n1304 585
R20956 GNDA.n1307 GNDA.n1306 585
R20957 GNDA.n1333 GNDA.n1308 585
R20958 GNDA.n4594 GNDA.n847 585
R20959 GNDA.n4594 GNDA.n1218 585
R20960 GNDA.n4819 GNDA.n4818 585
R20961 GNDA.n4816 GNDA.n4815 585
R20962 GNDA.n4814 GNDA.n4813 585
R20963 GNDA.n4727 GNDA.n1195 585
R20964 GNDA.n4747 GNDA.n4746 585
R20965 GNDA.n4743 GNDA.n4726 585
R20966 GNDA.n4730 GNDA.n4729 585
R20967 GNDA.n4738 GNDA.n4737 585
R20968 GNDA.n4736 GNDA.n4735 585
R20969 GNDA.n1216 GNDA.n1215 585
R20970 GNDA.n4752 GNDA.n4751 585
R20971 GNDA.n1232 GNDA.n1217 585
R20972 GNDA.n1231 GNDA.n847 585
R20973 GNDA.n1231 GNDA.n1218 585
R20974 GNDA.n4722 GNDA.n4721 585
R20975 GNDA.n4719 GNDA.n1230 585
R20976 GNDA.n1236 GNDA.n1235 585
R20977 GNDA.n4714 GNDA.n4713 585
R20978 GNDA.n4712 GNDA.n4711 585
R20979 GNDA.n4637 GNDA.n1240 585
R20980 GNDA.n4639 GNDA.n4638 585
R20981 GNDA.n4644 GNDA.n4643 585
R20982 GNDA.n4642 GNDA.n4635 585
R20983 GNDA.n4650 GNDA.n4649 585
R20984 GNDA.n4652 GNDA.n4651 585
R20985 GNDA.n4633 GNDA.n4632 585
R20986 GNDA.n1782 GNDA.n1378 585
R20987 GNDA.n1806 GNDA.n1784 585
R20988 GNDA.n1808 GNDA.n1807 585
R20989 GNDA.n1804 GNDA.n1803 585
R20990 GNDA.n1802 GNDA.n1801 585
R20991 GNDA.n1797 GNDA.n1796 585
R20992 GNDA.n1795 GNDA.n1794 585
R20993 GNDA.n1790 GNDA.n1789 585
R20994 GNDA.n1788 GNDA.n1709 585
R20995 GNDA.n1817 GNDA.n1816 585
R20996 GNDA.n1819 GNDA.n1818 585
R20997 GNDA.n1822 GNDA.n1821 585
R20998 GNDA.n5328 GNDA.n761 585
R20999 GNDA.n5331 GNDA.n5330 585
R21000 GNDA.n5330 GNDA.n5329 585
R21001 GNDA.n760 GNDA.n759 585
R21002 GNDA.n762 GNDA.n760 585
R21003 GNDA.n1271 GNDA.n1270 585
R21004 GNDA.n1270 GNDA.n1269 585
R21005 GNDA.n1272 GNDA.n1267 585
R21006 GNDA.n1268 GNDA.n1267 585
R21007 GNDA.n1274 GNDA.n1273 585
R21008 GNDA.n1274 GNDA.n774 585
R21009 GNDA.n1275 GNDA.n1266 585
R21010 GNDA.n1275 GNDA.n773 585
R21011 GNDA.n1278 GNDA.n1277 585
R21012 GNDA.n1277 GNDA.n1276 585
R21013 GNDA.n1279 GNDA.n1264 585
R21014 GNDA.n1264 GNDA.n1263 585
R21015 GNDA.n1281 GNDA.n1280 585
R21016 GNDA.n1282 GNDA.n1281 585
R21017 GNDA.n1265 GNDA.n1262 585
R21018 GNDA.n1283 GNDA.n1262 585
R21019 GNDA.n1285 GNDA.n1261 585
R21020 GNDA.n1285 GNDA.n1284 585
R21021 GNDA.n5327 GNDA.n5326 585
R21022 GNDA.n1826 GNDA.n1706 585
R21023 GNDA.n1829 GNDA.n1828 585
R21024 GNDA.n1828 GNDA.n1827 585
R21025 GNDA.n1830 GNDA.n1703 585
R21026 GNDA.n1703 GNDA.n1702 585
R21027 GNDA.n1832 GNDA.n1831 585
R21028 GNDA.n1833 GNDA.n1832 585
R21029 GNDA.n1704 GNDA.n1701 585
R21030 GNDA.n1834 GNDA.n1701 585
R21031 GNDA.n1836 GNDA.n1700 585
R21032 GNDA.n1836 GNDA.n1835 585
R21033 GNDA.n1839 GNDA.n1838 585
R21034 GNDA.n1838 GNDA.n1837 585
R21035 GNDA.n1840 GNDA.n1698 585
R21036 GNDA.n1698 GNDA.n1697 585
R21037 GNDA.n1842 GNDA.n1841 585
R21038 GNDA.n1843 GNDA.n1842 585
R21039 GNDA.n1699 GNDA.n1695 585
R21040 GNDA.n1844 GNDA.n1695 585
R21041 GNDA.n1846 GNDA.n1696 585
R21042 GNDA.n1846 GNDA.n1845 585
R21043 GNDA.n1847 GNDA.n1693 585
R21044 GNDA.n1847 GNDA.n1171 585
R21045 GNDA.n1825 GNDA.n1824 585
R21046 GNDA.n4348 GNDA.n4347 585
R21047 GNDA.n4350 GNDA.n1172 585
R21048 GNDA.n4446 GNDA.n4445 585
R21049 GNDA.n4443 GNDA.n4442 585
R21050 GNDA.n4441 GNDA.n4440 585
R21051 GNDA.n4356 GNDA.n1938 585
R21052 GNDA.n4358 GNDA.n4357 585
R21053 GNDA.n4362 GNDA.n4361 585
R21054 GNDA.n4364 GNDA.n4363 585
R21055 GNDA.n4371 GNDA.n4370 585
R21056 GNDA.n4369 GNDA.n4354 585
R21057 GNDA.n4377 GNDA.n4376 585
R21058 GNDA.n4379 GNDA.n4378 585
R21059 GNDA.n4352 GNDA.n4351 585
R21060 GNDA.n4342 GNDA.n1958 585
R21061 GNDA.n4346 GNDA.n1958 585
R21062 GNDA.n4344 GNDA.n4343 585
R21063 GNDA.n4345 GNDA.n4344 585
R21064 GNDA.n4341 GNDA.n1960 585
R21065 GNDA.n1960 GNDA.n1959 585
R21066 GNDA.n4340 GNDA.n4339 585
R21067 GNDA.n4339 GNDA.n4338 585
R21068 GNDA.n4337 GNDA.n1961 585
R21069 GNDA.n4337 GNDA.n1140 585
R21070 GNDA.n4336 GNDA.n4335 585
R21071 GNDA.n4336 GNDA.n1139 585
R21072 GNDA.n4334 GNDA.n1962 585
R21073 GNDA.n4330 GNDA.n1962 585
R21074 GNDA.n4333 GNDA.n4332 585
R21075 GNDA.n4332 GNDA.n4331 585
R21076 GNDA.n1964 GNDA.n1963 585
R21077 GNDA.n4329 GNDA.n1964 585
R21078 GNDA.n4326 GNDA.n4325 585
R21079 GNDA.n4327 GNDA.n4326 585
R21080 GNDA.n4324 GNDA.n4288 585
R21081 GNDA.n4288 GNDA.n4287 585
R21082 GNDA.n4323 GNDA.n4322 585
R21083 GNDA.n4322 GNDA.n4321 585
R21084 GNDA.n4290 GNDA.n4289 585
R21085 GNDA.n4320 GNDA.n4290 585
R21086 GNDA.n4318 GNDA.n4317 585
R21087 GNDA.n4319 GNDA.n4318 585
R21088 GNDA.n4316 GNDA.n4292 585
R21089 GNDA.n4292 GNDA.n4291 585
R21090 GNDA.n4315 GNDA.n4314 585
R21091 GNDA.n4314 GNDA.n4313 585
R21092 GNDA.n4294 GNDA.n4293 585
R21093 GNDA.n4312 GNDA.n4294 585
R21094 GNDA.n4309 GNDA.n4308 585
R21095 GNDA.n4310 GNDA.n4309 585
R21096 GNDA.n4307 GNDA.n4296 585
R21097 GNDA.n4296 GNDA.n4295 585
R21098 GNDA.n4306 GNDA.n4305 585
R21099 GNDA.n4305 GNDA.n4304 585
R21100 GNDA.n4298 GNDA.n4297 585
R21101 GNDA.n4303 GNDA.n4298 585
R21102 GNDA.n4301 GNDA.n4300 585
R21103 GNDA.n4302 GNDA.n4301 585
R21104 GNDA.n1127 GNDA.n1124 585
R21105 GNDA.n4299 GNDA.n1127 585
R21106 GNDA.n4869 GNDA.n1123 585
R21107 GNDA.n1123 GNDA.n1122 585
R21108 GNDA.n4871 GNDA.n4870 585
R21109 GNDA.n4872 GNDA.n4871 585
R21110 GNDA.n1121 GNDA.n1120 585
R21111 GNDA.n4873 GNDA.n1121 585
R21112 GNDA.n4876 GNDA.n4875 585
R21113 GNDA.n4875 GNDA.n4874 585
R21114 GNDA.n4877 GNDA.n1119 585
R21115 GNDA.n1119 GNDA.n1117 585
R21116 GNDA.n4879 GNDA.n4878 585
R21117 GNDA.n4880 GNDA.n4879 585
R21118 GNDA.n1584 GNDA.n1118 585
R21119 GNDA.n1118 GNDA.n1114 585
R21120 GNDA.n1587 GNDA.n1586 585
R21121 GNDA.n1586 GNDA.n1585 585
R21122 GNDA.n1588 GNDA.n1582 585
R21123 GNDA.n1582 GNDA.n1581 585
R21124 GNDA.n1590 GNDA.n1589 585
R21125 GNDA.n1591 GNDA.n1590 585
R21126 GNDA.n1583 GNDA.n1526 585
R21127 GNDA.n1592 GNDA.n1526 585
R21128 GNDA.n1594 GNDA.n1527 585
R21129 GNDA.n1594 GNDA.n1593 585
R21130 GNDA.n1934 GNDA.n1654 585
R21131 GNDA.n1933 GNDA.n1930 585
R21132 GNDA.n1928 GNDA.n1900 585
R21133 GNDA.n1926 GNDA.n1925 585
R21134 GNDA.n1922 GNDA.n1901 585
R21135 GNDA.n1921 GNDA.n1918 585
R21136 GNDA.n1916 GNDA.n1902 585
R21137 GNDA.n1914 GNDA.n1913 585
R21138 GNDA.n1910 GNDA.n1903 585
R21139 GNDA.n1909 GNDA.n1907 585
R21140 GNDA.n1905 GNDA.n1126 585
R21141 GNDA.n4867 GNDA.n1125 585
R21142 GNDA.n4449 GNDA.n4448 585
R21143 GNDA.n4449 GNDA.n1138 585
R21144 GNDA.n4867 GNDA.n4866 585
R21145 GNDA.n1128 GNDA.n1126 585
R21146 GNDA.n1909 GNDA.n1908 585
R21147 GNDA.n1911 GNDA.n1910 585
R21148 GNDA.n1913 GNDA.n1912 585
R21149 GNDA.n1919 GNDA.n1902 585
R21150 GNDA.n1921 GNDA.n1920 585
R21151 GNDA.n1923 GNDA.n1922 585
R21152 GNDA.n1925 GNDA.n1924 585
R21153 GNDA.n1931 GNDA.n1900 585
R21154 GNDA.n1933 GNDA.n1932 585
R21155 GNDA.n1935 GNDA.n1934 585
R21156 GNDA.n4448 GNDA.n4447 585
R21157 GNDA.n4447 GNDA.n1138 585
R21158 GNDA.n1379 GNDA.n1260 585
R21159 GNDA.n4625 GNDA.n4624 585
R21160 GNDA.n1383 GNDA.n1382 585
R21161 GNDA.n1880 GNDA.n1879 585
R21162 GNDA.n1885 GNDA.n1878 585
R21163 GNDA.n1886 GNDA.n1877 585
R21164 GNDA.n1887 GNDA.n1876 585
R21165 GNDA.n1874 GNDA.n1873 585
R21166 GNDA.n1892 GNDA.n1872 585
R21167 GNDA.n1893 GNDA.n1871 585
R21168 GNDA.n1870 GNDA.n1685 585
R21169 GNDA.n1898 GNDA.n1684 585
R21170 GNDA.n4631 GNDA.n4630 585
R21171 GNDA.n4631 GNDA.n1218 585
R21172 GNDA.n1898 GNDA.n1897 585
R21173 GNDA.n1895 GNDA.n1685 585
R21174 GNDA.n1894 GNDA.n1893 585
R21175 GNDA.n1892 GNDA.n1891 585
R21176 GNDA.n1890 GNDA.n1874 585
R21177 GNDA.n1888 GNDA.n1887 585
R21178 GNDA.n1886 GNDA.n1875 585
R21179 GNDA.n1885 GNDA.n1884 585
R21180 GNDA.n1882 GNDA.n1880 585
R21181 GNDA.n1382 GNDA.n1381 585
R21182 GNDA.n4626 GNDA.n4625 585
R21183 GNDA.n4628 GNDA.n1379 585
R21184 GNDA.n4630 GNDA.n4629 585
R21185 GNDA.n4629 GNDA.n1218 585
R21186 GNDA.n817 GNDA.n816 585
R21187 GNDA.n1355 GNDA.n1354 585
R21188 GNDA.n1352 GNDA.n1349 585
R21189 GNDA.n1361 GNDA.n1348 585
R21190 GNDA.n1362 GNDA.n1347 585
R21191 GNDA.n1363 GNDA.n1345 585
R21192 GNDA.n1344 GNDA.n1341 585
R21193 GNDA.n1369 GNDA.n1340 585
R21194 GNDA.n1370 GNDA.n1339 585
R21195 GNDA.n1371 GNDA.n1337 585
R21196 GNDA.n1336 GNDA.n1332 585
R21197 GNDA.n1376 GNDA.n1331 585
R21198 GNDA.n1376 GNDA.n1375 585
R21199 GNDA.n1373 GNDA.n1332 585
R21200 GNDA.n1372 GNDA.n1371 585
R21201 GNDA.n1372 GNDA.n775 585
R21202 GNDA.n1370 GNDA.n1334 585
R21203 GNDA.n1369 GNDA.n1368 585
R21204 GNDA.n1366 GNDA.n1341 585
R21205 GNDA.n1364 GNDA.n1363 585
R21206 GNDA.n1362 GNDA.n1342 585
R21207 GNDA.n1361 GNDA.n1360 585
R21208 GNDA.n1358 GNDA.n1349 585
R21209 GNDA.n1356 GNDA.n1355 585
R21210 GNDA.n1350 GNDA.n816 585
R21211 GNDA.n1350 GNDA.n775 585
R21212 GNDA.n5059 GNDA.n5056 585
R21213 GNDA.n5061 GNDA.n5060 585
R21214 GNDA.n5060 GNDA.n743 585
R21215 GNDA.n5070 GNDA.n5069 585
R21216 GNDA.n5145 GNDA.n5144 585
R21217 GNDA.n5144 GNDA.n5143 585
R21218 GNDA.n5164 GNDA.n5045 585
R21219 GNDA.n5155 GNDA.n5044 585
R21220 GNDA.n5167 GNDA.n5044 585
R21221 GNDA.n5160 GNDA.n5159 585
R21222 GNDA.n5306 GNDA.n770 585
R21223 GNDA.n5314 GNDA.n5313 585
R21224 GNDA.n5315 GNDA.n5314 585
R21225 GNDA.n5308 GNDA.n5305 585
R21226 GNDA.n884 GNDA.n881 585
R21227 GNDA.n884 GNDA.n824 585
R21228 GNDA.n5029 GNDA.n5028 585
R21229 GNDA.n5028 GNDA.n5027 585
R21230 GNDA.n5005 GNDA.n943 585
R21231 GNDA.n5026 GNDA.n943 585
R21232 GNDA.n5006 GNDA.n4927 585
R21233 GNDA.n4927 GNDA.n945 585
R21234 GNDA.n5014 GNDA.n5013 585
R21235 GNDA.n5015 GNDA.n5014 585
R21236 GNDA.n4930 GNDA.n4928 585
R21237 GNDA.n4928 GNDA.n4926 585
R21238 GNDA.n4935 GNDA.n4934 585
R21239 GNDA.n4934 GNDA.n895 585
R21240 GNDA.n4932 GNDA.n894 585
R21241 GNDA.n5168 GNDA.n894 585
R21242 GNDA.n5171 GNDA.n5170 585
R21243 GNDA.n5170 GNDA.n5169 585
R21244 GNDA.n891 GNDA.n886 585
R21245 GNDA.n886 GNDA.n885 585
R21246 GNDA.n5181 GNDA.n5180 585
R21247 GNDA.n5182 GNDA.n5181 585
R21248 GNDA.n888 GNDA.n883 585
R21249 GNDA.n5183 GNDA.n883 585
R21250 GNDA.n5186 GNDA.n5185 585
R21251 GNDA.n5185 GNDA.n5184 585
R21252 GNDA.n5222 GNDA.n5221 585
R21253 GNDA.n5221 GNDA.n5220 585
R21254 GNDA.n881 GNDA.n880 585
R21255 GNDA.n880 GNDA.n823 585
R21256 GNDA.n879 GNDA.n872 585
R21257 GNDA.n879 GNDA.n878 585
R21258 GNDA.n741 GNDA.n739 585
R21259 GNDA.n5350 GNDA.n741 585
R21260 GNDA.n5364 GNDA.n5363 585
R21261 GNDA.n5363 GNDA.n5362 585
R21262 GNDA.n5351 GNDA.n742 585
R21263 GNDA.n5361 GNDA.n742 585
R21264 GNDA.n5359 GNDA.n5358 585
R21265 GNDA.n5360 GNDA.n5359 585
R21266 GNDA.n5354 GNDA.n716 585
R21267 GNDA.n716 GNDA.n714 585
R21268 GNDA.n5373 GNDA.n5372 585
R21269 GNDA.n5374 GNDA.n5373 585
R21270 GNDA.n718 GNDA.n717 585
R21271 GNDA.n717 GNDA.n715 585
R21272 GNDA.n5076 GNDA.n5075 585
R21273 GNDA.n5075 GNDA.n5074 585
R21274 GNDA.n5079 GNDA.n5072 585
R21275 GNDA.n5072 GNDA.n5071 585
R21276 GNDA.n5138 GNDA.n5137 585
R21277 GNDA.n5139 GNDA.n5138 585
R21278 GNDA.n818 GNDA.n815 585
R21279 GNDA.n5140 GNDA.n818 585
R21280 GNDA.n5222 GNDA.n814 585
R21281 GNDA.n814 GNDA.n813 585
R21282 GNDA.n5277 GNDA.n5276 585
R21283 GNDA.n5278 GNDA.n5277 585
R21284 GNDA.n811 GNDA.n809 585
R21285 GNDA.n5279 GNDA.n811 585
R21286 GNDA.n5293 GNDA.n5292 585
R21287 GNDA.n5292 GNDA.n5291 585
R21288 GNDA.n5280 GNDA.n812 585
R21289 GNDA.n5290 GNDA.n812 585
R21290 GNDA.n5288 GNDA.n5287 585
R21291 GNDA.n5289 GNDA.n5288 585
R21292 GNDA.n5283 GNDA.n777 585
R21293 GNDA.n777 GNDA.n771 585
R21294 GNDA.n5302 GNDA.n5301 585
R21295 GNDA.n5303 GNDA.n5302 585
R21296 GNDA.n779 GNDA.n778 585
R21297 GNDA.n778 GNDA.n776 585
R21298 GNDA.n789 GNDA.n788 585
R21299 GNDA.n788 GNDA.n787 585
R21300 GNDA.n790 GNDA.n754 585
R21301 GNDA.n754 GNDA.n752 585
R21302 GNDA.n5336 GNDA.n5335 585
R21303 GNDA.n5337 GNDA.n5336 585
R21304 GNDA.n5333 GNDA.n755 585
R21305 GNDA.n755 GNDA.n753 585
R21306 GNDA.n926 GNDA.n925 585
R21307 GNDA.n925 GNDA.n924 585
R21308 GNDA.n927 GNDA.n903 585
R21309 GNDA.n903 GNDA.n902 585
R21310 GNDA.n929 GNDA.n928 585
R21311 GNDA.n930 GNDA.n929 585
R21312 GNDA.n901 GNDA.n900 585
R21313 GNDA.n931 GNDA.n901 585
R21314 GNDA.n934 GNDA.n933 585
R21315 GNDA.n933 GNDA.n932 585
R21316 GNDA.n935 GNDA.n898 585
R21317 GNDA.n898 GNDA.n896 585
R21318 GNDA.n5040 GNDA.n5039 585
R21319 GNDA.n5041 GNDA.n5040 585
R21320 GNDA.n5038 GNDA.n899 585
R21321 GNDA.n899 GNDA.n897 585
R21322 GNDA.n5037 GNDA.n5036 585
R21323 GNDA.n5036 GNDA.n5035 585
R21324 GNDA.n937 GNDA.n936 585
R21325 GNDA.n5034 GNDA.n937 585
R21326 GNDA.n5032 GNDA.n5031 585
R21327 GNDA.n5033 GNDA.n5032 585
R21328 GNDA.n939 GNDA.n938 585
R21329 GNDA.n4914 GNDA.n942 585
R21330 GNDA.n4844 GNDA.n4843 585
R21331 GNDA.n4845 GNDA.n4844 585
R21332 GNDA.n4842 GNDA.n1177 585
R21333 GNDA.n1177 GNDA.n1175 585
R21334 GNDA.n4841 GNDA.n4840 585
R21335 GNDA.n4840 GNDA.n4839 585
R21336 GNDA.n1180 GNDA.n1179 585
R21337 GNDA.n4838 GNDA.n1180 585
R21338 GNDA.n4836 GNDA.n4835 585
R21339 GNDA.n4837 GNDA.n4836 585
R21340 GNDA.n4834 GNDA.n1182 585
R21341 GNDA.n1182 GNDA.n1181 585
R21342 GNDA.n4833 GNDA.n4832 585
R21343 GNDA.n4832 GNDA.n4831 585
R21344 GNDA.n1184 GNDA.n1183 585
R21345 GNDA.n4830 GNDA.n1184 585
R21346 GNDA.n4828 GNDA.n4827 585
R21347 GNDA.n4829 GNDA.n4828 585
R21348 GNDA.n4826 GNDA.n1187 585
R21349 GNDA.n1187 GNDA.n1186 585
R21350 GNDA.n4825 GNDA.n4824 585
R21351 GNDA.n4824 GNDA.n4823 585
R21352 GNDA.n4822 GNDA.n1189 585
R21353 GNDA.n4821 GNDA.n4820 585
R21354 GNDA.n1539 GNDA.n1538 585
R21355 GNDA.n1553 GNDA.n1539 585
R21356 GNDA.n1551 GNDA.n1550 585
R21357 GNDA.n1552 GNDA.n1551 585
R21358 GNDA.n1549 GNDA.n1541 585
R21359 GNDA.n1544 GNDA.n1541 585
R21360 GNDA.n1548 GNDA.n1547 585
R21361 GNDA.n1547 GNDA.n1546 585
R21362 GNDA.n1543 GNDA.n1542 585
R21363 GNDA.n1545 GNDA.n1543 585
R21364 GNDA.n1145 GNDA.n1143 585
R21365 GNDA.n1143 GNDA.n1141 585
R21366 GNDA.n4861 GNDA.n4860 585
R21367 GNDA.n4862 GNDA.n4861 585
R21368 GNDA.n4859 GNDA.n1144 585
R21369 GNDA.n1144 GNDA.n1142 585
R21370 GNDA.n4858 GNDA.n4857 585
R21371 GNDA.n4857 GNDA.n4856 585
R21372 GNDA.n1147 GNDA.n1146 585
R21373 GNDA.n4855 GNDA.n1147 585
R21374 GNDA.n4853 GNDA.n4852 585
R21375 GNDA.n4854 GNDA.n4853 585
R21376 GNDA.n1149 GNDA.n1148 585
R21377 GNDA.n1174 GNDA.n1152 585
R21378 GNDA.n4916 GNDA.n4915 585
R21379 GNDA.n4919 GNDA.n4913 585
R21380 GNDA.n4913 GNDA.n944 585
R21381 GNDA.n5508 GNDA.n641 582.4
R21382 GNDA.n5408 GNDA.n5407 582.4
R21383 GNDA.n644 GNDA.n643 548.082
R21384 GNDA.n699 GNDA.n698 546.375
R21385 GNDA.n662 GNDA.n661 546.375
R21386 GNDA.n5451 GNDA.n5450 546.375
R21387 GNDA.n3298 GNDA.n3297 524.808
R21388 GNDA.n3304 GNDA.n3303 524.808
R21389 GNDA.n4277 GNDA.n4276 524.808
R21390 GNDA.n4182 GNDA.n4181 524.808
R21391 GNDA.n5325 GNDA.n5324 511.728
R21392 GNDA.n5425 GNDA.n5424 509.2
R21393 GNDA.n5421 GNDA.n5420 509.2
R21394 GNDA.n617 GNDA.n616 509.034
R21395 GNDA.n614 GNDA.n613 509.034
R21396 GNDA.n5399 GNDA.n5398 492.675
R21397 GNDA.n5405 GNDA.n5404 492.675
R21398 GNDA.n633 GNDA.n632 492.675
R21399 GNDA.n639 GNDA.n638 492.675
R21400 GNDA.n4846 GNDA.n1172 486.94
R21401 GNDA.n1825 GNDA.n825 486.94
R21402 GNDA.n4846 GNDA.n1174 486.94
R21403 GNDA.n4821 GNDA.n825 486.94
R21404 GNDA.n5525 GNDA.n5524 483.2
R21405 GNDA.n5524 GNDA.n37 476.8
R21406 GNDA.n4915 GNDA.n944 438.685
R21407 GNDA.n748 GNDA.n747 425.134
R21408 GNDA.n5023 GNDA.n5022 425.134
R21409 GNDA.n624 GNDA.n620 415.557
R21410 GNDA.n4921 GNDA.n4920 409.067
R21411 GNDA.n5341 GNDA.n5340 409.067
R21412 GNDA.n750 GNDA.n749 409.067
R21413 GNDA.n5347 GNDA.n5346 409.067
R21414 GNDA.n875 GNDA.n874 409.067
R21415 GNDA.n5019 GNDA.n5018 409.067
R21416 GNDA.n4327 GNDA.n4287 394.817
R21417 GNDA.n4331 GNDA.n4329 394.817
R21418 GNDA.n4331 GNDA.n4330 394.817
R21419 GNDA.n4330 GNDA.n1139 394.817
R21420 GNDA.n4338 GNDA.n1140 394.817
R21421 GNDA.n4338 GNDA.n1959 394.817
R21422 GNDA.n4345 GNDA.n1959 394.817
R21423 GNDA.n4346 GNDA.n4345 394.817
R21424 GNDA.n4347 GNDA.n4346 394.817
R21425 GNDA.n4347 GNDA.n1172 394.817
R21426 GNDA.n1845 GNDA.n1171 394.817
R21427 GNDA.n1845 GNDA.n1844 394.817
R21428 GNDA.n1844 GNDA.n1843 394.817
R21429 GNDA.n1843 GNDA.n1697 394.817
R21430 GNDA.n1837 GNDA.n1697 394.817
R21431 GNDA.n1835 GNDA.n1834 394.817
R21432 GNDA.n1834 GNDA.n1833 394.817
R21433 GNDA.n1833 GNDA.n1702 394.817
R21434 GNDA.n1827 GNDA.n1702 394.817
R21435 GNDA.n1827 GNDA.n1826 394.817
R21436 GNDA.n1826 GNDA.n1825 394.817
R21437 GNDA.n1284 GNDA.n1283 394.817
R21438 GNDA.n1283 GNDA.n1282 394.817
R21439 GNDA.n1282 GNDA.n1263 394.817
R21440 GNDA.n1276 GNDA.n1263 394.817
R21441 GNDA.n1276 GNDA.n773 394.817
R21442 GNDA.n1268 GNDA.n774 394.817
R21443 GNDA.n1269 GNDA.n1268 394.817
R21444 GNDA.n1269 GNDA.n762 394.817
R21445 GNDA.n5329 GNDA.n762 394.817
R21446 GNDA.n5329 GNDA.n5328 394.817
R21447 GNDA.n5328 GNDA.n5327 394.817
R21448 GNDA.n1553 GNDA.n1552 394.817
R21449 GNDA.n1546 GNDA.n1544 394.817
R21450 GNDA.n1546 GNDA.n1545 394.817
R21451 GNDA.n1545 GNDA.n1141 394.817
R21452 GNDA.n4862 GNDA.n1142 394.817
R21453 GNDA.n4856 GNDA.n1142 394.817
R21454 GNDA.n4856 GNDA.n4855 394.817
R21455 GNDA.n4855 GNDA.n4854 394.817
R21456 GNDA.n4854 GNDA.n1148 394.817
R21457 GNDA.n1174 GNDA.n1148 394.817
R21458 GNDA.n4845 GNDA.n1175 394.817
R21459 GNDA.n4839 GNDA.n1175 394.817
R21460 GNDA.n4839 GNDA.n4838 394.817
R21461 GNDA.n4838 GNDA.n4837 394.817
R21462 GNDA.n4837 GNDA.n1181 394.817
R21463 GNDA.n4831 GNDA.n4830 394.817
R21464 GNDA.n4830 GNDA.n4829 394.817
R21465 GNDA.n4829 GNDA.n1186 394.817
R21466 GNDA.n4823 GNDA.n1186 394.817
R21467 GNDA.n4823 GNDA.n4822 394.817
R21468 GNDA.n4822 GNDA.n4821 394.817
R21469 GNDA.n924 GNDA.n902 394.817
R21470 GNDA.n930 GNDA.n902 394.817
R21471 GNDA.n931 GNDA.n930 394.817
R21472 GNDA.n932 GNDA.n931 394.817
R21473 GNDA.n932 GNDA.n896 394.817
R21474 GNDA.n5041 GNDA.n897 394.817
R21475 GNDA.n5035 GNDA.n897 394.817
R21476 GNDA.n5035 GNDA.n5034 394.817
R21477 GNDA.n5034 GNDA.n5033 394.817
R21478 GNDA.n5033 GNDA.n938 394.817
R21479 GNDA.n4914 GNDA.n938 394.817
R21480 GNDA.n5518 GNDA.n5517 384
R21481 GNDA.n4328 GNDA.n4327 377.269
R21482 GNDA.n1552 GNDA.n1540 377.269
R21483 GNDA.n5216 GNDA.n712 370.214
R21484 GNDA.n4864 GNDA.n1129 370.214
R21485 GNDA.n1580 GNDA.n1137 370.214
R21486 GNDA.n4621 GNDA.n4620 370.214
R21487 GNDA.n4621 GNDA.n1380 370.214
R21488 GNDA.n5216 GNDA.n775 370.214
R21489 GNDA.n5216 GNDA.n822 365.957
R21490 GNDA.n1135 GNDA.n1129 365.957
R21491 GNDA.n1580 GNDA.n1136 365.957
R21492 GNDA.n4621 GNDA.n1389 365.957
R21493 GNDA.n4622 GNDA.n4621 365.957
R21494 GNDA.n5216 GNDA.n713 365.957
R21495 GNDA.n5519 GNDA.n5518 355.2
R21496 GNDA.n5517 GNDA.n623 345.601
R21497 GNDA.n5317 GNDA.n768 335
R21498 GNDA.n5310 GNDA.n5309 335
R21499 GNDA.n5158 GNDA.n5156 335
R21500 GNDA.n5042 GNDA.n822 327.661
R21501 GNDA.n4863 GNDA.n1135 327.661
R21502 GNDA.n4863 GNDA.n1136 327.661
R21503 GNDA.n1389 GNDA.n1185 327.661
R21504 GNDA.n4622 GNDA.n1185 327.661
R21505 GNDA.n5375 GNDA.n713 327.661
R21506 GNDA.n5375 GNDA.n712 323.404
R21507 GNDA.n4864 GNDA.n4863 323.404
R21508 GNDA.n4863 GNDA.n1137 323.404
R21509 GNDA.n4620 GNDA.n1185 323.404
R21510 GNDA.n1380 GNDA.n1185 323.404
R21511 GNDA.n5304 GNDA.n775 323.404
R21512 GNDA.n5519 GNDA.n623 316.8
R21513 GNDA.n620 GNDA.n619 293.651
R21514 GNDA.n620 GNDA.n615 293.651
R21515 GNDA.n5518 GNDA.n622 292.5
R21516 GNDA.n624 GNDA.n622 292.5
R21517 GNDA.n5517 GNDA.n5516 292.5
R21518 GNDA.n5516 GNDA.n5515 292.5
R21519 GNDA.n623 GNDA.n621 292.5
R21520 GNDA.n624 GNDA.n621 292.5
R21521 GNDA.n5520 GNDA.n5519 292.5
R21522 GNDA.n5521 GNDA.n5520 292.5
R21523 GNDA.n5524 GNDA.n5523 292.5
R21524 GNDA.n5523 GNDA.n5522 292.5
R21525 GNDA.n593 GNDA.n592 292.5
R21526 GNDA.n592 GNDA.n40 292.5
R21527 GNDA.n5397 GNDA.n629 292.5
R21528 GNDA.n670 GNDA.n629 292.5
R21529 GNDA.n702 GNDA.n628 292.5
R21530 GNDA.n671 GNDA.n628 292.5
R21531 GNDA.n5457 GNDA.n5456 292.5
R21532 GNDA.n5456 GNDA.n672 292.5
R21533 GNDA.n5464 GNDA.n5463 292.5
R21534 GNDA.n5465 GNDA.n5464 292.5
R21535 GNDA.n5477 GNDA.n5476 292.5
R21536 GNDA.n668 GNDA.n666 292.5
R21537 GNDA.n5466 GNDA.n668 292.5
R21538 GNDA.n5473 GNDA.n5472 292.5
R21539 GNDA.n5474 GNDA.n5473 292.5
R21540 GNDA.n669 GNDA.n667 292.5
R21541 GNDA.n591 GNDA.n39 292.5
R21542 GNDA.n5512 GNDA.n39 292.5
R21543 GNDA.n5510 GNDA.n5509 292.5
R21544 GNDA.n5511 GNDA.n5510 292.5
R21545 GNDA.n676 GNDA.n674 292.5
R21546 GNDA.n674 GNDA.n627 292.5
R21547 GNDA.n594 GNDA.n38 292.5
R21548 GNDA.n5393 GNDA.n38 292.5
R21549 GNDA.n5396 GNDA.n5395 292.5
R21550 GNDA.n5395 GNDA.n5394 292.5
R21551 GNDA.n677 GNDA.n673 292.5
R21552 GNDA.n5392 GNDA.n673 292.5
R21553 GNDA.n5154 GNDA.n5153 288.277
R21554 GNDA.n5163 GNDA.n5153 288.277
R21555 GNDA.n5312 GNDA.n769 267.865
R21556 GNDA.n5312 GNDA.n5311 267.865
R21557 GNDA.n5162 GNDA.n5161 267.865
R21558 GNDA.n4863 GNDA.n1139 267.598
R21559 GNDA.n1837 GNDA.n1185 267.598
R21560 GNDA.n5304 GNDA.n773 267.598
R21561 GNDA.n4863 GNDA.n1141 267.598
R21562 GNDA.n1185 GNDA.n1181 267.598
R21563 GNDA.n5042 GNDA.n896 267.598
R21564 GNDA.n5332 GNDA.n758 264.301
R21565 GNDA.n1823 GNDA.n1705 264.301
R21566 GNDA.n4349 GNDA.n1957 264.301
R21567 GNDA.n5030 GNDA.n940 264.301
R21568 GNDA.n1190 GNDA.n1188 264.301
R21569 GNDA.n4851 GNDA.n1150 264.301
R21570 GNDA.n1286 GNDA.n1285 259.416
R21571 GNDA.n1331 GNDA.n1330 259.416
R21572 GNDA.n5213 GNDA.n844 259.416
R21573 GNDA.n1125 GNDA.n1123 259.416
R21574 GNDA.n1598 GNDA.n1524 259.416
R21575 GNDA.n1848 GNDA.n1847 259.416
R21576 GNDA.n1684 GNDA.n1683 259.416
R21577 GNDA.n4577 GNDA.n4576 259.416
R21578 GNDA.n4322 GNDA.n4288 259.416
R21579 GNDA.n5258 GNDA.n5257 258.334
R21580 GNDA.n5099 GNDA.n5098 258.334
R21581 GNDA.n4689 GNDA.n1257 258.334
R21582 GNDA.n1456 GNDA.n1455 258.334
R21583 GNDA.n1765 GNDA.n1764 258.334
R21584 GNDA.n4791 GNDA.n4790 258.334
R21585 GNDA.n4517 GNDA.n4516 258.334
R21586 GNDA.n4987 GNDA.n4942 258.334
R21587 GNDA.n4418 GNDA.n4417 258.334
R21588 GNDA.n4881 GNDA.n1116 257.779
R21589 GNDA.n4549 GNDA.n1173 254.34
R21590 GNDA.n4571 GNDA.n1173 254.34
R21591 GNDA.n4565 GNDA.n1173 254.34
R21592 GNDA.n4563 GNDA.n1173 254.34
R21593 GNDA.n4557 GNDA.n1173 254.34
R21594 GNDA.n4555 GNDA.n1173 254.34
R21595 GNDA.n1682 GNDA.n1173 254.34
R21596 GNDA.n1676 GNDA.n1173 254.34
R21597 GNDA.n1674 GNDA.n1173 254.34
R21598 GNDA.n1668 GNDA.n1173 254.34
R21599 GNDA.n1666 GNDA.n1173 254.34
R21600 GNDA.n1661 GNDA.n1173 254.34
R21601 GNDA.n1694 GNDA.n1173 254.34
R21602 GNDA.n1853 GNDA.n1173 254.34
R21603 GNDA.n1691 GNDA.n1173 254.34
R21604 GNDA.n1860 GNDA.n1173 254.34
R21605 GNDA.n1688 GNDA.n1173 254.34
R21606 GNDA.n1867 GNDA.n1173 254.34
R21607 GNDA.n4847 GNDA.n1170 254.34
R21608 GNDA.n4847 GNDA.n1169 254.34
R21609 GNDA.n4847 GNDA.n1168 254.34
R21610 GNDA.n4847 GNDA.n1167 254.34
R21611 GNDA.n4847 GNDA.n1166 254.34
R21612 GNDA.n4847 GNDA.n1165 254.34
R21613 GNDA.n4848 GNDA.n4847 254.34
R21614 GNDA.n4847 GNDA.n1164 254.34
R21615 GNDA.n4847 GNDA.n1163 254.34
R21616 GNDA.n4847 GNDA.n1162 254.34
R21617 GNDA.n4847 GNDA.n1161 254.34
R21618 GNDA.n4847 GNDA.n1160 254.34
R21619 GNDA.n1626 GNDA.n1136 254.34
R21620 GNDA.n1623 GNDA.n1136 254.34
R21621 GNDA.n1613 GNDA.n1136 254.34
R21622 GNDA.n1611 GNDA.n1136 254.34
R21623 GNDA.n1601 GNDA.n1136 254.34
R21624 GNDA.n1599 GNDA.n1136 254.34
R21625 GNDA.n1595 GNDA.n1137 254.34
R21626 GNDA.n1605 GNDA.n1137 254.34
R21627 GNDA.n1607 GNDA.n1137 254.34
R21628 GNDA.n1617 GNDA.n1137 254.34
R21629 GNDA.n1619 GNDA.n1137 254.34
R21630 GNDA.n1630 GNDA.n1137 254.34
R21631 GNDA.n4593 GNDA.n1389 254.34
R21632 GNDA.n4590 GNDA.n1389 254.34
R21633 GNDA.n4587 GNDA.n1389 254.34
R21634 GNDA.n4584 GNDA.n1389 254.34
R21635 GNDA.n4581 GNDA.n1389 254.34
R21636 GNDA.n4578 GNDA.n1389 254.34
R21637 GNDA.n4620 GNDA.n4619 254.34
R21638 GNDA.n4620 GNDA.n1394 254.34
R21639 GNDA.n4620 GNDA.n1393 254.34
R21640 GNDA.n4620 GNDA.n1392 254.34
R21641 GNDA.n4620 GNDA.n1391 254.34
R21642 GNDA.n4620 GNDA.n1390 254.34
R21643 GNDA.n870 GNDA.n822 254.34
R21644 GNDA.n867 GNDA.n822 254.34
R21645 GNDA.n862 GNDA.n822 254.34
R21646 GNDA.n859 GNDA.n822 254.34
R21647 GNDA.n854 GNDA.n822 254.34
R21648 GNDA.n851 GNDA.n822 254.34
R21649 GNDA.n5208 GNDA.n712 254.34
R21650 GNDA.n5201 GNDA.n712 254.34
R21651 GNDA.n5199 GNDA.n712 254.34
R21652 GNDA.n5193 GNDA.n712 254.34
R21653 GNDA.n5191 GNDA.n712 254.34
R21654 GNDA.n5215 GNDA.n5214 254.34
R21655 GNDA.n5215 GNDA.n842 254.34
R21656 GNDA.n5215 GNDA.n841 254.34
R21657 GNDA.n5215 GNDA.n840 254.34
R21658 GNDA.n5215 GNDA.n839 254.34
R21659 GNDA.n5215 GNDA.n838 254.34
R21660 GNDA.n5215 GNDA.n837 254.34
R21661 GNDA.n5215 GNDA.n836 254.34
R21662 GNDA.n5215 GNDA.n835 254.34
R21663 GNDA.n5215 GNDA.n834 254.34
R21664 GNDA.n5215 GNDA.n833 254.34
R21665 GNDA.n5215 GNDA.n832 254.34
R21666 GNDA.n5215 GNDA.n831 254.34
R21667 GNDA.n5215 GNDA.n830 254.34
R21668 GNDA.n5215 GNDA.n829 254.34
R21669 GNDA.n5215 GNDA.n828 254.34
R21670 GNDA.n5215 GNDA.n827 254.34
R21671 GNDA.n5215 GNDA.n826 254.34
R21672 GNDA.n4749 GNDA.n1191 254.34
R21673 GNDA.n4749 GNDA.n1194 254.34
R21674 GNDA.n4749 GNDA.n4748 254.34
R21675 GNDA.n4749 GNDA.n4725 254.34
R21676 GNDA.n4749 GNDA.n4724 254.34
R21677 GNDA.n4750 GNDA.n4749 254.34
R21678 GNDA.n4749 GNDA.n4723 254.34
R21679 GNDA.n4749 GNDA.n1229 254.34
R21680 GNDA.n4749 GNDA.n1228 254.34
R21681 GNDA.n4749 GNDA.n1227 254.34
R21682 GNDA.n4749 GNDA.n1226 254.34
R21683 GNDA.n4749 GNDA.n1225 254.34
R21684 GNDA.n4749 GNDA.n1224 254.34
R21685 GNDA.n4749 GNDA.n1223 254.34
R21686 GNDA.n4749 GNDA.n1222 254.34
R21687 GNDA.n4749 GNDA.n1221 254.34
R21688 GNDA.n4749 GNDA.n1220 254.34
R21689 GNDA.n4749 GNDA.n1219 254.34
R21690 GNDA.n4847 GNDA.n1159 254.34
R21691 GNDA.n4847 GNDA.n1158 254.34
R21692 GNDA.n4847 GNDA.n1157 254.34
R21693 GNDA.n4847 GNDA.n1156 254.34
R21694 GNDA.n4847 GNDA.n1155 254.34
R21695 GNDA.n4847 GNDA.n1154 254.34
R21696 GNDA.n1929 GNDA.n1135 254.34
R21697 GNDA.n1927 GNDA.n1135 254.34
R21698 GNDA.n1917 GNDA.n1135 254.34
R21699 GNDA.n1915 GNDA.n1135 254.34
R21700 GNDA.n1906 GNDA.n1135 254.34
R21701 GNDA.n1904 GNDA.n1135 254.34
R21702 GNDA.n4865 GNDA.n4864 254.34
R21703 GNDA.n4864 GNDA.n1134 254.34
R21704 GNDA.n4864 GNDA.n1133 254.34
R21705 GNDA.n4864 GNDA.n1132 254.34
R21706 GNDA.n4864 GNDA.n1131 254.34
R21707 GNDA.n4864 GNDA.n1130 254.34
R21708 GNDA.n4623 GNDA.n4622 254.34
R21709 GNDA.n4622 GNDA.n1388 254.34
R21710 GNDA.n4622 GNDA.n1387 254.34
R21711 GNDA.n4622 GNDA.n1386 254.34
R21712 GNDA.n4622 GNDA.n1385 254.34
R21713 GNDA.n4622 GNDA.n1384 254.34
R21714 GNDA.n1896 GNDA.n1380 254.34
R21715 GNDA.n1869 GNDA.n1380 254.34
R21716 GNDA.n1889 GNDA.n1380 254.34
R21717 GNDA.n1883 GNDA.n1380 254.34
R21718 GNDA.n1881 GNDA.n1380 254.34
R21719 GNDA.n4627 GNDA.n1380 254.34
R21720 GNDA.n1353 GNDA.n713 254.34
R21721 GNDA.n1351 GNDA.n713 254.34
R21722 GNDA.n1346 GNDA.n713 254.34
R21723 GNDA.n1343 GNDA.n713 254.34
R21724 GNDA.n1338 GNDA.n713 254.34
R21725 GNDA.n1335 GNDA.n713 254.34
R21726 GNDA.n1374 GNDA.n775 254.34
R21727 GNDA.n1367 GNDA.n775 254.34
R21728 GNDA.n1365 GNDA.n775 254.34
R21729 GNDA.n1359 GNDA.n775 254.34
R21730 GNDA.n1357 GNDA.n775 254.34
R21731 GNDA.n5058 GNDA.n743 250.349
R21732 GNDA.n5143 GNDA.n5142 250.349
R21733 GNDA.n1375 GNDA.n1333 249.663
R21734 GNDA.n5209 GNDA.n849 249.663
R21735 GNDA.n925 GNDA.n923 249.663
R21736 GNDA.n1596 GNDA.n1594 249.663
R21737 GNDA.n1555 GNDA.n1539 249.663
R21738 GNDA.n1897 GNDA.n1868 249.663
R21739 GNDA.n4618 GNDA.n1396 249.663
R21740 GNDA.n4844 GNDA.n1176 249.663
R21741 GNDA.n4866 GNDA.n1127 249.663
R21742 GNDA.n5477 GNDA.n667 249.601
R21743 GNDA.n5472 GNDA.n667 249.601
R21744 GNDA.n5314 GNDA.n770 246.25
R21745 GNDA.n5314 GNDA.n5305 246.25
R21746 GNDA.n5045 GNDA.n5044 246.25
R21747 GNDA.n5159 GNDA.n5044 246.25
R21748 GNDA.n4916 GNDA.n4913 246.25
R21749 GNDA.n5167 GNDA.n5166 241.643
R21750 GNDA.n5167 GNDA.n5043 241.643
R21751 GNDA.n5316 GNDA.n5315 241.643
R21752 GNDA.n5315 GNDA.n772 241.643
R21753 GNDA.n5515 GNDA.n5514 207.779
R21754 GNDA.n5476 GNDA.n5475 202.423
R21755 GNDA.n5144 GNDA.n5070 197
R21756 GNDA.n5060 GNDA.n5059 197
R21757 GNDA.n5326 GNDA.n755 197
R21758 GNDA.n5221 GNDA.n818 197
R21759 GNDA.n5185 GNDA.n884 197
R21760 GNDA.n1512 GNDA.n1511 197
R21761 GNDA.n1824 GNDA.n1822 197
R21762 GNDA.n4632 GNDA.n4631 197
R21763 GNDA.n4594 GNDA.n1217 197
R21764 GNDA.n4450 GNDA.n4449 197
R21765 GNDA.n4351 GNDA.n4350 197
R21766 GNDA.n5277 GNDA.n814 187.249
R21767 GNDA.n880 GNDA.n879 187.249
R21768 GNDA.n5028 GNDA.n942 187.249
R21769 GNDA.n4849 GNDA.n1152 187.249
R21770 GNDA.n4629 GNDA.n1378 187.249
R21771 GNDA.n4722 GNDA.n1231 187.249
R21772 GNDA.n4820 GNDA.n4819 187.249
R21773 GNDA.n4546 GNDA.n4545 187.249
R21774 GNDA.n4447 GNDA.n4446 187.249
R21775 GNDA.n5259 GNDA.n5258 185
R21776 GNDA.n5261 GNDA.n5260 185
R21777 GNDA.n5263 GNDA.n5262 185
R21778 GNDA.n5265 GNDA.n5264 185
R21779 GNDA.n5267 GNDA.n5266 185
R21780 GNDA.n5269 GNDA.n5268 185
R21781 GNDA.n5271 GNDA.n5270 185
R21782 GNDA.n5273 GNDA.n5272 185
R21783 GNDA.n5274 GNDA.n807 185
R21784 GNDA.n5241 GNDA.n5240 185
R21785 GNDA.n5243 GNDA.n5242 185
R21786 GNDA.n5245 GNDA.n5244 185
R21787 GNDA.n5247 GNDA.n5246 185
R21788 GNDA.n5249 GNDA.n5248 185
R21789 GNDA.n5251 GNDA.n5250 185
R21790 GNDA.n5253 GNDA.n5252 185
R21791 GNDA.n5255 GNDA.n5254 185
R21792 GNDA.n5257 GNDA.n5256 185
R21793 GNDA.n799 GNDA.n757 185
R21794 GNDA.n5225 GNDA.n5224 185
R21795 GNDA.n5227 GNDA.n5226 185
R21796 GNDA.n5229 GNDA.n5228 185
R21797 GNDA.n5231 GNDA.n5230 185
R21798 GNDA.n5233 GNDA.n5232 185
R21799 GNDA.n5235 GNDA.n5234 185
R21800 GNDA.n5237 GNDA.n5236 185
R21801 GNDA.n5239 GNDA.n5238 185
R21802 GNDA.n798 GNDA.n756 185
R21803 GNDA.n792 GNDA.n791 185
R21804 GNDA.n786 GNDA.n781 185
R21805 GNDA.n5300 GNDA.n5299 185
R21806 GNDA.n5282 GNDA.n780 185
R21807 GNDA.n5286 GNDA.n5285 185
R21808 GNDA.n5284 GNDA.n5281 185
R21809 GNDA.n810 GNDA.n808 185
R21810 GNDA.n5295 GNDA.n5294 185
R21811 GNDA.n5098 GNDA.n5097 185
R21812 GNDA.n5096 GNDA.n5095 185
R21813 GNDA.n5094 GNDA.n5093 185
R21814 GNDA.n5092 GNDA.n5091 185
R21815 GNDA.n5090 GNDA.n5089 185
R21816 GNDA.n5088 GNDA.n5087 185
R21817 GNDA.n5086 GNDA.n5085 185
R21818 GNDA.n5084 GNDA.n5083 185
R21819 GNDA.n5082 GNDA.n737 185
R21820 GNDA.n5116 GNDA.n5115 185
R21821 GNDA.n5114 GNDA.n5113 185
R21822 GNDA.n5112 GNDA.n5111 185
R21823 GNDA.n5110 GNDA.n5109 185
R21824 GNDA.n5108 GNDA.n5107 185
R21825 GNDA.n5106 GNDA.n5105 185
R21826 GNDA.n5104 GNDA.n5103 185
R21827 GNDA.n5102 GNDA.n5101 185
R21828 GNDA.n5100 GNDA.n5099 185
R21829 GNDA.n5135 GNDA.n5134 185
R21830 GNDA.n5132 GNDA.n5131 185
R21831 GNDA.n5130 GNDA.n5129 185
R21832 GNDA.n5128 GNDA.n5127 185
R21833 GNDA.n5126 GNDA.n5125 185
R21834 GNDA.n5124 GNDA.n5123 185
R21835 GNDA.n5122 GNDA.n5121 185
R21836 GNDA.n5120 GNDA.n5119 185
R21837 GNDA.n5118 GNDA.n5117 185
R21838 GNDA.n5133 GNDA.n5080 185
R21839 GNDA.n5078 GNDA.n5077 185
R21840 GNDA.n5073 GNDA.n720 185
R21841 GNDA.n5371 GNDA.n5370 185
R21842 GNDA.n5353 GNDA.n719 185
R21843 GNDA.n5357 GNDA.n5356 185
R21844 GNDA.n5355 GNDA.n5352 185
R21845 GNDA.n740 GNDA.n738 185
R21846 GNDA.n5366 GNDA.n5365 185
R21847 GNDA.n4691 GNDA.n1257 185
R21848 GNDA.n4705 GNDA.n4704 185
R21849 GNDA.n4703 GNDA.n1258 185
R21850 GNDA.n4702 GNDA.n4701 185
R21851 GNDA.n4700 GNDA.n4699 185
R21852 GNDA.n4698 GNDA.n4697 185
R21853 GNDA.n4696 GNDA.n4695 185
R21854 GNDA.n4694 GNDA.n4693 185
R21855 GNDA.n4692 GNDA.n1234 185
R21856 GNDA.n4674 GNDA.n4673 185
R21857 GNDA.n4676 GNDA.n4675 185
R21858 GNDA.n4678 GNDA.n4677 185
R21859 GNDA.n4680 GNDA.n4679 185
R21860 GNDA.n4682 GNDA.n4681 185
R21861 GNDA.n4684 GNDA.n4683 185
R21862 GNDA.n4686 GNDA.n4685 185
R21863 GNDA.n4688 GNDA.n4687 185
R21864 GNDA.n4690 GNDA.n4689 185
R21865 GNDA.n4656 GNDA.n4655 185
R21866 GNDA.n4658 GNDA.n4657 185
R21867 GNDA.n4660 GNDA.n4659 185
R21868 GNDA.n4662 GNDA.n4661 185
R21869 GNDA.n4664 GNDA.n4663 185
R21870 GNDA.n4666 GNDA.n4665 185
R21871 GNDA.n4668 GNDA.n4667 185
R21872 GNDA.n4670 GNDA.n4669 185
R21873 GNDA.n4672 GNDA.n4671 185
R21874 GNDA.n4654 GNDA.n4653 185
R21875 GNDA.n4648 GNDA.n4647 185
R21876 GNDA.n4646 GNDA.n4645 185
R21877 GNDA.n4641 GNDA.n4640 185
R21878 GNDA.n4636 GNDA.n1242 185
R21879 GNDA.n4710 GNDA.n4709 185
R21880 GNDA.n1241 GNDA.n1239 185
R21881 GNDA.n4716 GNDA.n4715 185
R21882 GNDA.n4718 GNDA.n4717 185
R21883 GNDA.n5313 GNDA.n5312 185
R21884 GNDA.n5306 GNDA.n768 185
R21885 GNDA.n5313 GNDA.n5307 185
R21886 GNDA.n5309 GNDA.n5308 185
R21887 GNDA.n5164 GNDA.n5163 185
R21888 GNDA.n5162 GNDA.n5155 185
R21889 GNDA.n5164 GNDA.n5154 185
R21890 GNDA.n5157 GNDA.n5155 185
R21891 GNDA.n5160 GNDA.n5158 185
R21892 GNDA.n1457 GNDA.n1456 185
R21893 GNDA.n1459 GNDA.n1458 185
R21894 GNDA.n1461 GNDA.n1460 185
R21895 GNDA.n1463 GNDA.n1462 185
R21896 GNDA.n1465 GNDA.n1464 185
R21897 GNDA.n1467 GNDA.n1466 185
R21898 GNDA.n1469 GNDA.n1468 185
R21899 GNDA.n1470 GNDA.n1421 185
R21900 GNDA.n1472 GNDA.n1471 185
R21901 GNDA.n1439 GNDA.n1438 185
R21902 GNDA.n1441 GNDA.n1440 185
R21903 GNDA.n1443 GNDA.n1442 185
R21904 GNDA.n1445 GNDA.n1444 185
R21905 GNDA.n1447 GNDA.n1446 185
R21906 GNDA.n1449 GNDA.n1448 185
R21907 GNDA.n1451 GNDA.n1450 185
R21908 GNDA.n1453 GNDA.n1452 185
R21909 GNDA.n1455 GNDA.n1454 185
R21910 GNDA.n1413 GNDA.n1399 185
R21911 GNDA.n1423 GNDA.n1422 185
R21912 GNDA.n1425 GNDA.n1424 185
R21913 GNDA.n1427 GNDA.n1426 185
R21914 GNDA.n1429 GNDA.n1428 185
R21915 GNDA.n1431 GNDA.n1430 185
R21916 GNDA.n1433 GNDA.n1432 185
R21917 GNDA.n1435 GNDA.n1434 185
R21918 GNDA.n1437 GNDA.n1436 185
R21919 GNDA.n1766 GNDA.n1765 185
R21920 GNDA.n1768 GNDA.n1767 185
R21921 GNDA.n1770 GNDA.n1769 185
R21922 GNDA.n1772 GNDA.n1771 185
R21923 GNDA.n1774 GNDA.n1773 185
R21924 GNDA.n1776 GNDA.n1775 185
R21925 GNDA.n1778 GNDA.n1777 185
R21926 GNDA.n1780 GNDA.n1779 185
R21927 GNDA.n1781 GNDA.n1729 185
R21928 GNDA.n1748 GNDA.n1747 185
R21929 GNDA.n1750 GNDA.n1749 185
R21930 GNDA.n1752 GNDA.n1751 185
R21931 GNDA.n1754 GNDA.n1753 185
R21932 GNDA.n1756 GNDA.n1755 185
R21933 GNDA.n1758 GNDA.n1757 185
R21934 GNDA.n1760 GNDA.n1759 185
R21935 GNDA.n1762 GNDA.n1761 185
R21936 GNDA.n1764 GNDA.n1763 185
R21937 GNDA.n1721 GNDA.n1707 185
R21938 GNDA.n1732 GNDA.n1731 185
R21939 GNDA.n1734 GNDA.n1733 185
R21940 GNDA.n1736 GNDA.n1735 185
R21941 GNDA.n1738 GNDA.n1737 185
R21942 GNDA.n1740 GNDA.n1739 185
R21943 GNDA.n1742 GNDA.n1741 185
R21944 GNDA.n1744 GNDA.n1743 185
R21945 GNDA.n1746 GNDA.n1745 185
R21946 GNDA.n1711 GNDA.n1708 185
R21947 GNDA.n1815 GNDA.n1814 185
R21948 GNDA.n1787 GNDA.n1710 185
R21949 GNDA.n1793 GNDA.n1792 185
R21950 GNDA.n1791 GNDA.n1786 185
R21951 GNDA.n1800 GNDA.n1799 185
R21952 GNDA.n1798 GNDA.n1785 185
R21953 GNDA.n1805 GNDA.n1730 185
R21954 GNDA.n1810 GNDA.n1809 185
R21955 GNDA.n4792 GNDA.n4791 185
R21956 GNDA.n4794 GNDA.n4793 185
R21957 GNDA.n4796 GNDA.n4795 185
R21958 GNDA.n4798 GNDA.n4797 185
R21959 GNDA.n4800 GNDA.n4799 185
R21960 GNDA.n4802 GNDA.n4801 185
R21961 GNDA.n4804 GNDA.n4803 185
R21962 GNDA.n4806 GNDA.n4805 185
R21963 GNDA.n4807 GNDA.n1192 185
R21964 GNDA.n4774 GNDA.n4773 185
R21965 GNDA.n4776 GNDA.n4775 185
R21966 GNDA.n4778 GNDA.n4777 185
R21967 GNDA.n4780 GNDA.n4779 185
R21968 GNDA.n4782 GNDA.n4781 185
R21969 GNDA.n4784 GNDA.n4783 185
R21970 GNDA.n4786 GNDA.n4785 185
R21971 GNDA.n4788 GNDA.n4787 185
R21972 GNDA.n4790 GNDA.n4789 185
R21973 GNDA.n4756 GNDA.n4755 185
R21974 GNDA.n4758 GNDA.n4757 185
R21975 GNDA.n4760 GNDA.n4759 185
R21976 GNDA.n4762 GNDA.n4761 185
R21977 GNDA.n4764 GNDA.n4763 185
R21978 GNDA.n4766 GNDA.n4765 185
R21979 GNDA.n4768 GNDA.n4767 185
R21980 GNDA.n4770 GNDA.n4769 185
R21981 GNDA.n4772 GNDA.n4771 185
R21982 GNDA.n4754 GNDA.n4753 185
R21983 GNDA.n4734 GNDA.n4733 185
R21984 GNDA.n4732 GNDA.n4731 185
R21985 GNDA.n4740 GNDA.n4739 185
R21986 GNDA.n4742 GNDA.n4741 185
R21987 GNDA.n4745 GNDA.n4744 185
R21988 GNDA.n4728 GNDA.n1197 185
R21989 GNDA.n4812 GNDA.n4811 185
R21990 GNDA.n1196 GNDA.n1193 185
R21991 GNDA.n4518 GNDA.n4517 185
R21992 GNDA.n4520 GNDA.n4519 185
R21993 GNDA.n4522 GNDA.n4521 185
R21994 GNDA.n4524 GNDA.n4523 185
R21995 GNDA.n4526 GNDA.n4525 185
R21996 GNDA.n4528 GNDA.n4527 185
R21997 GNDA.n4530 GNDA.n4529 185
R21998 GNDA.n4532 GNDA.n4531 185
R21999 GNDA.n4533 GNDA.n1632 185
R22000 GNDA.n4500 GNDA.n4499 185
R22001 GNDA.n4502 GNDA.n4501 185
R22002 GNDA.n4504 GNDA.n4503 185
R22003 GNDA.n4506 GNDA.n4505 185
R22004 GNDA.n4508 GNDA.n4507 185
R22005 GNDA.n4510 GNDA.n4509 185
R22006 GNDA.n4512 GNDA.n4511 185
R22007 GNDA.n4514 GNDA.n4513 185
R22008 GNDA.n4516 GNDA.n4515 185
R22009 GNDA.n4482 GNDA.n4481 185
R22010 GNDA.n4484 GNDA.n4483 185
R22011 GNDA.n4486 GNDA.n4485 185
R22012 GNDA.n4488 GNDA.n4487 185
R22013 GNDA.n4490 GNDA.n4489 185
R22014 GNDA.n4492 GNDA.n4491 185
R22015 GNDA.n4494 GNDA.n4493 185
R22016 GNDA.n4496 GNDA.n4495 185
R22017 GNDA.n4498 GNDA.n4497 185
R22018 GNDA.n4480 GNDA.n4479 185
R22019 GNDA.n4474 GNDA.n4473 185
R22020 GNDA.n4472 GNDA.n4471 185
R22021 GNDA.n4467 GNDA.n4466 185
R22022 GNDA.n4465 GNDA.n4464 185
R22023 GNDA.n4459 GNDA.n4458 185
R22024 GNDA.n4454 GNDA.n1636 185
R22025 GNDA.n4538 GNDA.n4537 185
R22026 GNDA.n1635 GNDA.n1633 185
R22027 GNDA.n1403 GNDA.n1400 185
R22028 GNDA.n1504 GNDA.n1503 185
R22029 GNDA.n1477 GNDA.n1402 185
R22030 GNDA.n1483 GNDA.n1482 185
R22031 GNDA.n1481 GNDA.n1476 185
R22032 GNDA.n1490 GNDA.n1489 185
R22033 GNDA.n1488 GNDA.n1475 185
R22034 GNDA.n1495 GNDA.n1473 185
R22035 GNDA.n1499 GNDA.n1498 185
R22036 GNDA.n4987 GNDA.n4986 185
R22037 GNDA.n4989 GNDA.n4941 185
R22038 GNDA.n4992 GNDA.n4991 185
R22039 GNDA.n4993 GNDA.n4940 185
R22040 GNDA.n4995 GNDA.n4994 185
R22041 GNDA.n4997 GNDA.n4939 185
R22042 GNDA.n5000 GNDA.n4999 185
R22043 GNDA.n5001 GNDA.n4938 185
R22044 GNDA.n5003 GNDA.n5002 185
R22045 GNDA.n4969 GNDA.n4946 185
R22046 GNDA.n4971 GNDA.n4970 185
R22047 GNDA.n4973 GNDA.n4945 185
R22048 GNDA.n4976 GNDA.n4975 185
R22049 GNDA.n4977 GNDA.n4944 185
R22050 GNDA.n4979 GNDA.n4978 185
R22051 GNDA.n4981 GNDA.n4943 185
R22052 GNDA.n4984 GNDA.n4983 185
R22053 GNDA.n4985 GNDA.n4942 185
R22054 GNDA.n4953 GNDA.n889 185
R22055 GNDA.n4954 GNDA.n4952 185
R22056 GNDA.n4956 GNDA.n4955 185
R22057 GNDA.n4958 GNDA.n4949 185
R22058 GNDA.n4960 GNDA.n4959 185
R22059 GNDA.n4961 GNDA.n4948 185
R22060 GNDA.n4963 GNDA.n4962 185
R22061 GNDA.n4965 GNDA.n4947 185
R22062 GNDA.n4968 GNDA.n4967 185
R22063 GNDA.n5179 GNDA.n5178 185
R22064 GNDA.n5176 GNDA.n887 185
R22065 GNDA.n5175 GNDA.n892 185
R22066 GNDA.n5173 GNDA.n5172 185
R22067 GNDA.n4933 GNDA.n893 185
R22068 GNDA.n4937 GNDA.n4936 185
R22069 GNDA.n5012 GNDA.n5011 185
R22070 GNDA.n5009 GNDA.n4929 185
R22071 GNDA.n5008 GNDA.n5007 185
R22072 GNDA.n4419 GNDA.n4418 185
R22073 GNDA.n4421 GNDA.n4420 185
R22074 GNDA.n4423 GNDA.n4422 185
R22075 GNDA.n4425 GNDA.n4424 185
R22076 GNDA.n4427 GNDA.n4426 185
R22077 GNDA.n4429 GNDA.n4428 185
R22078 GNDA.n4431 GNDA.n4430 185
R22079 GNDA.n4433 GNDA.n4432 185
R22080 GNDA.n4434 GNDA.n1936 185
R22081 GNDA.n4401 GNDA.n4400 185
R22082 GNDA.n4403 GNDA.n4402 185
R22083 GNDA.n4405 GNDA.n4404 185
R22084 GNDA.n4407 GNDA.n4406 185
R22085 GNDA.n4409 GNDA.n4408 185
R22086 GNDA.n4411 GNDA.n4410 185
R22087 GNDA.n4413 GNDA.n4412 185
R22088 GNDA.n4415 GNDA.n4414 185
R22089 GNDA.n4417 GNDA.n4416 185
R22090 GNDA.n4383 GNDA.n4382 185
R22091 GNDA.n4385 GNDA.n4384 185
R22092 GNDA.n4387 GNDA.n4386 185
R22093 GNDA.n4389 GNDA.n4388 185
R22094 GNDA.n4391 GNDA.n4390 185
R22095 GNDA.n4393 GNDA.n4392 185
R22096 GNDA.n4395 GNDA.n4394 185
R22097 GNDA.n4397 GNDA.n4396 185
R22098 GNDA.n4399 GNDA.n4398 185
R22099 GNDA.n4381 GNDA.n4380 185
R22100 GNDA.n4375 GNDA.n4374 185
R22101 GNDA.n4373 GNDA.n4372 185
R22102 GNDA.n4368 GNDA.n4367 185
R22103 GNDA.n4366 GNDA.n4365 185
R22104 GNDA.n4360 GNDA.n4359 185
R22105 GNDA.n4355 GNDA.n1940 185
R22106 GNDA.n4439 GNDA.n4438 185
R22107 GNDA.n1939 GNDA.n1937 185
R22108 GNDA.n1285 GNDA.n1262 175.546
R22109 GNDA.n1281 GNDA.n1262 175.546
R22110 GNDA.n1281 GNDA.n1264 175.546
R22111 GNDA.n1277 GNDA.n1264 175.546
R22112 GNDA.n1277 GNDA.n1275 175.546
R22113 GNDA.n1275 GNDA.n1274 175.546
R22114 GNDA.n1274 GNDA.n1267 175.546
R22115 GNDA.n1270 GNDA.n1267 175.546
R22116 GNDA.n1270 GNDA.n760 175.546
R22117 GNDA.n5330 GNDA.n760 175.546
R22118 GNDA.n5330 GNDA.n761 175.546
R22119 GNDA.n5277 GNDA.n811 175.546
R22120 GNDA.n5292 GNDA.n811 175.546
R22121 GNDA.n5292 GNDA.n812 175.546
R22122 GNDA.n5288 GNDA.n812 175.546
R22123 GNDA.n5288 GNDA.n777 175.546
R22124 GNDA.n5302 GNDA.n777 175.546
R22125 GNDA.n5302 GNDA.n778 175.546
R22126 GNDA.n788 GNDA.n778 175.546
R22127 GNDA.n788 GNDA.n754 175.546
R22128 GNDA.n5336 GNDA.n754 175.546
R22129 GNDA.n5336 GNDA.n755 175.546
R22130 GNDA.n1373 GNDA.n1372 175.546
R22131 GNDA.n1372 GNDA.n1334 175.546
R22132 GNDA.n1368 GNDA.n1366 175.546
R22133 GNDA.n1364 GNDA.n1342 175.546
R22134 GNDA.n1360 GNDA.n1358 175.546
R22135 GNDA.n1356 GNDA.n1350 175.546
R22136 GNDA.n1306 GNDA.n1305 175.546
R22137 GNDA.n1302 GNDA.n1301 175.546
R22138 GNDA.n1298 GNDA.n1297 175.546
R22139 GNDA.n1294 GNDA.n1293 175.546
R22140 GNDA.n1290 GNDA.n1289 175.546
R22141 GNDA.n1337 GNDA.n1336 175.546
R22142 GNDA.n1340 GNDA.n1339 175.546
R22143 GNDA.n1345 GNDA.n1344 175.546
R22144 GNDA.n1348 GNDA.n1347 175.546
R22145 GNDA.n1354 GNDA.n1352 175.546
R22146 GNDA.n1311 GNDA.n1310 175.546
R22147 GNDA.n1315 GNDA.n1314 175.546
R22148 GNDA.n1319 GNDA.n1318 175.546
R22149 GNDA.n1323 GNDA.n1322 175.546
R22150 GNDA.n1327 GNDA.n1326 175.546
R22151 GNDA.n879 GNDA.n741 175.546
R22152 GNDA.n5363 GNDA.n741 175.546
R22153 GNDA.n5363 GNDA.n742 175.546
R22154 GNDA.n5359 GNDA.n742 175.546
R22155 GNDA.n5359 GNDA.n716 175.546
R22156 GNDA.n5373 GNDA.n716 175.546
R22157 GNDA.n5373 GNDA.n717 175.546
R22158 GNDA.n5075 GNDA.n717 175.546
R22159 GNDA.n5075 GNDA.n5072 175.546
R22160 GNDA.n5138 GNDA.n5072 175.546
R22161 GNDA.n5138 GNDA.n818 175.546
R22162 GNDA.n5207 GNDA.n5206 175.546
R22163 GNDA.n5206 GNDA.n850 175.546
R22164 GNDA.n5202 GNDA.n5200 175.546
R22165 GNDA.n5198 GNDA.n858 175.546
R22166 GNDA.n5194 GNDA.n5192 175.546
R22167 GNDA.n5190 GNDA.n866 175.546
R22168 GNDA.n925 GNDA.n903 175.546
R22169 GNDA.n929 GNDA.n903 175.546
R22170 GNDA.n929 GNDA.n901 175.546
R22171 GNDA.n933 GNDA.n901 175.546
R22172 GNDA.n933 GNDA.n898 175.546
R22173 GNDA.n5040 GNDA.n898 175.546
R22174 GNDA.n5040 GNDA.n899 175.546
R22175 GNDA.n5036 GNDA.n899 175.546
R22176 GNDA.n5036 GNDA.n937 175.546
R22177 GNDA.n5032 GNDA.n937 175.546
R22178 GNDA.n5032 GNDA.n939 175.546
R22179 GNDA.n920 GNDA.n919 175.546
R22180 GNDA.n916 GNDA.n915 175.546
R22181 GNDA.n912 GNDA.n911 175.546
R22182 GNDA.n908 GNDA.n907 175.546
R22183 GNDA.n904 GNDA.n843 175.546
R22184 GNDA.n5028 GNDA.n943 175.546
R22185 GNDA.n4927 GNDA.n943 175.546
R22186 GNDA.n5014 GNDA.n4927 175.546
R22187 GNDA.n5014 GNDA.n4928 175.546
R22188 GNDA.n4934 GNDA.n4928 175.546
R22189 GNDA.n4934 GNDA.n894 175.546
R22190 GNDA.n5170 GNDA.n894 175.546
R22191 GNDA.n5170 GNDA.n886 175.546
R22192 GNDA.n5181 GNDA.n886 175.546
R22193 GNDA.n5181 GNDA.n883 175.546
R22194 GNDA.n5185 GNDA.n883 175.546
R22195 GNDA.n853 GNDA.n852 175.546
R22196 GNDA.n856 GNDA.n855 175.546
R22197 GNDA.n861 GNDA.n860 175.546
R22198 GNDA.n864 GNDA.n863 175.546
R22199 GNDA.n869 GNDA.n868 175.546
R22200 GNDA.n1907 GNDA.n1905 175.546
R22201 GNDA.n1914 GNDA.n1903 175.546
R22202 GNDA.n1918 GNDA.n1916 175.546
R22203 GNDA.n1926 GNDA.n1901 175.546
R22204 GNDA.n1930 GNDA.n1928 175.546
R22205 GNDA.n1594 GNDA.n1526 175.546
R22206 GNDA.n1590 GNDA.n1526 175.546
R22207 GNDA.n1590 GNDA.n1582 175.546
R22208 GNDA.n1586 GNDA.n1582 175.546
R22209 GNDA.n1586 GNDA.n1118 175.546
R22210 GNDA.n4879 GNDA.n1118 175.546
R22211 GNDA.n4879 GNDA.n1119 175.546
R22212 GNDA.n4875 GNDA.n1119 175.546
R22213 GNDA.n4875 GNDA.n1121 175.546
R22214 GNDA.n4871 GNDA.n1121 175.546
R22215 GNDA.n4871 GNDA.n1123 175.546
R22216 GNDA.n1604 GNDA.n1522 175.546
R22217 GNDA.n1608 GNDA.n1606 175.546
R22218 GNDA.n1616 GNDA.n1518 175.546
R22219 GNDA.n1620 GNDA.n1618 175.546
R22220 GNDA.n1629 GNDA.n1514 175.546
R22221 GNDA.n1602 GNDA.n1600 175.546
R22222 GNDA.n1610 GNDA.n1520 175.546
R22223 GNDA.n1614 GNDA.n1612 175.546
R22224 GNDA.n1622 GNDA.n1516 175.546
R22225 GNDA.n1627 GNDA.n1624 175.546
R22226 GNDA.n1496 GNDA.n1153 175.546
R22227 GNDA.n1493 GNDA.n1492 175.546
R22228 GNDA.n1486 GNDA.n1485 175.546
R22229 GNDA.n1479 GNDA.n1478 175.546
R22230 GNDA.n1507 GNDA.n1506 175.546
R22231 GNDA.n1551 GNDA.n1539 175.546
R22232 GNDA.n1551 GNDA.n1541 175.546
R22233 GNDA.n1547 GNDA.n1541 175.546
R22234 GNDA.n1547 GNDA.n1543 175.546
R22235 GNDA.n1543 GNDA.n1143 175.546
R22236 GNDA.n4861 GNDA.n1143 175.546
R22237 GNDA.n4861 GNDA.n1144 175.546
R22238 GNDA.n4857 GNDA.n1144 175.546
R22239 GNDA.n4857 GNDA.n1147 175.546
R22240 GNDA.n4853 GNDA.n1147 175.546
R22241 GNDA.n4853 GNDA.n1149 175.546
R22242 GNDA.n1555 GNDA.n1537 175.546
R22243 GNDA.n1559 GNDA.n1537 175.546
R22244 GNDA.n1559 GNDA.n1535 175.546
R22245 GNDA.n1564 GNDA.n1535 175.546
R22246 GNDA.n1564 GNDA.n1533 175.546
R22247 GNDA.n1568 GNDA.n1533 175.546
R22248 GNDA.n1568 GNDA.n1531 175.546
R22249 GNDA.n1572 GNDA.n1531 175.546
R22250 GNDA.n1572 GNDA.n1529 175.546
R22251 GNDA.n1577 GNDA.n1529 175.546
R22252 GNDA.n1577 GNDA.n1524 175.546
R22253 GNDA.n1847 GNDA.n1846 175.546
R22254 GNDA.n1846 GNDA.n1695 175.546
R22255 GNDA.n1842 GNDA.n1695 175.546
R22256 GNDA.n1842 GNDA.n1698 175.546
R22257 GNDA.n1838 GNDA.n1698 175.546
R22258 GNDA.n1838 GNDA.n1836 175.546
R22259 GNDA.n1836 GNDA.n1701 175.546
R22260 GNDA.n1832 GNDA.n1701 175.546
R22261 GNDA.n1832 GNDA.n1703 175.546
R22262 GNDA.n1828 GNDA.n1703 175.546
R22263 GNDA.n1828 GNDA.n1706 175.546
R22264 GNDA.n1807 GNDA.n1806 175.546
R22265 GNDA.n1803 GNDA.n1802 175.546
R22266 GNDA.n1796 GNDA.n1795 175.546
R22267 GNDA.n1789 GNDA.n1788 175.546
R22268 GNDA.n1818 GNDA.n1817 175.546
R22269 GNDA.n1895 GNDA.n1894 175.546
R22270 GNDA.n1891 GNDA.n1890 175.546
R22271 GNDA.n1888 GNDA.n1875 175.546
R22272 GNDA.n1884 GNDA.n1882 175.546
R22273 GNDA.n4626 GNDA.n1381 175.546
R22274 GNDA.n1866 GNDA.n1686 175.546
R22275 GNDA.n1862 GNDA.n1861 175.546
R22276 GNDA.n1859 GNDA.n1689 175.546
R22277 GNDA.n1855 GNDA.n1854 175.546
R22278 GNDA.n1852 GNDA.n1692 175.546
R22279 GNDA.n1871 GNDA.n1870 175.546
R22280 GNDA.n1873 GNDA.n1872 175.546
R22281 GNDA.n1877 GNDA.n1876 175.546
R22282 GNDA.n1879 GNDA.n1878 175.546
R22283 GNDA.n4624 GNDA.n1383 175.546
R22284 GNDA.n1235 GNDA.n1230 175.546
R22285 GNDA.n4713 GNDA.n4712 175.546
R22286 GNDA.n4638 GNDA.n4637 175.546
R22287 GNDA.n4643 GNDA.n4642 175.546
R22288 GNDA.n4651 GNDA.n4650 175.546
R22289 GNDA.n4614 GNDA.n1395 175.546
R22290 GNDA.n4612 GNDA.n4611 175.546
R22291 GNDA.n4608 GNDA.n4607 175.546
R22292 GNDA.n4604 GNDA.n4603 175.546
R22293 GNDA.n4600 GNDA.n4599 175.546
R22294 GNDA.n1665 GNDA.n1662 175.546
R22295 GNDA.n1669 GNDA.n1667 175.546
R22296 GNDA.n1673 GNDA.n1659 175.546
R22297 GNDA.n1677 GNDA.n1675 175.546
R22298 GNDA.n1681 GNDA.n1657 175.546
R22299 GNDA.n4580 GNDA.n4579 175.546
R22300 GNDA.n4583 GNDA.n4582 175.546
R22301 GNDA.n4586 GNDA.n4585 175.546
R22302 GNDA.n4589 GNDA.n4588 175.546
R22303 GNDA.n4592 GNDA.n4591 175.546
R22304 GNDA.n4815 GNDA.n4814 175.546
R22305 GNDA.n4747 GNDA.n4727 175.546
R22306 GNDA.n4729 GNDA.n4726 175.546
R22307 GNDA.n4737 GNDA.n4736 175.546
R22308 GNDA.n4751 GNDA.n1216 175.546
R22309 GNDA.n4844 GNDA.n1177 175.546
R22310 GNDA.n4840 GNDA.n1177 175.546
R22311 GNDA.n4840 GNDA.n1180 175.546
R22312 GNDA.n4836 GNDA.n1180 175.546
R22313 GNDA.n4836 GNDA.n1182 175.546
R22314 GNDA.n4832 GNDA.n1182 175.546
R22315 GNDA.n4832 GNDA.n1184 175.546
R22316 GNDA.n4828 GNDA.n1184 175.546
R22317 GNDA.n4828 GNDA.n1187 175.546
R22318 GNDA.n4824 GNDA.n1187 175.546
R22319 GNDA.n4824 GNDA.n1189 175.546
R22320 GNDA.n4558 GNDA.n4556 175.546
R22321 GNDA.n4562 GNDA.n4553 175.546
R22322 GNDA.n4566 GNDA.n4564 175.546
R22323 GNDA.n4570 GNDA.n4551 175.546
R22324 GNDA.n4573 GNDA.n4572 175.546
R22325 GNDA.n4541 GNDA.n4540 175.546
R22326 GNDA.n4456 GNDA.n4455 175.546
R22327 GNDA.n4462 GNDA.n4461 175.546
R22328 GNDA.n4469 GNDA.n4468 175.546
R22329 GNDA.n4477 GNDA.n4476 175.546
R22330 GNDA.n1908 GNDA.n1128 175.546
R22331 GNDA.n1912 GNDA.n1911 175.546
R22332 GNDA.n1920 GNDA.n1919 175.546
R22333 GNDA.n1924 GNDA.n1923 175.546
R22334 GNDA.n1932 GNDA.n1931 175.546
R22335 GNDA.n4301 GNDA.n1127 175.546
R22336 GNDA.n4301 GNDA.n4298 175.546
R22337 GNDA.n4305 GNDA.n4298 175.546
R22338 GNDA.n4305 GNDA.n4296 175.546
R22339 GNDA.n4309 GNDA.n4296 175.546
R22340 GNDA.n4309 GNDA.n4294 175.546
R22341 GNDA.n4314 GNDA.n4294 175.546
R22342 GNDA.n4314 GNDA.n4292 175.546
R22343 GNDA.n4318 GNDA.n4292 175.546
R22344 GNDA.n4318 GNDA.n4290 175.546
R22345 GNDA.n4322 GNDA.n4290 175.546
R22346 GNDA.n4442 GNDA.n4441 175.546
R22347 GNDA.n4357 GNDA.n4356 175.546
R22348 GNDA.n4363 GNDA.n4362 175.546
R22349 GNDA.n4370 GNDA.n4369 175.546
R22350 GNDA.n4378 GNDA.n4377 175.546
R22351 GNDA.n4326 GNDA.n4288 175.546
R22352 GNDA.n4326 GNDA.n1964 175.546
R22353 GNDA.n4332 GNDA.n1964 175.546
R22354 GNDA.n4332 GNDA.n1962 175.546
R22355 GNDA.n4336 GNDA.n1962 175.546
R22356 GNDA.n4337 GNDA.n4336 175.546
R22357 GNDA.n4339 GNDA.n4337 175.546
R22358 GNDA.n4339 GNDA.n1960 175.546
R22359 GNDA.n4344 GNDA.n1960 175.546
R22360 GNDA.n4344 GNDA.n1958 175.546
R22361 GNDA.n4348 GNDA.n1958 175.546
R22362 GNDA.n5344 GNDA.n746 173.727
R22363 GNDA.n4924 GNDA.n4923 173.727
R22364 GNDA.n5478 GNDA.n5477 166.4
R22365 GNDA.n5472 GNDA.n5471 166.4
R22366 GNDA.n799 GNDA.n798 163.333
R22367 GNDA.n5134 GNDA.n5133 163.333
R22368 GNDA.n4655 GNDA.n4654 163.333
R22369 GNDA.n1413 GNDA.n1403 163.333
R22370 GNDA.n1721 GNDA.n1711 163.333
R22371 GNDA.n4755 GNDA.n4754 163.333
R22372 GNDA.n4481 GNDA.n4480 163.333
R22373 GNDA.n5178 GNDA.n889 163.333
R22374 GNDA.n4382 GNDA.n4381 163.333
R22375 GNDA.n4882 GNDA.n1113 157.601
R22376 GNDA.n5254 GNDA.n5253 150
R22377 GNDA.n5250 GNDA.n5249 150
R22378 GNDA.n5246 GNDA.n5245 150
R22379 GNDA.n5242 GNDA.n5241 150
R22380 GNDA.n5238 GNDA.n5237 150
R22381 GNDA.n5234 GNDA.n5233 150
R22382 GNDA.n5230 GNDA.n5229 150
R22383 GNDA.n5226 GNDA.n5225 150
R22384 GNDA.n5295 GNDA.n808 150
R22385 GNDA.n5285 GNDA.n5284 150
R22386 GNDA.n5299 GNDA.n780 150
R22387 GNDA.n792 GNDA.n781 150
R22388 GNDA.n5262 GNDA.n5261 150
R22389 GNDA.n5266 GNDA.n5265 150
R22390 GNDA.n5270 GNDA.n5269 150
R22391 GNDA.n5272 GNDA.n807 150
R22392 GNDA.n5103 GNDA.n5102 150
R22393 GNDA.n5107 GNDA.n5106 150
R22394 GNDA.n5111 GNDA.n5110 150
R22395 GNDA.n5115 GNDA.n5114 150
R22396 GNDA.n5119 GNDA.n5118 150
R22397 GNDA.n5123 GNDA.n5122 150
R22398 GNDA.n5127 GNDA.n5126 150
R22399 GNDA.n5131 GNDA.n5130 150
R22400 GNDA.n5366 GNDA.n738 150
R22401 GNDA.n5356 GNDA.n5355 150
R22402 GNDA.n5370 GNDA.n719 150
R22403 GNDA.n5077 GNDA.n720 150
R22404 GNDA.n5095 GNDA.n5094 150
R22405 GNDA.n5091 GNDA.n5090 150
R22406 GNDA.n5087 GNDA.n5086 150
R22407 GNDA.n5083 GNDA.n737 150
R22408 GNDA.n4687 GNDA.n4686 150
R22409 GNDA.n4683 GNDA.n4682 150
R22410 GNDA.n4679 GNDA.n4678 150
R22411 GNDA.n4675 GNDA.n4674 150
R22412 GNDA.n4671 GNDA.n4670 150
R22413 GNDA.n4667 GNDA.n4666 150
R22414 GNDA.n4663 GNDA.n4662 150
R22415 GNDA.n4659 GNDA.n4658 150
R22416 GNDA.n4717 GNDA.n4716 150
R22417 GNDA.n4709 GNDA.n1241 150
R22418 GNDA.n4640 GNDA.n1242 150
R22419 GNDA.n4647 GNDA.n4646 150
R22420 GNDA.n4705 GNDA.n1258 150
R22421 GNDA.n4701 GNDA.n4700 150
R22422 GNDA.n4697 GNDA.n4696 150
R22423 GNDA.n4693 GNDA.n4692 150
R22424 GNDA.n5307 GNDA.n768 150
R22425 GNDA.n5309 GNDA.n5307 150
R22426 GNDA.n5157 GNDA.n5154 150
R22427 GNDA.n5158 GNDA.n5157 150
R22428 GNDA.n5163 GNDA.n5162 150
R22429 GNDA.n1452 GNDA.n1451 150
R22430 GNDA.n1448 GNDA.n1447 150
R22431 GNDA.n1444 GNDA.n1443 150
R22432 GNDA.n1440 GNDA.n1439 150
R22433 GNDA.n1436 GNDA.n1435 150
R22434 GNDA.n1432 GNDA.n1431 150
R22435 GNDA.n1428 GNDA.n1427 150
R22436 GNDA.n1424 GNDA.n1423 150
R22437 GNDA.n1499 GNDA.n1473 150
R22438 GNDA.n1489 GNDA.n1488 150
R22439 GNDA.n1482 GNDA.n1481 150
R22440 GNDA.n1503 GNDA.n1402 150
R22441 GNDA.n1460 GNDA.n1459 150
R22442 GNDA.n1464 GNDA.n1463 150
R22443 GNDA.n1468 GNDA.n1467 150
R22444 GNDA.n1472 GNDA.n1421 150
R22445 GNDA.n1761 GNDA.n1760 150
R22446 GNDA.n1757 GNDA.n1756 150
R22447 GNDA.n1753 GNDA.n1752 150
R22448 GNDA.n1749 GNDA.n1748 150
R22449 GNDA.n1745 GNDA.n1744 150
R22450 GNDA.n1741 GNDA.n1740 150
R22451 GNDA.n1737 GNDA.n1736 150
R22452 GNDA.n1733 GNDA.n1732 150
R22453 GNDA.n1810 GNDA.n1730 150
R22454 GNDA.n1799 GNDA.n1798 150
R22455 GNDA.n1792 GNDA.n1791 150
R22456 GNDA.n1814 GNDA.n1710 150
R22457 GNDA.n1769 GNDA.n1768 150
R22458 GNDA.n1773 GNDA.n1772 150
R22459 GNDA.n1777 GNDA.n1776 150
R22460 GNDA.n1779 GNDA.n1729 150
R22461 GNDA.n4787 GNDA.n4786 150
R22462 GNDA.n4783 GNDA.n4782 150
R22463 GNDA.n4779 GNDA.n4778 150
R22464 GNDA.n4775 GNDA.n4774 150
R22465 GNDA.n4771 GNDA.n4770 150
R22466 GNDA.n4767 GNDA.n4766 150
R22467 GNDA.n4763 GNDA.n4762 150
R22468 GNDA.n4759 GNDA.n4758 150
R22469 GNDA.n4811 GNDA.n1196 150
R22470 GNDA.n4744 GNDA.n1197 150
R22471 GNDA.n4741 GNDA.n4740 150
R22472 GNDA.n4733 GNDA.n4732 150
R22473 GNDA.n4795 GNDA.n4794 150
R22474 GNDA.n4799 GNDA.n4798 150
R22475 GNDA.n4803 GNDA.n4802 150
R22476 GNDA.n4807 GNDA.n4806 150
R22477 GNDA.n4513 GNDA.n4512 150
R22478 GNDA.n4509 GNDA.n4508 150
R22479 GNDA.n4505 GNDA.n4504 150
R22480 GNDA.n4501 GNDA.n4500 150
R22481 GNDA.n4497 GNDA.n4496 150
R22482 GNDA.n4493 GNDA.n4492 150
R22483 GNDA.n4489 GNDA.n4488 150
R22484 GNDA.n4485 GNDA.n4484 150
R22485 GNDA.n4537 GNDA.n1635 150
R22486 GNDA.n4458 GNDA.n1636 150
R22487 GNDA.n4466 GNDA.n4465 150
R22488 GNDA.n4473 GNDA.n4472 150
R22489 GNDA.n4521 GNDA.n4520 150
R22490 GNDA.n4525 GNDA.n4524 150
R22491 GNDA.n4529 GNDA.n4528 150
R22492 GNDA.n4533 GNDA.n4532 150
R22493 GNDA.n4983 GNDA.n4981 150
R22494 GNDA.n4979 GNDA.n4944 150
R22495 GNDA.n4975 GNDA.n4973 150
R22496 GNDA.n4971 GNDA.n4946 150
R22497 GNDA.n4967 GNDA.n4965 150
R22498 GNDA.n4963 GNDA.n4948 150
R22499 GNDA.n4959 GNDA.n4958 150
R22500 GNDA.n4956 GNDA.n4952 150
R22501 GNDA.n5009 GNDA.n5008 150
R22502 GNDA.n5011 GNDA.n4937 150
R22503 GNDA.n5173 GNDA.n893 150
R22504 GNDA.n5176 GNDA.n5175 150
R22505 GNDA.n4991 GNDA.n4989 150
R22506 GNDA.n4995 GNDA.n4940 150
R22507 GNDA.n4999 GNDA.n4997 150
R22508 GNDA.n5003 GNDA.n4938 150
R22509 GNDA.n4414 GNDA.n4413 150
R22510 GNDA.n4410 GNDA.n4409 150
R22511 GNDA.n4406 GNDA.n4405 150
R22512 GNDA.n4402 GNDA.n4401 150
R22513 GNDA.n4398 GNDA.n4397 150
R22514 GNDA.n4394 GNDA.n4393 150
R22515 GNDA.n4390 GNDA.n4389 150
R22516 GNDA.n4386 GNDA.n4385 150
R22517 GNDA.n4438 GNDA.n1939 150
R22518 GNDA.n4359 GNDA.n1940 150
R22519 GNDA.n4367 GNDA.n4366 150
R22520 GNDA.n4374 GNDA.n4373 150
R22521 GNDA.n4422 GNDA.n4421 150
R22522 GNDA.n4426 GNDA.n4425 150
R22523 GNDA.n4430 GNDA.n4429 150
R22524 GNDA.n4434 GNDA.n4433 150
R22525 GNDA.n2200 GNDA.n2115 148.017
R22526 GNDA.n3622 GNDA.n1968 148.017
R22527 GNDA.n3617 GNDA.n1968 148.017
R22528 GNDA.n2205 GNDA.n2115 148.017
R22529 GNDA.n5339 GNDA.n751 130.001
R22530 GNDA.n5218 GNDA.n5217 130.001
R22531 GNDA.n820 GNDA.n819 130.001
R22532 GNDA.n5348 GNDA.n744 130.001
R22533 GNDA.n876 GNDA.n873 130.001
R22534 GNDA.n5017 GNDA.n4925 130.001
R22535 GNDA.n5024 GNDA.n946 130.001
R22536 GNDA.n4918 GNDA.n4917 127.754
R22537 GNDA.n4863 GNDA.n1140 127.219
R22538 GNDA.n1835 GNDA.n1185 127.219
R22539 GNDA.n5304 GNDA.n774 127.219
R22540 GNDA.n4863 GNDA.n4862 127.219
R22541 GNDA.n4831 GNDA.n1185 127.219
R22542 GNDA.n5042 GNDA.n5041 127.219
R22543 GNDA.n1350 GNDA.n814 124.832
R22544 GNDA.n5221 GNDA.n817 124.832
R22545 GNDA.n880 GNDA.n866 124.832
R22546 GNDA.n884 GNDA.n871 124.832
R22547 GNDA.n4449 GNDA.n1654 124.832
R22548 GNDA.n4546 GNDA.n1631 124.832
R22549 GNDA.n1625 GNDA.n1512 124.832
R22550 GNDA.n4629 GNDA.n4628 124.832
R22551 GNDA.n4631 GNDA.n1260 124.832
R22552 GNDA.n4596 GNDA.n1231 124.832
R22553 GNDA.n4595 GNDA.n4594 124.832
R22554 GNDA.n4447 GNDA.n1935 124.832
R22555 GNDA.n1580 GNDA.n1579 105.719
R22556 GNDA.n1129 GNDA.n1122 105.719
R22557 GNDA.n1593 GNDA.n1580 103.457
R22558 GNDA.n4299 GNDA.n1129 103.457
R22559 GNDA.n4847 GNDA.n4846 103.144
R22560 GNDA.n4749 GNDA.n825 103.144
R22561 GNDA.n5305 GNDA.n772 101.718
R22562 GNDA.n5159 GNDA.n5043 101.718
R22563 GNDA.n5166 GNDA.n5045 101.718
R22564 GNDA.n5316 GNDA.n770 101.718
R22565 GNDA.n5184 GNDA.n824 101.162
R22566 GNDA.n4846 GNDA.n1173 99.6276
R22567 GNDA.n5215 GNDA.n825 99.6276
R22568 GNDA.n5278 GNDA.n813 96.1535
R22569 GNDA.n595 GNDA.n594 92.8005
R22570 GNDA.n591 GNDA.n590 92.8005
R22571 GNDA.n4621 GNDA.n1173 91.423
R22572 GNDA.n5216 GNDA.n5215 91.423
R22573 GNDA.n5027 GNDA.n5026 90.1439
R22574 GNDA.n5015 GNDA.n4926 90.1439
R22575 GNDA.n4926 GNDA.n895 90.1439
R22576 GNDA.n5169 GNDA.n5168 90.1439
R22577 GNDA.n5169 GNDA.n885 90.1439
R22578 GNDA.n5182 GNDA.n885 90.1439
R22579 GNDA.n5183 GNDA.n5182 90.1439
R22580 GNDA.n5184 GNDA.n5183 90.1439
R22581 GNDA.n5362 GNDA.n5350 90.1439
R22582 GNDA.n5362 GNDA.n5361 90.1439
R22583 GNDA.n5361 GNDA.n5360 90.1439
R22584 GNDA.n5360 GNDA.n714 90.1439
R22585 GNDA.n5374 GNDA.n715 90.1439
R22586 GNDA.n5074 GNDA.n715 90.1439
R22587 GNDA.n5074 GNDA.n5071 90.1439
R22588 GNDA.n5139 GNDA.n5071 90.1439
R22589 GNDA.n5279 GNDA.n5278 90.1439
R22590 GNDA.n5291 GNDA.n5279 90.1439
R22591 GNDA.n5291 GNDA.n5290 90.1439
R22592 GNDA.n5290 GNDA.n5289 90.1439
R22593 GNDA.n5289 GNDA.n771 90.1439
R22594 GNDA.n5303 GNDA.n776 90.1439
R22595 GNDA.n787 GNDA.n776 90.1439
R22596 GNDA.n787 GNDA.n752 90.1439
R22597 GNDA.n5337 GNDA.n753 90.1439
R22598 GNDA.n5397 GNDA.n641 89.6005
R22599 GNDA.n5407 GNDA.n5397 89.6005
R22600 GNDA.n5016 GNDA.n945 87.1391
R22601 GNDA.n5216 GNDA.n823 87.1391
R22602 GNDA.n5216 GNDA.n813 87.1391
R22603 GNDA.n5216 GNDA.n824 86.1375
R22604 GNDA.n5059 GNDA.n5058 84.306
R22605 GNDA.n5142 GNDA.n5070 84.306
R22606 GNDA.n1375 GNDA.n1374 76.3222
R22607 GNDA.n1367 GNDA.n1334 76.3222
R22608 GNDA.n1366 GNDA.n1365 76.3222
R22609 GNDA.n1359 GNDA.n1342 76.3222
R22610 GNDA.n1358 GNDA.n1357 76.3222
R22611 GNDA.n1306 GNDA.n826 76.3222
R22612 GNDA.n1302 GNDA.n827 76.3222
R22613 GNDA.n1298 GNDA.n828 76.3222
R22614 GNDA.n1294 GNDA.n829 76.3222
R22615 GNDA.n1290 GNDA.n830 76.3222
R22616 GNDA.n1286 GNDA.n831 76.3222
R22617 GNDA.n1336 GNDA.n1335 76.3222
R22618 GNDA.n1339 GNDA.n1338 76.3222
R22619 GNDA.n1344 GNDA.n1343 76.3222
R22620 GNDA.n1347 GNDA.n1346 76.3222
R22621 GNDA.n1352 GNDA.n1351 76.3222
R22622 GNDA.n1353 GNDA.n817 76.3222
R22623 GNDA.n1310 GNDA.n832 76.3222
R22624 GNDA.n1314 GNDA.n833 76.3222
R22625 GNDA.n1318 GNDA.n834 76.3222
R22626 GNDA.n1322 GNDA.n835 76.3222
R22627 GNDA.n1326 GNDA.n836 76.3222
R22628 GNDA.n1330 GNDA.n837 76.3222
R22629 GNDA.n5209 GNDA.n5208 76.3222
R22630 GNDA.n5201 GNDA.n850 76.3222
R22631 GNDA.n5200 GNDA.n5199 76.3222
R22632 GNDA.n5193 GNDA.n858 76.3222
R22633 GNDA.n5192 GNDA.n5191 76.3222
R22634 GNDA.n920 GNDA.n838 76.3222
R22635 GNDA.n916 GNDA.n839 76.3222
R22636 GNDA.n912 GNDA.n840 76.3222
R22637 GNDA.n908 GNDA.n841 76.3222
R22638 GNDA.n904 GNDA.n842 76.3222
R22639 GNDA.n5214 GNDA.n5213 76.3222
R22640 GNDA.n851 GNDA.n844 76.3222
R22641 GNDA.n854 GNDA.n853 76.3222
R22642 GNDA.n859 GNDA.n856 76.3222
R22643 GNDA.n862 GNDA.n861 76.3222
R22644 GNDA.n867 GNDA.n864 76.3222
R22645 GNDA.n870 GNDA.n869 76.3222
R22646 GNDA.n1905 GNDA.n1904 76.3222
R22647 GNDA.n1906 GNDA.n1903 76.3222
R22648 GNDA.n1916 GNDA.n1915 76.3222
R22649 GNDA.n1917 GNDA.n1901 76.3222
R22650 GNDA.n1928 GNDA.n1927 76.3222
R22651 GNDA.n1929 GNDA.n1654 76.3222
R22652 GNDA.n1596 GNDA.n1595 76.3222
R22653 GNDA.n1605 GNDA.n1604 76.3222
R22654 GNDA.n1608 GNDA.n1607 76.3222
R22655 GNDA.n1617 GNDA.n1616 76.3222
R22656 GNDA.n1620 GNDA.n1619 76.3222
R22657 GNDA.n1630 GNDA.n1629 76.3222
R22658 GNDA.n1600 GNDA.n1599 76.3222
R22659 GNDA.n1601 GNDA.n1520 76.3222
R22660 GNDA.n1612 GNDA.n1611 76.3222
R22661 GNDA.n1613 GNDA.n1516 76.3222
R22662 GNDA.n1624 GNDA.n1623 76.3222
R22663 GNDA.n1626 GNDA.n1625 76.3222
R22664 GNDA.n4849 GNDA.n4848 76.3222
R22665 GNDA.n1493 GNDA.n1164 76.3222
R22666 GNDA.n1486 GNDA.n1163 76.3222
R22667 GNDA.n1479 GNDA.n1162 76.3222
R22668 GNDA.n1506 GNDA.n1161 76.3222
R22669 GNDA.n1511 GNDA.n1160 76.3222
R22670 GNDA.n1378 GNDA.n1224 76.3222
R22671 GNDA.n1807 GNDA.n1223 76.3222
R22672 GNDA.n1802 GNDA.n1222 76.3222
R22673 GNDA.n1795 GNDA.n1221 76.3222
R22674 GNDA.n1788 GNDA.n1220 76.3222
R22675 GNDA.n1818 GNDA.n1219 76.3222
R22676 GNDA.n1897 GNDA.n1896 76.3222
R22677 GNDA.n1894 GNDA.n1869 76.3222
R22678 GNDA.n1890 GNDA.n1889 76.3222
R22679 GNDA.n1883 GNDA.n1875 76.3222
R22680 GNDA.n1882 GNDA.n1881 76.3222
R22681 GNDA.n4627 GNDA.n4626 76.3222
R22682 GNDA.n1867 GNDA.n1866 76.3222
R22683 GNDA.n1862 GNDA.n1688 76.3222
R22684 GNDA.n1860 GNDA.n1859 76.3222
R22685 GNDA.n1855 GNDA.n1691 76.3222
R22686 GNDA.n1853 GNDA.n1852 76.3222
R22687 GNDA.n1848 GNDA.n1694 76.3222
R22688 GNDA.n1870 GNDA.n1384 76.3222
R22689 GNDA.n1872 GNDA.n1385 76.3222
R22690 GNDA.n1876 GNDA.n1386 76.3222
R22691 GNDA.n1878 GNDA.n1387 76.3222
R22692 GNDA.n1388 GNDA.n1383 76.3222
R22693 GNDA.n4623 GNDA.n1260 76.3222
R22694 GNDA.n4723 GNDA.n4722 76.3222
R22695 GNDA.n1235 GNDA.n1229 76.3222
R22696 GNDA.n4712 GNDA.n1228 76.3222
R22697 GNDA.n4638 GNDA.n1227 76.3222
R22698 GNDA.n4642 GNDA.n1226 76.3222
R22699 GNDA.n4651 GNDA.n1225 76.3222
R22700 GNDA.n4619 GNDA.n4618 76.3222
R22701 GNDA.n4614 GNDA.n1394 76.3222
R22702 GNDA.n4611 GNDA.n1393 76.3222
R22703 GNDA.n4607 GNDA.n1392 76.3222
R22704 GNDA.n4603 GNDA.n1391 76.3222
R22705 GNDA.n4599 GNDA.n1390 76.3222
R22706 GNDA.n1662 GNDA.n1661 76.3222
R22707 GNDA.n1667 GNDA.n1666 76.3222
R22708 GNDA.n1668 GNDA.n1659 76.3222
R22709 GNDA.n1675 GNDA.n1674 76.3222
R22710 GNDA.n1676 GNDA.n1657 76.3222
R22711 GNDA.n1683 GNDA.n1682 76.3222
R22712 GNDA.n4579 GNDA.n4578 76.3222
R22713 GNDA.n4582 GNDA.n4581 76.3222
R22714 GNDA.n4585 GNDA.n4584 76.3222
R22715 GNDA.n4588 GNDA.n4587 76.3222
R22716 GNDA.n4591 GNDA.n4590 76.3222
R22717 GNDA.n4595 GNDA.n4593 76.3222
R22718 GNDA.n4819 GNDA.n1191 76.3222
R22719 GNDA.n4814 GNDA.n1194 76.3222
R22720 GNDA.n4748 GNDA.n4747 76.3222
R22721 GNDA.n4729 GNDA.n4725 76.3222
R22722 GNDA.n4736 GNDA.n4724 76.3222
R22723 GNDA.n4751 GNDA.n4750 76.3222
R22724 GNDA.n4556 GNDA.n4555 76.3222
R22725 GNDA.n4557 GNDA.n4553 76.3222
R22726 GNDA.n4564 GNDA.n4563 76.3222
R22727 GNDA.n4565 GNDA.n4551 76.3222
R22728 GNDA.n4572 GNDA.n4571 76.3222
R22729 GNDA.n4576 GNDA.n4549 76.3222
R22730 GNDA.n4573 GNDA.n4549 76.3222
R22731 GNDA.n4571 GNDA.n4570 76.3222
R22732 GNDA.n4566 GNDA.n4565 76.3222
R22733 GNDA.n4563 GNDA.n4562 76.3222
R22734 GNDA.n4558 GNDA.n4557 76.3222
R22735 GNDA.n4555 GNDA.n1176 76.3222
R22736 GNDA.n1682 GNDA.n1681 76.3222
R22737 GNDA.n1677 GNDA.n1676 76.3222
R22738 GNDA.n1674 GNDA.n1673 76.3222
R22739 GNDA.n1669 GNDA.n1668 76.3222
R22740 GNDA.n1666 GNDA.n1665 76.3222
R22741 GNDA.n1661 GNDA.n1396 76.3222
R22742 GNDA.n1694 GNDA.n1692 76.3222
R22743 GNDA.n1854 GNDA.n1853 76.3222
R22744 GNDA.n1691 GNDA.n1689 76.3222
R22745 GNDA.n1861 GNDA.n1860 76.3222
R22746 GNDA.n1688 GNDA.n1686 76.3222
R22747 GNDA.n1868 GNDA.n1867 76.3222
R22748 GNDA.n4541 GNDA.n1170 76.3222
R22749 GNDA.n4455 GNDA.n1169 76.3222
R22750 GNDA.n4461 GNDA.n1168 76.3222
R22751 GNDA.n4469 GNDA.n1167 76.3222
R22752 GNDA.n4476 GNDA.n1166 76.3222
R22753 GNDA.n4450 GNDA.n1165 76.3222
R22754 GNDA.n4545 GNDA.n1170 76.3222
R22755 GNDA.n4540 GNDA.n1169 76.3222
R22756 GNDA.n4456 GNDA.n1168 76.3222
R22757 GNDA.n4462 GNDA.n1167 76.3222
R22758 GNDA.n4468 GNDA.n1166 76.3222
R22759 GNDA.n4477 GNDA.n1165 76.3222
R22760 GNDA.n4848 GNDA.n1153 76.3222
R22761 GNDA.n1496 GNDA.n1164 76.3222
R22762 GNDA.n1492 GNDA.n1163 76.3222
R22763 GNDA.n1485 GNDA.n1162 76.3222
R22764 GNDA.n1478 GNDA.n1161 76.3222
R22765 GNDA.n1507 GNDA.n1160 76.3222
R22766 GNDA.n1627 GNDA.n1626 76.3222
R22767 GNDA.n1623 GNDA.n1622 76.3222
R22768 GNDA.n1614 GNDA.n1613 76.3222
R22769 GNDA.n1611 GNDA.n1610 76.3222
R22770 GNDA.n1602 GNDA.n1601 76.3222
R22771 GNDA.n1599 GNDA.n1598 76.3222
R22772 GNDA.n1595 GNDA.n1522 76.3222
R22773 GNDA.n1606 GNDA.n1605 76.3222
R22774 GNDA.n1607 GNDA.n1518 76.3222
R22775 GNDA.n1618 GNDA.n1617 76.3222
R22776 GNDA.n1619 GNDA.n1514 76.3222
R22777 GNDA.n1631 GNDA.n1630 76.3222
R22778 GNDA.n4593 GNDA.n4592 76.3222
R22779 GNDA.n4590 GNDA.n4589 76.3222
R22780 GNDA.n4587 GNDA.n4586 76.3222
R22781 GNDA.n4584 GNDA.n4583 76.3222
R22782 GNDA.n4581 GNDA.n4580 76.3222
R22783 GNDA.n4578 GNDA.n4577 76.3222
R22784 GNDA.n4619 GNDA.n1395 76.3222
R22785 GNDA.n4612 GNDA.n1394 76.3222
R22786 GNDA.n4608 GNDA.n1393 76.3222
R22787 GNDA.n4604 GNDA.n1392 76.3222
R22788 GNDA.n4600 GNDA.n1391 76.3222
R22789 GNDA.n4596 GNDA.n1390 76.3222
R22790 GNDA.n871 GNDA.n870 76.3222
R22791 GNDA.n868 GNDA.n867 76.3222
R22792 GNDA.n863 GNDA.n862 76.3222
R22793 GNDA.n860 GNDA.n859 76.3222
R22794 GNDA.n855 GNDA.n854 76.3222
R22795 GNDA.n852 GNDA.n851 76.3222
R22796 GNDA.n5208 GNDA.n5207 76.3222
R22797 GNDA.n5202 GNDA.n5201 76.3222
R22798 GNDA.n5199 GNDA.n5198 76.3222
R22799 GNDA.n5194 GNDA.n5193 76.3222
R22800 GNDA.n5191 GNDA.n5190 76.3222
R22801 GNDA.n5214 GNDA.n843 76.3222
R22802 GNDA.n907 GNDA.n842 76.3222
R22803 GNDA.n911 GNDA.n841 76.3222
R22804 GNDA.n915 GNDA.n840 76.3222
R22805 GNDA.n919 GNDA.n839 76.3222
R22806 GNDA.n923 GNDA.n838 76.3222
R22807 GNDA.n1327 GNDA.n837 76.3222
R22808 GNDA.n1323 GNDA.n836 76.3222
R22809 GNDA.n1319 GNDA.n835 76.3222
R22810 GNDA.n1315 GNDA.n834 76.3222
R22811 GNDA.n1311 GNDA.n833 76.3222
R22812 GNDA.n849 GNDA.n832 76.3222
R22813 GNDA.n1289 GNDA.n831 76.3222
R22814 GNDA.n1293 GNDA.n830 76.3222
R22815 GNDA.n1297 GNDA.n829 76.3222
R22816 GNDA.n1301 GNDA.n828 76.3222
R22817 GNDA.n1305 GNDA.n827 76.3222
R22818 GNDA.n1333 GNDA.n826 76.3222
R22819 GNDA.n4815 GNDA.n1191 76.3222
R22820 GNDA.n4727 GNDA.n1194 76.3222
R22821 GNDA.n4748 GNDA.n4726 76.3222
R22822 GNDA.n4737 GNDA.n4725 76.3222
R22823 GNDA.n4724 GNDA.n1216 76.3222
R22824 GNDA.n4750 GNDA.n1217 76.3222
R22825 GNDA.n4723 GNDA.n1230 76.3222
R22826 GNDA.n4713 GNDA.n1229 76.3222
R22827 GNDA.n4637 GNDA.n1228 76.3222
R22828 GNDA.n4643 GNDA.n1227 76.3222
R22829 GNDA.n4650 GNDA.n1226 76.3222
R22830 GNDA.n4632 GNDA.n1225 76.3222
R22831 GNDA.n1806 GNDA.n1224 76.3222
R22832 GNDA.n1803 GNDA.n1223 76.3222
R22833 GNDA.n1796 GNDA.n1222 76.3222
R22834 GNDA.n1789 GNDA.n1221 76.3222
R22835 GNDA.n1817 GNDA.n1220 76.3222
R22836 GNDA.n1822 GNDA.n1219 76.3222
R22837 GNDA.n4866 GNDA.n4865 76.3222
R22838 GNDA.n1908 GNDA.n1134 76.3222
R22839 GNDA.n1912 GNDA.n1133 76.3222
R22840 GNDA.n1920 GNDA.n1132 76.3222
R22841 GNDA.n1924 GNDA.n1131 76.3222
R22842 GNDA.n1932 GNDA.n1130 76.3222
R22843 GNDA.n4442 GNDA.n1159 76.3222
R22844 GNDA.n4356 GNDA.n1158 76.3222
R22845 GNDA.n4362 GNDA.n1157 76.3222
R22846 GNDA.n4370 GNDA.n1156 76.3222
R22847 GNDA.n4377 GNDA.n1155 76.3222
R22848 GNDA.n4351 GNDA.n1154 76.3222
R22849 GNDA.n4446 GNDA.n1159 76.3222
R22850 GNDA.n4441 GNDA.n1158 76.3222
R22851 GNDA.n4357 GNDA.n1157 76.3222
R22852 GNDA.n4363 GNDA.n1156 76.3222
R22853 GNDA.n4369 GNDA.n1155 76.3222
R22854 GNDA.n4378 GNDA.n1154 76.3222
R22855 GNDA.n1930 GNDA.n1929 76.3222
R22856 GNDA.n1927 GNDA.n1926 76.3222
R22857 GNDA.n1918 GNDA.n1917 76.3222
R22858 GNDA.n1915 GNDA.n1914 76.3222
R22859 GNDA.n1907 GNDA.n1906 76.3222
R22860 GNDA.n1904 GNDA.n1125 76.3222
R22861 GNDA.n4865 GNDA.n1128 76.3222
R22862 GNDA.n1911 GNDA.n1134 76.3222
R22863 GNDA.n1919 GNDA.n1133 76.3222
R22864 GNDA.n1923 GNDA.n1132 76.3222
R22865 GNDA.n1931 GNDA.n1131 76.3222
R22866 GNDA.n1935 GNDA.n1130 76.3222
R22867 GNDA.n4624 GNDA.n4623 76.3222
R22868 GNDA.n1879 GNDA.n1388 76.3222
R22869 GNDA.n1877 GNDA.n1387 76.3222
R22870 GNDA.n1873 GNDA.n1386 76.3222
R22871 GNDA.n1871 GNDA.n1385 76.3222
R22872 GNDA.n1684 GNDA.n1384 76.3222
R22873 GNDA.n1896 GNDA.n1895 76.3222
R22874 GNDA.n1891 GNDA.n1869 76.3222
R22875 GNDA.n1889 GNDA.n1888 76.3222
R22876 GNDA.n1884 GNDA.n1883 76.3222
R22877 GNDA.n1881 GNDA.n1381 76.3222
R22878 GNDA.n4628 GNDA.n4627 76.3222
R22879 GNDA.n1354 GNDA.n1353 76.3222
R22880 GNDA.n1351 GNDA.n1348 76.3222
R22881 GNDA.n1346 GNDA.n1345 76.3222
R22882 GNDA.n1343 GNDA.n1340 76.3222
R22883 GNDA.n1338 GNDA.n1337 76.3222
R22884 GNDA.n1335 GNDA.n1331 76.3222
R22885 GNDA.n1374 GNDA.n1373 76.3222
R22886 GNDA.n1368 GNDA.n1367 76.3222
R22887 GNDA.n1365 GNDA.n1364 76.3222
R22888 GNDA.n1360 GNDA.n1359 76.3222
R22889 GNDA.n1357 GNDA.n1356 76.3222
R22890 GNDA.n5475 GNDA.n5474 74.6651
R22891 GNDA.n5241 GNDA.n794 74.5978
R22892 GNDA.n5238 GNDA.n794 74.5978
R22893 GNDA.n5115 GNDA.n726 74.5978
R22894 GNDA.n5118 GNDA.n726 74.5978
R22895 GNDA.n4674 GNDA.n1247 74.5978
R22896 GNDA.n4671 GNDA.n1247 74.5978
R22897 GNDA.n1439 GNDA.n1409 74.5978
R22898 GNDA.n1436 GNDA.n1409 74.5978
R22899 GNDA.n1748 GNDA.n1717 74.5978
R22900 GNDA.n1745 GNDA.n1717 74.5978
R22901 GNDA.n4774 GNDA.n1203 74.5978
R22902 GNDA.n4771 GNDA.n1203 74.5978
R22903 GNDA.n4500 GNDA.n1642 74.5978
R22904 GNDA.n4497 GNDA.n1642 74.5978
R22905 GNDA.n4966 GNDA.n4946 74.5978
R22906 GNDA.n4967 GNDA.n4966 74.5978
R22907 GNDA.n4401 GNDA.n1946 74.5978
R22908 GNDA.n4398 GNDA.n1946 74.5978
R22909 GNDA.n5220 GNDA.n821 74.1184
R22910 GNDA.n1116 GNDA.n1113 69.4466
R22911 GNDA.n5296 GNDA.n5295 69.3109
R22912 GNDA.n5296 GNDA.n807 69.3109
R22913 GNDA.n5367 GNDA.n5366 69.3109
R22914 GNDA.n5367 GNDA.n737 69.3109
R22915 GNDA.n4717 GNDA.n1237 69.3109
R22916 GNDA.n4692 GNDA.n1237 69.3109
R22917 GNDA.n1500 GNDA.n1499 69.3109
R22918 GNDA.n1500 GNDA.n1472 69.3109
R22919 GNDA.n1811 GNDA.n1810 69.3109
R22920 GNDA.n1811 GNDA.n1729 69.3109
R22921 GNDA.n4808 GNDA.n1196 69.3109
R22922 GNDA.n4808 GNDA.n4807 69.3109
R22923 GNDA.n4534 GNDA.n1635 69.3109
R22924 GNDA.n4534 GNDA.n4533 69.3109
R22925 GNDA.n5008 GNDA.n5004 69.3109
R22926 GNDA.n5004 GNDA.n5003 69.3109
R22927 GNDA.n4435 GNDA.n1939 69.3109
R22928 GNDA.n4435 GNDA.n4434 69.3109
R22929 GNDA.n5220 GNDA.n5219 66.1057
R22930 GNDA.n5297 GNDA.n806 65.8183
R22931 GNDA.n5297 GNDA.n805 65.8183
R22932 GNDA.n5297 GNDA.n804 65.8183
R22933 GNDA.n5297 GNDA.n803 65.8183
R22934 GNDA.n5297 GNDA.n785 65.8183
R22935 GNDA.n5297 GNDA.n801 65.8183
R22936 GNDA.n5297 GNDA.n783 65.8183
R22937 GNDA.n5297 GNDA.n802 65.8183
R22938 GNDA.n5297 GNDA.n800 65.8183
R22939 GNDA.n5297 GNDA.n797 65.8183
R22940 GNDA.n5297 GNDA.n796 65.8183
R22941 GNDA.n5297 GNDA.n795 65.8183
R22942 GNDA.n5297 GNDA.n793 65.8183
R22943 GNDA.n5298 GNDA.n5297 65.8183
R22944 GNDA.n5297 GNDA.n784 65.8183
R22945 GNDA.n5297 GNDA.n782 65.8183
R22946 GNDA.n5368 GNDA.n736 65.8183
R22947 GNDA.n5368 GNDA.n735 65.8183
R22948 GNDA.n5368 GNDA.n734 65.8183
R22949 GNDA.n5368 GNDA.n733 65.8183
R22950 GNDA.n5368 GNDA.n724 65.8183
R22951 GNDA.n5368 GNDA.n731 65.8183
R22952 GNDA.n5368 GNDA.n722 65.8183
R22953 GNDA.n5368 GNDA.n732 65.8183
R22954 GNDA.n5368 GNDA.n730 65.8183
R22955 GNDA.n5368 GNDA.n729 65.8183
R22956 GNDA.n5368 GNDA.n728 65.8183
R22957 GNDA.n5368 GNDA.n727 65.8183
R22958 GNDA.n5368 GNDA.n725 65.8183
R22959 GNDA.n5369 GNDA.n5368 65.8183
R22960 GNDA.n5368 GNDA.n723 65.8183
R22961 GNDA.n5368 GNDA.n721 65.8183
R22962 GNDA.n4707 GNDA.n4706 65.8183
R22963 GNDA.n4707 GNDA.n1256 65.8183
R22964 GNDA.n4707 GNDA.n1255 65.8183
R22965 GNDA.n4707 GNDA.n1254 65.8183
R22966 GNDA.n4707 GNDA.n1245 65.8183
R22967 GNDA.n4707 GNDA.n1252 65.8183
R22968 GNDA.n4707 GNDA.n1243 65.8183
R22969 GNDA.n4707 GNDA.n1253 65.8183
R22970 GNDA.n4707 GNDA.n1251 65.8183
R22971 GNDA.n4707 GNDA.n1250 65.8183
R22972 GNDA.n4707 GNDA.n1249 65.8183
R22973 GNDA.n4707 GNDA.n1248 65.8183
R22974 GNDA.n4707 GNDA.n1246 65.8183
R22975 GNDA.n4707 GNDA.n1244 65.8183
R22976 GNDA.n4708 GNDA.n4707 65.8183
R22977 GNDA.n4707 GNDA.n1238 65.8183
R22978 GNDA.n1501 GNDA.n1420 65.8183
R22979 GNDA.n1501 GNDA.n1419 65.8183
R22980 GNDA.n1501 GNDA.n1418 65.8183
R22981 GNDA.n1501 GNDA.n1417 65.8183
R22982 GNDA.n1501 GNDA.n1408 65.8183
R22983 GNDA.n1501 GNDA.n1415 65.8183
R22984 GNDA.n1501 GNDA.n1405 65.8183
R22985 GNDA.n1501 GNDA.n1416 65.8183
R22986 GNDA.n1501 GNDA.n1414 65.8183
R22987 GNDA.n1501 GNDA.n1412 65.8183
R22988 GNDA.n1501 GNDA.n1411 65.8183
R22989 GNDA.n1501 GNDA.n1410 65.8183
R22990 GNDA.n1812 GNDA.n1728 65.8183
R22991 GNDA.n1812 GNDA.n1727 65.8183
R22992 GNDA.n1812 GNDA.n1726 65.8183
R22993 GNDA.n1812 GNDA.n1725 65.8183
R22994 GNDA.n1812 GNDA.n1716 65.8183
R22995 GNDA.n1812 GNDA.n1723 65.8183
R22996 GNDA.n1812 GNDA.n1713 65.8183
R22997 GNDA.n1812 GNDA.n1724 65.8183
R22998 GNDA.n1812 GNDA.n1722 65.8183
R22999 GNDA.n1812 GNDA.n1720 65.8183
R23000 GNDA.n1812 GNDA.n1719 65.8183
R23001 GNDA.n1812 GNDA.n1718 65.8183
R23002 GNDA.n1813 GNDA.n1812 65.8183
R23003 GNDA.n1812 GNDA.n1715 65.8183
R23004 GNDA.n1812 GNDA.n1714 65.8183
R23005 GNDA.n1812 GNDA.n1712 65.8183
R23006 GNDA.n4809 GNDA.n1213 65.8183
R23007 GNDA.n4809 GNDA.n1212 65.8183
R23008 GNDA.n4809 GNDA.n1211 65.8183
R23009 GNDA.n4809 GNDA.n1210 65.8183
R23010 GNDA.n4809 GNDA.n1201 65.8183
R23011 GNDA.n4809 GNDA.n1208 65.8183
R23012 GNDA.n4809 GNDA.n1198 65.8183
R23013 GNDA.n4809 GNDA.n1209 65.8183
R23014 GNDA.n4809 GNDA.n1207 65.8183
R23015 GNDA.n4809 GNDA.n1206 65.8183
R23016 GNDA.n4809 GNDA.n1205 65.8183
R23017 GNDA.n4809 GNDA.n1204 65.8183
R23018 GNDA.n4809 GNDA.n1202 65.8183
R23019 GNDA.n4809 GNDA.n1200 65.8183
R23020 GNDA.n4809 GNDA.n1199 65.8183
R23021 GNDA.n4810 GNDA.n4809 65.8183
R23022 GNDA.n4535 GNDA.n1652 65.8183
R23023 GNDA.n4535 GNDA.n1651 65.8183
R23024 GNDA.n4535 GNDA.n1650 65.8183
R23025 GNDA.n4535 GNDA.n1649 65.8183
R23026 GNDA.n4535 GNDA.n1640 65.8183
R23027 GNDA.n4535 GNDA.n1647 65.8183
R23028 GNDA.n4535 GNDA.n1637 65.8183
R23029 GNDA.n4535 GNDA.n1648 65.8183
R23030 GNDA.n4535 GNDA.n1646 65.8183
R23031 GNDA.n4535 GNDA.n1645 65.8183
R23032 GNDA.n4535 GNDA.n1644 65.8183
R23033 GNDA.n4535 GNDA.n1643 65.8183
R23034 GNDA.n4535 GNDA.n1641 65.8183
R23035 GNDA.n4535 GNDA.n1639 65.8183
R23036 GNDA.n4535 GNDA.n1638 65.8183
R23037 GNDA.n4536 GNDA.n4535 65.8183
R23038 GNDA.n1502 GNDA.n1501 65.8183
R23039 GNDA.n1501 GNDA.n1407 65.8183
R23040 GNDA.n1501 GNDA.n1406 65.8183
R23041 GNDA.n1501 GNDA.n1404 65.8183
R23042 GNDA.n4988 GNDA.n890 65.8183
R23043 GNDA.n4990 GNDA.n890 65.8183
R23044 GNDA.n4996 GNDA.n890 65.8183
R23045 GNDA.n4998 GNDA.n890 65.8183
R23046 GNDA.n4972 GNDA.n890 65.8183
R23047 GNDA.n4974 GNDA.n890 65.8183
R23048 GNDA.n4980 GNDA.n890 65.8183
R23049 GNDA.n4982 GNDA.n890 65.8183
R23050 GNDA.n4951 GNDA.n890 65.8183
R23051 GNDA.n4957 GNDA.n890 65.8183
R23052 GNDA.n4950 GNDA.n890 65.8183
R23053 GNDA.n4964 GNDA.n890 65.8183
R23054 GNDA.n5177 GNDA.n890 65.8183
R23055 GNDA.n5174 GNDA.n890 65.8183
R23056 GNDA.n4931 GNDA.n890 65.8183
R23057 GNDA.n5010 GNDA.n890 65.8183
R23058 GNDA.n4436 GNDA.n1956 65.8183
R23059 GNDA.n4436 GNDA.n1955 65.8183
R23060 GNDA.n4436 GNDA.n1954 65.8183
R23061 GNDA.n4436 GNDA.n1953 65.8183
R23062 GNDA.n4436 GNDA.n1944 65.8183
R23063 GNDA.n4436 GNDA.n1951 65.8183
R23064 GNDA.n4436 GNDA.n1941 65.8183
R23065 GNDA.n4436 GNDA.n1952 65.8183
R23066 GNDA.n4436 GNDA.n1950 65.8183
R23067 GNDA.n4436 GNDA.n1949 65.8183
R23068 GNDA.n4436 GNDA.n1948 65.8183
R23069 GNDA.n4436 GNDA.n1947 65.8183
R23070 GNDA.n4436 GNDA.n1945 65.8183
R23071 GNDA.n4436 GNDA.n1943 65.8183
R23072 GNDA.n4436 GNDA.n1942 65.8183
R23073 GNDA.n4437 GNDA.n4436 65.8183
R23074 GNDA.n5403 GNDA.n5400 65.3505
R23075 GNDA.n5402 GNDA.n5401 65.3505
R23076 GNDA.n5425 GNDA.n5423 65.3505
R23077 GNDA.n5421 GNDA.n5419 65.3505
R23078 GNDA.n637 GNDA.n634 65.3505
R23079 GNDA.n636 GNDA.n635 65.3505
R23080 GNDA.n5471 GNDA.n666 64.0005
R23081 GNDA.n5478 GNDA.n666 64.0005
R23082 GNDA.n615 GNDA.n41 63.4011
R23083 GNDA.n619 GNDA.n618 63.4011
R23084 GNDA.n5338 GNDA.n5337 63.1009
R23085 GNDA.n644 GNDA.n642 62.2505
R23086 GNDA.n699 GNDA.n697 62.2505
R23087 GNDA.n662 GNDA.n660 62.2505
R23088 GNDA.n5451 GNDA.n5449 62.2505
R23089 GNDA.n4863 GNDA.n1138 60.9488
R23090 GNDA.n1218 GNDA.n1185 60.9488
R23091 GNDA.n3302 GNDA.n3301 59.2425
R23092 GNDA.n4279 GNDA.n1970 59.2425
R23093 GNDA.n4279 GNDA.n4278 59.2425
R23094 GNDA.n3301 GNDA.n3300 59.2425
R23095 GNDA.n5297 GNDA.n5296 57.8461
R23096 GNDA.n5368 GNDA.n5367 57.8461
R23097 GNDA.n4707 GNDA.n1237 57.8461
R23098 GNDA.n1812 GNDA.n1811 57.8461
R23099 GNDA.n4809 GNDA.n4808 57.8461
R23100 GNDA.n4535 GNDA.n4534 57.8461
R23101 GNDA.n1501 GNDA.n1500 57.8461
R23102 GNDA.n5004 GNDA.n890 57.8461
R23103 GNDA.n4436 GNDA.n4435 57.8461
R23104 GNDA.n878 GNDA.n743 57.0913
R23105 GNDA.n761 GNDA.n758 56.3995
R23106 GNDA.n940 GNDA.n939 56.3995
R23107 GNDA.n1150 GNDA.n1149 56.3995
R23108 GNDA.n1823 GNDA.n1706 56.3995
R23109 GNDA.n1190 GNDA.n1189 56.3995
R23110 GNDA.n5326 GNDA.n758 56.3995
R23111 GNDA.n1824 GNDA.n1823 56.3995
R23112 GNDA.n4349 GNDA.n4348 56.3995
R23113 GNDA.n4350 GNDA.n4349 56.3995
R23114 GNDA.n942 GNDA.n940 56.3995
R23115 GNDA.n4820 GNDA.n1190 56.3995
R23116 GNDA.n1152 GNDA.n1150 56.3995
R23117 GNDA.n5297 GNDA.n794 55.2026
R23118 GNDA.n5368 GNDA.n726 55.2026
R23119 GNDA.n4707 GNDA.n1247 55.2026
R23120 GNDA.n1501 GNDA.n1409 55.2026
R23121 GNDA.n1812 GNDA.n1717 55.2026
R23122 GNDA.n4809 GNDA.n1203 55.2026
R23123 GNDA.n4535 GNDA.n1642 55.2026
R23124 GNDA.n4966 GNDA.n890 55.2026
R23125 GNDA.n4436 GNDA.n1946 55.2026
R23126 GNDA.n5257 GNDA.n802 53.3664
R23127 GNDA.n5253 GNDA.n783 53.3664
R23128 GNDA.n5249 GNDA.n801 53.3664
R23129 GNDA.n5245 GNDA.n785 53.3664
R23130 GNDA.n5234 GNDA.n795 53.3664
R23131 GNDA.n5230 GNDA.n796 53.3664
R23132 GNDA.n5226 GNDA.n797 53.3664
R23133 GNDA.n800 GNDA.n799 53.3664
R23134 GNDA.n808 GNDA.n782 53.3664
R23135 GNDA.n5285 GNDA.n784 53.3664
R23136 GNDA.n5299 GNDA.n5298 53.3664
R23137 GNDA.n793 GNDA.n792 53.3664
R23138 GNDA.n5261 GNDA.n806 53.3664
R23139 GNDA.n5262 GNDA.n805 53.3664
R23140 GNDA.n5266 GNDA.n804 53.3664
R23141 GNDA.n5270 GNDA.n803 53.3664
R23142 GNDA.n5258 GNDA.n806 53.3664
R23143 GNDA.n5265 GNDA.n805 53.3664
R23144 GNDA.n5269 GNDA.n804 53.3664
R23145 GNDA.n5272 GNDA.n803 53.3664
R23146 GNDA.n5242 GNDA.n785 53.3664
R23147 GNDA.n5246 GNDA.n801 53.3664
R23148 GNDA.n5250 GNDA.n783 53.3664
R23149 GNDA.n5254 GNDA.n802 53.3664
R23150 GNDA.n5225 GNDA.n800 53.3664
R23151 GNDA.n5229 GNDA.n797 53.3664
R23152 GNDA.n5233 GNDA.n796 53.3664
R23153 GNDA.n5237 GNDA.n795 53.3664
R23154 GNDA.n798 GNDA.n793 53.3664
R23155 GNDA.n5298 GNDA.n781 53.3664
R23156 GNDA.n784 GNDA.n780 53.3664
R23157 GNDA.n5284 GNDA.n782 53.3664
R23158 GNDA.n5099 GNDA.n732 53.3664
R23159 GNDA.n5103 GNDA.n722 53.3664
R23160 GNDA.n5107 GNDA.n731 53.3664
R23161 GNDA.n5111 GNDA.n724 53.3664
R23162 GNDA.n5122 GNDA.n727 53.3664
R23163 GNDA.n5126 GNDA.n728 53.3664
R23164 GNDA.n5130 GNDA.n729 53.3664
R23165 GNDA.n5134 GNDA.n730 53.3664
R23166 GNDA.n738 GNDA.n721 53.3664
R23167 GNDA.n5356 GNDA.n723 53.3664
R23168 GNDA.n5370 GNDA.n5369 53.3664
R23169 GNDA.n5077 GNDA.n725 53.3664
R23170 GNDA.n5095 GNDA.n736 53.3664
R23171 GNDA.n5094 GNDA.n735 53.3664
R23172 GNDA.n5090 GNDA.n734 53.3664
R23173 GNDA.n5086 GNDA.n733 53.3664
R23174 GNDA.n5098 GNDA.n736 53.3664
R23175 GNDA.n5091 GNDA.n735 53.3664
R23176 GNDA.n5087 GNDA.n734 53.3664
R23177 GNDA.n5083 GNDA.n733 53.3664
R23178 GNDA.n5114 GNDA.n724 53.3664
R23179 GNDA.n5110 GNDA.n731 53.3664
R23180 GNDA.n5106 GNDA.n722 53.3664
R23181 GNDA.n5102 GNDA.n732 53.3664
R23182 GNDA.n5131 GNDA.n730 53.3664
R23183 GNDA.n5127 GNDA.n729 53.3664
R23184 GNDA.n5123 GNDA.n728 53.3664
R23185 GNDA.n5119 GNDA.n727 53.3664
R23186 GNDA.n5133 GNDA.n725 53.3664
R23187 GNDA.n5369 GNDA.n720 53.3664
R23188 GNDA.n723 GNDA.n719 53.3664
R23189 GNDA.n5355 GNDA.n721 53.3664
R23190 GNDA.n4689 GNDA.n1253 53.3664
R23191 GNDA.n4686 GNDA.n1243 53.3664
R23192 GNDA.n4682 GNDA.n1252 53.3664
R23193 GNDA.n4678 GNDA.n1245 53.3664
R23194 GNDA.n4667 GNDA.n1248 53.3664
R23195 GNDA.n4663 GNDA.n1249 53.3664
R23196 GNDA.n4659 GNDA.n1250 53.3664
R23197 GNDA.n4655 GNDA.n1251 53.3664
R23198 GNDA.n4716 GNDA.n1238 53.3664
R23199 GNDA.n4709 GNDA.n4708 53.3664
R23200 GNDA.n4640 GNDA.n1244 53.3664
R23201 GNDA.n4647 GNDA.n1246 53.3664
R23202 GNDA.n4706 GNDA.n4705 53.3664
R23203 GNDA.n1258 GNDA.n1256 53.3664
R23204 GNDA.n4700 GNDA.n1255 53.3664
R23205 GNDA.n4696 GNDA.n1254 53.3664
R23206 GNDA.n4706 GNDA.n1257 53.3664
R23207 GNDA.n4701 GNDA.n1256 53.3664
R23208 GNDA.n4697 GNDA.n1255 53.3664
R23209 GNDA.n4693 GNDA.n1254 53.3664
R23210 GNDA.n4675 GNDA.n1245 53.3664
R23211 GNDA.n4679 GNDA.n1252 53.3664
R23212 GNDA.n4683 GNDA.n1243 53.3664
R23213 GNDA.n4687 GNDA.n1253 53.3664
R23214 GNDA.n4658 GNDA.n1251 53.3664
R23215 GNDA.n4662 GNDA.n1250 53.3664
R23216 GNDA.n4666 GNDA.n1249 53.3664
R23217 GNDA.n4670 GNDA.n1248 53.3664
R23218 GNDA.n4654 GNDA.n1246 53.3664
R23219 GNDA.n4646 GNDA.n1244 53.3664
R23220 GNDA.n4708 GNDA.n1242 53.3664
R23221 GNDA.n1241 GNDA.n1238 53.3664
R23222 GNDA.n1455 GNDA.n1416 53.3664
R23223 GNDA.n1451 GNDA.n1405 53.3664
R23224 GNDA.n1447 GNDA.n1415 53.3664
R23225 GNDA.n1443 GNDA.n1408 53.3664
R23226 GNDA.n1432 GNDA.n1410 53.3664
R23227 GNDA.n1428 GNDA.n1411 53.3664
R23228 GNDA.n1424 GNDA.n1412 53.3664
R23229 GNDA.n1414 GNDA.n1413 53.3664
R23230 GNDA.n1473 GNDA.n1404 53.3664
R23231 GNDA.n1489 GNDA.n1406 53.3664
R23232 GNDA.n1482 GNDA.n1407 53.3664
R23233 GNDA.n1503 GNDA.n1502 53.3664
R23234 GNDA.n1459 GNDA.n1420 53.3664
R23235 GNDA.n1460 GNDA.n1419 53.3664
R23236 GNDA.n1464 GNDA.n1418 53.3664
R23237 GNDA.n1468 GNDA.n1417 53.3664
R23238 GNDA.n1456 GNDA.n1420 53.3664
R23239 GNDA.n1463 GNDA.n1419 53.3664
R23240 GNDA.n1467 GNDA.n1418 53.3664
R23241 GNDA.n1421 GNDA.n1417 53.3664
R23242 GNDA.n1440 GNDA.n1408 53.3664
R23243 GNDA.n1444 GNDA.n1415 53.3664
R23244 GNDA.n1448 GNDA.n1405 53.3664
R23245 GNDA.n1452 GNDA.n1416 53.3664
R23246 GNDA.n1423 GNDA.n1414 53.3664
R23247 GNDA.n1427 GNDA.n1412 53.3664
R23248 GNDA.n1431 GNDA.n1411 53.3664
R23249 GNDA.n1435 GNDA.n1410 53.3664
R23250 GNDA.n1764 GNDA.n1724 53.3664
R23251 GNDA.n1760 GNDA.n1713 53.3664
R23252 GNDA.n1756 GNDA.n1723 53.3664
R23253 GNDA.n1752 GNDA.n1716 53.3664
R23254 GNDA.n1741 GNDA.n1718 53.3664
R23255 GNDA.n1737 GNDA.n1719 53.3664
R23256 GNDA.n1733 GNDA.n1720 53.3664
R23257 GNDA.n1722 GNDA.n1721 53.3664
R23258 GNDA.n1730 GNDA.n1712 53.3664
R23259 GNDA.n1799 GNDA.n1714 53.3664
R23260 GNDA.n1792 GNDA.n1715 53.3664
R23261 GNDA.n1814 GNDA.n1813 53.3664
R23262 GNDA.n1768 GNDA.n1728 53.3664
R23263 GNDA.n1769 GNDA.n1727 53.3664
R23264 GNDA.n1773 GNDA.n1726 53.3664
R23265 GNDA.n1777 GNDA.n1725 53.3664
R23266 GNDA.n1765 GNDA.n1728 53.3664
R23267 GNDA.n1772 GNDA.n1727 53.3664
R23268 GNDA.n1776 GNDA.n1726 53.3664
R23269 GNDA.n1779 GNDA.n1725 53.3664
R23270 GNDA.n1749 GNDA.n1716 53.3664
R23271 GNDA.n1753 GNDA.n1723 53.3664
R23272 GNDA.n1757 GNDA.n1713 53.3664
R23273 GNDA.n1761 GNDA.n1724 53.3664
R23274 GNDA.n1732 GNDA.n1722 53.3664
R23275 GNDA.n1736 GNDA.n1720 53.3664
R23276 GNDA.n1740 GNDA.n1719 53.3664
R23277 GNDA.n1744 GNDA.n1718 53.3664
R23278 GNDA.n1813 GNDA.n1711 53.3664
R23279 GNDA.n1715 GNDA.n1710 53.3664
R23280 GNDA.n1791 GNDA.n1714 53.3664
R23281 GNDA.n1798 GNDA.n1712 53.3664
R23282 GNDA.n4790 GNDA.n1209 53.3664
R23283 GNDA.n4786 GNDA.n1198 53.3664
R23284 GNDA.n4782 GNDA.n1208 53.3664
R23285 GNDA.n4778 GNDA.n1201 53.3664
R23286 GNDA.n4767 GNDA.n1204 53.3664
R23287 GNDA.n4763 GNDA.n1205 53.3664
R23288 GNDA.n4759 GNDA.n1206 53.3664
R23289 GNDA.n4755 GNDA.n1207 53.3664
R23290 GNDA.n4811 GNDA.n4810 53.3664
R23291 GNDA.n4744 GNDA.n1199 53.3664
R23292 GNDA.n4740 GNDA.n1200 53.3664
R23293 GNDA.n4733 GNDA.n1202 53.3664
R23294 GNDA.n4794 GNDA.n1213 53.3664
R23295 GNDA.n4795 GNDA.n1212 53.3664
R23296 GNDA.n4799 GNDA.n1211 53.3664
R23297 GNDA.n4803 GNDA.n1210 53.3664
R23298 GNDA.n4791 GNDA.n1213 53.3664
R23299 GNDA.n4798 GNDA.n1212 53.3664
R23300 GNDA.n4802 GNDA.n1211 53.3664
R23301 GNDA.n4806 GNDA.n1210 53.3664
R23302 GNDA.n4775 GNDA.n1201 53.3664
R23303 GNDA.n4779 GNDA.n1208 53.3664
R23304 GNDA.n4783 GNDA.n1198 53.3664
R23305 GNDA.n4787 GNDA.n1209 53.3664
R23306 GNDA.n4758 GNDA.n1207 53.3664
R23307 GNDA.n4762 GNDA.n1206 53.3664
R23308 GNDA.n4766 GNDA.n1205 53.3664
R23309 GNDA.n4770 GNDA.n1204 53.3664
R23310 GNDA.n4754 GNDA.n1202 53.3664
R23311 GNDA.n4732 GNDA.n1200 53.3664
R23312 GNDA.n4741 GNDA.n1199 53.3664
R23313 GNDA.n4810 GNDA.n1197 53.3664
R23314 GNDA.n4516 GNDA.n1648 53.3664
R23315 GNDA.n4512 GNDA.n1637 53.3664
R23316 GNDA.n4508 GNDA.n1647 53.3664
R23317 GNDA.n4504 GNDA.n1640 53.3664
R23318 GNDA.n4493 GNDA.n1643 53.3664
R23319 GNDA.n4489 GNDA.n1644 53.3664
R23320 GNDA.n4485 GNDA.n1645 53.3664
R23321 GNDA.n4481 GNDA.n1646 53.3664
R23322 GNDA.n4537 GNDA.n4536 53.3664
R23323 GNDA.n4458 GNDA.n1638 53.3664
R23324 GNDA.n4466 GNDA.n1639 53.3664
R23325 GNDA.n4473 GNDA.n1641 53.3664
R23326 GNDA.n4520 GNDA.n1652 53.3664
R23327 GNDA.n4521 GNDA.n1651 53.3664
R23328 GNDA.n4525 GNDA.n1650 53.3664
R23329 GNDA.n4529 GNDA.n1649 53.3664
R23330 GNDA.n4517 GNDA.n1652 53.3664
R23331 GNDA.n4524 GNDA.n1651 53.3664
R23332 GNDA.n4528 GNDA.n1650 53.3664
R23333 GNDA.n4532 GNDA.n1649 53.3664
R23334 GNDA.n4501 GNDA.n1640 53.3664
R23335 GNDA.n4505 GNDA.n1647 53.3664
R23336 GNDA.n4509 GNDA.n1637 53.3664
R23337 GNDA.n4513 GNDA.n1648 53.3664
R23338 GNDA.n4484 GNDA.n1646 53.3664
R23339 GNDA.n4488 GNDA.n1645 53.3664
R23340 GNDA.n4492 GNDA.n1644 53.3664
R23341 GNDA.n4496 GNDA.n1643 53.3664
R23342 GNDA.n4480 GNDA.n1641 53.3664
R23343 GNDA.n4472 GNDA.n1639 53.3664
R23344 GNDA.n4465 GNDA.n1638 53.3664
R23345 GNDA.n4536 GNDA.n1636 53.3664
R23346 GNDA.n1502 GNDA.n1403 53.3664
R23347 GNDA.n1407 GNDA.n1402 53.3664
R23348 GNDA.n1481 GNDA.n1406 53.3664
R23349 GNDA.n1488 GNDA.n1404 53.3664
R23350 GNDA.n4982 GNDA.n4942 53.3664
R23351 GNDA.n4981 GNDA.n4980 53.3664
R23352 GNDA.n4974 GNDA.n4944 53.3664
R23353 GNDA.n4973 GNDA.n4972 53.3664
R23354 GNDA.n4964 GNDA.n4963 53.3664
R23355 GNDA.n4959 GNDA.n4950 53.3664
R23356 GNDA.n4957 GNDA.n4956 53.3664
R23357 GNDA.n4951 GNDA.n889 53.3664
R23358 GNDA.n5010 GNDA.n5009 53.3664
R23359 GNDA.n4937 GNDA.n4931 53.3664
R23360 GNDA.n5174 GNDA.n5173 53.3664
R23361 GNDA.n5177 GNDA.n5176 53.3664
R23362 GNDA.n4989 GNDA.n4988 53.3664
R23363 GNDA.n4991 GNDA.n4990 53.3664
R23364 GNDA.n4996 GNDA.n4995 53.3664
R23365 GNDA.n4999 GNDA.n4998 53.3664
R23366 GNDA.n4988 GNDA.n4987 53.3664
R23367 GNDA.n4990 GNDA.n4940 53.3664
R23368 GNDA.n4997 GNDA.n4996 53.3664
R23369 GNDA.n4998 GNDA.n4938 53.3664
R23370 GNDA.n4972 GNDA.n4971 53.3664
R23371 GNDA.n4975 GNDA.n4974 53.3664
R23372 GNDA.n4980 GNDA.n4979 53.3664
R23373 GNDA.n4983 GNDA.n4982 53.3664
R23374 GNDA.n4952 GNDA.n4951 53.3664
R23375 GNDA.n4958 GNDA.n4957 53.3664
R23376 GNDA.n4950 GNDA.n4948 53.3664
R23377 GNDA.n4965 GNDA.n4964 53.3664
R23378 GNDA.n5178 GNDA.n5177 53.3664
R23379 GNDA.n5175 GNDA.n5174 53.3664
R23380 GNDA.n4931 GNDA.n893 53.3664
R23381 GNDA.n5011 GNDA.n5010 53.3664
R23382 GNDA.n4417 GNDA.n1952 53.3664
R23383 GNDA.n4413 GNDA.n1941 53.3664
R23384 GNDA.n4409 GNDA.n1951 53.3664
R23385 GNDA.n4405 GNDA.n1944 53.3664
R23386 GNDA.n4394 GNDA.n1947 53.3664
R23387 GNDA.n4390 GNDA.n1948 53.3664
R23388 GNDA.n4386 GNDA.n1949 53.3664
R23389 GNDA.n4382 GNDA.n1950 53.3664
R23390 GNDA.n4438 GNDA.n4437 53.3664
R23391 GNDA.n4359 GNDA.n1942 53.3664
R23392 GNDA.n4367 GNDA.n1943 53.3664
R23393 GNDA.n4374 GNDA.n1945 53.3664
R23394 GNDA.n4421 GNDA.n1956 53.3664
R23395 GNDA.n4422 GNDA.n1955 53.3664
R23396 GNDA.n4426 GNDA.n1954 53.3664
R23397 GNDA.n4430 GNDA.n1953 53.3664
R23398 GNDA.n4418 GNDA.n1956 53.3664
R23399 GNDA.n4425 GNDA.n1955 53.3664
R23400 GNDA.n4429 GNDA.n1954 53.3664
R23401 GNDA.n4433 GNDA.n1953 53.3664
R23402 GNDA.n4402 GNDA.n1944 53.3664
R23403 GNDA.n4406 GNDA.n1951 53.3664
R23404 GNDA.n4410 GNDA.n1941 53.3664
R23405 GNDA.n4414 GNDA.n1952 53.3664
R23406 GNDA.n4385 GNDA.n1950 53.3664
R23407 GNDA.n4389 GNDA.n1949 53.3664
R23408 GNDA.n4393 GNDA.n1948 53.3664
R23409 GNDA.n4397 GNDA.n1947 53.3664
R23410 GNDA.n4381 GNDA.n1945 53.3664
R23411 GNDA.n4373 GNDA.n1943 53.3664
R23412 GNDA.n4366 GNDA.n1942 53.3664
R23413 GNDA.n4437 GNDA.n1940 53.3664
R23414 GNDA.n5025 GNDA.n945 53.085
R23415 GNDA.n878 GNDA.n877 53.085
R23416 GNDA.n5143 GNDA.n5140 53.085
R23417 GNDA.n1554 GNDA.n1536 50.8806
R23418 GNDA.n1560 GNDA.n1536 50.8806
R23419 GNDA.n1561 GNDA.n1560 50.8806
R23420 GNDA.n1563 GNDA.n1561 50.8806
R23421 GNDA.n1563 GNDA.n1562 50.8806
R23422 GNDA.n1570 GNDA.n1569 50.8806
R23423 GNDA.n1571 GNDA.n1570 50.8806
R23424 GNDA.n1571 GNDA.n1528 50.8806
R23425 GNDA.n1578 GNDA.n1528 50.8806
R23426 GNDA.n1579 GNDA.n1578 50.8806
R23427 GNDA.n1593 GNDA.n1592 50.8806
R23428 GNDA.n1592 GNDA.n1591 50.8806
R23429 GNDA.n1591 GNDA.n1581 50.8806
R23430 GNDA.n1585 GNDA.n1581 50.8806
R23431 GNDA.n1585 GNDA.n1114 50.8806
R23432 GNDA.n4880 GNDA.n1117 50.8806
R23433 GNDA.n4874 GNDA.n1117 50.8806
R23434 GNDA.n4874 GNDA.n4873 50.8806
R23435 GNDA.n4873 GNDA.n4872 50.8806
R23436 GNDA.n4872 GNDA.n1122 50.8806
R23437 GNDA.n4302 GNDA.n4299 50.8806
R23438 GNDA.n4303 GNDA.n4302 50.8806
R23439 GNDA.n4304 GNDA.n4303 50.8806
R23440 GNDA.n4304 GNDA.n4295 50.8806
R23441 GNDA.n4310 GNDA.n4295 50.8806
R23442 GNDA.n4313 GNDA.n4312 50.8806
R23443 GNDA.n4313 GNDA.n4291 50.8806
R23444 GNDA.n4319 GNDA.n4291 50.8806
R23445 GNDA.n4320 GNDA.n4319 50.8806
R23446 GNDA.n4321 GNDA.n4320 50.8806
R23447 GNDA.n5042 GNDA.n895 47.0754
R23448 GNDA.n5375 GNDA.n714 47.0754
R23449 GNDA.n585 GNDA.n584 44.1991
R23450 GNDA.n587 GNDA.n586 44.1991
R23451 GNDA.n877 GNDA.n823 43.069
R23452 GNDA.n5375 GNDA.n5374 43.069
R23453 GNDA.n5304 GNDA.n5303 43.069
R23454 GNDA.n5481 GNDA.n5479 42.6297
R23455 GNDA.n5469 GNDA.n5467 42.6297
R23456 GNDA.n32 GNDA.n30 42.6297
R23457 GNDA.n583 GNDA.n581 42.6297
R23458 GNDA.n5026 GNDA.n5025 37.0595
R23459 GNDA.n5143 GNDA.n5139 37.0595
R23460 GNDA.n5165 GNDA.n5152 33.0531
R23461 GNDA.n5318 GNDA.n5317 32.3969
R23462 GNDA.n4883 GNDA.n1112 31.3605
R23463 GNDA.n2205 GNDA.n2204 31.1255
R23464 GNDA.n2200 GNDA.n2199 31.1255
R23465 GNDA.n3617 GNDA.n3616 31.1255
R23466 GNDA.n3622 GNDA.n3621 31.1255
R23467 GNDA.n5349 GNDA.n743 30.0483
R23468 GNDA.n5259 GNDA.n5256 27.5561
R23469 GNDA.n5100 GNDA.n5097 27.5561
R23470 GNDA.n4691 GNDA.n4690 27.5561
R23471 GNDA.n1457 GNDA.n1454 27.5561
R23472 GNDA.n1766 GNDA.n1763 27.5561
R23473 GNDA.n4792 GNDA.n4789 27.5561
R23474 GNDA.n4518 GNDA.n4515 27.5561
R23475 GNDA.n4986 GNDA.n4985 27.5561
R23476 GNDA.n4419 GNDA.n4416 27.5561
R23477 GNDA.n5140 GNDA.n821 27.0435
R23478 GNDA.n5315 GNDA.n771 27.0435
R23479 GNDA.n5338 GNDA.n752 27.0435
R23480 GNDA.n4847 GNDA.n1138 26.9584
R23481 GNDA.n4749 GNDA.n1218 26.9584
R23482 GNDA.n5240 GNDA.n5239 26.6672
R23483 GNDA.n5117 GNDA.n5116 26.6672
R23484 GNDA.n4673 GNDA.n4672 26.6672
R23485 GNDA.n1438 GNDA.n1437 26.6672
R23486 GNDA.n1747 GNDA.n1746 26.6672
R23487 GNDA.n4773 GNDA.n4772 26.6672
R23488 GNDA.n4499 GNDA.n4498 26.6672
R23489 GNDA.n4969 GNDA.n4968 26.6672
R23490 GNDA.n4400 GNDA.n4399 26.6672
R23491 GNDA.n1562 GNDA.n1532 26.5712
R23492 GNDA.n4881 GNDA.n1114 26.5712
R23493 GNDA.n4311 GNDA.n4310 26.5712
R23494 GNDA.n1569 GNDA.n1532 24.3099
R23495 GNDA.n4881 GNDA.n4880 24.3099
R23496 GNDA.n4312 GNDA.n4311 24.3099
R23497 GNDA.n5165 GNDA.n5153 23.3628
R23498 GNDA.n5168 GNDA.n5167 23.0371
R23499 GNDA.n820 GNDA.n748 22.53
R23500 GNDA.n5514 GNDA.n625 20.9529
R23501 GNDA.n5341 GNDA.n5339 20.8233
R23502 GNDA.n5218 GNDA.n750 20.8233
R23503 GNDA.n5348 GNDA.n5347 20.8233
R23504 GNDA.n876 GNDA.n875 20.8233
R23505 GNDA.n5019 GNDA.n5017 20.8233
R23506 GNDA.n5024 GNDA.n5023 20.8233
R23507 GNDA.n5167 GNDA.n5042 20.0324
R23508 GNDA.n5219 GNDA.n5216 20.0324
R23509 GNDA.n5315 GNDA.n5304 20.0324
R23510 GNDA.n4921 GNDA.n4919 18.591
R23511 GNDA.n1287 GNDA.n1261 17.5843
R23512 GNDA.n1849 GNDA.n1693 17.5843
R23513 GNDA.n4324 GNDA.n4323 17.5843
R23514 GNDA.n4329 GNDA.n4328 17.5479
R23515 GNDA.n1544 GNDA.n1540 17.5479
R23516 GNDA.n1556 GNDA.n1538 16.9379
R23517 GNDA.n4843 GNDA.n1178 16.9379
R23518 GNDA.n926 GNDA.n922 16.9379
R23519 GNDA.n4548 GNDA.n4547 16.7709
R23520 GNDA.n5211 GNDA.n847 16.7709
R23521 GNDA.n4448 GNDA.n1899 16.7709
R23522 GNDA.n4630 GNDA.n1377 16.7709
R23523 GNDA.n5260 GNDA.n5259 16.0005
R23524 GNDA.n5263 GNDA.n5260 16.0005
R23525 GNDA.n5264 GNDA.n5263 16.0005
R23526 GNDA.n5267 GNDA.n5264 16.0005
R23527 GNDA.n5268 GNDA.n5267 16.0005
R23528 GNDA.n5271 GNDA.n5268 16.0005
R23529 GNDA.n5273 GNDA.n5271 16.0005
R23530 GNDA.n5274 GNDA.n5273 16.0005
R23531 GNDA.n5256 GNDA.n5255 16.0005
R23532 GNDA.n5255 GNDA.n5252 16.0005
R23533 GNDA.n5252 GNDA.n5251 16.0005
R23534 GNDA.n5251 GNDA.n5248 16.0005
R23535 GNDA.n5248 GNDA.n5247 16.0005
R23536 GNDA.n5247 GNDA.n5244 16.0005
R23537 GNDA.n5244 GNDA.n5243 16.0005
R23538 GNDA.n5243 GNDA.n5240 16.0005
R23539 GNDA.n5239 GNDA.n5236 16.0005
R23540 GNDA.n5236 GNDA.n5235 16.0005
R23541 GNDA.n5235 GNDA.n5232 16.0005
R23542 GNDA.n5232 GNDA.n5231 16.0005
R23543 GNDA.n5231 GNDA.n5228 16.0005
R23544 GNDA.n5228 GNDA.n5227 16.0005
R23545 GNDA.n5227 GNDA.n5224 16.0005
R23546 GNDA.n5224 GNDA.n757 16.0005
R23547 GNDA.n5097 GNDA.n5096 16.0005
R23548 GNDA.n5096 GNDA.n5093 16.0005
R23549 GNDA.n5093 GNDA.n5092 16.0005
R23550 GNDA.n5092 GNDA.n5089 16.0005
R23551 GNDA.n5089 GNDA.n5088 16.0005
R23552 GNDA.n5088 GNDA.n5085 16.0005
R23553 GNDA.n5085 GNDA.n5084 16.0005
R23554 GNDA.n5084 GNDA.n5082 16.0005
R23555 GNDA.n5101 GNDA.n5100 16.0005
R23556 GNDA.n5104 GNDA.n5101 16.0005
R23557 GNDA.n5105 GNDA.n5104 16.0005
R23558 GNDA.n5108 GNDA.n5105 16.0005
R23559 GNDA.n5109 GNDA.n5108 16.0005
R23560 GNDA.n5112 GNDA.n5109 16.0005
R23561 GNDA.n5113 GNDA.n5112 16.0005
R23562 GNDA.n5116 GNDA.n5113 16.0005
R23563 GNDA.n5120 GNDA.n5117 16.0005
R23564 GNDA.n5121 GNDA.n5120 16.0005
R23565 GNDA.n5124 GNDA.n5121 16.0005
R23566 GNDA.n5125 GNDA.n5124 16.0005
R23567 GNDA.n5128 GNDA.n5125 16.0005
R23568 GNDA.n5129 GNDA.n5128 16.0005
R23569 GNDA.n5132 GNDA.n5129 16.0005
R23570 GNDA.n5135 GNDA.n5132 16.0005
R23571 GNDA.n4704 GNDA.n4691 16.0005
R23572 GNDA.n4704 GNDA.n4703 16.0005
R23573 GNDA.n4703 GNDA.n4702 16.0005
R23574 GNDA.n4702 GNDA.n4699 16.0005
R23575 GNDA.n4699 GNDA.n4698 16.0005
R23576 GNDA.n4698 GNDA.n4695 16.0005
R23577 GNDA.n4695 GNDA.n4694 16.0005
R23578 GNDA.n4694 GNDA.n1234 16.0005
R23579 GNDA.n4690 GNDA.n4688 16.0005
R23580 GNDA.n4688 GNDA.n4685 16.0005
R23581 GNDA.n4685 GNDA.n4684 16.0005
R23582 GNDA.n4684 GNDA.n4681 16.0005
R23583 GNDA.n4681 GNDA.n4680 16.0005
R23584 GNDA.n4680 GNDA.n4677 16.0005
R23585 GNDA.n4677 GNDA.n4676 16.0005
R23586 GNDA.n4676 GNDA.n4673 16.0005
R23587 GNDA.n4672 GNDA.n4669 16.0005
R23588 GNDA.n4669 GNDA.n4668 16.0005
R23589 GNDA.n4668 GNDA.n4665 16.0005
R23590 GNDA.n4665 GNDA.n4664 16.0005
R23591 GNDA.n4664 GNDA.n4661 16.0005
R23592 GNDA.n4661 GNDA.n4660 16.0005
R23593 GNDA.n4660 GNDA.n4657 16.0005
R23594 GNDA.n4657 GNDA.n4656 16.0005
R23595 GNDA.n1458 GNDA.n1457 16.0005
R23596 GNDA.n1461 GNDA.n1458 16.0005
R23597 GNDA.n1462 GNDA.n1461 16.0005
R23598 GNDA.n1465 GNDA.n1462 16.0005
R23599 GNDA.n1466 GNDA.n1465 16.0005
R23600 GNDA.n1469 GNDA.n1466 16.0005
R23601 GNDA.n1470 GNDA.n1469 16.0005
R23602 GNDA.n1471 GNDA.n1470 16.0005
R23603 GNDA.n1454 GNDA.n1453 16.0005
R23604 GNDA.n1453 GNDA.n1450 16.0005
R23605 GNDA.n1450 GNDA.n1449 16.0005
R23606 GNDA.n1449 GNDA.n1446 16.0005
R23607 GNDA.n1446 GNDA.n1445 16.0005
R23608 GNDA.n1445 GNDA.n1442 16.0005
R23609 GNDA.n1442 GNDA.n1441 16.0005
R23610 GNDA.n1441 GNDA.n1438 16.0005
R23611 GNDA.n1437 GNDA.n1434 16.0005
R23612 GNDA.n1434 GNDA.n1433 16.0005
R23613 GNDA.n1433 GNDA.n1430 16.0005
R23614 GNDA.n1430 GNDA.n1429 16.0005
R23615 GNDA.n1429 GNDA.n1426 16.0005
R23616 GNDA.n1426 GNDA.n1425 16.0005
R23617 GNDA.n1425 GNDA.n1422 16.0005
R23618 GNDA.n1422 GNDA.n1399 16.0005
R23619 GNDA.n1767 GNDA.n1766 16.0005
R23620 GNDA.n1770 GNDA.n1767 16.0005
R23621 GNDA.n1771 GNDA.n1770 16.0005
R23622 GNDA.n1774 GNDA.n1771 16.0005
R23623 GNDA.n1775 GNDA.n1774 16.0005
R23624 GNDA.n1778 GNDA.n1775 16.0005
R23625 GNDA.n1780 GNDA.n1778 16.0005
R23626 GNDA.n1781 GNDA.n1780 16.0005
R23627 GNDA.n1763 GNDA.n1762 16.0005
R23628 GNDA.n1762 GNDA.n1759 16.0005
R23629 GNDA.n1759 GNDA.n1758 16.0005
R23630 GNDA.n1758 GNDA.n1755 16.0005
R23631 GNDA.n1755 GNDA.n1754 16.0005
R23632 GNDA.n1754 GNDA.n1751 16.0005
R23633 GNDA.n1751 GNDA.n1750 16.0005
R23634 GNDA.n1750 GNDA.n1747 16.0005
R23635 GNDA.n1746 GNDA.n1743 16.0005
R23636 GNDA.n1743 GNDA.n1742 16.0005
R23637 GNDA.n1742 GNDA.n1739 16.0005
R23638 GNDA.n1739 GNDA.n1738 16.0005
R23639 GNDA.n1738 GNDA.n1735 16.0005
R23640 GNDA.n1735 GNDA.n1734 16.0005
R23641 GNDA.n1734 GNDA.n1731 16.0005
R23642 GNDA.n1731 GNDA.n1707 16.0005
R23643 GNDA.n4793 GNDA.n4792 16.0005
R23644 GNDA.n4796 GNDA.n4793 16.0005
R23645 GNDA.n4797 GNDA.n4796 16.0005
R23646 GNDA.n4800 GNDA.n4797 16.0005
R23647 GNDA.n4801 GNDA.n4800 16.0005
R23648 GNDA.n4804 GNDA.n4801 16.0005
R23649 GNDA.n4805 GNDA.n4804 16.0005
R23650 GNDA.n4805 GNDA.n1192 16.0005
R23651 GNDA.n4789 GNDA.n4788 16.0005
R23652 GNDA.n4788 GNDA.n4785 16.0005
R23653 GNDA.n4785 GNDA.n4784 16.0005
R23654 GNDA.n4784 GNDA.n4781 16.0005
R23655 GNDA.n4781 GNDA.n4780 16.0005
R23656 GNDA.n4780 GNDA.n4777 16.0005
R23657 GNDA.n4777 GNDA.n4776 16.0005
R23658 GNDA.n4776 GNDA.n4773 16.0005
R23659 GNDA.n4772 GNDA.n4769 16.0005
R23660 GNDA.n4769 GNDA.n4768 16.0005
R23661 GNDA.n4768 GNDA.n4765 16.0005
R23662 GNDA.n4765 GNDA.n4764 16.0005
R23663 GNDA.n4764 GNDA.n4761 16.0005
R23664 GNDA.n4761 GNDA.n4760 16.0005
R23665 GNDA.n4760 GNDA.n4757 16.0005
R23666 GNDA.n4757 GNDA.n4756 16.0005
R23667 GNDA.n4519 GNDA.n4518 16.0005
R23668 GNDA.n4522 GNDA.n4519 16.0005
R23669 GNDA.n4523 GNDA.n4522 16.0005
R23670 GNDA.n4526 GNDA.n4523 16.0005
R23671 GNDA.n4527 GNDA.n4526 16.0005
R23672 GNDA.n4530 GNDA.n4527 16.0005
R23673 GNDA.n4531 GNDA.n4530 16.0005
R23674 GNDA.n4531 GNDA.n1632 16.0005
R23675 GNDA.n4515 GNDA.n4514 16.0005
R23676 GNDA.n4514 GNDA.n4511 16.0005
R23677 GNDA.n4511 GNDA.n4510 16.0005
R23678 GNDA.n4510 GNDA.n4507 16.0005
R23679 GNDA.n4507 GNDA.n4506 16.0005
R23680 GNDA.n4506 GNDA.n4503 16.0005
R23681 GNDA.n4503 GNDA.n4502 16.0005
R23682 GNDA.n4502 GNDA.n4499 16.0005
R23683 GNDA.n4498 GNDA.n4495 16.0005
R23684 GNDA.n4495 GNDA.n4494 16.0005
R23685 GNDA.n4494 GNDA.n4491 16.0005
R23686 GNDA.n4491 GNDA.n4490 16.0005
R23687 GNDA.n4490 GNDA.n4487 16.0005
R23688 GNDA.n4487 GNDA.n4486 16.0005
R23689 GNDA.n4486 GNDA.n4483 16.0005
R23690 GNDA.n4483 GNDA.n4482 16.0005
R23691 GNDA.n4986 GNDA.n4941 16.0005
R23692 GNDA.n4992 GNDA.n4941 16.0005
R23693 GNDA.n4993 GNDA.n4992 16.0005
R23694 GNDA.n4994 GNDA.n4993 16.0005
R23695 GNDA.n4994 GNDA.n4939 16.0005
R23696 GNDA.n5000 GNDA.n4939 16.0005
R23697 GNDA.n5001 GNDA.n5000 16.0005
R23698 GNDA.n5002 GNDA.n5001 16.0005
R23699 GNDA.n4985 GNDA.n4984 16.0005
R23700 GNDA.n4984 GNDA.n4943 16.0005
R23701 GNDA.n4978 GNDA.n4943 16.0005
R23702 GNDA.n4978 GNDA.n4977 16.0005
R23703 GNDA.n4977 GNDA.n4976 16.0005
R23704 GNDA.n4976 GNDA.n4945 16.0005
R23705 GNDA.n4970 GNDA.n4945 16.0005
R23706 GNDA.n4970 GNDA.n4969 16.0005
R23707 GNDA.n4968 GNDA.n4947 16.0005
R23708 GNDA.n4962 GNDA.n4947 16.0005
R23709 GNDA.n4962 GNDA.n4961 16.0005
R23710 GNDA.n4961 GNDA.n4960 16.0005
R23711 GNDA.n4960 GNDA.n4949 16.0005
R23712 GNDA.n4955 GNDA.n4949 16.0005
R23713 GNDA.n4955 GNDA.n4954 16.0005
R23714 GNDA.n4954 GNDA.n4953 16.0005
R23715 GNDA.n4420 GNDA.n4419 16.0005
R23716 GNDA.n4423 GNDA.n4420 16.0005
R23717 GNDA.n4424 GNDA.n4423 16.0005
R23718 GNDA.n4427 GNDA.n4424 16.0005
R23719 GNDA.n4428 GNDA.n4427 16.0005
R23720 GNDA.n4431 GNDA.n4428 16.0005
R23721 GNDA.n4432 GNDA.n4431 16.0005
R23722 GNDA.n4432 GNDA.n1936 16.0005
R23723 GNDA.n4416 GNDA.n4415 16.0005
R23724 GNDA.n4415 GNDA.n4412 16.0005
R23725 GNDA.n4412 GNDA.n4411 16.0005
R23726 GNDA.n4411 GNDA.n4408 16.0005
R23727 GNDA.n4408 GNDA.n4407 16.0005
R23728 GNDA.n4407 GNDA.n4404 16.0005
R23729 GNDA.n4404 GNDA.n4403 16.0005
R23730 GNDA.n4403 GNDA.n4400 16.0005
R23731 GNDA.n4399 GNDA.n4396 16.0005
R23732 GNDA.n4396 GNDA.n4395 16.0005
R23733 GNDA.n4395 GNDA.n4392 16.0005
R23734 GNDA.n4392 GNDA.n4391 16.0005
R23735 GNDA.n4391 GNDA.n4388 16.0005
R23736 GNDA.n4388 GNDA.n4387 16.0005
R23737 GNDA.n4387 GNDA.n4384 16.0005
R23738 GNDA.n4384 GNDA.n4383 16.0005
R23739 GNDA.n5407 GNDA.n5406 14.238
R23740 GNDA.n641 GNDA.n640 14.238
R23741 GNDA.n5141 GNDA.n5069 12.8005
R23742 GNDA.n5145 GNDA.n5069 12.8005
R23743 GNDA.n5057 GNDA.n5056 12.8005
R23744 GNDA.n5061 GNDA.n5056 12.8005
R23745 GNDA.n1115 GNDA.n1111 12.8005
R23746 GNDA.n4883 GNDA.n1111 12.8005
R23747 GNDA.n5462 GNDA.n676 12.8005
R23748 GNDA.n5458 GNDA.n676 12.8005
R23749 GNDA.n677 GNDA.n675 12.8005
R23750 GNDA.n5455 GNDA.n677 12.8005
R23751 GNDA.n5509 GNDA.n630 12.8005
R23752 GNDA.n5509 GNDA.n5508 12.8005
R23753 GNDA.n5396 GNDA.n703 12.8005
R23754 GNDA.n5408 GNDA.n5396 12.8005
R23755 GNDA.n590 GNDA.n36 12.8005
R23756 GNDA.n5525 GNDA.n36 12.8005
R23757 GNDA.n596 GNDA.n595 12.8005
R23758 GNDA.n596 GNDA.n37 12.8005
R23759 GNDA.n3300 GNDA.n3299 12.6791
R23760 GNDA.n3302 GNDA.n2114 12.6791
R23761 GNDA.n4278 GNDA.n1971 12.6791
R23762 GNDA.n1970 GNDA.n1969 12.6791
R23763 GNDA.n1265 GNDA.n1261 11.6369
R23764 GNDA.n1280 GNDA.n1265 11.6369
R23765 GNDA.n1280 GNDA.n1279 11.6369
R23766 GNDA.n1279 GNDA.n1278 11.6369
R23767 GNDA.n1278 GNDA.n1266 11.6369
R23768 GNDA.n1273 GNDA.n1266 11.6369
R23769 GNDA.n1273 GNDA.n1272 11.6369
R23770 GNDA.n1272 GNDA.n1271 11.6369
R23771 GNDA.n1271 GNDA.n759 11.6369
R23772 GNDA.n5331 GNDA.n759 11.6369
R23773 GNDA.n1308 GNDA.n1307 11.6369
R23774 GNDA.n1307 GNDA.n1304 11.6369
R23775 GNDA.n1304 GNDA.n1303 11.6369
R23776 GNDA.n1303 GNDA.n1300 11.6369
R23777 GNDA.n1300 GNDA.n1299 11.6369
R23778 GNDA.n1299 GNDA.n1296 11.6369
R23779 GNDA.n1296 GNDA.n1295 11.6369
R23780 GNDA.n1295 GNDA.n1292 11.6369
R23781 GNDA.n1292 GNDA.n1291 11.6369
R23782 GNDA.n1291 GNDA.n1288 11.6369
R23783 GNDA.n1288 GNDA.n1287 11.6369
R23784 GNDA.n1309 GNDA.n846 11.6369
R23785 GNDA.n1312 GNDA.n1309 11.6369
R23786 GNDA.n1313 GNDA.n1312 11.6369
R23787 GNDA.n1316 GNDA.n1313 11.6369
R23788 GNDA.n1317 GNDA.n1316 11.6369
R23789 GNDA.n1320 GNDA.n1317 11.6369
R23790 GNDA.n1321 GNDA.n1320 11.6369
R23791 GNDA.n1324 GNDA.n1321 11.6369
R23792 GNDA.n1325 GNDA.n1324 11.6369
R23793 GNDA.n1328 GNDA.n1325 11.6369
R23794 GNDA.n1329 GNDA.n1328 11.6369
R23795 GNDA.n1557 GNDA.n1556 11.6369
R23796 GNDA.n1558 GNDA.n1557 11.6369
R23797 GNDA.n1558 GNDA.n1534 11.6369
R23798 GNDA.n1565 GNDA.n1534 11.6369
R23799 GNDA.n1566 GNDA.n1565 11.6369
R23800 GNDA.n1567 GNDA.n1566 11.6369
R23801 GNDA.n1567 GNDA.n1530 11.6369
R23802 GNDA.n1573 GNDA.n1530 11.6369
R23803 GNDA.n1574 GNDA.n1573 11.6369
R23804 GNDA.n1576 GNDA.n1574 11.6369
R23805 GNDA.n1576 GNDA.n1575 11.6369
R23806 GNDA.n1550 GNDA.n1538 11.6369
R23807 GNDA.n1550 GNDA.n1549 11.6369
R23808 GNDA.n1549 GNDA.n1548 11.6369
R23809 GNDA.n1548 GNDA.n1542 11.6369
R23810 GNDA.n1542 GNDA.n1145 11.6369
R23811 GNDA.n4860 GNDA.n1145 11.6369
R23812 GNDA.n4860 GNDA.n4859 11.6369
R23813 GNDA.n4859 GNDA.n4858 11.6369
R23814 GNDA.n4858 GNDA.n1146 11.6369
R23815 GNDA.n4852 GNDA.n1146 11.6369
R23816 GNDA.n1696 GNDA.n1693 11.6369
R23817 GNDA.n1699 GNDA.n1696 11.6369
R23818 GNDA.n1841 GNDA.n1699 11.6369
R23819 GNDA.n1841 GNDA.n1840 11.6369
R23820 GNDA.n1840 GNDA.n1839 11.6369
R23821 GNDA.n1839 GNDA.n1700 11.6369
R23822 GNDA.n1704 GNDA.n1700 11.6369
R23823 GNDA.n1831 GNDA.n1704 11.6369
R23824 GNDA.n1831 GNDA.n1830 11.6369
R23825 GNDA.n1830 GNDA.n1829 11.6369
R23826 GNDA.n1865 GNDA.n1655 11.6369
R23827 GNDA.n1865 GNDA.n1864 11.6369
R23828 GNDA.n1864 GNDA.n1863 11.6369
R23829 GNDA.n1863 GNDA.n1687 11.6369
R23830 GNDA.n1858 GNDA.n1687 11.6369
R23831 GNDA.n1858 GNDA.n1857 11.6369
R23832 GNDA.n1857 GNDA.n1856 11.6369
R23833 GNDA.n1856 GNDA.n1690 11.6369
R23834 GNDA.n1851 GNDA.n1690 11.6369
R23835 GNDA.n1851 GNDA.n1850 11.6369
R23836 GNDA.n1850 GNDA.n1849 11.6369
R23837 GNDA.n1663 GNDA.n1397 11.6369
R23838 GNDA.n1664 GNDA.n1663 11.6369
R23839 GNDA.n1664 GNDA.n1660 11.6369
R23840 GNDA.n1670 GNDA.n1660 11.6369
R23841 GNDA.n1671 GNDA.n1670 11.6369
R23842 GNDA.n1672 GNDA.n1671 11.6369
R23843 GNDA.n1672 GNDA.n1658 11.6369
R23844 GNDA.n1678 GNDA.n1658 11.6369
R23845 GNDA.n1679 GNDA.n1678 11.6369
R23846 GNDA.n1680 GNDA.n1679 11.6369
R23847 GNDA.n1680 GNDA.n1656 11.6369
R23848 GNDA.n4843 GNDA.n4842 11.6369
R23849 GNDA.n4842 GNDA.n4841 11.6369
R23850 GNDA.n4841 GNDA.n1179 11.6369
R23851 GNDA.n4835 GNDA.n1179 11.6369
R23852 GNDA.n4835 GNDA.n4834 11.6369
R23853 GNDA.n4834 GNDA.n4833 11.6369
R23854 GNDA.n4833 GNDA.n1183 11.6369
R23855 GNDA.n4827 GNDA.n1183 11.6369
R23856 GNDA.n4827 GNDA.n4826 11.6369
R23857 GNDA.n4826 GNDA.n4825 11.6369
R23858 GNDA.n4554 GNDA.n1178 11.6369
R23859 GNDA.n4559 GNDA.n4554 11.6369
R23860 GNDA.n4560 GNDA.n4559 11.6369
R23861 GNDA.n4561 GNDA.n4560 11.6369
R23862 GNDA.n4561 GNDA.n4552 11.6369
R23863 GNDA.n4567 GNDA.n4552 11.6369
R23864 GNDA.n4568 GNDA.n4567 11.6369
R23865 GNDA.n4569 GNDA.n4568 11.6369
R23866 GNDA.n4569 GNDA.n4550 11.6369
R23867 GNDA.n4574 GNDA.n4550 11.6369
R23868 GNDA.n4575 GNDA.n4574 11.6369
R23869 GNDA.n927 GNDA.n926 11.6369
R23870 GNDA.n928 GNDA.n927 11.6369
R23871 GNDA.n928 GNDA.n900 11.6369
R23872 GNDA.n934 GNDA.n900 11.6369
R23873 GNDA.n935 GNDA.n934 11.6369
R23874 GNDA.n5039 GNDA.n935 11.6369
R23875 GNDA.n5039 GNDA.n5038 11.6369
R23876 GNDA.n5038 GNDA.n5037 11.6369
R23877 GNDA.n5037 GNDA.n936 11.6369
R23878 GNDA.n5031 GNDA.n936 11.6369
R23879 GNDA.n922 GNDA.n921 11.6369
R23880 GNDA.n921 GNDA.n918 11.6369
R23881 GNDA.n918 GNDA.n917 11.6369
R23882 GNDA.n917 GNDA.n914 11.6369
R23883 GNDA.n914 GNDA.n913 11.6369
R23884 GNDA.n913 GNDA.n910 11.6369
R23885 GNDA.n910 GNDA.n909 11.6369
R23886 GNDA.n909 GNDA.n906 11.6369
R23887 GNDA.n906 GNDA.n905 11.6369
R23888 GNDA.n905 GNDA.n845 11.6369
R23889 GNDA.n5212 GNDA.n845 11.6369
R23890 GNDA.n4325 GNDA.n4324 11.6369
R23891 GNDA.n4325 GNDA.n1963 11.6369
R23892 GNDA.n4333 GNDA.n1963 11.6369
R23893 GNDA.n4334 GNDA.n4333 11.6369
R23894 GNDA.n4335 GNDA.n4334 11.6369
R23895 GNDA.n4335 GNDA.n1961 11.6369
R23896 GNDA.n4340 GNDA.n1961 11.6369
R23897 GNDA.n4341 GNDA.n4340 11.6369
R23898 GNDA.n4343 GNDA.n4341 11.6369
R23899 GNDA.n4343 GNDA.n4342 11.6369
R23900 GNDA.n4300 GNDA.n1124 11.6369
R23901 GNDA.n4300 GNDA.n4297 11.6369
R23902 GNDA.n4306 GNDA.n4297 11.6369
R23903 GNDA.n4307 GNDA.n4306 11.6369
R23904 GNDA.n4308 GNDA.n4307 11.6369
R23905 GNDA.n4308 GNDA.n4293 11.6369
R23906 GNDA.n4315 GNDA.n4293 11.6369
R23907 GNDA.n4316 GNDA.n4315 11.6369
R23908 GNDA.n4317 GNDA.n4316 11.6369
R23909 GNDA.n4317 GNDA.n4289 11.6369
R23910 GNDA.n4323 GNDA.n4289 11.6369
R23911 GNDA.n1583 GNDA.n1527 11.6369
R23912 GNDA.n1589 GNDA.n1583 11.6369
R23913 GNDA.n1589 GNDA.n1588 11.6369
R23914 GNDA.n1588 GNDA.n1587 11.6369
R23915 GNDA.n1587 GNDA.n1584 11.6369
R23916 GNDA.n4878 GNDA.n4877 11.6369
R23917 GNDA.n4877 GNDA.n4876 11.6369
R23918 GNDA.n4876 GNDA.n1120 11.6369
R23919 GNDA.n4870 GNDA.n1120 11.6369
R23920 GNDA.n4870 GNDA.n4869 11.6369
R23921 GNDA.n5342 GNDA.n5341 11.3283
R23922 GNDA.n4922 GNDA.n4921 10.87
R23923 GNDA.n5023 GNDA.n5021 10.87
R23924 GNDA.n5020 GNDA.n5019 10.87
R23925 GNDA.n875 GNDA.n745 10.87
R23926 GNDA.n5347 GNDA.n5345 10.87
R23927 GNDA.n5343 GNDA.n748 10.87
R23928 GNDA.n5342 GNDA.n750 10.87
R23929 GNDA.n5482 GNDA.n5478 9.42329
R23930 GNDA.n5471 GNDA.n5470 9.42293
R23931 GNDA.n5141 GNDA.n5067 9.36264
R23932 GNDA.n5057 GNDA.n5054 9.36264
R23933 GNDA.n1115 GNDA.n1109 9.36264
R23934 GNDA.n703 GNDA.n700 9.36264
R23935 GNDA.n5459 GNDA.n5458 9.36264
R23936 GNDA.n5452 GNDA.n675 9.36264
R23937 GNDA.n5508 GNDA.n5507 9.36264
R23938 GNDA.n595 GNDA.n589 9.36264
R23939 GNDA.n590 GNDA.n34 9.36264
R23940 GNDA.n5069 GNDA.n5068 9.3005
R23941 GNDA.n5146 GNDA.n5145 9.3005
R23942 GNDA.n5056 GNDA.n5055 9.3005
R23943 GNDA.n5062 GNDA.n5061 9.3005
R23944 GNDA.n1111 GNDA.n1110 9.3005
R23945 GNDA.n4884 GNDA.n4883 9.3005
R23946 GNDA.n5460 GNDA.n676 9.3005
R23947 GNDA.n5462 GNDA.n5461 9.3005
R23948 GNDA.n678 GNDA.n677 9.3005
R23949 GNDA.n5455 GNDA.n5454 9.3005
R23950 GNDA.n5509 GNDA.n631 9.3005
R23951 GNDA.n645 GNDA.n630 9.3005
R23952 GNDA.n5396 GNDA.n701 9.3005
R23953 GNDA.n5409 GNDA.n5408 9.3005
R23954 GNDA.n36 GNDA.n35 9.3005
R23955 GNDA.n5526 GNDA.n5525 9.3005
R23956 GNDA.n597 GNDA.n596 9.3005
R23957 GNDA.n598 GNDA.n37 9.3005
R23958 GNDA.n1377 GNDA.n1329 6.72373
R23959 GNDA.n1575 GNDA.n1525 6.72373
R23960 GNDA.n1899 GNDA.n1656 6.72373
R23961 GNDA.n4575 GNDA.n4548 6.72373
R23962 GNDA.n5212 GNDA.n5211 6.72373
R23963 GNDA.n4869 GNDA.n4868 6.72373
R23964 GNDA.n1377 GNDA.n1308 6.20656
R23965 GNDA.n5211 GNDA.n846 6.20656
R23966 GNDA.n1899 GNDA.n1655 6.20656
R23967 GNDA.n4548 GNDA.n1397 6.20656
R23968 GNDA.n4868 GNDA.n1124 6.20656
R23969 GNDA.n1527 GNDA.n1525 6.20656
R23970 GNDA.n1584 GNDA.n1112 6.07727
R23971 GNDA.n5313 GNDA.n5306 5.81868
R23972 GNDA.n5313 GNDA.n5308 5.81868
R23973 GNDA.n5165 GNDA.n5164 5.81868
R23974 GNDA.n5164 GNDA.n5155 5.81868
R23975 GNDA.n5160 GNDA.n5155 5.81868
R23976 GNDA.n4878 GNDA.n1112 5.5601
R23977 GNDA.n5334 GNDA.n757 5.51161
R23978 GNDA.n5136 GNDA.n5135 5.51161
R23979 GNDA.n4656 GNDA.n4634 5.51161
R23980 GNDA.n1509 GNDA.n1399 5.51161
R23981 GNDA.n1820 GNDA.n1707 5.51161
R23982 GNDA.n4756 GNDA.n1214 5.51161
R23983 GNDA.n4482 GNDA.n4452 5.51161
R23984 GNDA.n4953 GNDA.n882 5.51161
R23985 GNDA.n4383 GNDA.n4353 5.51161
R23986 GNDA.n5333 GNDA.n5332 5.1717
R23987 GNDA.n1821 GNDA.n1705 5.1717
R23988 GNDA.n4352 GNDA.n1957 5.1717
R23989 GNDA.n4818 GNDA.n1188 4.9157
R23990 GNDA.n4851 GNDA.n4850 4.9157
R23991 GNDA.n5030 GNDA.n5029 4.9157
R23992 GNDA.n5506 GNDA.n644 4.663
R23993 GNDA.n5410 GNDA.n699 4.663
R23994 GNDA.n663 GNDA.n662 4.663
R23995 GNDA.n5453 GNDA.n5451 4.663
R23996 GNDA.n5406 GNDA.n5399 4.64112
R23997 GNDA.n5406 GNDA.n5405 4.64112
R23998 GNDA.n640 GNDA.n633 4.64112
R23999 GNDA.n640 GNDA.n639 4.64112
R24000 GNDA.n2216 GNDA.n2215 4.5005
R24001 GNDA.n2112 GNDA.n2111 4.5005
R24002 GNDA.n2033 GNDA.n2032 4.5005
R24003 GNDA.n2055 GNDA.n2034 4.5005
R24004 GNDA.n2056 GNDA.n2035 4.5005
R24005 GNDA.n2057 GNDA.n2036 4.5005
R24006 GNDA.n2058 GNDA.n2037 4.5005
R24007 GNDA.n2059 GNDA.n2038 4.5005
R24008 GNDA.n2060 GNDA.n2039 4.5005
R24009 GNDA.n2061 GNDA.n2040 4.5005
R24010 GNDA.n2062 GNDA.n2041 4.5005
R24011 GNDA.n2063 GNDA.n2042 4.5005
R24012 GNDA.n2064 GNDA.n2043 4.5005
R24013 GNDA.n2065 GNDA.n2044 4.5005
R24014 GNDA.n2066 GNDA.n2045 4.5005
R24015 GNDA.n2067 GNDA.n2046 4.5005
R24016 GNDA.n2068 GNDA.n2047 4.5005
R24017 GNDA.n2069 GNDA.n2048 4.5005
R24018 GNDA.n2070 GNDA.n2049 4.5005
R24019 GNDA.n2071 GNDA.n2050 4.5005
R24020 GNDA.n2072 GNDA.n2051 4.5005
R24021 GNDA.n2073 GNDA.n2052 4.5005
R24022 GNDA.n2074 GNDA.n2053 4.5005
R24023 GNDA.n4147 GNDA.n4146 4.5005
R24024 GNDA.n4145 GNDA.n3661 4.5005
R24025 GNDA.n4144 GNDA.n4143 4.5005
R24026 GNDA.n4142 GNDA.n3665 4.5005
R24027 GNDA.n4141 GNDA.n4140 4.5005
R24028 GNDA.n4139 GNDA.n3666 4.5005
R24029 GNDA.n4138 GNDA.n4137 4.5005
R24030 GNDA.n4136 GNDA.n3670 4.5005
R24031 GNDA.n4135 GNDA.n4134 4.5005
R24032 GNDA.n4133 GNDA.n3671 4.5005
R24033 GNDA.n4132 GNDA.n4131 4.5005
R24034 GNDA.n4130 GNDA.n3675 4.5005
R24035 GNDA.n4129 GNDA.n4128 4.5005
R24036 GNDA.n4127 GNDA.n3676 4.5005
R24037 GNDA.n4126 GNDA.n4125 4.5005
R24038 GNDA.n4124 GNDA.n3680 4.5005
R24039 GNDA.n4123 GNDA.n4122 4.5005
R24040 GNDA.n4121 GNDA.n3681 4.5005
R24041 GNDA.n4120 GNDA.n4119 4.5005
R24042 GNDA.n4118 GNDA.n3685 4.5005
R24043 GNDA.n4117 GNDA.n4116 4.5005
R24044 GNDA.n4115 GNDA.n3686 4.5005
R24045 GNDA.n4048 GNDA.n3656 4.5005
R24046 GNDA.n4051 GNDA.n4050 4.5005
R24047 GNDA.n4052 GNDA.n4045 4.5005
R24048 GNDA.n4054 GNDA.n4053 4.5005
R24049 GNDA.n4055 GNDA.n4044 4.5005
R24050 GNDA.n4059 GNDA.n4058 4.5005
R24051 GNDA.n4060 GNDA.n4041 4.5005
R24052 GNDA.n4062 GNDA.n4061 4.5005
R24053 GNDA.n4063 GNDA.n4040 4.5005
R24054 GNDA.n4067 GNDA.n4066 4.5005
R24055 GNDA.n4068 GNDA.n4037 4.5005
R24056 GNDA.n4070 GNDA.n4069 4.5005
R24057 GNDA.n4071 GNDA.n4036 4.5005
R24058 GNDA.n4075 GNDA.n4074 4.5005
R24059 GNDA.n4076 GNDA.n4033 4.5005
R24060 GNDA.n4078 GNDA.n4077 4.5005
R24061 GNDA.n4079 GNDA.n4032 4.5005
R24062 GNDA.n4083 GNDA.n4082 4.5005
R24063 GNDA.n4084 GNDA.n4029 4.5005
R24064 GNDA.n4086 GNDA.n4085 4.5005
R24065 GNDA.n4087 GNDA.n4028 4.5005
R24066 GNDA.n4091 GNDA.n4090 4.5005
R24067 GNDA.n3967 GNDA.n3651 4.5005
R24068 GNDA.n3970 GNDA.n3969 4.5005
R24069 GNDA.n3971 GNDA.n3964 4.5005
R24070 GNDA.n3973 GNDA.n3972 4.5005
R24071 GNDA.n3974 GNDA.n3963 4.5005
R24072 GNDA.n3978 GNDA.n3977 4.5005
R24073 GNDA.n3979 GNDA.n3960 4.5005
R24074 GNDA.n3981 GNDA.n3980 4.5005
R24075 GNDA.n3982 GNDA.n3959 4.5005
R24076 GNDA.n3986 GNDA.n3985 4.5005
R24077 GNDA.n3987 GNDA.n3956 4.5005
R24078 GNDA.n3989 GNDA.n3988 4.5005
R24079 GNDA.n3990 GNDA.n3955 4.5005
R24080 GNDA.n3994 GNDA.n3993 4.5005
R24081 GNDA.n3995 GNDA.n3952 4.5005
R24082 GNDA.n3997 GNDA.n3996 4.5005
R24083 GNDA.n3998 GNDA.n3951 4.5005
R24084 GNDA.n4002 GNDA.n4001 4.5005
R24085 GNDA.n4003 GNDA.n3948 4.5005
R24086 GNDA.n4005 GNDA.n4004 4.5005
R24087 GNDA.n4006 GNDA.n3947 4.5005
R24088 GNDA.n4010 GNDA.n4009 4.5005
R24089 GNDA.n3886 GNDA.n3646 4.5005
R24090 GNDA.n3889 GNDA.n3888 4.5005
R24091 GNDA.n3890 GNDA.n3883 4.5005
R24092 GNDA.n3892 GNDA.n3891 4.5005
R24093 GNDA.n3893 GNDA.n3882 4.5005
R24094 GNDA.n3897 GNDA.n3896 4.5005
R24095 GNDA.n3898 GNDA.n3879 4.5005
R24096 GNDA.n3900 GNDA.n3899 4.5005
R24097 GNDA.n3901 GNDA.n3878 4.5005
R24098 GNDA.n3905 GNDA.n3904 4.5005
R24099 GNDA.n3906 GNDA.n3875 4.5005
R24100 GNDA.n3908 GNDA.n3907 4.5005
R24101 GNDA.n3909 GNDA.n3874 4.5005
R24102 GNDA.n3913 GNDA.n3912 4.5005
R24103 GNDA.n3914 GNDA.n3871 4.5005
R24104 GNDA.n3916 GNDA.n3915 4.5005
R24105 GNDA.n3917 GNDA.n3870 4.5005
R24106 GNDA.n3921 GNDA.n3920 4.5005
R24107 GNDA.n3922 GNDA.n3867 4.5005
R24108 GNDA.n3924 GNDA.n3923 4.5005
R24109 GNDA.n3925 GNDA.n3866 4.5005
R24110 GNDA.n3929 GNDA.n3928 4.5005
R24111 GNDA.n4190 GNDA.n4189 4.5005
R24112 GNDA.n4193 GNDA.n4192 4.5005
R24113 GNDA.n4194 GNDA.n3506 4.5005
R24114 GNDA.n4196 GNDA.n4195 4.5005
R24115 GNDA.n4197 GNDA.n3505 4.5005
R24116 GNDA.n4201 GNDA.n4200 4.5005
R24117 GNDA.n4202 GNDA.n3502 4.5005
R24118 GNDA.n4204 GNDA.n4203 4.5005
R24119 GNDA.n4205 GNDA.n3501 4.5005
R24120 GNDA.n4209 GNDA.n4208 4.5005
R24121 GNDA.n4210 GNDA.n3498 4.5005
R24122 GNDA.n4212 GNDA.n4211 4.5005
R24123 GNDA.n4213 GNDA.n3497 4.5005
R24124 GNDA.n4217 GNDA.n4216 4.5005
R24125 GNDA.n4218 GNDA.n3494 4.5005
R24126 GNDA.n4220 GNDA.n4219 4.5005
R24127 GNDA.n4221 GNDA.n3493 4.5005
R24128 GNDA.n4225 GNDA.n4224 4.5005
R24129 GNDA.n4226 GNDA.n3490 4.5005
R24130 GNDA.n4228 GNDA.n4227 4.5005
R24131 GNDA.n4229 GNDA.n3489 4.5005
R24132 GNDA.n4233 GNDA.n4232 4.5005
R24133 GNDA.n3805 GNDA.n3604 4.5005
R24134 GNDA.n3808 GNDA.n3807 4.5005
R24135 GNDA.n3809 GNDA.n3802 4.5005
R24136 GNDA.n3811 GNDA.n3810 4.5005
R24137 GNDA.n3812 GNDA.n3801 4.5005
R24138 GNDA.n3816 GNDA.n3815 4.5005
R24139 GNDA.n3817 GNDA.n3798 4.5005
R24140 GNDA.n3819 GNDA.n3818 4.5005
R24141 GNDA.n3820 GNDA.n3797 4.5005
R24142 GNDA.n3824 GNDA.n3823 4.5005
R24143 GNDA.n3825 GNDA.n3794 4.5005
R24144 GNDA.n3827 GNDA.n3826 4.5005
R24145 GNDA.n3828 GNDA.n3793 4.5005
R24146 GNDA.n3832 GNDA.n3831 4.5005
R24147 GNDA.n3833 GNDA.n3790 4.5005
R24148 GNDA.n3835 GNDA.n3834 4.5005
R24149 GNDA.n3836 GNDA.n3789 4.5005
R24150 GNDA.n3840 GNDA.n3839 4.5005
R24151 GNDA.n3841 GNDA.n3786 4.5005
R24152 GNDA.n3843 GNDA.n3842 4.5005
R24153 GNDA.n3844 GNDA.n3785 4.5005
R24154 GNDA.n3848 GNDA.n3847 4.5005
R24155 GNDA.n3724 GNDA.n3599 4.5005
R24156 GNDA.n3727 GNDA.n3726 4.5005
R24157 GNDA.n3728 GNDA.n3721 4.5005
R24158 GNDA.n3730 GNDA.n3729 4.5005
R24159 GNDA.n3731 GNDA.n3720 4.5005
R24160 GNDA.n3735 GNDA.n3734 4.5005
R24161 GNDA.n3736 GNDA.n3717 4.5005
R24162 GNDA.n3738 GNDA.n3737 4.5005
R24163 GNDA.n3739 GNDA.n3716 4.5005
R24164 GNDA.n3743 GNDA.n3742 4.5005
R24165 GNDA.n3744 GNDA.n3713 4.5005
R24166 GNDA.n3746 GNDA.n3745 4.5005
R24167 GNDA.n3747 GNDA.n3712 4.5005
R24168 GNDA.n3751 GNDA.n3750 4.5005
R24169 GNDA.n3752 GNDA.n3709 4.5005
R24170 GNDA.n3754 GNDA.n3753 4.5005
R24171 GNDA.n3755 GNDA.n3708 4.5005
R24172 GNDA.n3759 GNDA.n3758 4.5005
R24173 GNDA.n3760 GNDA.n3705 4.5005
R24174 GNDA.n3762 GNDA.n3761 4.5005
R24175 GNDA.n3763 GNDA.n3704 4.5005
R24176 GNDA.n3767 GNDA.n3766 4.5005
R24177 GNDA.n3594 GNDA.n3593 4.5005
R24178 GNDA.n3592 GNDA.n3514 4.5005
R24179 GNDA.n3591 GNDA.n3590 4.5005
R24180 GNDA.n3589 GNDA.n3519 4.5005
R24181 GNDA.n3588 GNDA.n3587 4.5005
R24182 GNDA.n3586 GNDA.n3520 4.5005
R24183 GNDA.n3585 GNDA.n3584 4.5005
R24184 GNDA.n3583 GNDA.n3527 4.5005
R24185 GNDA.n3582 GNDA.n3581 4.5005
R24186 GNDA.n3580 GNDA.n3528 4.5005
R24187 GNDA.n3579 GNDA.n3578 4.5005
R24188 GNDA.n3577 GNDA.n3535 4.5005
R24189 GNDA.n3576 GNDA.n3575 4.5005
R24190 GNDA.n3574 GNDA.n3536 4.5005
R24191 GNDA.n3573 GNDA.n3572 4.5005
R24192 GNDA.n3571 GNDA.n3543 4.5005
R24193 GNDA.n3570 GNDA.n3569 4.5005
R24194 GNDA.n3568 GNDA.n3544 4.5005
R24195 GNDA.n3567 GNDA.n3566 4.5005
R24196 GNDA.n3565 GNDA.n3551 4.5005
R24197 GNDA.n3564 GNDA.n3563 4.5005
R24198 GNDA.n3562 GNDA.n3552 4.5005
R24199 GNDA.n4273 GNDA.n4272 4.5005
R24200 GNDA.n4271 GNDA.n1974 4.5005
R24201 GNDA.n4270 GNDA.n4269 4.5005
R24202 GNDA.n4268 GNDA.n1978 4.5005
R24203 GNDA.n4267 GNDA.n4266 4.5005
R24204 GNDA.n4265 GNDA.n1979 4.5005
R24205 GNDA.n4264 GNDA.n4263 4.5005
R24206 GNDA.n4262 GNDA.n1983 4.5005
R24207 GNDA.n4261 GNDA.n4260 4.5005
R24208 GNDA.n4259 GNDA.n1984 4.5005
R24209 GNDA.n4258 GNDA.n4257 4.5005
R24210 GNDA.n4256 GNDA.n1988 4.5005
R24211 GNDA.n4255 GNDA.n4254 4.5005
R24212 GNDA.n4253 GNDA.n1989 4.5005
R24213 GNDA.n4252 GNDA.n4251 4.5005
R24214 GNDA.n4250 GNDA.n1993 4.5005
R24215 GNDA.n4249 GNDA.n4248 4.5005
R24216 GNDA.n4247 GNDA.n1994 4.5005
R24217 GNDA.n4246 GNDA.n4245 4.5005
R24218 GNDA.n4244 GNDA.n1998 4.5005
R24219 GNDA.n4243 GNDA.n4242 4.5005
R24220 GNDA.n4241 GNDA.n1999 4.5005
R24221 GNDA.n3632 GNDA.n3631 4.5005
R24222 GNDA.n3638 GNDA.n3626 4.5005
R24223 GNDA.n3639 GNDA.n3608 4.5005
R24224 GNDA.n3639 GNDA.n3638 4.5005
R24225 GNDA.n5063 GNDA.n5062 4.5005
R24226 GNDA.n5147 GNDA.n5146 4.5005
R24227 GNDA.n5053 GNDA.n5052 4.5005
R24228 GNDA.n5152 GNDA.n5046 4.5005
R24229 GNDA.n5151 GNDA.n767 4.5005
R24230 GNDA.n5152 GNDA.n5151 4.5005
R24231 GNDA.n1067 GNDA.n1061 4.5005
R24232 GNDA.n1069 GNDA.n1068 4.5005
R24233 GNDA.n1070 GNDA.n1060 4.5005
R24234 GNDA.n1074 GNDA.n1073 4.5005
R24235 GNDA.n1075 GNDA.n1057 4.5005
R24236 GNDA.n1077 GNDA.n1076 4.5005
R24237 GNDA.n1078 GNDA.n1056 4.5005
R24238 GNDA.n1082 GNDA.n1081 4.5005
R24239 GNDA.n1083 GNDA.n1053 4.5005
R24240 GNDA.n1085 GNDA.n1084 4.5005
R24241 GNDA.n1086 GNDA.n1052 4.5005
R24242 GNDA.n1090 GNDA.n1089 4.5005
R24243 GNDA.n1091 GNDA.n1049 4.5005
R24244 GNDA.n1093 GNDA.n1092 4.5005
R24245 GNDA.n1094 GNDA.n1048 4.5005
R24246 GNDA.n1098 GNDA.n1097 4.5005
R24247 GNDA.n1099 GNDA.n1045 4.5005
R24248 GNDA.n1101 GNDA.n1100 4.5005
R24249 GNDA.n1102 GNDA.n1044 4.5005
R24250 GNDA.n1106 GNDA.n1105 4.5005
R24251 GNDA.n1107 GNDA.n1043 4.5005
R24252 GNDA.n4894 GNDA.n4893 4.5005
R24253 GNDA.n766 GNDA.n765 4.5005
R24254 GNDA.n4887 GNDA.n4886 4.5005
R24255 GNDA.n4890 GNDA.n763 4.5005
R24256 GNDA.n4886 GNDA.n763 4.5005
R24257 GNDA.n4885 GNDA.n4884 4.5005
R24258 GNDA.n4180 GNDA.n3511 4.5005
R24259 GNDA.n4179 GNDA.n4178 4.5005
R24260 GNDA.n4180 GNDA.n4179 4.5005
R24261 GNDA.n4176 GNDA.n3596 4.5005
R24262 GNDA.n4175 GNDA.n4174 4.5005
R24263 GNDA.n4176 GNDA.n4175 4.5005
R24264 GNDA.n4172 GNDA.n3601 4.5005
R24265 GNDA.n4171 GNDA.n4170 4.5005
R24266 GNDA.n4172 GNDA.n4171 4.5005
R24267 GNDA.n4184 GNDA.n1973 4.5005
R24268 GNDA.n4188 GNDA.n4187 4.5005
R24269 GNDA.n4188 GNDA.n1973 4.5005
R24270 GNDA.n4164 GNDA.n3643 4.5005
R24271 GNDA.n4163 GNDA.n4162 4.5005
R24272 GNDA.n4164 GNDA.n4163 4.5005
R24273 GNDA.n4160 GNDA.n3648 4.5005
R24274 GNDA.n4159 GNDA.n4158 4.5005
R24275 GNDA.n4160 GNDA.n4159 4.5005
R24276 GNDA.n4156 GNDA.n3653 4.5005
R24277 GNDA.n4155 GNDA.n4154 4.5005
R24278 GNDA.n4156 GNDA.n4155 4.5005
R24279 GNDA.n4152 GNDA.n3658 4.5005
R24280 GNDA.n4151 GNDA.n4150 4.5005
R24281 GNDA.n4152 GNDA.n4151 4.5005
R24282 GNDA.n4165 GNDA.n3640 4.5005
R24283 GNDA.n4168 GNDA.n3640 4.5005
R24284 GNDA.n4168 GNDA.n3606 4.5005
R24285 GNDA.n3397 GNDA.n3396 4.5005
R24286 GNDA.n3401 GNDA.n3400 4.5005
R24287 GNDA.n3404 GNDA.n3403 4.5005
R24288 GNDA.n3405 GNDA.n3392 4.5005
R24289 GNDA.n3409 GNDA.n3406 4.5005
R24290 GNDA.n3410 GNDA.n3391 4.5005
R24291 GNDA.n3414 GNDA.n3413 4.5005
R24292 GNDA.n3415 GNDA.n3390 4.5005
R24293 GNDA.n3419 GNDA.n3416 4.5005
R24294 GNDA.n3420 GNDA.n3389 4.5005
R24295 GNDA.n3424 GNDA.n3423 4.5005
R24296 GNDA.n3425 GNDA.n3388 4.5005
R24297 GNDA.n3429 GNDA.n3426 4.5005
R24298 GNDA.n3430 GNDA.n3387 4.5005
R24299 GNDA.n3434 GNDA.n3433 4.5005
R24300 GNDA.n3435 GNDA.n3386 4.5005
R24301 GNDA.n3439 GNDA.n3436 4.5005
R24302 GNDA.n3440 GNDA.n3385 4.5005
R24303 GNDA.n3444 GNDA.n3443 4.5005
R24304 GNDA.n3445 GNDA.n3384 4.5005
R24305 GNDA.n3449 GNDA.n3446 4.5005
R24306 GNDA.n3450 GNDA.n3383 4.5005
R24307 GNDA.n3454 GNDA.n3453 4.5005
R24308 GNDA.n3312 GNDA.n3311 4.5005
R24309 GNDA.n3315 GNDA.n3314 4.5005
R24310 GNDA.n3316 GNDA.n2027 4.5005
R24311 GNDA.n3320 GNDA.n3317 4.5005
R24312 GNDA.n3321 GNDA.n2026 4.5005
R24313 GNDA.n3325 GNDA.n3324 4.5005
R24314 GNDA.n3326 GNDA.n2025 4.5005
R24315 GNDA.n3330 GNDA.n3327 4.5005
R24316 GNDA.n3331 GNDA.n2024 4.5005
R24317 GNDA.n3335 GNDA.n3334 4.5005
R24318 GNDA.n3336 GNDA.n2023 4.5005
R24319 GNDA.n3340 GNDA.n3337 4.5005
R24320 GNDA.n3341 GNDA.n2022 4.5005
R24321 GNDA.n3345 GNDA.n3344 4.5005
R24322 GNDA.n3346 GNDA.n2021 4.5005
R24323 GNDA.n3350 GNDA.n3347 4.5005
R24324 GNDA.n3351 GNDA.n2020 4.5005
R24325 GNDA.n3355 GNDA.n3354 4.5005
R24326 GNDA.n3356 GNDA.n2019 4.5005
R24327 GNDA.n3360 GNDA.n3357 4.5005
R24328 GNDA.n3361 GNDA.n2018 4.5005
R24329 GNDA.n3365 GNDA.n3364 4.5005
R24330 GNDA.n3288 GNDA.n3287 4.5005
R24331 GNDA.n2120 GNDA.n2119 4.5005
R24332 GNDA.n3233 GNDA.n3232 4.5005
R24333 GNDA.n3237 GNDA.n3234 4.5005
R24334 GNDA.n3238 GNDA.n3231 4.5005
R24335 GNDA.n3242 GNDA.n3241 4.5005
R24336 GNDA.n3243 GNDA.n3230 4.5005
R24337 GNDA.n3247 GNDA.n3244 4.5005
R24338 GNDA.n3248 GNDA.n3229 4.5005
R24339 GNDA.n3252 GNDA.n3251 4.5005
R24340 GNDA.n3253 GNDA.n3228 4.5005
R24341 GNDA.n3257 GNDA.n3254 4.5005
R24342 GNDA.n3258 GNDA.n3227 4.5005
R24343 GNDA.n3262 GNDA.n3261 4.5005
R24344 GNDA.n3263 GNDA.n3226 4.5005
R24345 GNDA.n3267 GNDA.n3264 4.5005
R24346 GNDA.n3268 GNDA.n3225 4.5005
R24347 GNDA.n3272 GNDA.n3271 4.5005
R24348 GNDA.n3273 GNDA.n3224 4.5005
R24349 GNDA.n3277 GNDA.n3274 4.5005
R24350 GNDA.n3278 GNDA.n3223 4.5005
R24351 GNDA.n3282 GNDA.n3281 4.5005
R24352 GNDA.n3153 GNDA.n3152 4.5005
R24353 GNDA.n3156 GNDA.n3155 4.5005
R24354 GNDA.n3157 GNDA.n2146 4.5005
R24355 GNDA.n3161 GNDA.n3158 4.5005
R24356 GNDA.n3162 GNDA.n2145 4.5005
R24357 GNDA.n3166 GNDA.n3165 4.5005
R24358 GNDA.n3167 GNDA.n2144 4.5005
R24359 GNDA.n3171 GNDA.n3168 4.5005
R24360 GNDA.n3172 GNDA.n2143 4.5005
R24361 GNDA.n3176 GNDA.n3175 4.5005
R24362 GNDA.n3177 GNDA.n2142 4.5005
R24363 GNDA.n3181 GNDA.n3178 4.5005
R24364 GNDA.n3182 GNDA.n2141 4.5005
R24365 GNDA.n3186 GNDA.n3185 4.5005
R24366 GNDA.n3187 GNDA.n2140 4.5005
R24367 GNDA.n3191 GNDA.n3188 4.5005
R24368 GNDA.n3192 GNDA.n2139 4.5005
R24369 GNDA.n3196 GNDA.n3195 4.5005
R24370 GNDA.n3197 GNDA.n2138 4.5005
R24371 GNDA.n3201 GNDA.n3198 4.5005
R24372 GNDA.n3202 GNDA.n2137 4.5005
R24373 GNDA.n3206 GNDA.n3205 4.5005
R24374 GNDA.n3141 GNDA.n3140 4.5005
R24375 GNDA.n3062 GNDA.n3061 4.5005
R24376 GNDA.n3084 GNDA.n3063 4.5005
R24377 GNDA.n3085 GNDA.n3064 4.5005
R24378 GNDA.n3086 GNDA.n3065 4.5005
R24379 GNDA.n3087 GNDA.n3066 4.5005
R24380 GNDA.n3088 GNDA.n3067 4.5005
R24381 GNDA.n3089 GNDA.n3068 4.5005
R24382 GNDA.n3090 GNDA.n3069 4.5005
R24383 GNDA.n3091 GNDA.n3070 4.5005
R24384 GNDA.n3092 GNDA.n3071 4.5005
R24385 GNDA.n3093 GNDA.n3072 4.5005
R24386 GNDA.n3094 GNDA.n3073 4.5005
R24387 GNDA.n3095 GNDA.n3074 4.5005
R24388 GNDA.n3096 GNDA.n3075 4.5005
R24389 GNDA.n3097 GNDA.n3076 4.5005
R24390 GNDA.n3098 GNDA.n3077 4.5005
R24391 GNDA.n3099 GNDA.n3078 4.5005
R24392 GNDA.n3100 GNDA.n3079 4.5005
R24393 GNDA.n3101 GNDA.n3080 4.5005
R24394 GNDA.n3102 GNDA.n3081 4.5005
R24395 GNDA.n3103 GNDA.n3082 4.5005
R24396 GNDA.n3054 GNDA.n3053 4.5005
R24397 GNDA.n2159 GNDA.n2158 4.5005
R24398 GNDA.n2999 GNDA.n2998 4.5005
R24399 GNDA.n3003 GNDA.n3000 4.5005
R24400 GNDA.n3004 GNDA.n2997 4.5005
R24401 GNDA.n3008 GNDA.n3007 4.5005
R24402 GNDA.n3009 GNDA.n2996 4.5005
R24403 GNDA.n3013 GNDA.n3010 4.5005
R24404 GNDA.n3014 GNDA.n2995 4.5005
R24405 GNDA.n3018 GNDA.n3017 4.5005
R24406 GNDA.n3019 GNDA.n2994 4.5005
R24407 GNDA.n3023 GNDA.n3020 4.5005
R24408 GNDA.n3024 GNDA.n2993 4.5005
R24409 GNDA.n3028 GNDA.n3027 4.5005
R24410 GNDA.n3029 GNDA.n2992 4.5005
R24411 GNDA.n3033 GNDA.n3030 4.5005
R24412 GNDA.n3034 GNDA.n2991 4.5005
R24413 GNDA.n3038 GNDA.n3037 4.5005
R24414 GNDA.n3039 GNDA.n2990 4.5005
R24415 GNDA.n3043 GNDA.n3040 4.5005
R24416 GNDA.n3044 GNDA.n2989 4.5005
R24417 GNDA.n3048 GNDA.n3047 4.5005
R24418 GNDA.n2919 GNDA.n2918 4.5005
R24419 GNDA.n2922 GNDA.n2921 4.5005
R24420 GNDA.n2923 GNDA.n2185 4.5005
R24421 GNDA.n2927 GNDA.n2924 4.5005
R24422 GNDA.n2928 GNDA.n2184 4.5005
R24423 GNDA.n2932 GNDA.n2931 4.5005
R24424 GNDA.n2933 GNDA.n2183 4.5005
R24425 GNDA.n2937 GNDA.n2934 4.5005
R24426 GNDA.n2938 GNDA.n2182 4.5005
R24427 GNDA.n2942 GNDA.n2941 4.5005
R24428 GNDA.n2943 GNDA.n2181 4.5005
R24429 GNDA.n2947 GNDA.n2944 4.5005
R24430 GNDA.n2948 GNDA.n2180 4.5005
R24431 GNDA.n2952 GNDA.n2951 4.5005
R24432 GNDA.n2953 GNDA.n2179 4.5005
R24433 GNDA.n2957 GNDA.n2954 4.5005
R24434 GNDA.n2958 GNDA.n2178 4.5005
R24435 GNDA.n2962 GNDA.n2961 4.5005
R24436 GNDA.n2963 GNDA.n2177 4.5005
R24437 GNDA.n2967 GNDA.n2964 4.5005
R24438 GNDA.n2968 GNDA.n2176 4.5005
R24439 GNDA.n2972 GNDA.n2971 4.5005
R24440 GNDA.n2907 GNDA.n2906 4.5005
R24441 GNDA.n2828 GNDA.n2827 4.5005
R24442 GNDA.n2850 GNDA.n2829 4.5005
R24443 GNDA.n2851 GNDA.n2830 4.5005
R24444 GNDA.n2852 GNDA.n2831 4.5005
R24445 GNDA.n2853 GNDA.n2832 4.5005
R24446 GNDA.n2854 GNDA.n2833 4.5005
R24447 GNDA.n2855 GNDA.n2834 4.5005
R24448 GNDA.n2856 GNDA.n2835 4.5005
R24449 GNDA.n2857 GNDA.n2836 4.5005
R24450 GNDA.n2858 GNDA.n2837 4.5005
R24451 GNDA.n2859 GNDA.n2838 4.5005
R24452 GNDA.n2860 GNDA.n2839 4.5005
R24453 GNDA.n2861 GNDA.n2840 4.5005
R24454 GNDA.n2862 GNDA.n2841 4.5005
R24455 GNDA.n2863 GNDA.n2842 4.5005
R24456 GNDA.n2864 GNDA.n2843 4.5005
R24457 GNDA.n2865 GNDA.n2844 4.5005
R24458 GNDA.n2866 GNDA.n2845 4.5005
R24459 GNDA.n2867 GNDA.n2846 4.5005
R24460 GNDA.n2868 GNDA.n2847 4.5005
R24461 GNDA.n2869 GNDA.n2848 4.5005
R24462 GNDA.n2820 GNDA.n2819 4.5005
R24463 GNDA.n2243 GNDA.n2242 4.5005
R24464 GNDA.n2765 GNDA.n2764 4.5005
R24465 GNDA.n2769 GNDA.n2766 4.5005
R24466 GNDA.n2770 GNDA.n2763 4.5005
R24467 GNDA.n2774 GNDA.n2773 4.5005
R24468 GNDA.n2775 GNDA.n2762 4.5005
R24469 GNDA.n2779 GNDA.n2776 4.5005
R24470 GNDA.n2780 GNDA.n2761 4.5005
R24471 GNDA.n2784 GNDA.n2783 4.5005
R24472 GNDA.n2785 GNDA.n2760 4.5005
R24473 GNDA.n2789 GNDA.n2786 4.5005
R24474 GNDA.n2790 GNDA.n2759 4.5005
R24475 GNDA.n2794 GNDA.n2793 4.5005
R24476 GNDA.n2795 GNDA.n2758 4.5005
R24477 GNDA.n2799 GNDA.n2796 4.5005
R24478 GNDA.n2800 GNDA.n2757 4.5005
R24479 GNDA.n2804 GNDA.n2803 4.5005
R24480 GNDA.n2805 GNDA.n2756 4.5005
R24481 GNDA.n2809 GNDA.n2806 4.5005
R24482 GNDA.n2810 GNDA.n2755 4.5005
R24483 GNDA.n2814 GNDA.n2813 4.5005
R24484 GNDA.n2686 GNDA.n2678 4.5005
R24485 GNDA.n2688 GNDA.n2687 4.5005
R24486 GNDA.n2691 GNDA.n2677 4.5005
R24487 GNDA.n2695 GNDA.n2694 4.5005
R24488 GNDA.n2696 GNDA.n2676 4.5005
R24489 GNDA.n2698 GNDA.n2697 4.5005
R24490 GNDA.n2701 GNDA.n2675 4.5005
R24491 GNDA.n2705 GNDA.n2704 4.5005
R24492 GNDA.n2706 GNDA.n2674 4.5005
R24493 GNDA.n2708 GNDA.n2707 4.5005
R24494 GNDA.n2711 GNDA.n2673 4.5005
R24495 GNDA.n2715 GNDA.n2714 4.5005
R24496 GNDA.n2716 GNDA.n2672 4.5005
R24497 GNDA.n2718 GNDA.n2717 4.5005
R24498 GNDA.n2721 GNDA.n2671 4.5005
R24499 GNDA.n2725 GNDA.n2724 4.5005
R24500 GNDA.n2726 GNDA.n2670 4.5005
R24501 GNDA.n2728 GNDA.n2727 4.5005
R24502 GNDA.n2731 GNDA.n2669 4.5005
R24503 GNDA.n2734 GNDA.n2733 4.5005
R24504 GNDA.n2735 GNDA.n2667 4.5005
R24505 GNDA.n2738 GNDA.n2737 4.5005
R24506 GNDA.n2684 GNDA.n2680 4.5005
R24507 GNDA.n2685 GNDA.n2240 4.5005
R24508 GNDA.n2685 GNDA.n2684 4.5005
R24509 GNDA.n2825 GNDA.n2824 4.5005
R24510 GNDA.n2824 GNDA.n2823 4.5005
R24511 GNDA.n2823 GNDA.n2241 4.5005
R24512 GNDA.n2912 GNDA.n2911 4.5005
R24513 GNDA.n2911 GNDA.n2910 4.5005
R24514 GNDA.n2910 GNDA.n2826 4.5005
R24515 GNDA.n2913 GNDA.n2231 4.5005
R24516 GNDA.n2914 GNDA.n2913 4.5005
R24517 GNDA.n2915 GNDA.n2914 4.5005
R24518 GNDA.n3059 GNDA.n3058 4.5005
R24519 GNDA.n3058 GNDA.n3057 4.5005
R24520 GNDA.n3057 GNDA.n2157 4.5005
R24521 GNDA.n3146 GNDA.n3145 4.5005
R24522 GNDA.n3145 GNDA.n3144 4.5005
R24523 GNDA.n3144 GNDA.n3060 4.5005
R24524 GNDA.n3147 GNDA.n2116 4.5005
R24525 GNDA.n3148 GNDA.n3147 4.5005
R24526 GNDA.n3149 GNDA.n3148 4.5005
R24527 GNDA.n3292 GNDA.n2118 4.5005
R24528 GNDA.n3295 GNDA.n2118 4.5005
R24529 GNDA.n3295 GNDA.n2117 4.5005
R24530 GNDA.n3306 GNDA.n2029 4.5005
R24531 GNDA.n3307 GNDA.n3306 4.5005
R24532 GNDA.n3308 GNDA.n3307 4.5005
R24533 GNDA.n2230 GNDA.n2187 4.5005
R24534 GNDA.n2229 GNDA.n2156 4.5005
R24535 GNDA.n2230 GNDA.n2229 4.5005
R24536 GNDA.n2219 GNDA.n2209 4.5005
R24537 GNDA.n2220 GNDA.n2219 4.5005
R24538 GNDA.n2221 GNDA.n2220 4.5005
R24539 GNDA.n5410 GNDA.n5409 4.5005
R24540 GNDA.n5430 GNDA.n5429 4.5005
R24541 GNDA.n5439 GNDA.n5417 4.5005
R24542 GNDA.n5438 GNDA.n655 4.5005
R24543 GNDA.n5439 GNDA.n5438 4.5005
R24544 GNDA.n5461 GNDA.n663 4.5005
R24545 GNDA.n5454 GNDA.n5453 4.5005
R24546 GNDA.n689 GNDA.n680 4.5005
R24547 GNDA.n692 GNDA.n691 4.5005
R24548 GNDA.n695 GNDA.n694 4.5005
R24549 GNDA.n2193 GNDA.n2190 4.5005
R24550 GNDA.n687 GNDA.n683 4.5005
R24551 GNDA.n688 GNDA.n682 4.5005
R24552 GNDA.n688 GNDA.n687 4.5005
R24553 GNDA.n5488 GNDA.n5487 4.5005
R24554 GNDA.n5491 GNDA.n657 4.5005
R24555 GNDA.n5492 GNDA.n5491 4.5005
R24556 GNDA.n5493 GNDA.n5492 4.5005
R24557 GNDA.n5496 GNDA.n652 4.5005
R24558 GNDA.n5497 GNDA.n5496 4.5005
R24559 GNDA.n5498 GNDA.n5497 4.5005
R24560 GNDA.n3615 GNDA.n649 4.5005
R24561 GNDA.n3612 GNDA.n649 4.5005
R24562 GNDA.n3613 GNDA.n3612 4.5005
R24563 GNDA.n5505 GNDA.n646 4.5005
R24564 GNDA.n5504 GNDA.n5503 4.5005
R24565 GNDA.n5505 GNDA.n5504 4.5005
R24566 GNDA.n5506 GNDA.n645 4.5005
R24567 GNDA.n599 GNDA.n598 4.5005
R24568 GNDA.n5527 GNDA.n5526 4.5005
R24569 GNDA.n5532 GNDA.n5531 4.5005
R24570 GNDA.n5538 GNDA.n5537 4.5005
R24571 GNDA.n5543 GNDA.n5542 4.5005
R24572 GNDA.n5546 GNDA.n5545 4.5005
R24573 GNDA.n5547 GNDA.n24 4.5005
R24574 GNDA.n5551 GNDA.n5548 4.5005
R24575 GNDA.n5552 GNDA.n23 4.5005
R24576 GNDA.n5556 GNDA.n5555 4.5005
R24577 GNDA.n5557 GNDA.n22 4.5005
R24578 GNDA.n5561 GNDA.n5558 4.5005
R24579 GNDA.n5562 GNDA.n21 4.5005
R24580 GNDA.n5566 GNDA.n5565 4.5005
R24581 GNDA.n5567 GNDA.n20 4.5005
R24582 GNDA.n5571 GNDA.n5568 4.5005
R24583 GNDA.n5572 GNDA.n19 4.5005
R24584 GNDA.n5576 GNDA.n5575 4.5005
R24585 GNDA.n5577 GNDA.n18 4.5005
R24586 GNDA.n5581 GNDA.n5578 4.5005
R24587 GNDA.n5582 GNDA.n17 4.5005
R24588 GNDA.n5586 GNDA.n5585 4.5005
R24589 GNDA.n5587 GNDA.n16 4.5005
R24590 GNDA.n5591 GNDA.n5588 4.5005
R24591 GNDA.n5592 GNDA.n15 4.5005
R24592 GNDA.n5596 GNDA.n5595 4.5005
R24593 GNDA.n577 GNDA.n576 4.5005
R24594 GNDA.n47 GNDA.n46 4.5005
R24595 GNDA.n522 GNDA.n521 4.5005
R24596 GNDA.n526 GNDA.n523 4.5005
R24597 GNDA.n527 GNDA.n520 4.5005
R24598 GNDA.n531 GNDA.n530 4.5005
R24599 GNDA.n532 GNDA.n519 4.5005
R24600 GNDA.n536 GNDA.n533 4.5005
R24601 GNDA.n537 GNDA.n518 4.5005
R24602 GNDA.n541 GNDA.n540 4.5005
R24603 GNDA.n542 GNDA.n517 4.5005
R24604 GNDA.n546 GNDA.n543 4.5005
R24605 GNDA.n547 GNDA.n516 4.5005
R24606 GNDA.n551 GNDA.n550 4.5005
R24607 GNDA.n552 GNDA.n515 4.5005
R24608 GNDA.n556 GNDA.n553 4.5005
R24609 GNDA.n557 GNDA.n514 4.5005
R24610 GNDA.n561 GNDA.n560 4.5005
R24611 GNDA.n562 GNDA.n513 4.5005
R24612 GNDA.n566 GNDA.n563 4.5005
R24613 GNDA.n567 GNDA.n512 4.5005
R24614 GNDA.n571 GNDA.n570 4.5005
R24615 GNDA.n353 GNDA.n352 4.5005
R24616 GNDA.n274 GNDA.n273 4.5005
R24617 GNDA.n296 GNDA.n275 4.5005
R24618 GNDA.n297 GNDA.n276 4.5005
R24619 GNDA.n298 GNDA.n277 4.5005
R24620 GNDA.n299 GNDA.n278 4.5005
R24621 GNDA.n300 GNDA.n279 4.5005
R24622 GNDA.n301 GNDA.n280 4.5005
R24623 GNDA.n302 GNDA.n281 4.5005
R24624 GNDA.n303 GNDA.n282 4.5005
R24625 GNDA.n304 GNDA.n283 4.5005
R24626 GNDA.n305 GNDA.n284 4.5005
R24627 GNDA.n306 GNDA.n285 4.5005
R24628 GNDA.n307 GNDA.n286 4.5005
R24629 GNDA.n308 GNDA.n287 4.5005
R24630 GNDA.n309 GNDA.n288 4.5005
R24631 GNDA.n310 GNDA.n289 4.5005
R24632 GNDA.n311 GNDA.n290 4.5005
R24633 GNDA.n312 GNDA.n291 4.5005
R24634 GNDA.n313 GNDA.n292 4.5005
R24635 GNDA.n314 GNDA.n293 4.5005
R24636 GNDA.n315 GNDA.n294 4.5005
R24637 GNDA.n267 GNDA.n266 4.5005
R24638 GNDA.n187 GNDA.n186 4.5005
R24639 GNDA.n212 GNDA.n211 4.5005
R24640 GNDA.n216 GNDA.n213 4.5005
R24641 GNDA.n217 GNDA.n210 4.5005
R24642 GNDA.n221 GNDA.n220 4.5005
R24643 GNDA.n222 GNDA.n209 4.5005
R24644 GNDA.n226 GNDA.n223 4.5005
R24645 GNDA.n227 GNDA.n208 4.5005
R24646 GNDA.n231 GNDA.n230 4.5005
R24647 GNDA.n232 GNDA.n207 4.5005
R24648 GNDA.n236 GNDA.n233 4.5005
R24649 GNDA.n237 GNDA.n206 4.5005
R24650 GNDA.n241 GNDA.n240 4.5005
R24651 GNDA.n242 GNDA.n205 4.5005
R24652 GNDA.n246 GNDA.n243 4.5005
R24653 GNDA.n247 GNDA.n204 4.5005
R24654 GNDA.n251 GNDA.n250 4.5005
R24655 GNDA.n252 GNDA.n203 4.5005
R24656 GNDA.n256 GNDA.n253 4.5005
R24657 GNDA.n257 GNDA.n202 4.5005
R24658 GNDA.n261 GNDA.n260 4.5005
R24659 GNDA.n180 GNDA.n179 4.5005
R24660 GNDA.n101 GNDA.n100 4.5005
R24661 GNDA.n123 GNDA.n102 4.5005
R24662 GNDA.n124 GNDA.n103 4.5005
R24663 GNDA.n125 GNDA.n104 4.5005
R24664 GNDA.n126 GNDA.n105 4.5005
R24665 GNDA.n127 GNDA.n106 4.5005
R24666 GNDA.n128 GNDA.n107 4.5005
R24667 GNDA.n129 GNDA.n108 4.5005
R24668 GNDA.n130 GNDA.n109 4.5005
R24669 GNDA.n131 GNDA.n110 4.5005
R24670 GNDA.n132 GNDA.n111 4.5005
R24671 GNDA.n133 GNDA.n112 4.5005
R24672 GNDA.n134 GNDA.n113 4.5005
R24673 GNDA.n135 GNDA.n114 4.5005
R24674 GNDA.n136 GNDA.n115 4.5005
R24675 GNDA.n137 GNDA.n116 4.5005
R24676 GNDA.n138 GNDA.n117 4.5005
R24677 GNDA.n139 GNDA.n118 4.5005
R24678 GNDA.n140 GNDA.n119 4.5005
R24679 GNDA.n141 GNDA.n120 4.5005
R24680 GNDA.n142 GNDA.n121 4.5005
R24681 GNDA.n452 GNDA.n451 4.5005
R24682 GNDA.n455 GNDA.n454 4.5005
R24683 GNDA.n456 GNDA.n96 4.5005
R24684 GNDA.n460 GNDA.n457 4.5005
R24685 GNDA.n461 GNDA.n95 4.5005
R24686 GNDA.n465 GNDA.n464 4.5005
R24687 GNDA.n466 GNDA.n94 4.5005
R24688 GNDA.n470 GNDA.n467 4.5005
R24689 GNDA.n471 GNDA.n93 4.5005
R24690 GNDA.n475 GNDA.n474 4.5005
R24691 GNDA.n476 GNDA.n92 4.5005
R24692 GNDA.n480 GNDA.n477 4.5005
R24693 GNDA.n481 GNDA.n91 4.5005
R24694 GNDA.n485 GNDA.n484 4.5005
R24695 GNDA.n486 GNDA.n90 4.5005
R24696 GNDA.n490 GNDA.n487 4.5005
R24697 GNDA.n491 GNDA.n89 4.5005
R24698 GNDA.n495 GNDA.n494 4.5005
R24699 GNDA.n496 GNDA.n88 4.5005
R24700 GNDA.n500 GNDA.n497 4.5005
R24701 GNDA.n501 GNDA.n87 4.5005
R24702 GNDA.n505 GNDA.n504 4.5005
R24703 GNDA.n443 GNDA.n442 4.5005
R24704 GNDA.n441 GNDA.n376 4.5005
R24705 GNDA.n440 GNDA.n439 4.5005
R24706 GNDA.n438 GNDA.n379 4.5005
R24707 GNDA.n437 GNDA.n436 4.5005
R24708 GNDA.n435 GNDA.n380 4.5005
R24709 GNDA.n434 GNDA.n433 4.5005
R24710 GNDA.n432 GNDA.n385 4.5005
R24711 GNDA.n431 GNDA.n430 4.5005
R24712 GNDA.n429 GNDA.n386 4.5005
R24713 GNDA.n428 GNDA.n427 4.5005
R24714 GNDA.n426 GNDA.n391 4.5005
R24715 GNDA.n425 GNDA.n424 4.5005
R24716 GNDA.n423 GNDA.n392 4.5005
R24717 GNDA.n422 GNDA.n421 4.5005
R24718 GNDA.n420 GNDA.n397 4.5005
R24719 GNDA.n419 GNDA.n418 4.5005
R24720 GNDA.n417 GNDA.n398 4.5005
R24721 GNDA.n416 GNDA.n415 4.5005
R24722 GNDA.n414 GNDA.n403 4.5005
R24723 GNDA.n413 GNDA.n412 4.5005
R24724 GNDA.n411 GNDA.n404 4.5005
R24725 GNDA.n374 GNDA.n45 4.5005
R24726 GNDA.n445 GNDA.n444 4.5005
R24727 GNDA.n444 GNDA.n45 4.5005
R24728 GNDA.n446 GNDA.n368 4.5005
R24729 GNDA.n447 GNDA.n446 4.5005
R24730 GNDA.n448 GNDA.n447 4.5005
R24731 GNDA.n364 GNDA.n99 4.5005
R24732 GNDA.n367 GNDA.n99 4.5005
R24733 GNDA.n367 GNDA.n98 4.5005
R24734 GNDA.n360 GNDA.n185 4.5005
R24735 GNDA.n363 GNDA.n185 4.5005
R24736 GNDA.n363 GNDA.n184 4.5005
R24737 GNDA.n272 GNDA.n25 4.5005
R24738 GNDA.n359 GNDA.n272 4.5005
R24739 GNDA.n359 GNDA.n271 4.5005
R24740 GNDA.n603 GNDA.n600 4.5005
R24741 GNDA.n604 GNDA.n603 4.5005
R24742 GNDA.n605 GNDA.n604 4.5005
R24743 GNDA.n610 GNDA.n579 4.5005
R24744 GNDA.n612 GNDA.n611 4.5005
R24745 GNDA.n611 GNDA.n610 4.5005
R24746 GNDA.n4904 GNDA.n4903 4.5005
R24747 GNDA.n4907 GNDA.n948 4.5005
R24748 GNDA.n980 GNDA.n976 4.5005
R24749 GNDA.n984 GNDA.n983 4.5005
R24750 GNDA.n985 GNDA.n975 4.5005
R24751 GNDA.n989 GNDA.n986 4.5005
R24752 GNDA.n990 GNDA.n974 4.5005
R24753 GNDA.n994 GNDA.n993 4.5005
R24754 GNDA.n995 GNDA.n973 4.5005
R24755 GNDA.n999 GNDA.n996 4.5005
R24756 GNDA.n1000 GNDA.n972 4.5005
R24757 GNDA.n1004 GNDA.n1003 4.5005
R24758 GNDA.n1005 GNDA.n971 4.5005
R24759 GNDA.n1009 GNDA.n1006 4.5005
R24760 GNDA.n1010 GNDA.n970 4.5005
R24761 GNDA.n1014 GNDA.n1013 4.5005
R24762 GNDA.n1015 GNDA.n969 4.5005
R24763 GNDA.n1019 GNDA.n1016 4.5005
R24764 GNDA.n1020 GNDA.n968 4.5005
R24765 GNDA.n1024 GNDA.n1023 4.5005
R24766 GNDA.n1025 GNDA.n967 4.5005
R24767 GNDA.n1027 GNDA.n1026 4.5005
R24768 GNDA.n952 GNDA.n951 4.5005
R24769 GNDA.n4900 GNDA.n4899 4.5005
R24770 GNDA.n4919 GNDA.n4918 4.49344
R24771 GNDA.n1597 GNDA.n1523 4.26717
R24772 GNDA.n1603 GNDA.n1523 4.26717
R24773 GNDA.n1603 GNDA.n1521 4.26717
R24774 GNDA.n1609 GNDA.n1521 4.26717
R24775 GNDA.n1609 GNDA.n1519 4.26717
R24776 GNDA.n1615 GNDA.n1519 4.26717
R24777 GNDA.n1615 GNDA.n1517 4.26717
R24778 GNDA.n1621 GNDA.n1517 4.26717
R24779 GNDA.n1621 GNDA.n1515 4.26717
R24780 GNDA.n1628 GNDA.n1515 4.26717
R24781 GNDA.n1628 GNDA.n1513 4.26717
R24782 GNDA.n4617 GNDA.n4616 4.26717
R24783 GNDA.n4616 GNDA.n4615 4.26717
R24784 GNDA.n4615 GNDA.n4613 4.26717
R24785 GNDA.n4613 GNDA.n4610 4.26717
R24786 GNDA.n4610 GNDA.n4609 4.26717
R24787 GNDA.n4609 GNDA.n4606 4.26717
R24788 GNDA.n4606 GNDA.n4605 4.26717
R24789 GNDA.n4605 GNDA.n4602 4.26717
R24790 GNDA.n4602 GNDA.n4601 4.26717
R24791 GNDA.n4601 GNDA.n4598 4.26717
R24792 GNDA.n4598 GNDA.n4597 4.26717
R24793 GNDA.n5210 GNDA.n848 4.26717
R24794 GNDA.n5205 GNDA.n848 4.26717
R24795 GNDA.n5205 GNDA.n5204 4.26717
R24796 GNDA.n5204 GNDA.n5203 4.26717
R24797 GNDA.n5203 GNDA.n857 4.26717
R24798 GNDA.n5197 GNDA.n857 4.26717
R24799 GNDA.n5197 GNDA.n5196 4.26717
R24800 GNDA.n5196 GNDA.n5195 4.26717
R24801 GNDA.n5195 GNDA.n865 4.26717
R24802 GNDA.n5189 GNDA.n865 4.26717
R24803 GNDA.n5189 GNDA.n5188 4.26717
R24804 GNDA.n4867 GNDA.n1126 4.26717
R24805 GNDA.n1909 GNDA.n1126 4.26717
R24806 GNDA.n1910 GNDA.n1909 4.26717
R24807 GNDA.n1913 GNDA.n1910 4.26717
R24808 GNDA.n1913 GNDA.n1902 4.26717
R24809 GNDA.n1921 GNDA.n1902 4.26717
R24810 GNDA.n1922 GNDA.n1921 4.26717
R24811 GNDA.n1925 GNDA.n1922 4.26717
R24812 GNDA.n1925 GNDA.n1900 4.26717
R24813 GNDA.n1933 GNDA.n1900 4.26717
R24814 GNDA.n1934 GNDA.n1933 4.26717
R24815 GNDA.n1898 GNDA.n1685 4.26717
R24816 GNDA.n1893 GNDA.n1685 4.26717
R24817 GNDA.n1893 GNDA.n1892 4.26717
R24818 GNDA.n1892 GNDA.n1874 4.26717
R24819 GNDA.n1887 GNDA.n1874 4.26717
R24820 GNDA.n1887 GNDA.n1886 4.26717
R24821 GNDA.n1886 GNDA.n1885 4.26717
R24822 GNDA.n1885 GNDA.n1880 4.26717
R24823 GNDA.n1880 GNDA.n1382 4.26717
R24824 GNDA.n4625 GNDA.n1382 4.26717
R24825 GNDA.n4625 GNDA.n1379 4.26717
R24826 GNDA.n1376 GNDA.n1332 4.26717
R24827 GNDA.n1371 GNDA.n1332 4.26717
R24828 GNDA.n1371 GNDA.n1370 4.26717
R24829 GNDA.n1370 GNDA.n1369 4.26717
R24830 GNDA.n1369 GNDA.n1341 4.26717
R24831 GNDA.n1363 GNDA.n1341 4.26717
R24832 GNDA.n1363 GNDA.n1362 4.26717
R24833 GNDA.n1362 GNDA.n1361 4.26717
R24834 GNDA.n1361 GNDA.n1349 4.26717
R24835 GNDA.n1355 GNDA.n1349 4.26717
R24836 GNDA.n1355 GNDA.n816 4.26717
R24837 GNDA.n1597 GNDA.n1525 3.93531
R24838 GNDA.n4617 GNDA.n4548 3.93531
R24839 GNDA.n5211 GNDA.n5210 3.93531
R24840 GNDA.n4868 GNDA.n4867 3.93531
R24841 GNDA.n1899 GNDA.n1898 3.93531
R24842 GNDA.n1377 GNDA.n1376 3.93531
R24843 GNDA.n3305 GNDA.n3304 3.84081
R24844 GNDA.n4183 GNDA.n4182 3.84081
R24845 GNDA.n4277 GNDA.n4275 3.84081
R24846 GNDA.n3298 GNDA.n3296 3.84045
R24847 GNDA.n5294 GNDA.n809 3.7893
R24848 GNDA.n5293 GNDA.n810 3.7893
R24849 GNDA.n5281 GNDA.n5280 3.7893
R24850 GNDA.n5287 GNDA.n5286 3.7893
R24851 GNDA.n5283 GNDA.n5282 3.7893
R24852 GNDA.n786 GNDA.n779 3.7893
R24853 GNDA.n791 GNDA.n789 3.7893
R24854 GNDA.n790 GNDA.n756 3.7893
R24855 GNDA.n5365 GNDA.n739 3.7893
R24856 GNDA.n5364 GNDA.n740 3.7893
R24857 GNDA.n5352 GNDA.n5351 3.7893
R24858 GNDA.n5358 GNDA.n5357 3.7893
R24859 GNDA.n5354 GNDA.n5353 3.7893
R24860 GNDA.n5073 GNDA.n718 3.7893
R24861 GNDA.n5078 GNDA.n5076 3.7893
R24862 GNDA.n5080 GNDA.n5079 3.7893
R24863 GNDA.n4719 GNDA.n4718 3.7893
R24864 GNDA.n4715 GNDA.n1236 3.7893
R24865 GNDA.n4714 GNDA.n1239 3.7893
R24866 GNDA.n4711 GNDA.n4710 3.7893
R24867 GNDA.n4636 GNDA.n1240 3.7893
R24868 GNDA.n4645 GNDA.n4644 3.7893
R24869 GNDA.n4648 GNDA.n4635 3.7893
R24870 GNDA.n4653 GNDA.n4649 3.7893
R24871 GNDA.n1809 GNDA.n1784 3.7893
R24872 GNDA.n1808 GNDA.n1805 3.7893
R24873 GNDA.n1804 GNDA.n1785 3.7893
R24874 GNDA.n1801 GNDA.n1800 3.7893
R24875 GNDA.n1797 GNDA.n1786 3.7893
R24876 GNDA.n1790 GNDA.n1787 3.7893
R24877 GNDA.n1815 GNDA.n1709 3.7893
R24878 GNDA.n1816 GNDA.n1708 3.7893
R24879 GNDA.n4816 GNDA.n1193 3.7893
R24880 GNDA.n4813 GNDA.n4812 3.7893
R24881 GNDA.n4728 GNDA.n1195 3.7893
R24882 GNDA.n4746 GNDA.n4745 3.7893
R24883 GNDA.n4743 GNDA.n4742 3.7893
R24884 GNDA.n4738 GNDA.n4731 3.7893
R24885 GNDA.n4735 GNDA.n4734 3.7893
R24886 GNDA.n4753 GNDA.n1215 3.7893
R24887 GNDA.n4542 GNDA.n1633 3.7893
R24888 GNDA.n4539 GNDA.n4538 3.7893
R24889 GNDA.n4454 GNDA.n1634 3.7893
R24890 GNDA.n4459 GNDA.n4457 3.7893
R24891 GNDA.n4464 GNDA.n4460 3.7893
R24892 GNDA.n4471 GNDA.n4470 3.7893
R24893 GNDA.n4474 GNDA.n4453 3.7893
R24894 GNDA.n4479 GNDA.n4475 3.7893
R24895 GNDA.n1498 GNDA.n1474 3.7893
R24896 GNDA.n1497 GNDA.n1495 3.7893
R24897 GNDA.n1494 GNDA.n1475 3.7893
R24898 GNDA.n1491 GNDA.n1490 3.7893
R24899 GNDA.n1487 GNDA.n1476 3.7893
R24900 GNDA.n1480 GNDA.n1477 3.7893
R24901 GNDA.n1504 GNDA.n1401 3.7893
R24902 GNDA.n1505 GNDA.n1400 3.7893
R24903 GNDA.n5007 GNDA.n5005 3.7893
R24904 GNDA.n5006 GNDA.n4929 3.7893
R24905 GNDA.n5013 GNDA.n5012 3.7893
R24906 GNDA.n4936 GNDA.n4930 3.7893
R24907 GNDA.n4935 GNDA.n4933 3.7893
R24908 GNDA.n5171 GNDA.n892 3.7893
R24909 GNDA.n891 GNDA.n887 3.7893
R24910 GNDA.n5180 GNDA.n5179 3.7893
R24911 GNDA.n4443 GNDA.n1937 3.7893
R24912 GNDA.n4440 GNDA.n4439 3.7893
R24913 GNDA.n4355 GNDA.n1938 3.7893
R24914 GNDA.n4360 GNDA.n4358 3.7893
R24915 GNDA.n4365 GNDA.n4361 3.7893
R24916 GNDA.n4372 GNDA.n4371 3.7893
R24917 GNDA.n4375 GNDA.n4354 3.7893
R24918 GNDA.n4380 GNDA.n4376 3.7893
R24919 GNDA_2 GNDA.n5300 3.7381
R24920 GNDA_2 GNDA.n5371 3.7381
R24921 GNDA.n4641 GNDA_2 3.7381
R24922 GNDA_2 GNDA.n1793 3.7381
R24923 GNDA.n4739 GNDA_2 3.7381
R24924 GNDA.n4467 GNDA_2 3.7381
R24925 GNDA_2 GNDA.n1483 3.7381
R24926 GNDA.n5172 GNDA_2 3.7381
R24927 GNDA.n4368 GNDA_2 3.7381
R24928 GNDA.n5317 GNDA.n769 3.70778
R24929 GNDA.n5311 GNDA.n5310 3.70778
R24930 GNDA.n5161 GNDA.n5156 3.70778
R24931 GNDA.n2736 GNDA.n2654 3.50398
R24932 GNDA.n409 GNDA.n60 3.50398
R24933 GNDA.n977 GNDA.n955 3.47871
R24934 GNDA.n2076 GNDA.n2075 3.47821
R24935 GNDA.n4113 GNDA.n4112 3.47821
R24936 GNDA.n4093 GNDA.n4092 3.47821
R24937 GNDA.n4012 GNDA.n4011 3.47821
R24938 GNDA.n3931 GNDA.n3930 3.47821
R24939 GNDA.n4235 GNDA.n4234 3.47821
R24940 GNDA.n3850 GNDA.n3849 3.47821
R24941 GNDA.n3769 GNDA.n3768 3.47821
R24942 GNDA.n3560 GNDA.n3559 3.47821
R24943 GNDA.n4239 GNDA.n4238 3.47821
R24944 GNDA.n1066 GNDA.n1030 3.47821
R24945 GNDA.n3456 GNDA.n3455 3.47821
R24946 GNDA.n3367 GNDA.n3366 3.47821
R24947 GNDA.n3284 GNDA.n3283 3.47821
R24948 GNDA.n3208 GNDA.n3207 3.47821
R24949 GNDA.n3105 GNDA.n3104 3.47821
R24950 GNDA.n3050 GNDA.n3049 3.47821
R24951 GNDA.n2974 GNDA.n2973 3.47821
R24952 GNDA.n2871 GNDA.n2870 3.47821
R24953 GNDA.n2816 GNDA.n2815 3.47821
R24954 GNDA.n5598 GNDA.n5597 3.47821
R24955 GNDA.n573 GNDA.n572 3.47821
R24956 GNDA.n317 GNDA.n316 3.47821
R24957 GNDA.n263 GNDA.n262 3.47821
R24958 GNDA.n144 GNDA.n143 3.47821
R24959 GNDA.n507 GNDA.n506 3.47821
R24960 GNDA.n2678 GNDA.n2655 3.43627
R24961 GNDA.n442 GNDA.n61 3.43627
R24962 GNDA.n2077 GNDA.n2054 3.4105
R24963 GNDA.n2079 GNDA.n2053 3.4105
R24964 GNDA.n2080 GNDA.n2052 3.4105
R24965 GNDA.n2082 GNDA.n2051 3.4105
R24966 GNDA.n2083 GNDA.n2050 3.4105
R24967 GNDA.n2085 GNDA.n2049 3.4105
R24968 GNDA.n2086 GNDA.n2048 3.4105
R24969 GNDA.n2088 GNDA.n2047 3.4105
R24970 GNDA.n2089 GNDA.n2046 3.4105
R24971 GNDA.n2091 GNDA.n2045 3.4105
R24972 GNDA.n2092 GNDA.n2044 3.4105
R24973 GNDA.n2094 GNDA.n2043 3.4105
R24974 GNDA.n2095 GNDA.n2042 3.4105
R24975 GNDA.n2097 GNDA.n2041 3.4105
R24976 GNDA.n2098 GNDA.n2040 3.4105
R24977 GNDA.n2100 GNDA.n2039 3.4105
R24978 GNDA.n2101 GNDA.n2038 3.4105
R24979 GNDA.n2103 GNDA.n2037 3.4105
R24980 GNDA.n2104 GNDA.n2036 3.4105
R24981 GNDA.n2106 GNDA.n2035 3.4105
R24982 GNDA.n2107 GNDA.n2034 3.4105
R24983 GNDA.n2109 GNDA.n2033 3.4105
R24984 GNDA.n2111 GNDA.n2110 3.4105
R24985 GNDA.n4114 GNDA.n3689 3.4105
R24986 GNDA.n4115 GNDA.n3688 3.4105
R24987 GNDA.n4116 GNDA.n3687 3.4105
R24988 GNDA.n4108 GNDA.n3685 3.4105
R24989 GNDA.n4120 GNDA.n3684 3.4105
R24990 GNDA.n4121 GNDA.n3683 3.4105
R24991 GNDA.n4122 GNDA.n3682 3.4105
R24992 GNDA.n4105 GNDA.n3680 3.4105
R24993 GNDA.n4126 GNDA.n3679 3.4105
R24994 GNDA.n4127 GNDA.n3678 3.4105
R24995 GNDA.n4128 GNDA.n3677 3.4105
R24996 GNDA.n4102 GNDA.n3675 3.4105
R24997 GNDA.n4132 GNDA.n3674 3.4105
R24998 GNDA.n4133 GNDA.n3673 3.4105
R24999 GNDA.n4134 GNDA.n3672 3.4105
R25000 GNDA.n4099 GNDA.n3670 3.4105
R25001 GNDA.n4138 GNDA.n3669 3.4105
R25002 GNDA.n4139 GNDA.n3668 3.4105
R25003 GNDA.n4140 GNDA.n3667 3.4105
R25004 GNDA.n4096 GNDA.n3665 3.4105
R25005 GNDA.n4144 GNDA.n3664 3.4105
R25006 GNDA.n4145 GNDA.n3663 3.4105
R25007 GNDA.n4146 GNDA.n3662 3.4105
R25008 GNDA.n4027 GNDA.n4026 3.4105
R25009 GNDA.n4090 GNDA.n4089 3.4105
R25010 GNDA.n4088 GNDA.n4087 3.4105
R25011 GNDA.n4086 GNDA.n4031 3.4105
R25012 GNDA.n4030 GNDA.n4029 3.4105
R25013 GNDA.n4082 GNDA.n4081 3.4105
R25014 GNDA.n4080 GNDA.n4079 3.4105
R25015 GNDA.n4078 GNDA.n4035 3.4105
R25016 GNDA.n4034 GNDA.n4033 3.4105
R25017 GNDA.n4074 GNDA.n4073 3.4105
R25018 GNDA.n4072 GNDA.n4071 3.4105
R25019 GNDA.n4070 GNDA.n4039 3.4105
R25020 GNDA.n4038 GNDA.n4037 3.4105
R25021 GNDA.n4066 GNDA.n4065 3.4105
R25022 GNDA.n4064 GNDA.n4063 3.4105
R25023 GNDA.n4062 GNDA.n4043 3.4105
R25024 GNDA.n4042 GNDA.n4041 3.4105
R25025 GNDA.n4058 GNDA.n4057 3.4105
R25026 GNDA.n4056 GNDA.n4055 3.4105
R25027 GNDA.n4054 GNDA.n4047 3.4105
R25028 GNDA.n4046 GNDA.n4045 3.4105
R25029 GNDA.n4050 GNDA.n4049 3.4105
R25030 GNDA.n4048 GNDA.n4014 3.4105
R25031 GNDA.n3946 GNDA.n3945 3.4105
R25032 GNDA.n4009 GNDA.n4008 3.4105
R25033 GNDA.n4007 GNDA.n4006 3.4105
R25034 GNDA.n4005 GNDA.n3950 3.4105
R25035 GNDA.n3949 GNDA.n3948 3.4105
R25036 GNDA.n4001 GNDA.n4000 3.4105
R25037 GNDA.n3999 GNDA.n3998 3.4105
R25038 GNDA.n3997 GNDA.n3954 3.4105
R25039 GNDA.n3953 GNDA.n3952 3.4105
R25040 GNDA.n3993 GNDA.n3992 3.4105
R25041 GNDA.n3991 GNDA.n3990 3.4105
R25042 GNDA.n3989 GNDA.n3958 3.4105
R25043 GNDA.n3957 GNDA.n3956 3.4105
R25044 GNDA.n3985 GNDA.n3984 3.4105
R25045 GNDA.n3983 GNDA.n3982 3.4105
R25046 GNDA.n3981 GNDA.n3962 3.4105
R25047 GNDA.n3961 GNDA.n3960 3.4105
R25048 GNDA.n3977 GNDA.n3976 3.4105
R25049 GNDA.n3975 GNDA.n3974 3.4105
R25050 GNDA.n3973 GNDA.n3966 3.4105
R25051 GNDA.n3965 GNDA.n3964 3.4105
R25052 GNDA.n3969 GNDA.n3968 3.4105
R25053 GNDA.n3967 GNDA.n3933 3.4105
R25054 GNDA.n3865 GNDA.n3864 3.4105
R25055 GNDA.n3928 GNDA.n3927 3.4105
R25056 GNDA.n3926 GNDA.n3925 3.4105
R25057 GNDA.n3924 GNDA.n3869 3.4105
R25058 GNDA.n3868 GNDA.n3867 3.4105
R25059 GNDA.n3920 GNDA.n3919 3.4105
R25060 GNDA.n3918 GNDA.n3917 3.4105
R25061 GNDA.n3916 GNDA.n3873 3.4105
R25062 GNDA.n3872 GNDA.n3871 3.4105
R25063 GNDA.n3912 GNDA.n3911 3.4105
R25064 GNDA.n3910 GNDA.n3909 3.4105
R25065 GNDA.n3908 GNDA.n3877 3.4105
R25066 GNDA.n3876 GNDA.n3875 3.4105
R25067 GNDA.n3904 GNDA.n3903 3.4105
R25068 GNDA.n3902 GNDA.n3901 3.4105
R25069 GNDA.n3900 GNDA.n3881 3.4105
R25070 GNDA.n3880 GNDA.n3879 3.4105
R25071 GNDA.n3896 GNDA.n3895 3.4105
R25072 GNDA.n3894 GNDA.n3893 3.4105
R25073 GNDA.n3892 GNDA.n3885 3.4105
R25074 GNDA.n3884 GNDA.n3883 3.4105
R25075 GNDA.n3888 GNDA.n3887 3.4105
R25076 GNDA.n3886 GNDA.n3852 3.4105
R25077 GNDA.n3488 GNDA.n3487 3.4105
R25078 GNDA.n4232 GNDA.n4231 3.4105
R25079 GNDA.n4230 GNDA.n4229 3.4105
R25080 GNDA.n4228 GNDA.n3492 3.4105
R25081 GNDA.n3491 GNDA.n3490 3.4105
R25082 GNDA.n4224 GNDA.n4223 3.4105
R25083 GNDA.n4222 GNDA.n4221 3.4105
R25084 GNDA.n4220 GNDA.n3496 3.4105
R25085 GNDA.n3495 GNDA.n3494 3.4105
R25086 GNDA.n4216 GNDA.n4215 3.4105
R25087 GNDA.n4214 GNDA.n4213 3.4105
R25088 GNDA.n4212 GNDA.n3500 3.4105
R25089 GNDA.n3499 GNDA.n3498 3.4105
R25090 GNDA.n4208 GNDA.n4207 3.4105
R25091 GNDA.n4206 GNDA.n4205 3.4105
R25092 GNDA.n4204 GNDA.n3504 3.4105
R25093 GNDA.n3503 GNDA.n3502 3.4105
R25094 GNDA.n4200 GNDA.n4199 3.4105
R25095 GNDA.n4198 GNDA.n4197 3.4105
R25096 GNDA.n4196 GNDA.n3508 3.4105
R25097 GNDA.n3507 GNDA.n3506 3.4105
R25098 GNDA.n4192 GNDA.n4191 3.4105
R25099 GNDA.n4190 GNDA.n3474 3.4105
R25100 GNDA.n3784 GNDA.n3783 3.4105
R25101 GNDA.n3847 GNDA.n3846 3.4105
R25102 GNDA.n3845 GNDA.n3844 3.4105
R25103 GNDA.n3843 GNDA.n3788 3.4105
R25104 GNDA.n3787 GNDA.n3786 3.4105
R25105 GNDA.n3839 GNDA.n3838 3.4105
R25106 GNDA.n3837 GNDA.n3836 3.4105
R25107 GNDA.n3835 GNDA.n3792 3.4105
R25108 GNDA.n3791 GNDA.n3790 3.4105
R25109 GNDA.n3831 GNDA.n3830 3.4105
R25110 GNDA.n3829 GNDA.n3828 3.4105
R25111 GNDA.n3827 GNDA.n3796 3.4105
R25112 GNDA.n3795 GNDA.n3794 3.4105
R25113 GNDA.n3823 GNDA.n3822 3.4105
R25114 GNDA.n3821 GNDA.n3820 3.4105
R25115 GNDA.n3819 GNDA.n3800 3.4105
R25116 GNDA.n3799 GNDA.n3798 3.4105
R25117 GNDA.n3815 GNDA.n3814 3.4105
R25118 GNDA.n3813 GNDA.n3812 3.4105
R25119 GNDA.n3811 GNDA.n3804 3.4105
R25120 GNDA.n3803 GNDA.n3802 3.4105
R25121 GNDA.n3807 GNDA.n3806 3.4105
R25122 GNDA.n3805 GNDA.n3771 3.4105
R25123 GNDA.n3703 GNDA.n3702 3.4105
R25124 GNDA.n3766 GNDA.n3765 3.4105
R25125 GNDA.n3764 GNDA.n3763 3.4105
R25126 GNDA.n3762 GNDA.n3707 3.4105
R25127 GNDA.n3706 GNDA.n3705 3.4105
R25128 GNDA.n3758 GNDA.n3757 3.4105
R25129 GNDA.n3756 GNDA.n3755 3.4105
R25130 GNDA.n3754 GNDA.n3711 3.4105
R25131 GNDA.n3710 GNDA.n3709 3.4105
R25132 GNDA.n3750 GNDA.n3749 3.4105
R25133 GNDA.n3748 GNDA.n3747 3.4105
R25134 GNDA.n3746 GNDA.n3715 3.4105
R25135 GNDA.n3714 GNDA.n3713 3.4105
R25136 GNDA.n3742 GNDA.n3741 3.4105
R25137 GNDA.n3740 GNDA.n3739 3.4105
R25138 GNDA.n3738 GNDA.n3719 3.4105
R25139 GNDA.n3718 GNDA.n3717 3.4105
R25140 GNDA.n3734 GNDA.n3733 3.4105
R25141 GNDA.n3732 GNDA.n3731 3.4105
R25142 GNDA.n3730 GNDA.n3723 3.4105
R25143 GNDA.n3722 GNDA.n3721 3.4105
R25144 GNDA.n3726 GNDA.n3725 3.4105
R25145 GNDA.n3724 GNDA.n3690 3.4105
R25146 GNDA.n3561 GNDA.n3558 3.4105
R25147 GNDA.n3562 GNDA.n3556 3.4105
R25148 GNDA.n3563 GNDA.n3555 3.4105
R25149 GNDA.n3553 GNDA.n3551 3.4105
R25150 GNDA.n3567 GNDA.n3550 3.4105
R25151 GNDA.n3568 GNDA.n3548 3.4105
R25152 GNDA.n3569 GNDA.n3547 3.4105
R25153 GNDA.n3545 GNDA.n3543 3.4105
R25154 GNDA.n3573 GNDA.n3542 3.4105
R25155 GNDA.n3574 GNDA.n3540 3.4105
R25156 GNDA.n3575 GNDA.n3539 3.4105
R25157 GNDA.n3537 GNDA.n3535 3.4105
R25158 GNDA.n3579 GNDA.n3534 3.4105
R25159 GNDA.n3580 GNDA.n3532 3.4105
R25160 GNDA.n3581 GNDA.n3531 3.4105
R25161 GNDA.n3529 GNDA.n3527 3.4105
R25162 GNDA.n3585 GNDA.n3526 3.4105
R25163 GNDA.n3586 GNDA.n3524 3.4105
R25164 GNDA.n3587 GNDA.n3523 3.4105
R25165 GNDA.n3521 GNDA.n3519 3.4105
R25166 GNDA.n3591 GNDA.n3518 3.4105
R25167 GNDA.n3592 GNDA.n3516 3.4105
R25168 GNDA.n3593 GNDA.n3515 3.4105
R25169 GNDA.n4240 GNDA.n2002 3.4105
R25170 GNDA.n4241 GNDA.n2001 3.4105
R25171 GNDA.n4242 GNDA.n2000 3.4105
R25172 GNDA.n3471 GNDA.n1998 3.4105
R25173 GNDA.n4246 GNDA.n1997 3.4105
R25174 GNDA.n4247 GNDA.n1996 3.4105
R25175 GNDA.n4248 GNDA.n1995 3.4105
R25176 GNDA.n3468 GNDA.n1993 3.4105
R25177 GNDA.n4252 GNDA.n1992 3.4105
R25178 GNDA.n4253 GNDA.n1991 3.4105
R25179 GNDA.n4254 GNDA.n1990 3.4105
R25180 GNDA.n3465 GNDA.n1988 3.4105
R25181 GNDA.n4258 GNDA.n1987 3.4105
R25182 GNDA.n4259 GNDA.n1986 3.4105
R25183 GNDA.n4260 GNDA.n1985 3.4105
R25184 GNDA.n3462 GNDA.n1983 3.4105
R25185 GNDA.n4264 GNDA.n1982 3.4105
R25186 GNDA.n4265 GNDA.n1981 3.4105
R25187 GNDA.n4266 GNDA.n1980 3.4105
R25188 GNDA.n3459 GNDA.n1978 3.4105
R25189 GNDA.n4270 GNDA.n1977 3.4105
R25190 GNDA.n4271 GNDA.n1976 3.4105
R25191 GNDA.n4272 GNDA.n1975 3.4105
R25192 GNDA.n1043 GNDA.n1042 3.4105
R25193 GNDA.n1105 GNDA.n1104 3.4105
R25194 GNDA.n1103 GNDA.n1102 3.4105
R25195 GNDA.n1101 GNDA.n1047 3.4105
R25196 GNDA.n1046 GNDA.n1045 3.4105
R25197 GNDA.n1097 GNDA.n1096 3.4105
R25198 GNDA.n1095 GNDA.n1094 3.4105
R25199 GNDA.n1093 GNDA.n1051 3.4105
R25200 GNDA.n1050 GNDA.n1049 3.4105
R25201 GNDA.n1089 GNDA.n1088 3.4105
R25202 GNDA.n1087 GNDA.n1086 3.4105
R25203 GNDA.n1085 GNDA.n1055 3.4105
R25204 GNDA.n1054 GNDA.n1053 3.4105
R25205 GNDA.n1081 GNDA.n1080 3.4105
R25206 GNDA.n1079 GNDA.n1078 3.4105
R25207 GNDA.n1077 GNDA.n1059 3.4105
R25208 GNDA.n1058 GNDA.n1057 3.4105
R25209 GNDA.n1073 GNDA.n1072 3.4105
R25210 GNDA.n1071 GNDA.n1070 3.4105
R25211 GNDA.n1069 GNDA.n1063 3.4105
R25212 GNDA.n1062 GNDA.n1061 3.4105
R25213 GNDA.n1065 GNDA.n1064 3.4105
R25214 GNDA.n4895 GNDA.n4894 3.4105
R25215 GNDA.n3382 GNDA.n3381 3.4105
R25216 GNDA.n3453 GNDA.n3452 3.4105
R25217 GNDA.n3451 GNDA.n3450 3.4105
R25218 GNDA.n3449 GNDA.n3448 3.4105
R25219 GNDA.n3447 GNDA.n3384 3.4105
R25220 GNDA.n3443 GNDA.n3442 3.4105
R25221 GNDA.n3441 GNDA.n3440 3.4105
R25222 GNDA.n3439 GNDA.n3438 3.4105
R25223 GNDA.n3437 GNDA.n3386 3.4105
R25224 GNDA.n3433 GNDA.n3432 3.4105
R25225 GNDA.n3431 GNDA.n3430 3.4105
R25226 GNDA.n3429 GNDA.n3428 3.4105
R25227 GNDA.n3427 GNDA.n3388 3.4105
R25228 GNDA.n3423 GNDA.n3422 3.4105
R25229 GNDA.n3421 GNDA.n3420 3.4105
R25230 GNDA.n3419 GNDA.n3418 3.4105
R25231 GNDA.n3417 GNDA.n3390 3.4105
R25232 GNDA.n3413 GNDA.n3412 3.4105
R25233 GNDA.n3411 GNDA.n3410 3.4105
R25234 GNDA.n3409 GNDA.n3408 3.4105
R25235 GNDA.n3407 GNDA.n3392 3.4105
R25236 GNDA.n3403 GNDA.n3402 3.4105
R25237 GNDA.n3401 GNDA.n3369 3.4105
R25238 GNDA.n2017 GNDA.n2016 3.4105
R25239 GNDA.n3364 GNDA.n3363 3.4105
R25240 GNDA.n3362 GNDA.n3361 3.4105
R25241 GNDA.n3360 GNDA.n3359 3.4105
R25242 GNDA.n3358 GNDA.n2019 3.4105
R25243 GNDA.n3354 GNDA.n3353 3.4105
R25244 GNDA.n3352 GNDA.n3351 3.4105
R25245 GNDA.n3350 GNDA.n3349 3.4105
R25246 GNDA.n3348 GNDA.n2021 3.4105
R25247 GNDA.n3344 GNDA.n3343 3.4105
R25248 GNDA.n3342 GNDA.n3341 3.4105
R25249 GNDA.n3340 GNDA.n3339 3.4105
R25250 GNDA.n3338 GNDA.n2023 3.4105
R25251 GNDA.n3334 GNDA.n3333 3.4105
R25252 GNDA.n3332 GNDA.n3331 3.4105
R25253 GNDA.n3330 GNDA.n3329 3.4105
R25254 GNDA.n3328 GNDA.n2025 3.4105
R25255 GNDA.n3324 GNDA.n3323 3.4105
R25256 GNDA.n3322 GNDA.n3321 3.4105
R25257 GNDA.n3320 GNDA.n3319 3.4105
R25258 GNDA.n3318 GNDA.n2027 3.4105
R25259 GNDA.n3314 GNDA.n3313 3.4105
R25260 GNDA.n3312 GNDA.n2004 3.4105
R25261 GNDA.n3222 GNDA.n3221 3.4105
R25262 GNDA.n3281 GNDA.n3280 3.4105
R25263 GNDA.n3279 GNDA.n3278 3.4105
R25264 GNDA.n3277 GNDA.n3276 3.4105
R25265 GNDA.n3275 GNDA.n3224 3.4105
R25266 GNDA.n3271 GNDA.n3270 3.4105
R25267 GNDA.n3269 GNDA.n3268 3.4105
R25268 GNDA.n3267 GNDA.n3266 3.4105
R25269 GNDA.n3265 GNDA.n3226 3.4105
R25270 GNDA.n3261 GNDA.n3260 3.4105
R25271 GNDA.n3259 GNDA.n3258 3.4105
R25272 GNDA.n3257 GNDA.n3256 3.4105
R25273 GNDA.n3255 GNDA.n3228 3.4105
R25274 GNDA.n3251 GNDA.n3250 3.4105
R25275 GNDA.n3249 GNDA.n3248 3.4105
R25276 GNDA.n3247 GNDA.n3246 3.4105
R25277 GNDA.n3245 GNDA.n3230 3.4105
R25278 GNDA.n3241 GNDA.n3240 3.4105
R25279 GNDA.n3239 GNDA.n3238 3.4105
R25280 GNDA.n3237 GNDA.n3236 3.4105
R25281 GNDA.n3235 GNDA.n3232 3.4105
R25282 GNDA.n2121 GNDA.n2120 3.4105
R25283 GNDA.n3287 GNDA.n3286 3.4105
R25284 GNDA.n2136 GNDA.n2135 3.4105
R25285 GNDA.n3205 GNDA.n3204 3.4105
R25286 GNDA.n3203 GNDA.n3202 3.4105
R25287 GNDA.n3201 GNDA.n3200 3.4105
R25288 GNDA.n3199 GNDA.n2138 3.4105
R25289 GNDA.n3195 GNDA.n3194 3.4105
R25290 GNDA.n3193 GNDA.n3192 3.4105
R25291 GNDA.n3191 GNDA.n3190 3.4105
R25292 GNDA.n3189 GNDA.n2140 3.4105
R25293 GNDA.n3185 GNDA.n3184 3.4105
R25294 GNDA.n3183 GNDA.n3182 3.4105
R25295 GNDA.n3181 GNDA.n3180 3.4105
R25296 GNDA.n3179 GNDA.n2142 3.4105
R25297 GNDA.n3175 GNDA.n3174 3.4105
R25298 GNDA.n3173 GNDA.n3172 3.4105
R25299 GNDA.n3171 GNDA.n3170 3.4105
R25300 GNDA.n3169 GNDA.n2144 3.4105
R25301 GNDA.n3165 GNDA.n3164 3.4105
R25302 GNDA.n3163 GNDA.n3162 3.4105
R25303 GNDA.n3161 GNDA.n3160 3.4105
R25304 GNDA.n3159 GNDA.n2146 3.4105
R25305 GNDA.n3155 GNDA.n3154 3.4105
R25306 GNDA.n3153 GNDA.n2123 3.4105
R25307 GNDA.n3106 GNDA.n3083 3.4105
R25308 GNDA.n3108 GNDA.n3082 3.4105
R25309 GNDA.n3109 GNDA.n3081 3.4105
R25310 GNDA.n3111 GNDA.n3080 3.4105
R25311 GNDA.n3112 GNDA.n3079 3.4105
R25312 GNDA.n3114 GNDA.n3078 3.4105
R25313 GNDA.n3115 GNDA.n3077 3.4105
R25314 GNDA.n3117 GNDA.n3076 3.4105
R25315 GNDA.n3118 GNDA.n3075 3.4105
R25316 GNDA.n3120 GNDA.n3074 3.4105
R25317 GNDA.n3121 GNDA.n3073 3.4105
R25318 GNDA.n3123 GNDA.n3072 3.4105
R25319 GNDA.n3124 GNDA.n3071 3.4105
R25320 GNDA.n3126 GNDA.n3070 3.4105
R25321 GNDA.n3127 GNDA.n3069 3.4105
R25322 GNDA.n3129 GNDA.n3068 3.4105
R25323 GNDA.n3130 GNDA.n3067 3.4105
R25324 GNDA.n3132 GNDA.n3066 3.4105
R25325 GNDA.n3133 GNDA.n3065 3.4105
R25326 GNDA.n3135 GNDA.n3064 3.4105
R25327 GNDA.n3136 GNDA.n3063 3.4105
R25328 GNDA.n3138 GNDA.n3062 3.4105
R25329 GNDA.n3140 GNDA.n3139 3.4105
R25330 GNDA.n2988 GNDA.n2987 3.4105
R25331 GNDA.n3047 GNDA.n3046 3.4105
R25332 GNDA.n3045 GNDA.n3044 3.4105
R25333 GNDA.n3043 GNDA.n3042 3.4105
R25334 GNDA.n3041 GNDA.n2990 3.4105
R25335 GNDA.n3037 GNDA.n3036 3.4105
R25336 GNDA.n3035 GNDA.n3034 3.4105
R25337 GNDA.n3033 GNDA.n3032 3.4105
R25338 GNDA.n3031 GNDA.n2992 3.4105
R25339 GNDA.n3027 GNDA.n3026 3.4105
R25340 GNDA.n3025 GNDA.n3024 3.4105
R25341 GNDA.n3023 GNDA.n3022 3.4105
R25342 GNDA.n3021 GNDA.n2994 3.4105
R25343 GNDA.n3017 GNDA.n3016 3.4105
R25344 GNDA.n3015 GNDA.n3014 3.4105
R25345 GNDA.n3013 GNDA.n3012 3.4105
R25346 GNDA.n3011 GNDA.n2996 3.4105
R25347 GNDA.n3007 GNDA.n3006 3.4105
R25348 GNDA.n3005 GNDA.n3004 3.4105
R25349 GNDA.n3003 GNDA.n3002 3.4105
R25350 GNDA.n3001 GNDA.n2998 3.4105
R25351 GNDA.n2160 GNDA.n2159 3.4105
R25352 GNDA.n3053 GNDA.n3052 3.4105
R25353 GNDA.n2175 GNDA.n2174 3.4105
R25354 GNDA.n2971 GNDA.n2970 3.4105
R25355 GNDA.n2969 GNDA.n2968 3.4105
R25356 GNDA.n2967 GNDA.n2966 3.4105
R25357 GNDA.n2965 GNDA.n2177 3.4105
R25358 GNDA.n2961 GNDA.n2960 3.4105
R25359 GNDA.n2959 GNDA.n2958 3.4105
R25360 GNDA.n2957 GNDA.n2956 3.4105
R25361 GNDA.n2955 GNDA.n2179 3.4105
R25362 GNDA.n2951 GNDA.n2950 3.4105
R25363 GNDA.n2949 GNDA.n2948 3.4105
R25364 GNDA.n2947 GNDA.n2946 3.4105
R25365 GNDA.n2945 GNDA.n2181 3.4105
R25366 GNDA.n2941 GNDA.n2940 3.4105
R25367 GNDA.n2939 GNDA.n2938 3.4105
R25368 GNDA.n2937 GNDA.n2936 3.4105
R25369 GNDA.n2935 GNDA.n2183 3.4105
R25370 GNDA.n2931 GNDA.n2930 3.4105
R25371 GNDA.n2929 GNDA.n2928 3.4105
R25372 GNDA.n2927 GNDA.n2926 3.4105
R25373 GNDA.n2925 GNDA.n2185 3.4105
R25374 GNDA.n2921 GNDA.n2920 3.4105
R25375 GNDA.n2919 GNDA.n2162 3.4105
R25376 GNDA.n2872 GNDA.n2849 3.4105
R25377 GNDA.n2874 GNDA.n2848 3.4105
R25378 GNDA.n2875 GNDA.n2847 3.4105
R25379 GNDA.n2877 GNDA.n2846 3.4105
R25380 GNDA.n2878 GNDA.n2845 3.4105
R25381 GNDA.n2880 GNDA.n2844 3.4105
R25382 GNDA.n2881 GNDA.n2843 3.4105
R25383 GNDA.n2883 GNDA.n2842 3.4105
R25384 GNDA.n2884 GNDA.n2841 3.4105
R25385 GNDA.n2886 GNDA.n2840 3.4105
R25386 GNDA.n2887 GNDA.n2839 3.4105
R25387 GNDA.n2889 GNDA.n2838 3.4105
R25388 GNDA.n2890 GNDA.n2837 3.4105
R25389 GNDA.n2892 GNDA.n2836 3.4105
R25390 GNDA.n2893 GNDA.n2835 3.4105
R25391 GNDA.n2895 GNDA.n2834 3.4105
R25392 GNDA.n2896 GNDA.n2833 3.4105
R25393 GNDA.n2898 GNDA.n2832 3.4105
R25394 GNDA.n2899 GNDA.n2831 3.4105
R25395 GNDA.n2901 GNDA.n2830 3.4105
R25396 GNDA.n2902 GNDA.n2829 3.4105
R25397 GNDA.n2904 GNDA.n2828 3.4105
R25398 GNDA.n2906 GNDA.n2905 3.4105
R25399 GNDA.n2754 GNDA.n2753 3.4105
R25400 GNDA.n2813 GNDA.n2812 3.4105
R25401 GNDA.n2811 GNDA.n2810 3.4105
R25402 GNDA.n2809 GNDA.n2808 3.4105
R25403 GNDA.n2807 GNDA.n2756 3.4105
R25404 GNDA.n2803 GNDA.n2802 3.4105
R25405 GNDA.n2801 GNDA.n2800 3.4105
R25406 GNDA.n2799 GNDA.n2798 3.4105
R25407 GNDA.n2797 GNDA.n2758 3.4105
R25408 GNDA.n2793 GNDA.n2792 3.4105
R25409 GNDA.n2791 GNDA.n2790 3.4105
R25410 GNDA.n2789 GNDA.n2788 3.4105
R25411 GNDA.n2787 GNDA.n2760 3.4105
R25412 GNDA.n2783 GNDA.n2782 3.4105
R25413 GNDA.n2781 GNDA.n2780 3.4105
R25414 GNDA.n2779 GNDA.n2778 3.4105
R25415 GNDA.n2777 GNDA.n2762 3.4105
R25416 GNDA.n2773 GNDA.n2772 3.4105
R25417 GNDA.n2771 GNDA.n2770 3.4105
R25418 GNDA.n2769 GNDA.n2768 3.4105
R25419 GNDA.n2767 GNDA.n2764 3.4105
R25420 GNDA.n2244 GNDA.n2243 3.4105
R25421 GNDA.n2819 GNDA.n2818 3.4105
R25422 GNDA.n2818 GNDA.n2817 3.4105
R25423 GNDA.n2817 GNDA.n2816 3.4105
R25424 GNDA.n2905 GNDA.n2161 3.4105
R25425 GNDA.n2871 GNDA.n2161 3.4105
R25426 GNDA.n2975 GNDA.n2162 3.4105
R25427 GNDA.n2975 GNDA.n2974 3.4105
R25428 GNDA.n3052 GNDA.n3051 3.4105
R25429 GNDA.n3051 GNDA.n3050 3.4105
R25430 GNDA.n3139 GNDA.n2122 3.4105
R25431 GNDA.n3105 GNDA.n2122 3.4105
R25432 GNDA.n3209 GNDA.n2123 3.4105
R25433 GNDA.n3209 GNDA.n3208 3.4105
R25434 GNDA.n3286 GNDA.n3285 3.4105
R25435 GNDA.n3285 GNDA.n3284 3.4105
R25436 GNDA.n3368 GNDA.n2004 3.4105
R25437 GNDA.n3368 GNDA.n3367 3.4105
R25438 GNDA.n3457 GNDA.n3369 3.4105
R25439 GNDA.n3457 GNDA.n3456 3.4105
R25440 GNDA.n2110 GNDA.n2003 3.4105
R25441 GNDA.n2076 GNDA.n2003 3.4105
R25442 GNDA.n4237 GNDA.n1975 3.4105
R25443 GNDA.n4238 GNDA.n4237 3.4105
R25444 GNDA.n3515 GNDA.n3486 3.4105
R25445 GNDA.n3559 GNDA.n3486 3.4105
R25446 GNDA.n3770 GNDA.n3690 3.4105
R25447 GNDA.n3770 GNDA.n3769 3.4105
R25448 GNDA.n3851 GNDA.n3771 3.4105
R25449 GNDA.n3851 GNDA.n3850 3.4105
R25450 GNDA.n4236 GNDA.n3474 3.4105
R25451 GNDA.n4236 GNDA.n4235 3.4105
R25452 GNDA.n3932 GNDA.n3852 3.4105
R25453 GNDA.n3932 GNDA.n3931 3.4105
R25454 GNDA.n4013 GNDA.n3933 3.4105
R25455 GNDA.n4013 GNDA.n4012 3.4105
R25456 GNDA.n4094 GNDA.n4014 3.4105
R25457 GNDA.n4094 GNDA.n4093 3.4105
R25458 GNDA.n4111 GNDA.n3662 3.4105
R25459 GNDA.n4112 GNDA.n4111 3.4105
R25460 GNDA.n2668 GNDA.n2666 3.4105
R25461 GNDA.n2739 GNDA.n2738 3.4105
R25462 GNDA.n2667 GNDA.n2665 3.4105
R25463 GNDA.n2733 GNDA.n2732 3.4105
R25464 GNDA.n2731 GNDA.n2730 3.4105
R25465 GNDA.n2729 GNDA.n2728 3.4105
R25466 GNDA.n2722 GNDA.n2670 3.4105
R25467 GNDA.n2724 GNDA.n2723 3.4105
R25468 GNDA.n2721 GNDA.n2720 3.4105
R25469 GNDA.n2719 GNDA.n2718 3.4105
R25470 GNDA.n2712 GNDA.n2672 3.4105
R25471 GNDA.n2714 GNDA.n2713 3.4105
R25472 GNDA.n2711 GNDA.n2710 3.4105
R25473 GNDA.n2709 GNDA.n2708 3.4105
R25474 GNDA.n2702 GNDA.n2674 3.4105
R25475 GNDA.n2704 GNDA.n2703 3.4105
R25476 GNDA.n2701 GNDA.n2700 3.4105
R25477 GNDA.n2699 GNDA.n2698 3.4105
R25478 GNDA.n2692 GNDA.n2676 3.4105
R25479 GNDA.n2694 GNDA.n2693 3.4105
R25480 GNDA.n2691 GNDA.n2690 3.4105
R25481 GNDA.n2689 GNDA.n2688 3.4105
R25482 GNDA.n14 GNDA.n13 3.4105
R25483 GNDA.n5595 GNDA.n5594 3.4105
R25484 GNDA.n5593 GNDA.n5592 3.4105
R25485 GNDA.n5591 GNDA.n5590 3.4105
R25486 GNDA.n5589 GNDA.n16 3.4105
R25487 GNDA.n5585 GNDA.n5584 3.4105
R25488 GNDA.n5583 GNDA.n5582 3.4105
R25489 GNDA.n5581 GNDA.n5580 3.4105
R25490 GNDA.n5579 GNDA.n18 3.4105
R25491 GNDA.n5575 GNDA.n5574 3.4105
R25492 GNDA.n5573 GNDA.n5572 3.4105
R25493 GNDA.n5571 GNDA.n5570 3.4105
R25494 GNDA.n5569 GNDA.n20 3.4105
R25495 GNDA.n5565 GNDA.n5564 3.4105
R25496 GNDA.n5563 GNDA.n5562 3.4105
R25497 GNDA.n5561 GNDA.n5560 3.4105
R25498 GNDA.n5559 GNDA.n22 3.4105
R25499 GNDA.n5555 GNDA.n5554 3.4105
R25500 GNDA.n5553 GNDA.n5552 3.4105
R25501 GNDA.n5551 GNDA.n5550 3.4105
R25502 GNDA.n5549 GNDA.n24 3.4105
R25503 GNDA.n5545 GNDA.n5544 3.4105
R25504 GNDA.n5543 GNDA.n1 3.4105
R25505 GNDA.n511 GNDA.n510 3.4105
R25506 GNDA.n570 GNDA.n569 3.4105
R25507 GNDA.n568 GNDA.n567 3.4105
R25508 GNDA.n566 GNDA.n565 3.4105
R25509 GNDA.n564 GNDA.n513 3.4105
R25510 GNDA.n560 GNDA.n559 3.4105
R25511 GNDA.n558 GNDA.n557 3.4105
R25512 GNDA.n556 GNDA.n555 3.4105
R25513 GNDA.n554 GNDA.n515 3.4105
R25514 GNDA.n550 GNDA.n549 3.4105
R25515 GNDA.n548 GNDA.n547 3.4105
R25516 GNDA.n546 GNDA.n545 3.4105
R25517 GNDA.n544 GNDA.n517 3.4105
R25518 GNDA.n540 GNDA.n539 3.4105
R25519 GNDA.n538 GNDA.n537 3.4105
R25520 GNDA.n536 GNDA.n535 3.4105
R25521 GNDA.n534 GNDA.n519 3.4105
R25522 GNDA.n530 GNDA.n529 3.4105
R25523 GNDA.n528 GNDA.n527 3.4105
R25524 GNDA.n526 GNDA.n525 3.4105
R25525 GNDA.n524 GNDA.n521 3.4105
R25526 GNDA.n48 GNDA.n47 3.4105
R25527 GNDA.n576 GNDA.n575 3.4105
R25528 GNDA.n318 GNDA.n295 3.4105
R25529 GNDA.n320 GNDA.n294 3.4105
R25530 GNDA.n321 GNDA.n293 3.4105
R25531 GNDA.n323 GNDA.n292 3.4105
R25532 GNDA.n324 GNDA.n291 3.4105
R25533 GNDA.n326 GNDA.n290 3.4105
R25534 GNDA.n327 GNDA.n289 3.4105
R25535 GNDA.n329 GNDA.n288 3.4105
R25536 GNDA.n330 GNDA.n287 3.4105
R25537 GNDA.n332 GNDA.n286 3.4105
R25538 GNDA.n333 GNDA.n285 3.4105
R25539 GNDA.n335 GNDA.n284 3.4105
R25540 GNDA.n336 GNDA.n283 3.4105
R25541 GNDA.n338 GNDA.n282 3.4105
R25542 GNDA.n339 GNDA.n281 3.4105
R25543 GNDA.n341 GNDA.n280 3.4105
R25544 GNDA.n342 GNDA.n279 3.4105
R25545 GNDA.n344 GNDA.n278 3.4105
R25546 GNDA.n345 GNDA.n277 3.4105
R25547 GNDA.n347 GNDA.n276 3.4105
R25548 GNDA.n348 GNDA.n275 3.4105
R25549 GNDA.n350 GNDA.n274 3.4105
R25550 GNDA.n352 GNDA.n351 3.4105
R25551 GNDA.n201 GNDA.n200 3.4105
R25552 GNDA.n260 GNDA.n259 3.4105
R25553 GNDA.n258 GNDA.n257 3.4105
R25554 GNDA.n256 GNDA.n255 3.4105
R25555 GNDA.n254 GNDA.n203 3.4105
R25556 GNDA.n250 GNDA.n249 3.4105
R25557 GNDA.n248 GNDA.n247 3.4105
R25558 GNDA.n246 GNDA.n245 3.4105
R25559 GNDA.n244 GNDA.n205 3.4105
R25560 GNDA.n240 GNDA.n239 3.4105
R25561 GNDA.n238 GNDA.n237 3.4105
R25562 GNDA.n236 GNDA.n235 3.4105
R25563 GNDA.n234 GNDA.n207 3.4105
R25564 GNDA.n230 GNDA.n229 3.4105
R25565 GNDA.n228 GNDA.n227 3.4105
R25566 GNDA.n226 GNDA.n225 3.4105
R25567 GNDA.n224 GNDA.n209 3.4105
R25568 GNDA.n220 GNDA.n219 3.4105
R25569 GNDA.n218 GNDA.n217 3.4105
R25570 GNDA.n216 GNDA.n215 3.4105
R25571 GNDA.n214 GNDA.n211 3.4105
R25572 GNDA.n188 GNDA.n187 3.4105
R25573 GNDA.n266 GNDA.n265 3.4105
R25574 GNDA.n145 GNDA.n122 3.4105
R25575 GNDA.n147 GNDA.n121 3.4105
R25576 GNDA.n148 GNDA.n120 3.4105
R25577 GNDA.n150 GNDA.n119 3.4105
R25578 GNDA.n151 GNDA.n118 3.4105
R25579 GNDA.n153 GNDA.n117 3.4105
R25580 GNDA.n154 GNDA.n116 3.4105
R25581 GNDA.n156 GNDA.n115 3.4105
R25582 GNDA.n157 GNDA.n114 3.4105
R25583 GNDA.n159 GNDA.n113 3.4105
R25584 GNDA.n160 GNDA.n112 3.4105
R25585 GNDA.n162 GNDA.n111 3.4105
R25586 GNDA.n163 GNDA.n110 3.4105
R25587 GNDA.n165 GNDA.n109 3.4105
R25588 GNDA.n166 GNDA.n108 3.4105
R25589 GNDA.n168 GNDA.n107 3.4105
R25590 GNDA.n169 GNDA.n106 3.4105
R25591 GNDA.n171 GNDA.n105 3.4105
R25592 GNDA.n172 GNDA.n104 3.4105
R25593 GNDA.n174 GNDA.n103 3.4105
R25594 GNDA.n175 GNDA.n102 3.4105
R25595 GNDA.n177 GNDA.n101 3.4105
R25596 GNDA.n179 GNDA.n178 3.4105
R25597 GNDA.n86 GNDA.n85 3.4105
R25598 GNDA.n504 GNDA.n503 3.4105
R25599 GNDA.n502 GNDA.n501 3.4105
R25600 GNDA.n500 GNDA.n499 3.4105
R25601 GNDA.n498 GNDA.n88 3.4105
R25602 GNDA.n494 GNDA.n493 3.4105
R25603 GNDA.n492 GNDA.n491 3.4105
R25604 GNDA.n490 GNDA.n489 3.4105
R25605 GNDA.n488 GNDA.n90 3.4105
R25606 GNDA.n484 GNDA.n483 3.4105
R25607 GNDA.n482 GNDA.n481 3.4105
R25608 GNDA.n480 GNDA.n479 3.4105
R25609 GNDA.n478 GNDA.n92 3.4105
R25610 GNDA.n474 GNDA.n473 3.4105
R25611 GNDA.n472 GNDA.n471 3.4105
R25612 GNDA.n470 GNDA.n469 3.4105
R25613 GNDA.n468 GNDA.n94 3.4105
R25614 GNDA.n464 GNDA.n463 3.4105
R25615 GNDA.n462 GNDA.n461 3.4105
R25616 GNDA.n460 GNDA.n459 3.4105
R25617 GNDA.n458 GNDA.n96 3.4105
R25618 GNDA.n454 GNDA.n453 3.4105
R25619 GNDA.n452 GNDA.n72 3.4105
R25620 GNDA.n508 GNDA.n72 3.4105
R25621 GNDA.n508 GNDA.n507 3.4105
R25622 GNDA.n178 GNDA.n84 3.4105
R25623 GNDA.n144 GNDA.n84 3.4105
R25624 GNDA.n265 GNDA.n264 3.4105
R25625 GNDA.n264 GNDA.n263 3.4105
R25626 GNDA.n351 GNDA.n0 3.4105
R25627 GNDA.n317 GNDA.n0 3.4105
R25628 GNDA.n575 GNDA.n574 3.4105
R25629 GNDA.n574 GNDA.n573 3.4105
R25630 GNDA.n5599 GNDA.n1 3.4105
R25631 GNDA.n5599 GNDA.n5598 3.4105
R25632 GNDA.n410 GNDA.n408 3.4105
R25633 GNDA.n411 GNDA.n407 3.4105
R25634 GNDA.n412 GNDA.n406 3.4105
R25635 GNDA.n405 GNDA.n403 3.4105
R25636 GNDA.n416 GNDA.n402 3.4105
R25637 GNDA.n417 GNDA.n401 3.4105
R25638 GNDA.n418 GNDA.n400 3.4105
R25639 GNDA.n399 GNDA.n397 3.4105
R25640 GNDA.n422 GNDA.n396 3.4105
R25641 GNDA.n423 GNDA.n395 3.4105
R25642 GNDA.n424 GNDA.n394 3.4105
R25643 GNDA.n393 GNDA.n391 3.4105
R25644 GNDA.n428 GNDA.n390 3.4105
R25645 GNDA.n429 GNDA.n389 3.4105
R25646 GNDA.n430 GNDA.n388 3.4105
R25647 GNDA.n387 GNDA.n385 3.4105
R25648 GNDA.n434 GNDA.n384 3.4105
R25649 GNDA.n435 GNDA.n383 3.4105
R25650 GNDA.n436 GNDA.n382 3.4105
R25651 GNDA.n381 GNDA.n379 3.4105
R25652 GNDA.n440 GNDA.n378 3.4105
R25653 GNDA.n441 GNDA.n377 3.4105
R25654 GNDA.n953 GNDA.n952 3.4105
R25655 GNDA.n1028 GNDA.n1027 3.4105
R25656 GNDA.n967 GNDA.n966 3.4105
R25657 GNDA.n1023 GNDA.n1022 3.4105
R25658 GNDA.n1021 GNDA.n1020 3.4105
R25659 GNDA.n1019 GNDA.n1018 3.4105
R25660 GNDA.n1017 GNDA.n969 3.4105
R25661 GNDA.n1013 GNDA.n1012 3.4105
R25662 GNDA.n1011 GNDA.n1010 3.4105
R25663 GNDA.n1009 GNDA.n1008 3.4105
R25664 GNDA.n1007 GNDA.n971 3.4105
R25665 GNDA.n1003 GNDA.n1002 3.4105
R25666 GNDA.n1001 GNDA.n1000 3.4105
R25667 GNDA.n999 GNDA.n998 3.4105
R25668 GNDA.n997 GNDA.n973 3.4105
R25669 GNDA.n993 GNDA.n992 3.4105
R25670 GNDA.n991 GNDA.n990 3.4105
R25671 GNDA.n989 GNDA.n988 3.4105
R25672 GNDA.n987 GNDA.n975 3.4105
R25673 GNDA.n983 GNDA.n982 3.4105
R25674 GNDA.n981 GNDA.n980 3.4105
R25675 GNDA.n979 GNDA.n978 3.4105
R25676 GNDA.n4899 GNDA.n4898 3.4105
R25677 GNDA.n4897 GNDA.n955 3.4105
R25678 GNDA.n4898 GNDA.n4897 3.4105
R25679 GNDA.n4896 GNDA.n1030 3.4105
R25680 GNDA.n4896 GNDA.n4895 3.4105
R25681 GNDA.n2540 GNDA.n2492 3.4105
R25682 GNDA.n2543 GNDA.n2492 3.4105
R25683 GNDA.n2543 GNDA.n2473 3.4105
R25684 GNDA.n2540 GNDA.n2495 3.4105
R25685 GNDA.n2495 GNDA.n2426 3.4105
R25686 GNDA.n2495 GNDA.n2424 3.4105
R25687 GNDA.n2495 GNDA.n2427 3.4105
R25688 GNDA.n2495 GNDA.n2423 3.4105
R25689 GNDA.n2495 GNDA.n2428 3.4105
R25690 GNDA.n2495 GNDA.n2422 3.4105
R25691 GNDA.n2495 GNDA.n2429 3.4105
R25692 GNDA.n2495 GNDA.n2421 3.4105
R25693 GNDA.n2495 GNDA.n2430 3.4105
R25694 GNDA.n2495 GNDA.n2420 3.4105
R25695 GNDA.n2495 GNDA.n2431 3.4105
R25696 GNDA.n2495 GNDA.n2419 3.4105
R25697 GNDA.n2495 GNDA.n2432 3.4105
R25698 GNDA.n2495 GNDA.n2418 3.4105
R25699 GNDA.n2495 GNDA.n2433 3.4105
R25700 GNDA.n2495 GNDA.n2417 3.4105
R25701 GNDA.n2495 GNDA.n2434 3.4105
R25702 GNDA.n2495 GNDA.n2416 3.4105
R25703 GNDA.n2495 GNDA.n2435 3.4105
R25704 GNDA.n2495 GNDA.n2415 3.4105
R25705 GNDA.n2495 GNDA.n2436 3.4105
R25706 GNDA.n2495 GNDA.n2414 3.4105
R25707 GNDA.n2495 GNDA.n2437 3.4105
R25708 GNDA.n2495 GNDA.n2413 3.4105
R25709 GNDA.n2495 GNDA.n2438 3.4105
R25710 GNDA.n2495 GNDA.n2412 3.4105
R25711 GNDA.n2495 GNDA.n2439 3.4105
R25712 GNDA.n2495 GNDA.n2411 3.4105
R25713 GNDA.n2495 GNDA.n2440 3.4105
R25714 GNDA.n2495 GNDA.n2410 3.4105
R25715 GNDA.n2495 GNDA.n2441 3.4105
R25716 GNDA.n2543 GNDA.n2495 3.4105
R25717 GNDA.n2540 GNDA.n2457 3.4105
R25718 GNDA.n2457 GNDA.n2426 3.4105
R25719 GNDA.n2457 GNDA.n2424 3.4105
R25720 GNDA.n2457 GNDA.n2427 3.4105
R25721 GNDA.n2457 GNDA.n2423 3.4105
R25722 GNDA.n2457 GNDA.n2428 3.4105
R25723 GNDA.n2457 GNDA.n2422 3.4105
R25724 GNDA.n2457 GNDA.n2429 3.4105
R25725 GNDA.n2457 GNDA.n2421 3.4105
R25726 GNDA.n2457 GNDA.n2430 3.4105
R25727 GNDA.n2457 GNDA.n2420 3.4105
R25728 GNDA.n2457 GNDA.n2431 3.4105
R25729 GNDA.n2457 GNDA.n2419 3.4105
R25730 GNDA.n2457 GNDA.n2432 3.4105
R25731 GNDA.n2457 GNDA.n2418 3.4105
R25732 GNDA.n2457 GNDA.n2433 3.4105
R25733 GNDA.n2457 GNDA.n2417 3.4105
R25734 GNDA.n2457 GNDA.n2434 3.4105
R25735 GNDA.n2457 GNDA.n2416 3.4105
R25736 GNDA.n2457 GNDA.n2435 3.4105
R25737 GNDA.n2457 GNDA.n2415 3.4105
R25738 GNDA.n2457 GNDA.n2436 3.4105
R25739 GNDA.n2457 GNDA.n2414 3.4105
R25740 GNDA.n2457 GNDA.n2437 3.4105
R25741 GNDA.n2457 GNDA.n2413 3.4105
R25742 GNDA.n2457 GNDA.n2438 3.4105
R25743 GNDA.n2457 GNDA.n2412 3.4105
R25744 GNDA.n2457 GNDA.n2439 3.4105
R25745 GNDA.n2457 GNDA.n2411 3.4105
R25746 GNDA.n2457 GNDA.n2440 3.4105
R25747 GNDA.n2457 GNDA.n2410 3.4105
R25748 GNDA.n2457 GNDA.n2441 3.4105
R25749 GNDA.n2543 GNDA.n2457 3.4105
R25750 GNDA.n2540 GNDA.n2498 3.4105
R25751 GNDA.n2498 GNDA.n2426 3.4105
R25752 GNDA.n2498 GNDA.n2424 3.4105
R25753 GNDA.n2498 GNDA.n2427 3.4105
R25754 GNDA.n2498 GNDA.n2423 3.4105
R25755 GNDA.n2498 GNDA.n2428 3.4105
R25756 GNDA.n2498 GNDA.n2422 3.4105
R25757 GNDA.n2498 GNDA.n2429 3.4105
R25758 GNDA.n2498 GNDA.n2421 3.4105
R25759 GNDA.n2498 GNDA.n2430 3.4105
R25760 GNDA.n2498 GNDA.n2420 3.4105
R25761 GNDA.n2498 GNDA.n2431 3.4105
R25762 GNDA.n2498 GNDA.n2419 3.4105
R25763 GNDA.n2498 GNDA.n2432 3.4105
R25764 GNDA.n2498 GNDA.n2418 3.4105
R25765 GNDA.n2498 GNDA.n2433 3.4105
R25766 GNDA.n2498 GNDA.n2417 3.4105
R25767 GNDA.n2498 GNDA.n2434 3.4105
R25768 GNDA.n2498 GNDA.n2416 3.4105
R25769 GNDA.n2498 GNDA.n2435 3.4105
R25770 GNDA.n2498 GNDA.n2415 3.4105
R25771 GNDA.n2498 GNDA.n2436 3.4105
R25772 GNDA.n2498 GNDA.n2414 3.4105
R25773 GNDA.n2498 GNDA.n2437 3.4105
R25774 GNDA.n2498 GNDA.n2413 3.4105
R25775 GNDA.n2498 GNDA.n2438 3.4105
R25776 GNDA.n2498 GNDA.n2412 3.4105
R25777 GNDA.n2498 GNDA.n2439 3.4105
R25778 GNDA.n2498 GNDA.n2411 3.4105
R25779 GNDA.n2498 GNDA.n2440 3.4105
R25780 GNDA.n2498 GNDA.n2410 3.4105
R25781 GNDA.n2498 GNDA.n2441 3.4105
R25782 GNDA.n2543 GNDA.n2498 3.4105
R25783 GNDA.n2540 GNDA.n2456 3.4105
R25784 GNDA.n2456 GNDA.n2426 3.4105
R25785 GNDA.n2456 GNDA.n2424 3.4105
R25786 GNDA.n2456 GNDA.n2427 3.4105
R25787 GNDA.n2456 GNDA.n2423 3.4105
R25788 GNDA.n2456 GNDA.n2428 3.4105
R25789 GNDA.n2456 GNDA.n2422 3.4105
R25790 GNDA.n2456 GNDA.n2429 3.4105
R25791 GNDA.n2456 GNDA.n2421 3.4105
R25792 GNDA.n2456 GNDA.n2430 3.4105
R25793 GNDA.n2456 GNDA.n2420 3.4105
R25794 GNDA.n2456 GNDA.n2431 3.4105
R25795 GNDA.n2456 GNDA.n2419 3.4105
R25796 GNDA.n2456 GNDA.n2432 3.4105
R25797 GNDA.n2456 GNDA.n2418 3.4105
R25798 GNDA.n2456 GNDA.n2433 3.4105
R25799 GNDA.n2456 GNDA.n2417 3.4105
R25800 GNDA.n2456 GNDA.n2434 3.4105
R25801 GNDA.n2456 GNDA.n2416 3.4105
R25802 GNDA.n2456 GNDA.n2435 3.4105
R25803 GNDA.n2456 GNDA.n2415 3.4105
R25804 GNDA.n2456 GNDA.n2436 3.4105
R25805 GNDA.n2456 GNDA.n2414 3.4105
R25806 GNDA.n2456 GNDA.n2437 3.4105
R25807 GNDA.n2456 GNDA.n2413 3.4105
R25808 GNDA.n2456 GNDA.n2438 3.4105
R25809 GNDA.n2456 GNDA.n2412 3.4105
R25810 GNDA.n2456 GNDA.n2439 3.4105
R25811 GNDA.n2456 GNDA.n2411 3.4105
R25812 GNDA.n2456 GNDA.n2440 3.4105
R25813 GNDA.n2456 GNDA.n2410 3.4105
R25814 GNDA.n2456 GNDA.n2441 3.4105
R25815 GNDA.n2543 GNDA.n2456 3.4105
R25816 GNDA.n2540 GNDA.n2501 3.4105
R25817 GNDA.n2501 GNDA.n2426 3.4105
R25818 GNDA.n2501 GNDA.n2424 3.4105
R25819 GNDA.n2501 GNDA.n2427 3.4105
R25820 GNDA.n2501 GNDA.n2423 3.4105
R25821 GNDA.n2501 GNDA.n2428 3.4105
R25822 GNDA.n2501 GNDA.n2422 3.4105
R25823 GNDA.n2501 GNDA.n2429 3.4105
R25824 GNDA.n2501 GNDA.n2421 3.4105
R25825 GNDA.n2501 GNDA.n2430 3.4105
R25826 GNDA.n2501 GNDA.n2420 3.4105
R25827 GNDA.n2501 GNDA.n2431 3.4105
R25828 GNDA.n2501 GNDA.n2419 3.4105
R25829 GNDA.n2501 GNDA.n2432 3.4105
R25830 GNDA.n2501 GNDA.n2418 3.4105
R25831 GNDA.n2501 GNDA.n2433 3.4105
R25832 GNDA.n2501 GNDA.n2417 3.4105
R25833 GNDA.n2501 GNDA.n2434 3.4105
R25834 GNDA.n2501 GNDA.n2416 3.4105
R25835 GNDA.n2501 GNDA.n2435 3.4105
R25836 GNDA.n2501 GNDA.n2415 3.4105
R25837 GNDA.n2501 GNDA.n2436 3.4105
R25838 GNDA.n2501 GNDA.n2414 3.4105
R25839 GNDA.n2501 GNDA.n2437 3.4105
R25840 GNDA.n2501 GNDA.n2413 3.4105
R25841 GNDA.n2501 GNDA.n2438 3.4105
R25842 GNDA.n2501 GNDA.n2412 3.4105
R25843 GNDA.n2501 GNDA.n2439 3.4105
R25844 GNDA.n2501 GNDA.n2411 3.4105
R25845 GNDA.n2501 GNDA.n2440 3.4105
R25846 GNDA.n2501 GNDA.n2410 3.4105
R25847 GNDA.n2501 GNDA.n2441 3.4105
R25848 GNDA.n2543 GNDA.n2501 3.4105
R25849 GNDA.n2540 GNDA.n2455 3.4105
R25850 GNDA.n2455 GNDA.n2426 3.4105
R25851 GNDA.n2455 GNDA.n2424 3.4105
R25852 GNDA.n2455 GNDA.n2427 3.4105
R25853 GNDA.n2455 GNDA.n2423 3.4105
R25854 GNDA.n2455 GNDA.n2428 3.4105
R25855 GNDA.n2455 GNDA.n2422 3.4105
R25856 GNDA.n2455 GNDA.n2429 3.4105
R25857 GNDA.n2455 GNDA.n2421 3.4105
R25858 GNDA.n2455 GNDA.n2430 3.4105
R25859 GNDA.n2455 GNDA.n2420 3.4105
R25860 GNDA.n2455 GNDA.n2431 3.4105
R25861 GNDA.n2455 GNDA.n2419 3.4105
R25862 GNDA.n2455 GNDA.n2432 3.4105
R25863 GNDA.n2455 GNDA.n2418 3.4105
R25864 GNDA.n2455 GNDA.n2433 3.4105
R25865 GNDA.n2455 GNDA.n2417 3.4105
R25866 GNDA.n2455 GNDA.n2434 3.4105
R25867 GNDA.n2455 GNDA.n2416 3.4105
R25868 GNDA.n2455 GNDA.n2435 3.4105
R25869 GNDA.n2455 GNDA.n2415 3.4105
R25870 GNDA.n2455 GNDA.n2436 3.4105
R25871 GNDA.n2455 GNDA.n2414 3.4105
R25872 GNDA.n2455 GNDA.n2437 3.4105
R25873 GNDA.n2455 GNDA.n2413 3.4105
R25874 GNDA.n2455 GNDA.n2438 3.4105
R25875 GNDA.n2455 GNDA.n2412 3.4105
R25876 GNDA.n2455 GNDA.n2439 3.4105
R25877 GNDA.n2455 GNDA.n2411 3.4105
R25878 GNDA.n2455 GNDA.n2440 3.4105
R25879 GNDA.n2455 GNDA.n2410 3.4105
R25880 GNDA.n2455 GNDA.n2441 3.4105
R25881 GNDA.n2543 GNDA.n2455 3.4105
R25882 GNDA.n2540 GNDA.n2504 3.4105
R25883 GNDA.n2504 GNDA.n2426 3.4105
R25884 GNDA.n2504 GNDA.n2424 3.4105
R25885 GNDA.n2504 GNDA.n2427 3.4105
R25886 GNDA.n2504 GNDA.n2423 3.4105
R25887 GNDA.n2504 GNDA.n2428 3.4105
R25888 GNDA.n2504 GNDA.n2422 3.4105
R25889 GNDA.n2504 GNDA.n2429 3.4105
R25890 GNDA.n2504 GNDA.n2421 3.4105
R25891 GNDA.n2504 GNDA.n2430 3.4105
R25892 GNDA.n2504 GNDA.n2420 3.4105
R25893 GNDA.n2504 GNDA.n2431 3.4105
R25894 GNDA.n2504 GNDA.n2419 3.4105
R25895 GNDA.n2504 GNDA.n2432 3.4105
R25896 GNDA.n2504 GNDA.n2418 3.4105
R25897 GNDA.n2504 GNDA.n2433 3.4105
R25898 GNDA.n2504 GNDA.n2417 3.4105
R25899 GNDA.n2504 GNDA.n2434 3.4105
R25900 GNDA.n2504 GNDA.n2416 3.4105
R25901 GNDA.n2504 GNDA.n2435 3.4105
R25902 GNDA.n2504 GNDA.n2415 3.4105
R25903 GNDA.n2504 GNDA.n2436 3.4105
R25904 GNDA.n2504 GNDA.n2414 3.4105
R25905 GNDA.n2504 GNDA.n2437 3.4105
R25906 GNDA.n2504 GNDA.n2413 3.4105
R25907 GNDA.n2504 GNDA.n2438 3.4105
R25908 GNDA.n2504 GNDA.n2412 3.4105
R25909 GNDA.n2504 GNDA.n2439 3.4105
R25910 GNDA.n2504 GNDA.n2411 3.4105
R25911 GNDA.n2504 GNDA.n2440 3.4105
R25912 GNDA.n2504 GNDA.n2410 3.4105
R25913 GNDA.n2504 GNDA.n2441 3.4105
R25914 GNDA.n2543 GNDA.n2504 3.4105
R25915 GNDA.n2540 GNDA.n2454 3.4105
R25916 GNDA.n2454 GNDA.n2426 3.4105
R25917 GNDA.n2454 GNDA.n2424 3.4105
R25918 GNDA.n2454 GNDA.n2427 3.4105
R25919 GNDA.n2454 GNDA.n2423 3.4105
R25920 GNDA.n2454 GNDA.n2428 3.4105
R25921 GNDA.n2454 GNDA.n2422 3.4105
R25922 GNDA.n2454 GNDA.n2429 3.4105
R25923 GNDA.n2454 GNDA.n2421 3.4105
R25924 GNDA.n2454 GNDA.n2430 3.4105
R25925 GNDA.n2454 GNDA.n2420 3.4105
R25926 GNDA.n2454 GNDA.n2431 3.4105
R25927 GNDA.n2454 GNDA.n2419 3.4105
R25928 GNDA.n2454 GNDA.n2432 3.4105
R25929 GNDA.n2454 GNDA.n2418 3.4105
R25930 GNDA.n2454 GNDA.n2433 3.4105
R25931 GNDA.n2454 GNDA.n2417 3.4105
R25932 GNDA.n2454 GNDA.n2434 3.4105
R25933 GNDA.n2454 GNDA.n2416 3.4105
R25934 GNDA.n2454 GNDA.n2435 3.4105
R25935 GNDA.n2454 GNDA.n2415 3.4105
R25936 GNDA.n2454 GNDA.n2436 3.4105
R25937 GNDA.n2454 GNDA.n2414 3.4105
R25938 GNDA.n2454 GNDA.n2437 3.4105
R25939 GNDA.n2454 GNDA.n2413 3.4105
R25940 GNDA.n2454 GNDA.n2438 3.4105
R25941 GNDA.n2454 GNDA.n2412 3.4105
R25942 GNDA.n2454 GNDA.n2439 3.4105
R25943 GNDA.n2454 GNDA.n2411 3.4105
R25944 GNDA.n2454 GNDA.n2440 3.4105
R25945 GNDA.n2454 GNDA.n2410 3.4105
R25946 GNDA.n2454 GNDA.n2441 3.4105
R25947 GNDA.n2543 GNDA.n2454 3.4105
R25948 GNDA.n2540 GNDA.n2507 3.4105
R25949 GNDA.n2507 GNDA.n2426 3.4105
R25950 GNDA.n2507 GNDA.n2424 3.4105
R25951 GNDA.n2507 GNDA.n2427 3.4105
R25952 GNDA.n2507 GNDA.n2423 3.4105
R25953 GNDA.n2507 GNDA.n2428 3.4105
R25954 GNDA.n2507 GNDA.n2422 3.4105
R25955 GNDA.n2507 GNDA.n2429 3.4105
R25956 GNDA.n2507 GNDA.n2421 3.4105
R25957 GNDA.n2507 GNDA.n2430 3.4105
R25958 GNDA.n2507 GNDA.n2420 3.4105
R25959 GNDA.n2507 GNDA.n2431 3.4105
R25960 GNDA.n2507 GNDA.n2419 3.4105
R25961 GNDA.n2507 GNDA.n2432 3.4105
R25962 GNDA.n2507 GNDA.n2418 3.4105
R25963 GNDA.n2507 GNDA.n2433 3.4105
R25964 GNDA.n2507 GNDA.n2417 3.4105
R25965 GNDA.n2507 GNDA.n2434 3.4105
R25966 GNDA.n2507 GNDA.n2416 3.4105
R25967 GNDA.n2507 GNDA.n2435 3.4105
R25968 GNDA.n2507 GNDA.n2415 3.4105
R25969 GNDA.n2507 GNDA.n2436 3.4105
R25970 GNDA.n2507 GNDA.n2414 3.4105
R25971 GNDA.n2507 GNDA.n2437 3.4105
R25972 GNDA.n2507 GNDA.n2413 3.4105
R25973 GNDA.n2507 GNDA.n2438 3.4105
R25974 GNDA.n2507 GNDA.n2412 3.4105
R25975 GNDA.n2507 GNDA.n2439 3.4105
R25976 GNDA.n2507 GNDA.n2411 3.4105
R25977 GNDA.n2507 GNDA.n2440 3.4105
R25978 GNDA.n2507 GNDA.n2410 3.4105
R25979 GNDA.n2507 GNDA.n2441 3.4105
R25980 GNDA.n2543 GNDA.n2507 3.4105
R25981 GNDA.n2540 GNDA.n2453 3.4105
R25982 GNDA.n2453 GNDA.n2426 3.4105
R25983 GNDA.n2453 GNDA.n2424 3.4105
R25984 GNDA.n2453 GNDA.n2427 3.4105
R25985 GNDA.n2453 GNDA.n2423 3.4105
R25986 GNDA.n2453 GNDA.n2428 3.4105
R25987 GNDA.n2453 GNDA.n2422 3.4105
R25988 GNDA.n2453 GNDA.n2429 3.4105
R25989 GNDA.n2453 GNDA.n2421 3.4105
R25990 GNDA.n2453 GNDA.n2430 3.4105
R25991 GNDA.n2453 GNDA.n2420 3.4105
R25992 GNDA.n2453 GNDA.n2431 3.4105
R25993 GNDA.n2453 GNDA.n2419 3.4105
R25994 GNDA.n2453 GNDA.n2432 3.4105
R25995 GNDA.n2453 GNDA.n2418 3.4105
R25996 GNDA.n2453 GNDA.n2433 3.4105
R25997 GNDA.n2453 GNDA.n2417 3.4105
R25998 GNDA.n2453 GNDA.n2434 3.4105
R25999 GNDA.n2453 GNDA.n2416 3.4105
R26000 GNDA.n2453 GNDA.n2435 3.4105
R26001 GNDA.n2453 GNDA.n2415 3.4105
R26002 GNDA.n2453 GNDA.n2436 3.4105
R26003 GNDA.n2453 GNDA.n2414 3.4105
R26004 GNDA.n2453 GNDA.n2437 3.4105
R26005 GNDA.n2453 GNDA.n2413 3.4105
R26006 GNDA.n2453 GNDA.n2438 3.4105
R26007 GNDA.n2453 GNDA.n2412 3.4105
R26008 GNDA.n2453 GNDA.n2439 3.4105
R26009 GNDA.n2453 GNDA.n2411 3.4105
R26010 GNDA.n2453 GNDA.n2440 3.4105
R26011 GNDA.n2453 GNDA.n2410 3.4105
R26012 GNDA.n2453 GNDA.n2441 3.4105
R26013 GNDA.n2543 GNDA.n2453 3.4105
R26014 GNDA.n2540 GNDA.n2510 3.4105
R26015 GNDA.n2510 GNDA.n2426 3.4105
R26016 GNDA.n2510 GNDA.n2424 3.4105
R26017 GNDA.n2510 GNDA.n2427 3.4105
R26018 GNDA.n2510 GNDA.n2423 3.4105
R26019 GNDA.n2510 GNDA.n2428 3.4105
R26020 GNDA.n2510 GNDA.n2422 3.4105
R26021 GNDA.n2510 GNDA.n2429 3.4105
R26022 GNDA.n2510 GNDA.n2421 3.4105
R26023 GNDA.n2510 GNDA.n2430 3.4105
R26024 GNDA.n2510 GNDA.n2420 3.4105
R26025 GNDA.n2510 GNDA.n2431 3.4105
R26026 GNDA.n2510 GNDA.n2419 3.4105
R26027 GNDA.n2510 GNDA.n2432 3.4105
R26028 GNDA.n2510 GNDA.n2418 3.4105
R26029 GNDA.n2510 GNDA.n2433 3.4105
R26030 GNDA.n2510 GNDA.n2417 3.4105
R26031 GNDA.n2510 GNDA.n2434 3.4105
R26032 GNDA.n2510 GNDA.n2416 3.4105
R26033 GNDA.n2510 GNDA.n2435 3.4105
R26034 GNDA.n2510 GNDA.n2415 3.4105
R26035 GNDA.n2510 GNDA.n2436 3.4105
R26036 GNDA.n2510 GNDA.n2414 3.4105
R26037 GNDA.n2510 GNDA.n2437 3.4105
R26038 GNDA.n2510 GNDA.n2413 3.4105
R26039 GNDA.n2510 GNDA.n2438 3.4105
R26040 GNDA.n2510 GNDA.n2412 3.4105
R26041 GNDA.n2510 GNDA.n2439 3.4105
R26042 GNDA.n2510 GNDA.n2411 3.4105
R26043 GNDA.n2510 GNDA.n2440 3.4105
R26044 GNDA.n2510 GNDA.n2410 3.4105
R26045 GNDA.n2510 GNDA.n2441 3.4105
R26046 GNDA.n2543 GNDA.n2510 3.4105
R26047 GNDA.n2540 GNDA.n2452 3.4105
R26048 GNDA.n2452 GNDA.n2426 3.4105
R26049 GNDA.n2452 GNDA.n2424 3.4105
R26050 GNDA.n2452 GNDA.n2427 3.4105
R26051 GNDA.n2452 GNDA.n2423 3.4105
R26052 GNDA.n2452 GNDA.n2428 3.4105
R26053 GNDA.n2452 GNDA.n2422 3.4105
R26054 GNDA.n2452 GNDA.n2429 3.4105
R26055 GNDA.n2452 GNDA.n2421 3.4105
R26056 GNDA.n2452 GNDA.n2430 3.4105
R26057 GNDA.n2452 GNDA.n2420 3.4105
R26058 GNDA.n2452 GNDA.n2431 3.4105
R26059 GNDA.n2452 GNDA.n2419 3.4105
R26060 GNDA.n2452 GNDA.n2432 3.4105
R26061 GNDA.n2452 GNDA.n2418 3.4105
R26062 GNDA.n2452 GNDA.n2433 3.4105
R26063 GNDA.n2452 GNDA.n2417 3.4105
R26064 GNDA.n2452 GNDA.n2434 3.4105
R26065 GNDA.n2452 GNDA.n2416 3.4105
R26066 GNDA.n2452 GNDA.n2435 3.4105
R26067 GNDA.n2452 GNDA.n2415 3.4105
R26068 GNDA.n2452 GNDA.n2436 3.4105
R26069 GNDA.n2452 GNDA.n2414 3.4105
R26070 GNDA.n2452 GNDA.n2437 3.4105
R26071 GNDA.n2452 GNDA.n2413 3.4105
R26072 GNDA.n2452 GNDA.n2438 3.4105
R26073 GNDA.n2452 GNDA.n2412 3.4105
R26074 GNDA.n2452 GNDA.n2439 3.4105
R26075 GNDA.n2452 GNDA.n2411 3.4105
R26076 GNDA.n2452 GNDA.n2440 3.4105
R26077 GNDA.n2452 GNDA.n2410 3.4105
R26078 GNDA.n2452 GNDA.n2441 3.4105
R26079 GNDA.n2543 GNDA.n2452 3.4105
R26080 GNDA.n2540 GNDA.n2513 3.4105
R26081 GNDA.n2513 GNDA.n2426 3.4105
R26082 GNDA.n2513 GNDA.n2424 3.4105
R26083 GNDA.n2513 GNDA.n2427 3.4105
R26084 GNDA.n2513 GNDA.n2423 3.4105
R26085 GNDA.n2513 GNDA.n2428 3.4105
R26086 GNDA.n2513 GNDA.n2422 3.4105
R26087 GNDA.n2513 GNDA.n2429 3.4105
R26088 GNDA.n2513 GNDA.n2421 3.4105
R26089 GNDA.n2513 GNDA.n2430 3.4105
R26090 GNDA.n2513 GNDA.n2420 3.4105
R26091 GNDA.n2513 GNDA.n2431 3.4105
R26092 GNDA.n2513 GNDA.n2419 3.4105
R26093 GNDA.n2513 GNDA.n2432 3.4105
R26094 GNDA.n2513 GNDA.n2418 3.4105
R26095 GNDA.n2513 GNDA.n2433 3.4105
R26096 GNDA.n2513 GNDA.n2417 3.4105
R26097 GNDA.n2513 GNDA.n2434 3.4105
R26098 GNDA.n2513 GNDA.n2416 3.4105
R26099 GNDA.n2513 GNDA.n2435 3.4105
R26100 GNDA.n2513 GNDA.n2415 3.4105
R26101 GNDA.n2513 GNDA.n2436 3.4105
R26102 GNDA.n2513 GNDA.n2414 3.4105
R26103 GNDA.n2513 GNDA.n2437 3.4105
R26104 GNDA.n2513 GNDA.n2413 3.4105
R26105 GNDA.n2513 GNDA.n2438 3.4105
R26106 GNDA.n2513 GNDA.n2412 3.4105
R26107 GNDA.n2513 GNDA.n2439 3.4105
R26108 GNDA.n2513 GNDA.n2411 3.4105
R26109 GNDA.n2513 GNDA.n2440 3.4105
R26110 GNDA.n2513 GNDA.n2410 3.4105
R26111 GNDA.n2513 GNDA.n2441 3.4105
R26112 GNDA.n2543 GNDA.n2513 3.4105
R26113 GNDA.n2540 GNDA.n2451 3.4105
R26114 GNDA.n2451 GNDA.n2426 3.4105
R26115 GNDA.n2451 GNDA.n2424 3.4105
R26116 GNDA.n2451 GNDA.n2427 3.4105
R26117 GNDA.n2451 GNDA.n2423 3.4105
R26118 GNDA.n2451 GNDA.n2428 3.4105
R26119 GNDA.n2451 GNDA.n2422 3.4105
R26120 GNDA.n2451 GNDA.n2429 3.4105
R26121 GNDA.n2451 GNDA.n2421 3.4105
R26122 GNDA.n2451 GNDA.n2430 3.4105
R26123 GNDA.n2451 GNDA.n2420 3.4105
R26124 GNDA.n2451 GNDA.n2431 3.4105
R26125 GNDA.n2451 GNDA.n2419 3.4105
R26126 GNDA.n2451 GNDA.n2432 3.4105
R26127 GNDA.n2451 GNDA.n2418 3.4105
R26128 GNDA.n2451 GNDA.n2433 3.4105
R26129 GNDA.n2451 GNDA.n2417 3.4105
R26130 GNDA.n2451 GNDA.n2434 3.4105
R26131 GNDA.n2451 GNDA.n2416 3.4105
R26132 GNDA.n2451 GNDA.n2435 3.4105
R26133 GNDA.n2451 GNDA.n2415 3.4105
R26134 GNDA.n2451 GNDA.n2436 3.4105
R26135 GNDA.n2451 GNDA.n2414 3.4105
R26136 GNDA.n2451 GNDA.n2437 3.4105
R26137 GNDA.n2451 GNDA.n2413 3.4105
R26138 GNDA.n2451 GNDA.n2438 3.4105
R26139 GNDA.n2451 GNDA.n2412 3.4105
R26140 GNDA.n2451 GNDA.n2439 3.4105
R26141 GNDA.n2451 GNDA.n2411 3.4105
R26142 GNDA.n2451 GNDA.n2440 3.4105
R26143 GNDA.n2451 GNDA.n2410 3.4105
R26144 GNDA.n2451 GNDA.n2441 3.4105
R26145 GNDA.n2543 GNDA.n2451 3.4105
R26146 GNDA.n2540 GNDA.n2516 3.4105
R26147 GNDA.n2516 GNDA.n2426 3.4105
R26148 GNDA.n2516 GNDA.n2424 3.4105
R26149 GNDA.n2516 GNDA.n2427 3.4105
R26150 GNDA.n2516 GNDA.n2423 3.4105
R26151 GNDA.n2516 GNDA.n2428 3.4105
R26152 GNDA.n2516 GNDA.n2422 3.4105
R26153 GNDA.n2516 GNDA.n2429 3.4105
R26154 GNDA.n2516 GNDA.n2421 3.4105
R26155 GNDA.n2516 GNDA.n2430 3.4105
R26156 GNDA.n2516 GNDA.n2420 3.4105
R26157 GNDA.n2516 GNDA.n2431 3.4105
R26158 GNDA.n2516 GNDA.n2419 3.4105
R26159 GNDA.n2516 GNDA.n2432 3.4105
R26160 GNDA.n2516 GNDA.n2418 3.4105
R26161 GNDA.n2516 GNDA.n2433 3.4105
R26162 GNDA.n2516 GNDA.n2417 3.4105
R26163 GNDA.n2516 GNDA.n2434 3.4105
R26164 GNDA.n2516 GNDA.n2416 3.4105
R26165 GNDA.n2516 GNDA.n2435 3.4105
R26166 GNDA.n2516 GNDA.n2415 3.4105
R26167 GNDA.n2516 GNDA.n2436 3.4105
R26168 GNDA.n2516 GNDA.n2414 3.4105
R26169 GNDA.n2516 GNDA.n2437 3.4105
R26170 GNDA.n2516 GNDA.n2413 3.4105
R26171 GNDA.n2516 GNDA.n2438 3.4105
R26172 GNDA.n2516 GNDA.n2412 3.4105
R26173 GNDA.n2516 GNDA.n2439 3.4105
R26174 GNDA.n2516 GNDA.n2411 3.4105
R26175 GNDA.n2516 GNDA.n2440 3.4105
R26176 GNDA.n2516 GNDA.n2410 3.4105
R26177 GNDA.n2516 GNDA.n2441 3.4105
R26178 GNDA.n2543 GNDA.n2516 3.4105
R26179 GNDA.n2540 GNDA.n2450 3.4105
R26180 GNDA.n2450 GNDA.n2426 3.4105
R26181 GNDA.n2450 GNDA.n2424 3.4105
R26182 GNDA.n2450 GNDA.n2427 3.4105
R26183 GNDA.n2450 GNDA.n2423 3.4105
R26184 GNDA.n2450 GNDA.n2428 3.4105
R26185 GNDA.n2450 GNDA.n2422 3.4105
R26186 GNDA.n2450 GNDA.n2429 3.4105
R26187 GNDA.n2450 GNDA.n2421 3.4105
R26188 GNDA.n2450 GNDA.n2430 3.4105
R26189 GNDA.n2450 GNDA.n2420 3.4105
R26190 GNDA.n2450 GNDA.n2431 3.4105
R26191 GNDA.n2450 GNDA.n2419 3.4105
R26192 GNDA.n2450 GNDA.n2432 3.4105
R26193 GNDA.n2450 GNDA.n2418 3.4105
R26194 GNDA.n2450 GNDA.n2433 3.4105
R26195 GNDA.n2450 GNDA.n2417 3.4105
R26196 GNDA.n2450 GNDA.n2434 3.4105
R26197 GNDA.n2450 GNDA.n2416 3.4105
R26198 GNDA.n2450 GNDA.n2435 3.4105
R26199 GNDA.n2450 GNDA.n2415 3.4105
R26200 GNDA.n2450 GNDA.n2436 3.4105
R26201 GNDA.n2450 GNDA.n2414 3.4105
R26202 GNDA.n2450 GNDA.n2437 3.4105
R26203 GNDA.n2450 GNDA.n2413 3.4105
R26204 GNDA.n2450 GNDA.n2438 3.4105
R26205 GNDA.n2450 GNDA.n2412 3.4105
R26206 GNDA.n2450 GNDA.n2439 3.4105
R26207 GNDA.n2450 GNDA.n2411 3.4105
R26208 GNDA.n2450 GNDA.n2440 3.4105
R26209 GNDA.n2450 GNDA.n2410 3.4105
R26210 GNDA.n2450 GNDA.n2441 3.4105
R26211 GNDA.n2543 GNDA.n2450 3.4105
R26212 GNDA.n2540 GNDA.n2519 3.4105
R26213 GNDA.n2519 GNDA.n2426 3.4105
R26214 GNDA.n2519 GNDA.n2424 3.4105
R26215 GNDA.n2519 GNDA.n2427 3.4105
R26216 GNDA.n2519 GNDA.n2423 3.4105
R26217 GNDA.n2519 GNDA.n2428 3.4105
R26218 GNDA.n2519 GNDA.n2422 3.4105
R26219 GNDA.n2519 GNDA.n2429 3.4105
R26220 GNDA.n2519 GNDA.n2421 3.4105
R26221 GNDA.n2519 GNDA.n2430 3.4105
R26222 GNDA.n2519 GNDA.n2420 3.4105
R26223 GNDA.n2519 GNDA.n2431 3.4105
R26224 GNDA.n2519 GNDA.n2419 3.4105
R26225 GNDA.n2519 GNDA.n2432 3.4105
R26226 GNDA.n2519 GNDA.n2418 3.4105
R26227 GNDA.n2519 GNDA.n2433 3.4105
R26228 GNDA.n2519 GNDA.n2417 3.4105
R26229 GNDA.n2519 GNDA.n2434 3.4105
R26230 GNDA.n2519 GNDA.n2416 3.4105
R26231 GNDA.n2519 GNDA.n2435 3.4105
R26232 GNDA.n2519 GNDA.n2415 3.4105
R26233 GNDA.n2519 GNDA.n2436 3.4105
R26234 GNDA.n2519 GNDA.n2414 3.4105
R26235 GNDA.n2519 GNDA.n2437 3.4105
R26236 GNDA.n2519 GNDA.n2413 3.4105
R26237 GNDA.n2519 GNDA.n2438 3.4105
R26238 GNDA.n2519 GNDA.n2412 3.4105
R26239 GNDA.n2519 GNDA.n2439 3.4105
R26240 GNDA.n2519 GNDA.n2411 3.4105
R26241 GNDA.n2519 GNDA.n2440 3.4105
R26242 GNDA.n2519 GNDA.n2410 3.4105
R26243 GNDA.n2519 GNDA.n2441 3.4105
R26244 GNDA.n2543 GNDA.n2519 3.4105
R26245 GNDA.n2540 GNDA.n2449 3.4105
R26246 GNDA.n2449 GNDA.n2426 3.4105
R26247 GNDA.n2449 GNDA.n2424 3.4105
R26248 GNDA.n2449 GNDA.n2427 3.4105
R26249 GNDA.n2449 GNDA.n2423 3.4105
R26250 GNDA.n2449 GNDA.n2428 3.4105
R26251 GNDA.n2449 GNDA.n2422 3.4105
R26252 GNDA.n2449 GNDA.n2429 3.4105
R26253 GNDA.n2449 GNDA.n2421 3.4105
R26254 GNDA.n2449 GNDA.n2430 3.4105
R26255 GNDA.n2449 GNDA.n2420 3.4105
R26256 GNDA.n2449 GNDA.n2431 3.4105
R26257 GNDA.n2449 GNDA.n2419 3.4105
R26258 GNDA.n2449 GNDA.n2432 3.4105
R26259 GNDA.n2449 GNDA.n2418 3.4105
R26260 GNDA.n2449 GNDA.n2433 3.4105
R26261 GNDA.n2449 GNDA.n2417 3.4105
R26262 GNDA.n2449 GNDA.n2434 3.4105
R26263 GNDA.n2449 GNDA.n2416 3.4105
R26264 GNDA.n2449 GNDA.n2435 3.4105
R26265 GNDA.n2449 GNDA.n2415 3.4105
R26266 GNDA.n2449 GNDA.n2436 3.4105
R26267 GNDA.n2449 GNDA.n2414 3.4105
R26268 GNDA.n2449 GNDA.n2437 3.4105
R26269 GNDA.n2449 GNDA.n2413 3.4105
R26270 GNDA.n2449 GNDA.n2438 3.4105
R26271 GNDA.n2449 GNDA.n2412 3.4105
R26272 GNDA.n2449 GNDA.n2439 3.4105
R26273 GNDA.n2449 GNDA.n2411 3.4105
R26274 GNDA.n2449 GNDA.n2440 3.4105
R26275 GNDA.n2449 GNDA.n2410 3.4105
R26276 GNDA.n2449 GNDA.n2441 3.4105
R26277 GNDA.n2543 GNDA.n2449 3.4105
R26278 GNDA.n2540 GNDA.n2522 3.4105
R26279 GNDA.n2522 GNDA.n2426 3.4105
R26280 GNDA.n2522 GNDA.n2424 3.4105
R26281 GNDA.n2522 GNDA.n2427 3.4105
R26282 GNDA.n2522 GNDA.n2423 3.4105
R26283 GNDA.n2522 GNDA.n2428 3.4105
R26284 GNDA.n2522 GNDA.n2422 3.4105
R26285 GNDA.n2522 GNDA.n2429 3.4105
R26286 GNDA.n2522 GNDA.n2421 3.4105
R26287 GNDA.n2522 GNDA.n2430 3.4105
R26288 GNDA.n2522 GNDA.n2420 3.4105
R26289 GNDA.n2522 GNDA.n2431 3.4105
R26290 GNDA.n2522 GNDA.n2419 3.4105
R26291 GNDA.n2522 GNDA.n2432 3.4105
R26292 GNDA.n2522 GNDA.n2418 3.4105
R26293 GNDA.n2522 GNDA.n2433 3.4105
R26294 GNDA.n2522 GNDA.n2417 3.4105
R26295 GNDA.n2522 GNDA.n2434 3.4105
R26296 GNDA.n2522 GNDA.n2416 3.4105
R26297 GNDA.n2522 GNDA.n2435 3.4105
R26298 GNDA.n2522 GNDA.n2415 3.4105
R26299 GNDA.n2522 GNDA.n2436 3.4105
R26300 GNDA.n2522 GNDA.n2414 3.4105
R26301 GNDA.n2522 GNDA.n2437 3.4105
R26302 GNDA.n2522 GNDA.n2413 3.4105
R26303 GNDA.n2522 GNDA.n2438 3.4105
R26304 GNDA.n2522 GNDA.n2412 3.4105
R26305 GNDA.n2522 GNDA.n2439 3.4105
R26306 GNDA.n2522 GNDA.n2411 3.4105
R26307 GNDA.n2522 GNDA.n2440 3.4105
R26308 GNDA.n2522 GNDA.n2410 3.4105
R26309 GNDA.n2522 GNDA.n2441 3.4105
R26310 GNDA.n2543 GNDA.n2522 3.4105
R26311 GNDA.n2540 GNDA.n2448 3.4105
R26312 GNDA.n2448 GNDA.n2426 3.4105
R26313 GNDA.n2448 GNDA.n2424 3.4105
R26314 GNDA.n2448 GNDA.n2427 3.4105
R26315 GNDA.n2448 GNDA.n2423 3.4105
R26316 GNDA.n2448 GNDA.n2428 3.4105
R26317 GNDA.n2448 GNDA.n2422 3.4105
R26318 GNDA.n2448 GNDA.n2429 3.4105
R26319 GNDA.n2448 GNDA.n2421 3.4105
R26320 GNDA.n2448 GNDA.n2430 3.4105
R26321 GNDA.n2448 GNDA.n2420 3.4105
R26322 GNDA.n2448 GNDA.n2431 3.4105
R26323 GNDA.n2448 GNDA.n2419 3.4105
R26324 GNDA.n2448 GNDA.n2432 3.4105
R26325 GNDA.n2448 GNDA.n2418 3.4105
R26326 GNDA.n2448 GNDA.n2433 3.4105
R26327 GNDA.n2448 GNDA.n2417 3.4105
R26328 GNDA.n2448 GNDA.n2434 3.4105
R26329 GNDA.n2448 GNDA.n2416 3.4105
R26330 GNDA.n2448 GNDA.n2435 3.4105
R26331 GNDA.n2448 GNDA.n2415 3.4105
R26332 GNDA.n2448 GNDA.n2436 3.4105
R26333 GNDA.n2448 GNDA.n2414 3.4105
R26334 GNDA.n2448 GNDA.n2437 3.4105
R26335 GNDA.n2448 GNDA.n2413 3.4105
R26336 GNDA.n2448 GNDA.n2438 3.4105
R26337 GNDA.n2448 GNDA.n2412 3.4105
R26338 GNDA.n2448 GNDA.n2439 3.4105
R26339 GNDA.n2448 GNDA.n2411 3.4105
R26340 GNDA.n2448 GNDA.n2440 3.4105
R26341 GNDA.n2448 GNDA.n2410 3.4105
R26342 GNDA.n2448 GNDA.n2441 3.4105
R26343 GNDA.n2543 GNDA.n2448 3.4105
R26344 GNDA.n2540 GNDA.n2525 3.4105
R26345 GNDA.n2525 GNDA.n2426 3.4105
R26346 GNDA.n2525 GNDA.n2424 3.4105
R26347 GNDA.n2525 GNDA.n2427 3.4105
R26348 GNDA.n2525 GNDA.n2423 3.4105
R26349 GNDA.n2525 GNDA.n2428 3.4105
R26350 GNDA.n2525 GNDA.n2422 3.4105
R26351 GNDA.n2525 GNDA.n2429 3.4105
R26352 GNDA.n2525 GNDA.n2421 3.4105
R26353 GNDA.n2525 GNDA.n2430 3.4105
R26354 GNDA.n2525 GNDA.n2420 3.4105
R26355 GNDA.n2525 GNDA.n2431 3.4105
R26356 GNDA.n2525 GNDA.n2419 3.4105
R26357 GNDA.n2525 GNDA.n2432 3.4105
R26358 GNDA.n2525 GNDA.n2418 3.4105
R26359 GNDA.n2525 GNDA.n2433 3.4105
R26360 GNDA.n2525 GNDA.n2417 3.4105
R26361 GNDA.n2525 GNDA.n2434 3.4105
R26362 GNDA.n2525 GNDA.n2416 3.4105
R26363 GNDA.n2525 GNDA.n2435 3.4105
R26364 GNDA.n2525 GNDA.n2415 3.4105
R26365 GNDA.n2525 GNDA.n2436 3.4105
R26366 GNDA.n2525 GNDA.n2414 3.4105
R26367 GNDA.n2525 GNDA.n2437 3.4105
R26368 GNDA.n2525 GNDA.n2413 3.4105
R26369 GNDA.n2525 GNDA.n2438 3.4105
R26370 GNDA.n2525 GNDA.n2412 3.4105
R26371 GNDA.n2525 GNDA.n2439 3.4105
R26372 GNDA.n2525 GNDA.n2411 3.4105
R26373 GNDA.n2525 GNDA.n2440 3.4105
R26374 GNDA.n2525 GNDA.n2410 3.4105
R26375 GNDA.n2525 GNDA.n2441 3.4105
R26376 GNDA.n2543 GNDA.n2525 3.4105
R26377 GNDA.n2540 GNDA.n2447 3.4105
R26378 GNDA.n2447 GNDA.n2426 3.4105
R26379 GNDA.n2447 GNDA.n2424 3.4105
R26380 GNDA.n2447 GNDA.n2427 3.4105
R26381 GNDA.n2447 GNDA.n2423 3.4105
R26382 GNDA.n2447 GNDA.n2428 3.4105
R26383 GNDA.n2447 GNDA.n2422 3.4105
R26384 GNDA.n2447 GNDA.n2429 3.4105
R26385 GNDA.n2447 GNDA.n2421 3.4105
R26386 GNDA.n2447 GNDA.n2430 3.4105
R26387 GNDA.n2447 GNDA.n2420 3.4105
R26388 GNDA.n2447 GNDA.n2431 3.4105
R26389 GNDA.n2447 GNDA.n2419 3.4105
R26390 GNDA.n2447 GNDA.n2432 3.4105
R26391 GNDA.n2447 GNDA.n2418 3.4105
R26392 GNDA.n2447 GNDA.n2433 3.4105
R26393 GNDA.n2447 GNDA.n2417 3.4105
R26394 GNDA.n2447 GNDA.n2434 3.4105
R26395 GNDA.n2447 GNDA.n2416 3.4105
R26396 GNDA.n2447 GNDA.n2435 3.4105
R26397 GNDA.n2447 GNDA.n2415 3.4105
R26398 GNDA.n2447 GNDA.n2436 3.4105
R26399 GNDA.n2447 GNDA.n2414 3.4105
R26400 GNDA.n2447 GNDA.n2437 3.4105
R26401 GNDA.n2447 GNDA.n2413 3.4105
R26402 GNDA.n2447 GNDA.n2438 3.4105
R26403 GNDA.n2447 GNDA.n2412 3.4105
R26404 GNDA.n2447 GNDA.n2439 3.4105
R26405 GNDA.n2447 GNDA.n2411 3.4105
R26406 GNDA.n2447 GNDA.n2440 3.4105
R26407 GNDA.n2447 GNDA.n2410 3.4105
R26408 GNDA.n2447 GNDA.n2441 3.4105
R26409 GNDA.n2543 GNDA.n2447 3.4105
R26410 GNDA.n2540 GNDA.n2528 3.4105
R26411 GNDA.n2528 GNDA.n2426 3.4105
R26412 GNDA.n2528 GNDA.n2424 3.4105
R26413 GNDA.n2528 GNDA.n2427 3.4105
R26414 GNDA.n2528 GNDA.n2423 3.4105
R26415 GNDA.n2528 GNDA.n2428 3.4105
R26416 GNDA.n2528 GNDA.n2422 3.4105
R26417 GNDA.n2528 GNDA.n2429 3.4105
R26418 GNDA.n2528 GNDA.n2421 3.4105
R26419 GNDA.n2528 GNDA.n2430 3.4105
R26420 GNDA.n2528 GNDA.n2420 3.4105
R26421 GNDA.n2528 GNDA.n2431 3.4105
R26422 GNDA.n2528 GNDA.n2419 3.4105
R26423 GNDA.n2528 GNDA.n2432 3.4105
R26424 GNDA.n2528 GNDA.n2418 3.4105
R26425 GNDA.n2528 GNDA.n2433 3.4105
R26426 GNDA.n2528 GNDA.n2417 3.4105
R26427 GNDA.n2528 GNDA.n2434 3.4105
R26428 GNDA.n2528 GNDA.n2416 3.4105
R26429 GNDA.n2528 GNDA.n2435 3.4105
R26430 GNDA.n2528 GNDA.n2415 3.4105
R26431 GNDA.n2528 GNDA.n2436 3.4105
R26432 GNDA.n2528 GNDA.n2414 3.4105
R26433 GNDA.n2528 GNDA.n2437 3.4105
R26434 GNDA.n2528 GNDA.n2413 3.4105
R26435 GNDA.n2528 GNDA.n2438 3.4105
R26436 GNDA.n2528 GNDA.n2412 3.4105
R26437 GNDA.n2528 GNDA.n2439 3.4105
R26438 GNDA.n2528 GNDA.n2411 3.4105
R26439 GNDA.n2528 GNDA.n2440 3.4105
R26440 GNDA.n2528 GNDA.n2410 3.4105
R26441 GNDA.n2528 GNDA.n2441 3.4105
R26442 GNDA.n2543 GNDA.n2528 3.4105
R26443 GNDA.n2540 GNDA.n2446 3.4105
R26444 GNDA.n2446 GNDA.n2426 3.4105
R26445 GNDA.n2446 GNDA.n2424 3.4105
R26446 GNDA.n2446 GNDA.n2427 3.4105
R26447 GNDA.n2446 GNDA.n2423 3.4105
R26448 GNDA.n2446 GNDA.n2428 3.4105
R26449 GNDA.n2446 GNDA.n2422 3.4105
R26450 GNDA.n2446 GNDA.n2429 3.4105
R26451 GNDA.n2446 GNDA.n2421 3.4105
R26452 GNDA.n2446 GNDA.n2430 3.4105
R26453 GNDA.n2446 GNDA.n2420 3.4105
R26454 GNDA.n2446 GNDA.n2431 3.4105
R26455 GNDA.n2446 GNDA.n2419 3.4105
R26456 GNDA.n2446 GNDA.n2432 3.4105
R26457 GNDA.n2446 GNDA.n2418 3.4105
R26458 GNDA.n2446 GNDA.n2433 3.4105
R26459 GNDA.n2446 GNDA.n2417 3.4105
R26460 GNDA.n2446 GNDA.n2434 3.4105
R26461 GNDA.n2446 GNDA.n2416 3.4105
R26462 GNDA.n2446 GNDA.n2435 3.4105
R26463 GNDA.n2446 GNDA.n2415 3.4105
R26464 GNDA.n2446 GNDA.n2436 3.4105
R26465 GNDA.n2446 GNDA.n2414 3.4105
R26466 GNDA.n2446 GNDA.n2437 3.4105
R26467 GNDA.n2446 GNDA.n2413 3.4105
R26468 GNDA.n2446 GNDA.n2438 3.4105
R26469 GNDA.n2446 GNDA.n2412 3.4105
R26470 GNDA.n2446 GNDA.n2439 3.4105
R26471 GNDA.n2446 GNDA.n2411 3.4105
R26472 GNDA.n2446 GNDA.n2440 3.4105
R26473 GNDA.n2446 GNDA.n2410 3.4105
R26474 GNDA.n2446 GNDA.n2441 3.4105
R26475 GNDA.n2543 GNDA.n2446 3.4105
R26476 GNDA.n2540 GNDA.n2531 3.4105
R26477 GNDA.n2531 GNDA.n2426 3.4105
R26478 GNDA.n2531 GNDA.n2424 3.4105
R26479 GNDA.n2531 GNDA.n2427 3.4105
R26480 GNDA.n2531 GNDA.n2423 3.4105
R26481 GNDA.n2531 GNDA.n2428 3.4105
R26482 GNDA.n2531 GNDA.n2422 3.4105
R26483 GNDA.n2531 GNDA.n2429 3.4105
R26484 GNDA.n2531 GNDA.n2421 3.4105
R26485 GNDA.n2531 GNDA.n2430 3.4105
R26486 GNDA.n2531 GNDA.n2420 3.4105
R26487 GNDA.n2531 GNDA.n2431 3.4105
R26488 GNDA.n2531 GNDA.n2419 3.4105
R26489 GNDA.n2531 GNDA.n2432 3.4105
R26490 GNDA.n2531 GNDA.n2418 3.4105
R26491 GNDA.n2531 GNDA.n2433 3.4105
R26492 GNDA.n2531 GNDA.n2417 3.4105
R26493 GNDA.n2531 GNDA.n2434 3.4105
R26494 GNDA.n2531 GNDA.n2416 3.4105
R26495 GNDA.n2531 GNDA.n2435 3.4105
R26496 GNDA.n2531 GNDA.n2415 3.4105
R26497 GNDA.n2531 GNDA.n2436 3.4105
R26498 GNDA.n2531 GNDA.n2414 3.4105
R26499 GNDA.n2531 GNDA.n2437 3.4105
R26500 GNDA.n2531 GNDA.n2413 3.4105
R26501 GNDA.n2531 GNDA.n2438 3.4105
R26502 GNDA.n2531 GNDA.n2412 3.4105
R26503 GNDA.n2531 GNDA.n2439 3.4105
R26504 GNDA.n2531 GNDA.n2411 3.4105
R26505 GNDA.n2531 GNDA.n2440 3.4105
R26506 GNDA.n2531 GNDA.n2410 3.4105
R26507 GNDA.n2531 GNDA.n2441 3.4105
R26508 GNDA.n2543 GNDA.n2531 3.4105
R26509 GNDA.n2540 GNDA.n2445 3.4105
R26510 GNDA.n2445 GNDA.n2426 3.4105
R26511 GNDA.n2445 GNDA.n2424 3.4105
R26512 GNDA.n2445 GNDA.n2427 3.4105
R26513 GNDA.n2445 GNDA.n2423 3.4105
R26514 GNDA.n2445 GNDA.n2428 3.4105
R26515 GNDA.n2445 GNDA.n2422 3.4105
R26516 GNDA.n2445 GNDA.n2429 3.4105
R26517 GNDA.n2445 GNDA.n2421 3.4105
R26518 GNDA.n2445 GNDA.n2430 3.4105
R26519 GNDA.n2445 GNDA.n2420 3.4105
R26520 GNDA.n2445 GNDA.n2431 3.4105
R26521 GNDA.n2445 GNDA.n2419 3.4105
R26522 GNDA.n2445 GNDA.n2432 3.4105
R26523 GNDA.n2445 GNDA.n2418 3.4105
R26524 GNDA.n2445 GNDA.n2433 3.4105
R26525 GNDA.n2445 GNDA.n2417 3.4105
R26526 GNDA.n2445 GNDA.n2434 3.4105
R26527 GNDA.n2445 GNDA.n2416 3.4105
R26528 GNDA.n2445 GNDA.n2435 3.4105
R26529 GNDA.n2445 GNDA.n2415 3.4105
R26530 GNDA.n2445 GNDA.n2436 3.4105
R26531 GNDA.n2445 GNDA.n2414 3.4105
R26532 GNDA.n2445 GNDA.n2437 3.4105
R26533 GNDA.n2445 GNDA.n2413 3.4105
R26534 GNDA.n2445 GNDA.n2438 3.4105
R26535 GNDA.n2445 GNDA.n2412 3.4105
R26536 GNDA.n2445 GNDA.n2439 3.4105
R26537 GNDA.n2445 GNDA.n2411 3.4105
R26538 GNDA.n2445 GNDA.n2440 3.4105
R26539 GNDA.n2445 GNDA.n2410 3.4105
R26540 GNDA.n2445 GNDA.n2441 3.4105
R26541 GNDA.n2543 GNDA.n2445 3.4105
R26542 GNDA.n2540 GNDA.n2534 3.4105
R26543 GNDA.n2534 GNDA.n2426 3.4105
R26544 GNDA.n2534 GNDA.n2424 3.4105
R26545 GNDA.n2534 GNDA.n2427 3.4105
R26546 GNDA.n2534 GNDA.n2423 3.4105
R26547 GNDA.n2534 GNDA.n2428 3.4105
R26548 GNDA.n2534 GNDA.n2422 3.4105
R26549 GNDA.n2534 GNDA.n2429 3.4105
R26550 GNDA.n2534 GNDA.n2421 3.4105
R26551 GNDA.n2534 GNDA.n2430 3.4105
R26552 GNDA.n2534 GNDA.n2420 3.4105
R26553 GNDA.n2534 GNDA.n2431 3.4105
R26554 GNDA.n2534 GNDA.n2419 3.4105
R26555 GNDA.n2534 GNDA.n2432 3.4105
R26556 GNDA.n2534 GNDA.n2418 3.4105
R26557 GNDA.n2534 GNDA.n2433 3.4105
R26558 GNDA.n2534 GNDA.n2417 3.4105
R26559 GNDA.n2534 GNDA.n2434 3.4105
R26560 GNDA.n2534 GNDA.n2416 3.4105
R26561 GNDA.n2534 GNDA.n2435 3.4105
R26562 GNDA.n2534 GNDA.n2415 3.4105
R26563 GNDA.n2534 GNDA.n2436 3.4105
R26564 GNDA.n2534 GNDA.n2414 3.4105
R26565 GNDA.n2534 GNDA.n2437 3.4105
R26566 GNDA.n2534 GNDA.n2413 3.4105
R26567 GNDA.n2534 GNDA.n2438 3.4105
R26568 GNDA.n2534 GNDA.n2412 3.4105
R26569 GNDA.n2534 GNDA.n2439 3.4105
R26570 GNDA.n2534 GNDA.n2411 3.4105
R26571 GNDA.n2534 GNDA.n2440 3.4105
R26572 GNDA.n2534 GNDA.n2410 3.4105
R26573 GNDA.n2534 GNDA.n2441 3.4105
R26574 GNDA.n2543 GNDA.n2534 3.4105
R26575 GNDA.n2540 GNDA.n2444 3.4105
R26576 GNDA.n2444 GNDA.n2426 3.4105
R26577 GNDA.n2444 GNDA.n2424 3.4105
R26578 GNDA.n2444 GNDA.n2427 3.4105
R26579 GNDA.n2444 GNDA.n2423 3.4105
R26580 GNDA.n2444 GNDA.n2428 3.4105
R26581 GNDA.n2444 GNDA.n2422 3.4105
R26582 GNDA.n2444 GNDA.n2429 3.4105
R26583 GNDA.n2444 GNDA.n2421 3.4105
R26584 GNDA.n2444 GNDA.n2430 3.4105
R26585 GNDA.n2444 GNDA.n2420 3.4105
R26586 GNDA.n2444 GNDA.n2431 3.4105
R26587 GNDA.n2444 GNDA.n2419 3.4105
R26588 GNDA.n2444 GNDA.n2432 3.4105
R26589 GNDA.n2444 GNDA.n2418 3.4105
R26590 GNDA.n2444 GNDA.n2433 3.4105
R26591 GNDA.n2444 GNDA.n2417 3.4105
R26592 GNDA.n2444 GNDA.n2434 3.4105
R26593 GNDA.n2444 GNDA.n2416 3.4105
R26594 GNDA.n2444 GNDA.n2435 3.4105
R26595 GNDA.n2444 GNDA.n2415 3.4105
R26596 GNDA.n2444 GNDA.n2436 3.4105
R26597 GNDA.n2444 GNDA.n2414 3.4105
R26598 GNDA.n2444 GNDA.n2437 3.4105
R26599 GNDA.n2444 GNDA.n2413 3.4105
R26600 GNDA.n2444 GNDA.n2438 3.4105
R26601 GNDA.n2444 GNDA.n2412 3.4105
R26602 GNDA.n2444 GNDA.n2439 3.4105
R26603 GNDA.n2444 GNDA.n2411 3.4105
R26604 GNDA.n2444 GNDA.n2440 3.4105
R26605 GNDA.n2444 GNDA.n2410 3.4105
R26606 GNDA.n2444 GNDA.n2441 3.4105
R26607 GNDA.n2543 GNDA.n2444 3.4105
R26608 GNDA.n2540 GNDA.n2537 3.4105
R26609 GNDA.n2537 GNDA.n2426 3.4105
R26610 GNDA.n2537 GNDA.n2424 3.4105
R26611 GNDA.n2537 GNDA.n2427 3.4105
R26612 GNDA.n2537 GNDA.n2423 3.4105
R26613 GNDA.n2537 GNDA.n2428 3.4105
R26614 GNDA.n2537 GNDA.n2422 3.4105
R26615 GNDA.n2537 GNDA.n2429 3.4105
R26616 GNDA.n2537 GNDA.n2421 3.4105
R26617 GNDA.n2537 GNDA.n2430 3.4105
R26618 GNDA.n2537 GNDA.n2420 3.4105
R26619 GNDA.n2537 GNDA.n2431 3.4105
R26620 GNDA.n2537 GNDA.n2419 3.4105
R26621 GNDA.n2537 GNDA.n2432 3.4105
R26622 GNDA.n2537 GNDA.n2418 3.4105
R26623 GNDA.n2537 GNDA.n2433 3.4105
R26624 GNDA.n2537 GNDA.n2417 3.4105
R26625 GNDA.n2537 GNDA.n2434 3.4105
R26626 GNDA.n2537 GNDA.n2416 3.4105
R26627 GNDA.n2537 GNDA.n2435 3.4105
R26628 GNDA.n2537 GNDA.n2415 3.4105
R26629 GNDA.n2537 GNDA.n2436 3.4105
R26630 GNDA.n2537 GNDA.n2414 3.4105
R26631 GNDA.n2537 GNDA.n2437 3.4105
R26632 GNDA.n2537 GNDA.n2413 3.4105
R26633 GNDA.n2537 GNDA.n2438 3.4105
R26634 GNDA.n2537 GNDA.n2412 3.4105
R26635 GNDA.n2537 GNDA.n2439 3.4105
R26636 GNDA.n2537 GNDA.n2411 3.4105
R26637 GNDA.n2537 GNDA.n2440 3.4105
R26638 GNDA.n2537 GNDA.n2410 3.4105
R26639 GNDA.n2537 GNDA.n2441 3.4105
R26640 GNDA.n2543 GNDA.n2537 3.4105
R26641 GNDA.n2540 GNDA.n2443 3.4105
R26642 GNDA.n2443 GNDA.n2426 3.4105
R26643 GNDA.n2443 GNDA.n2424 3.4105
R26644 GNDA.n2443 GNDA.n2427 3.4105
R26645 GNDA.n2443 GNDA.n2423 3.4105
R26646 GNDA.n2443 GNDA.n2428 3.4105
R26647 GNDA.n2443 GNDA.n2422 3.4105
R26648 GNDA.n2443 GNDA.n2429 3.4105
R26649 GNDA.n2443 GNDA.n2421 3.4105
R26650 GNDA.n2443 GNDA.n2430 3.4105
R26651 GNDA.n2443 GNDA.n2420 3.4105
R26652 GNDA.n2443 GNDA.n2431 3.4105
R26653 GNDA.n2443 GNDA.n2419 3.4105
R26654 GNDA.n2443 GNDA.n2432 3.4105
R26655 GNDA.n2443 GNDA.n2418 3.4105
R26656 GNDA.n2443 GNDA.n2433 3.4105
R26657 GNDA.n2443 GNDA.n2417 3.4105
R26658 GNDA.n2443 GNDA.n2434 3.4105
R26659 GNDA.n2443 GNDA.n2416 3.4105
R26660 GNDA.n2443 GNDA.n2435 3.4105
R26661 GNDA.n2443 GNDA.n2415 3.4105
R26662 GNDA.n2443 GNDA.n2436 3.4105
R26663 GNDA.n2443 GNDA.n2414 3.4105
R26664 GNDA.n2443 GNDA.n2437 3.4105
R26665 GNDA.n2443 GNDA.n2413 3.4105
R26666 GNDA.n2443 GNDA.n2438 3.4105
R26667 GNDA.n2443 GNDA.n2412 3.4105
R26668 GNDA.n2443 GNDA.n2439 3.4105
R26669 GNDA.n2443 GNDA.n2411 3.4105
R26670 GNDA.n2443 GNDA.n2440 3.4105
R26671 GNDA.n2443 GNDA.n2410 3.4105
R26672 GNDA.n2443 GNDA.n2441 3.4105
R26673 GNDA.n2543 GNDA.n2443 3.4105
R26674 GNDA.n2542 GNDA.n2540 3.4105
R26675 GNDA.n2542 GNDA.n2426 3.4105
R26676 GNDA.n2542 GNDA.n2424 3.4105
R26677 GNDA.n2542 GNDA.n2427 3.4105
R26678 GNDA.n2542 GNDA.n2423 3.4105
R26679 GNDA.n2542 GNDA.n2428 3.4105
R26680 GNDA.n2542 GNDA.n2422 3.4105
R26681 GNDA.n2542 GNDA.n2429 3.4105
R26682 GNDA.n2542 GNDA.n2421 3.4105
R26683 GNDA.n2542 GNDA.n2430 3.4105
R26684 GNDA.n2542 GNDA.n2420 3.4105
R26685 GNDA.n2542 GNDA.n2431 3.4105
R26686 GNDA.n2542 GNDA.n2419 3.4105
R26687 GNDA.n2542 GNDA.n2432 3.4105
R26688 GNDA.n2542 GNDA.n2418 3.4105
R26689 GNDA.n2542 GNDA.n2433 3.4105
R26690 GNDA.n2542 GNDA.n2417 3.4105
R26691 GNDA.n2542 GNDA.n2434 3.4105
R26692 GNDA.n2542 GNDA.n2416 3.4105
R26693 GNDA.n2542 GNDA.n2435 3.4105
R26694 GNDA.n2542 GNDA.n2415 3.4105
R26695 GNDA.n2542 GNDA.n2436 3.4105
R26696 GNDA.n2542 GNDA.n2414 3.4105
R26697 GNDA.n2542 GNDA.n2437 3.4105
R26698 GNDA.n2542 GNDA.n2413 3.4105
R26699 GNDA.n2542 GNDA.n2438 3.4105
R26700 GNDA.n2542 GNDA.n2412 3.4105
R26701 GNDA.n2542 GNDA.n2439 3.4105
R26702 GNDA.n2542 GNDA.n2411 3.4105
R26703 GNDA.n2542 GNDA.n2440 3.4105
R26704 GNDA.n2542 GNDA.n2410 3.4105
R26705 GNDA.n2542 GNDA.n2441 3.4105
R26706 GNDA.n2543 GNDA.n2542 3.4105
R26707 GNDA.n2540 GNDA.n2442 3.4105
R26708 GNDA.n2442 GNDA.n2426 3.4105
R26709 GNDA.n2442 GNDA.n2424 3.4105
R26710 GNDA.n2442 GNDA.n2427 3.4105
R26711 GNDA.n2442 GNDA.n2423 3.4105
R26712 GNDA.n2442 GNDA.n2428 3.4105
R26713 GNDA.n2442 GNDA.n2422 3.4105
R26714 GNDA.n2442 GNDA.n2429 3.4105
R26715 GNDA.n2442 GNDA.n2421 3.4105
R26716 GNDA.n2442 GNDA.n2430 3.4105
R26717 GNDA.n2442 GNDA.n2420 3.4105
R26718 GNDA.n2442 GNDA.n2431 3.4105
R26719 GNDA.n2442 GNDA.n2419 3.4105
R26720 GNDA.n2442 GNDA.n2432 3.4105
R26721 GNDA.n2442 GNDA.n2418 3.4105
R26722 GNDA.n2442 GNDA.n2433 3.4105
R26723 GNDA.n2442 GNDA.n2417 3.4105
R26724 GNDA.n2442 GNDA.n2434 3.4105
R26725 GNDA.n2442 GNDA.n2416 3.4105
R26726 GNDA.n2442 GNDA.n2435 3.4105
R26727 GNDA.n2442 GNDA.n2415 3.4105
R26728 GNDA.n2442 GNDA.n2436 3.4105
R26729 GNDA.n2442 GNDA.n2414 3.4105
R26730 GNDA.n2442 GNDA.n2437 3.4105
R26731 GNDA.n2442 GNDA.n2413 3.4105
R26732 GNDA.n2442 GNDA.n2438 3.4105
R26733 GNDA.n2442 GNDA.n2412 3.4105
R26734 GNDA.n2442 GNDA.n2439 3.4105
R26735 GNDA.n2442 GNDA.n2411 3.4105
R26736 GNDA.n2442 GNDA.n2440 3.4105
R26737 GNDA.n2442 GNDA.n2410 3.4105
R26738 GNDA.n2442 GNDA.n2441 3.4105
R26739 GNDA.n2543 GNDA.n2442 3.4105
R26740 GNDA.n2544 GNDA.n2426 3.4105
R26741 GNDA.n2544 GNDA.n2424 3.4105
R26742 GNDA.n2544 GNDA.n2427 3.4105
R26743 GNDA.n2544 GNDA.n2423 3.4105
R26744 GNDA.n2544 GNDA.n2428 3.4105
R26745 GNDA.n2544 GNDA.n2422 3.4105
R26746 GNDA.n2544 GNDA.n2429 3.4105
R26747 GNDA.n2544 GNDA.n2421 3.4105
R26748 GNDA.n2544 GNDA.n2430 3.4105
R26749 GNDA.n2544 GNDA.n2420 3.4105
R26750 GNDA.n2544 GNDA.n2431 3.4105
R26751 GNDA.n2544 GNDA.n2419 3.4105
R26752 GNDA.n2544 GNDA.n2432 3.4105
R26753 GNDA.n2544 GNDA.n2418 3.4105
R26754 GNDA.n2544 GNDA.n2433 3.4105
R26755 GNDA.n2544 GNDA.n2417 3.4105
R26756 GNDA.n2544 GNDA.n2434 3.4105
R26757 GNDA.n2544 GNDA.n2416 3.4105
R26758 GNDA.n2544 GNDA.n2435 3.4105
R26759 GNDA.n2544 GNDA.n2415 3.4105
R26760 GNDA.n2544 GNDA.n2436 3.4105
R26761 GNDA.n2544 GNDA.n2414 3.4105
R26762 GNDA.n2544 GNDA.n2437 3.4105
R26763 GNDA.n2544 GNDA.n2413 3.4105
R26764 GNDA.n2544 GNDA.n2438 3.4105
R26765 GNDA.n2544 GNDA.n2412 3.4105
R26766 GNDA.n2544 GNDA.n2439 3.4105
R26767 GNDA.n2544 GNDA.n2411 3.4105
R26768 GNDA.n2544 GNDA.n2440 3.4105
R26769 GNDA.n2544 GNDA.n2410 3.4105
R26770 GNDA.n2544 GNDA.n2441 3.4105
R26771 GNDA.n2544 GNDA.n2543 3.4105
R26772 GNDA.n2650 GNDA.n2649 3.4105
R26773 GNDA.n2651 GNDA.n2650 3.4105
R26774 GNDA.n2653 GNDA.n2261 3.4105
R26775 GNDA.n2649 GNDA.n2261 3.4105
R26776 GNDA.n2651 GNDA.n2261 3.4105
R26777 GNDA.n2653 GNDA.n2263 3.4105
R26778 GNDA.n2294 GNDA.n2263 3.4105
R26779 GNDA.n2296 GNDA.n2263 3.4105
R26780 GNDA.n2293 GNDA.n2263 3.4105
R26781 GNDA.n2298 GNDA.n2263 3.4105
R26782 GNDA.n2292 GNDA.n2263 3.4105
R26783 GNDA.n2300 GNDA.n2263 3.4105
R26784 GNDA.n2291 GNDA.n2263 3.4105
R26785 GNDA.n2302 GNDA.n2263 3.4105
R26786 GNDA.n2290 GNDA.n2263 3.4105
R26787 GNDA.n2304 GNDA.n2263 3.4105
R26788 GNDA.n2289 GNDA.n2263 3.4105
R26789 GNDA.n2306 GNDA.n2263 3.4105
R26790 GNDA.n2288 GNDA.n2263 3.4105
R26791 GNDA.n2308 GNDA.n2263 3.4105
R26792 GNDA.n2287 GNDA.n2263 3.4105
R26793 GNDA.n2310 GNDA.n2263 3.4105
R26794 GNDA.n2286 GNDA.n2263 3.4105
R26795 GNDA.n2312 GNDA.n2263 3.4105
R26796 GNDA.n2285 GNDA.n2263 3.4105
R26797 GNDA.n2314 GNDA.n2263 3.4105
R26798 GNDA.n2284 GNDA.n2263 3.4105
R26799 GNDA.n2316 GNDA.n2263 3.4105
R26800 GNDA.n2283 GNDA.n2263 3.4105
R26801 GNDA.n2318 GNDA.n2263 3.4105
R26802 GNDA.n2282 GNDA.n2263 3.4105
R26803 GNDA.n2320 GNDA.n2263 3.4105
R26804 GNDA.n2281 GNDA.n2263 3.4105
R26805 GNDA.n2322 GNDA.n2263 3.4105
R26806 GNDA.n2280 GNDA.n2263 3.4105
R26807 GNDA.n2324 GNDA.n2263 3.4105
R26808 GNDA.n2649 GNDA.n2263 3.4105
R26809 GNDA.n2651 GNDA.n2263 3.4105
R26810 GNDA.n2653 GNDA.n2260 3.4105
R26811 GNDA.n2294 GNDA.n2260 3.4105
R26812 GNDA.n2296 GNDA.n2260 3.4105
R26813 GNDA.n2293 GNDA.n2260 3.4105
R26814 GNDA.n2298 GNDA.n2260 3.4105
R26815 GNDA.n2292 GNDA.n2260 3.4105
R26816 GNDA.n2300 GNDA.n2260 3.4105
R26817 GNDA.n2291 GNDA.n2260 3.4105
R26818 GNDA.n2302 GNDA.n2260 3.4105
R26819 GNDA.n2290 GNDA.n2260 3.4105
R26820 GNDA.n2304 GNDA.n2260 3.4105
R26821 GNDA.n2289 GNDA.n2260 3.4105
R26822 GNDA.n2306 GNDA.n2260 3.4105
R26823 GNDA.n2288 GNDA.n2260 3.4105
R26824 GNDA.n2308 GNDA.n2260 3.4105
R26825 GNDA.n2287 GNDA.n2260 3.4105
R26826 GNDA.n2310 GNDA.n2260 3.4105
R26827 GNDA.n2286 GNDA.n2260 3.4105
R26828 GNDA.n2312 GNDA.n2260 3.4105
R26829 GNDA.n2285 GNDA.n2260 3.4105
R26830 GNDA.n2314 GNDA.n2260 3.4105
R26831 GNDA.n2284 GNDA.n2260 3.4105
R26832 GNDA.n2316 GNDA.n2260 3.4105
R26833 GNDA.n2283 GNDA.n2260 3.4105
R26834 GNDA.n2318 GNDA.n2260 3.4105
R26835 GNDA.n2282 GNDA.n2260 3.4105
R26836 GNDA.n2320 GNDA.n2260 3.4105
R26837 GNDA.n2281 GNDA.n2260 3.4105
R26838 GNDA.n2322 GNDA.n2260 3.4105
R26839 GNDA.n2280 GNDA.n2260 3.4105
R26840 GNDA.n2324 GNDA.n2260 3.4105
R26841 GNDA.n2649 GNDA.n2260 3.4105
R26842 GNDA.n2651 GNDA.n2260 3.4105
R26843 GNDA.n2653 GNDA.n2264 3.4105
R26844 GNDA.n2294 GNDA.n2264 3.4105
R26845 GNDA.n2296 GNDA.n2264 3.4105
R26846 GNDA.n2293 GNDA.n2264 3.4105
R26847 GNDA.n2298 GNDA.n2264 3.4105
R26848 GNDA.n2292 GNDA.n2264 3.4105
R26849 GNDA.n2300 GNDA.n2264 3.4105
R26850 GNDA.n2291 GNDA.n2264 3.4105
R26851 GNDA.n2302 GNDA.n2264 3.4105
R26852 GNDA.n2290 GNDA.n2264 3.4105
R26853 GNDA.n2304 GNDA.n2264 3.4105
R26854 GNDA.n2289 GNDA.n2264 3.4105
R26855 GNDA.n2306 GNDA.n2264 3.4105
R26856 GNDA.n2288 GNDA.n2264 3.4105
R26857 GNDA.n2308 GNDA.n2264 3.4105
R26858 GNDA.n2287 GNDA.n2264 3.4105
R26859 GNDA.n2310 GNDA.n2264 3.4105
R26860 GNDA.n2286 GNDA.n2264 3.4105
R26861 GNDA.n2312 GNDA.n2264 3.4105
R26862 GNDA.n2285 GNDA.n2264 3.4105
R26863 GNDA.n2314 GNDA.n2264 3.4105
R26864 GNDA.n2284 GNDA.n2264 3.4105
R26865 GNDA.n2316 GNDA.n2264 3.4105
R26866 GNDA.n2283 GNDA.n2264 3.4105
R26867 GNDA.n2318 GNDA.n2264 3.4105
R26868 GNDA.n2282 GNDA.n2264 3.4105
R26869 GNDA.n2320 GNDA.n2264 3.4105
R26870 GNDA.n2281 GNDA.n2264 3.4105
R26871 GNDA.n2322 GNDA.n2264 3.4105
R26872 GNDA.n2280 GNDA.n2264 3.4105
R26873 GNDA.n2324 GNDA.n2264 3.4105
R26874 GNDA.n2649 GNDA.n2264 3.4105
R26875 GNDA.n2651 GNDA.n2264 3.4105
R26876 GNDA.n2653 GNDA.n2259 3.4105
R26877 GNDA.n2294 GNDA.n2259 3.4105
R26878 GNDA.n2296 GNDA.n2259 3.4105
R26879 GNDA.n2293 GNDA.n2259 3.4105
R26880 GNDA.n2298 GNDA.n2259 3.4105
R26881 GNDA.n2292 GNDA.n2259 3.4105
R26882 GNDA.n2300 GNDA.n2259 3.4105
R26883 GNDA.n2291 GNDA.n2259 3.4105
R26884 GNDA.n2302 GNDA.n2259 3.4105
R26885 GNDA.n2290 GNDA.n2259 3.4105
R26886 GNDA.n2304 GNDA.n2259 3.4105
R26887 GNDA.n2289 GNDA.n2259 3.4105
R26888 GNDA.n2306 GNDA.n2259 3.4105
R26889 GNDA.n2288 GNDA.n2259 3.4105
R26890 GNDA.n2308 GNDA.n2259 3.4105
R26891 GNDA.n2287 GNDA.n2259 3.4105
R26892 GNDA.n2310 GNDA.n2259 3.4105
R26893 GNDA.n2286 GNDA.n2259 3.4105
R26894 GNDA.n2312 GNDA.n2259 3.4105
R26895 GNDA.n2285 GNDA.n2259 3.4105
R26896 GNDA.n2314 GNDA.n2259 3.4105
R26897 GNDA.n2284 GNDA.n2259 3.4105
R26898 GNDA.n2316 GNDA.n2259 3.4105
R26899 GNDA.n2283 GNDA.n2259 3.4105
R26900 GNDA.n2318 GNDA.n2259 3.4105
R26901 GNDA.n2282 GNDA.n2259 3.4105
R26902 GNDA.n2320 GNDA.n2259 3.4105
R26903 GNDA.n2281 GNDA.n2259 3.4105
R26904 GNDA.n2322 GNDA.n2259 3.4105
R26905 GNDA.n2280 GNDA.n2259 3.4105
R26906 GNDA.n2324 GNDA.n2259 3.4105
R26907 GNDA.n2649 GNDA.n2259 3.4105
R26908 GNDA.n2651 GNDA.n2259 3.4105
R26909 GNDA.n2653 GNDA.n2265 3.4105
R26910 GNDA.n2294 GNDA.n2265 3.4105
R26911 GNDA.n2296 GNDA.n2265 3.4105
R26912 GNDA.n2293 GNDA.n2265 3.4105
R26913 GNDA.n2298 GNDA.n2265 3.4105
R26914 GNDA.n2292 GNDA.n2265 3.4105
R26915 GNDA.n2300 GNDA.n2265 3.4105
R26916 GNDA.n2291 GNDA.n2265 3.4105
R26917 GNDA.n2302 GNDA.n2265 3.4105
R26918 GNDA.n2290 GNDA.n2265 3.4105
R26919 GNDA.n2304 GNDA.n2265 3.4105
R26920 GNDA.n2289 GNDA.n2265 3.4105
R26921 GNDA.n2306 GNDA.n2265 3.4105
R26922 GNDA.n2288 GNDA.n2265 3.4105
R26923 GNDA.n2308 GNDA.n2265 3.4105
R26924 GNDA.n2287 GNDA.n2265 3.4105
R26925 GNDA.n2310 GNDA.n2265 3.4105
R26926 GNDA.n2286 GNDA.n2265 3.4105
R26927 GNDA.n2312 GNDA.n2265 3.4105
R26928 GNDA.n2285 GNDA.n2265 3.4105
R26929 GNDA.n2314 GNDA.n2265 3.4105
R26930 GNDA.n2284 GNDA.n2265 3.4105
R26931 GNDA.n2316 GNDA.n2265 3.4105
R26932 GNDA.n2283 GNDA.n2265 3.4105
R26933 GNDA.n2318 GNDA.n2265 3.4105
R26934 GNDA.n2282 GNDA.n2265 3.4105
R26935 GNDA.n2320 GNDA.n2265 3.4105
R26936 GNDA.n2281 GNDA.n2265 3.4105
R26937 GNDA.n2322 GNDA.n2265 3.4105
R26938 GNDA.n2280 GNDA.n2265 3.4105
R26939 GNDA.n2324 GNDA.n2265 3.4105
R26940 GNDA.n2649 GNDA.n2265 3.4105
R26941 GNDA.n2651 GNDA.n2265 3.4105
R26942 GNDA.n2653 GNDA.n2258 3.4105
R26943 GNDA.n2294 GNDA.n2258 3.4105
R26944 GNDA.n2296 GNDA.n2258 3.4105
R26945 GNDA.n2293 GNDA.n2258 3.4105
R26946 GNDA.n2298 GNDA.n2258 3.4105
R26947 GNDA.n2292 GNDA.n2258 3.4105
R26948 GNDA.n2300 GNDA.n2258 3.4105
R26949 GNDA.n2291 GNDA.n2258 3.4105
R26950 GNDA.n2302 GNDA.n2258 3.4105
R26951 GNDA.n2290 GNDA.n2258 3.4105
R26952 GNDA.n2304 GNDA.n2258 3.4105
R26953 GNDA.n2289 GNDA.n2258 3.4105
R26954 GNDA.n2306 GNDA.n2258 3.4105
R26955 GNDA.n2288 GNDA.n2258 3.4105
R26956 GNDA.n2308 GNDA.n2258 3.4105
R26957 GNDA.n2287 GNDA.n2258 3.4105
R26958 GNDA.n2310 GNDA.n2258 3.4105
R26959 GNDA.n2286 GNDA.n2258 3.4105
R26960 GNDA.n2312 GNDA.n2258 3.4105
R26961 GNDA.n2285 GNDA.n2258 3.4105
R26962 GNDA.n2314 GNDA.n2258 3.4105
R26963 GNDA.n2284 GNDA.n2258 3.4105
R26964 GNDA.n2316 GNDA.n2258 3.4105
R26965 GNDA.n2283 GNDA.n2258 3.4105
R26966 GNDA.n2318 GNDA.n2258 3.4105
R26967 GNDA.n2282 GNDA.n2258 3.4105
R26968 GNDA.n2320 GNDA.n2258 3.4105
R26969 GNDA.n2281 GNDA.n2258 3.4105
R26970 GNDA.n2322 GNDA.n2258 3.4105
R26971 GNDA.n2280 GNDA.n2258 3.4105
R26972 GNDA.n2324 GNDA.n2258 3.4105
R26973 GNDA.n2649 GNDA.n2258 3.4105
R26974 GNDA.n2651 GNDA.n2258 3.4105
R26975 GNDA.n2653 GNDA.n2266 3.4105
R26976 GNDA.n2294 GNDA.n2266 3.4105
R26977 GNDA.n2296 GNDA.n2266 3.4105
R26978 GNDA.n2293 GNDA.n2266 3.4105
R26979 GNDA.n2298 GNDA.n2266 3.4105
R26980 GNDA.n2292 GNDA.n2266 3.4105
R26981 GNDA.n2300 GNDA.n2266 3.4105
R26982 GNDA.n2291 GNDA.n2266 3.4105
R26983 GNDA.n2302 GNDA.n2266 3.4105
R26984 GNDA.n2290 GNDA.n2266 3.4105
R26985 GNDA.n2304 GNDA.n2266 3.4105
R26986 GNDA.n2289 GNDA.n2266 3.4105
R26987 GNDA.n2306 GNDA.n2266 3.4105
R26988 GNDA.n2288 GNDA.n2266 3.4105
R26989 GNDA.n2308 GNDA.n2266 3.4105
R26990 GNDA.n2287 GNDA.n2266 3.4105
R26991 GNDA.n2310 GNDA.n2266 3.4105
R26992 GNDA.n2286 GNDA.n2266 3.4105
R26993 GNDA.n2312 GNDA.n2266 3.4105
R26994 GNDA.n2285 GNDA.n2266 3.4105
R26995 GNDA.n2314 GNDA.n2266 3.4105
R26996 GNDA.n2284 GNDA.n2266 3.4105
R26997 GNDA.n2316 GNDA.n2266 3.4105
R26998 GNDA.n2283 GNDA.n2266 3.4105
R26999 GNDA.n2318 GNDA.n2266 3.4105
R27000 GNDA.n2282 GNDA.n2266 3.4105
R27001 GNDA.n2320 GNDA.n2266 3.4105
R27002 GNDA.n2281 GNDA.n2266 3.4105
R27003 GNDA.n2322 GNDA.n2266 3.4105
R27004 GNDA.n2280 GNDA.n2266 3.4105
R27005 GNDA.n2324 GNDA.n2266 3.4105
R27006 GNDA.n2649 GNDA.n2266 3.4105
R27007 GNDA.n2651 GNDA.n2266 3.4105
R27008 GNDA.n2653 GNDA.n2257 3.4105
R27009 GNDA.n2294 GNDA.n2257 3.4105
R27010 GNDA.n2296 GNDA.n2257 3.4105
R27011 GNDA.n2293 GNDA.n2257 3.4105
R27012 GNDA.n2298 GNDA.n2257 3.4105
R27013 GNDA.n2292 GNDA.n2257 3.4105
R27014 GNDA.n2300 GNDA.n2257 3.4105
R27015 GNDA.n2291 GNDA.n2257 3.4105
R27016 GNDA.n2302 GNDA.n2257 3.4105
R27017 GNDA.n2290 GNDA.n2257 3.4105
R27018 GNDA.n2304 GNDA.n2257 3.4105
R27019 GNDA.n2289 GNDA.n2257 3.4105
R27020 GNDA.n2306 GNDA.n2257 3.4105
R27021 GNDA.n2288 GNDA.n2257 3.4105
R27022 GNDA.n2308 GNDA.n2257 3.4105
R27023 GNDA.n2287 GNDA.n2257 3.4105
R27024 GNDA.n2310 GNDA.n2257 3.4105
R27025 GNDA.n2286 GNDA.n2257 3.4105
R27026 GNDA.n2312 GNDA.n2257 3.4105
R27027 GNDA.n2285 GNDA.n2257 3.4105
R27028 GNDA.n2314 GNDA.n2257 3.4105
R27029 GNDA.n2284 GNDA.n2257 3.4105
R27030 GNDA.n2316 GNDA.n2257 3.4105
R27031 GNDA.n2283 GNDA.n2257 3.4105
R27032 GNDA.n2318 GNDA.n2257 3.4105
R27033 GNDA.n2282 GNDA.n2257 3.4105
R27034 GNDA.n2320 GNDA.n2257 3.4105
R27035 GNDA.n2281 GNDA.n2257 3.4105
R27036 GNDA.n2322 GNDA.n2257 3.4105
R27037 GNDA.n2280 GNDA.n2257 3.4105
R27038 GNDA.n2324 GNDA.n2257 3.4105
R27039 GNDA.n2649 GNDA.n2257 3.4105
R27040 GNDA.n2651 GNDA.n2257 3.4105
R27041 GNDA.n2653 GNDA.n2267 3.4105
R27042 GNDA.n2294 GNDA.n2267 3.4105
R27043 GNDA.n2296 GNDA.n2267 3.4105
R27044 GNDA.n2293 GNDA.n2267 3.4105
R27045 GNDA.n2298 GNDA.n2267 3.4105
R27046 GNDA.n2292 GNDA.n2267 3.4105
R27047 GNDA.n2300 GNDA.n2267 3.4105
R27048 GNDA.n2291 GNDA.n2267 3.4105
R27049 GNDA.n2302 GNDA.n2267 3.4105
R27050 GNDA.n2290 GNDA.n2267 3.4105
R27051 GNDA.n2304 GNDA.n2267 3.4105
R27052 GNDA.n2289 GNDA.n2267 3.4105
R27053 GNDA.n2306 GNDA.n2267 3.4105
R27054 GNDA.n2288 GNDA.n2267 3.4105
R27055 GNDA.n2308 GNDA.n2267 3.4105
R27056 GNDA.n2287 GNDA.n2267 3.4105
R27057 GNDA.n2310 GNDA.n2267 3.4105
R27058 GNDA.n2286 GNDA.n2267 3.4105
R27059 GNDA.n2312 GNDA.n2267 3.4105
R27060 GNDA.n2285 GNDA.n2267 3.4105
R27061 GNDA.n2314 GNDA.n2267 3.4105
R27062 GNDA.n2284 GNDA.n2267 3.4105
R27063 GNDA.n2316 GNDA.n2267 3.4105
R27064 GNDA.n2283 GNDA.n2267 3.4105
R27065 GNDA.n2318 GNDA.n2267 3.4105
R27066 GNDA.n2282 GNDA.n2267 3.4105
R27067 GNDA.n2320 GNDA.n2267 3.4105
R27068 GNDA.n2281 GNDA.n2267 3.4105
R27069 GNDA.n2322 GNDA.n2267 3.4105
R27070 GNDA.n2280 GNDA.n2267 3.4105
R27071 GNDA.n2324 GNDA.n2267 3.4105
R27072 GNDA.n2649 GNDA.n2267 3.4105
R27073 GNDA.n2651 GNDA.n2267 3.4105
R27074 GNDA.n2653 GNDA.n2256 3.4105
R27075 GNDA.n2294 GNDA.n2256 3.4105
R27076 GNDA.n2296 GNDA.n2256 3.4105
R27077 GNDA.n2293 GNDA.n2256 3.4105
R27078 GNDA.n2298 GNDA.n2256 3.4105
R27079 GNDA.n2292 GNDA.n2256 3.4105
R27080 GNDA.n2300 GNDA.n2256 3.4105
R27081 GNDA.n2291 GNDA.n2256 3.4105
R27082 GNDA.n2302 GNDA.n2256 3.4105
R27083 GNDA.n2290 GNDA.n2256 3.4105
R27084 GNDA.n2304 GNDA.n2256 3.4105
R27085 GNDA.n2289 GNDA.n2256 3.4105
R27086 GNDA.n2306 GNDA.n2256 3.4105
R27087 GNDA.n2288 GNDA.n2256 3.4105
R27088 GNDA.n2308 GNDA.n2256 3.4105
R27089 GNDA.n2287 GNDA.n2256 3.4105
R27090 GNDA.n2310 GNDA.n2256 3.4105
R27091 GNDA.n2286 GNDA.n2256 3.4105
R27092 GNDA.n2312 GNDA.n2256 3.4105
R27093 GNDA.n2285 GNDA.n2256 3.4105
R27094 GNDA.n2314 GNDA.n2256 3.4105
R27095 GNDA.n2284 GNDA.n2256 3.4105
R27096 GNDA.n2316 GNDA.n2256 3.4105
R27097 GNDA.n2283 GNDA.n2256 3.4105
R27098 GNDA.n2318 GNDA.n2256 3.4105
R27099 GNDA.n2282 GNDA.n2256 3.4105
R27100 GNDA.n2320 GNDA.n2256 3.4105
R27101 GNDA.n2281 GNDA.n2256 3.4105
R27102 GNDA.n2322 GNDA.n2256 3.4105
R27103 GNDA.n2280 GNDA.n2256 3.4105
R27104 GNDA.n2324 GNDA.n2256 3.4105
R27105 GNDA.n2649 GNDA.n2256 3.4105
R27106 GNDA.n2651 GNDA.n2256 3.4105
R27107 GNDA.n2653 GNDA.n2268 3.4105
R27108 GNDA.n2294 GNDA.n2268 3.4105
R27109 GNDA.n2296 GNDA.n2268 3.4105
R27110 GNDA.n2293 GNDA.n2268 3.4105
R27111 GNDA.n2298 GNDA.n2268 3.4105
R27112 GNDA.n2292 GNDA.n2268 3.4105
R27113 GNDA.n2300 GNDA.n2268 3.4105
R27114 GNDA.n2291 GNDA.n2268 3.4105
R27115 GNDA.n2302 GNDA.n2268 3.4105
R27116 GNDA.n2290 GNDA.n2268 3.4105
R27117 GNDA.n2304 GNDA.n2268 3.4105
R27118 GNDA.n2289 GNDA.n2268 3.4105
R27119 GNDA.n2306 GNDA.n2268 3.4105
R27120 GNDA.n2288 GNDA.n2268 3.4105
R27121 GNDA.n2308 GNDA.n2268 3.4105
R27122 GNDA.n2287 GNDA.n2268 3.4105
R27123 GNDA.n2310 GNDA.n2268 3.4105
R27124 GNDA.n2286 GNDA.n2268 3.4105
R27125 GNDA.n2312 GNDA.n2268 3.4105
R27126 GNDA.n2285 GNDA.n2268 3.4105
R27127 GNDA.n2314 GNDA.n2268 3.4105
R27128 GNDA.n2284 GNDA.n2268 3.4105
R27129 GNDA.n2316 GNDA.n2268 3.4105
R27130 GNDA.n2283 GNDA.n2268 3.4105
R27131 GNDA.n2318 GNDA.n2268 3.4105
R27132 GNDA.n2282 GNDA.n2268 3.4105
R27133 GNDA.n2320 GNDA.n2268 3.4105
R27134 GNDA.n2281 GNDA.n2268 3.4105
R27135 GNDA.n2322 GNDA.n2268 3.4105
R27136 GNDA.n2280 GNDA.n2268 3.4105
R27137 GNDA.n2324 GNDA.n2268 3.4105
R27138 GNDA.n2649 GNDA.n2268 3.4105
R27139 GNDA.n2651 GNDA.n2268 3.4105
R27140 GNDA.n2653 GNDA.n2255 3.4105
R27141 GNDA.n2294 GNDA.n2255 3.4105
R27142 GNDA.n2296 GNDA.n2255 3.4105
R27143 GNDA.n2293 GNDA.n2255 3.4105
R27144 GNDA.n2298 GNDA.n2255 3.4105
R27145 GNDA.n2292 GNDA.n2255 3.4105
R27146 GNDA.n2300 GNDA.n2255 3.4105
R27147 GNDA.n2291 GNDA.n2255 3.4105
R27148 GNDA.n2302 GNDA.n2255 3.4105
R27149 GNDA.n2290 GNDA.n2255 3.4105
R27150 GNDA.n2304 GNDA.n2255 3.4105
R27151 GNDA.n2289 GNDA.n2255 3.4105
R27152 GNDA.n2306 GNDA.n2255 3.4105
R27153 GNDA.n2288 GNDA.n2255 3.4105
R27154 GNDA.n2308 GNDA.n2255 3.4105
R27155 GNDA.n2287 GNDA.n2255 3.4105
R27156 GNDA.n2310 GNDA.n2255 3.4105
R27157 GNDA.n2286 GNDA.n2255 3.4105
R27158 GNDA.n2312 GNDA.n2255 3.4105
R27159 GNDA.n2285 GNDA.n2255 3.4105
R27160 GNDA.n2314 GNDA.n2255 3.4105
R27161 GNDA.n2284 GNDA.n2255 3.4105
R27162 GNDA.n2316 GNDA.n2255 3.4105
R27163 GNDA.n2283 GNDA.n2255 3.4105
R27164 GNDA.n2318 GNDA.n2255 3.4105
R27165 GNDA.n2282 GNDA.n2255 3.4105
R27166 GNDA.n2320 GNDA.n2255 3.4105
R27167 GNDA.n2281 GNDA.n2255 3.4105
R27168 GNDA.n2322 GNDA.n2255 3.4105
R27169 GNDA.n2280 GNDA.n2255 3.4105
R27170 GNDA.n2324 GNDA.n2255 3.4105
R27171 GNDA.n2649 GNDA.n2255 3.4105
R27172 GNDA.n2651 GNDA.n2255 3.4105
R27173 GNDA.n2653 GNDA.n2269 3.4105
R27174 GNDA.n2294 GNDA.n2269 3.4105
R27175 GNDA.n2296 GNDA.n2269 3.4105
R27176 GNDA.n2293 GNDA.n2269 3.4105
R27177 GNDA.n2298 GNDA.n2269 3.4105
R27178 GNDA.n2292 GNDA.n2269 3.4105
R27179 GNDA.n2300 GNDA.n2269 3.4105
R27180 GNDA.n2291 GNDA.n2269 3.4105
R27181 GNDA.n2302 GNDA.n2269 3.4105
R27182 GNDA.n2290 GNDA.n2269 3.4105
R27183 GNDA.n2304 GNDA.n2269 3.4105
R27184 GNDA.n2289 GNDA.n2269 3.4105
R27185 GNDA.n2306 GNDA.n2269 3.4105
R27186 GNDA.n2288 GNDA.n2269 3.4105
R27187 GNDA.n2308 GNDA.n2269 3.4105
R27188 GNDA.n2287 GNDA.n2269 3.4105
R27189 GNDA.n2310 GNDA.n2269 3.4105
R27190 GNDA.n2286 GNDA.n2269 3.4105
R27191 GNDA.n2312 GNDA.n2269 3.4105
R27192 GNDA.n2285 GNDA.n2269 3.4105
R27193 GNDA.n2314 GNDA.n2269 3.4105
R27194 GNDA.n2284 GNDA.n2269 3.4105
R27195 GNDA.n2316 GNDA.n2269 3.4105
R27196 GNDA.n2283 GNDA.n2269 3.4105
R27197 GNDA.n2318 GNDA.n2269 3.4105
R27198 GNDA.n2282 GNDA.n2269 3.4105
R27199 GNDA.n2320 GNDA.n2269 3.4105
R27200 GNDA.n2281 GNDA.n2269 3.4105
R27201 GNDA.n2322 GNDA.n2269 3.4105
R27202 GNDA.n2280 GNDA.n2269 3.4105
R27203 GNDA.n2324 GNDA.n2269 3.4105
R27204 GNDA.n2649 GNDA.n2269 3.4105
R27205 GNDA.n2651 GNDA.n2269 3.4105
R27206 GNDA.n2653 GNDA.n2254 3.4105
R27207 GNDA.n2294 GNDA.n2254 3.4105
R27208 GNDA.n2296 GNDA.n2254 3.4105
R27209 GNDA.n2293 GNDA.n2254 3.4105
R27210 GNDA.n2298 GNDA.n2254 3.4105
R27211 GNDA.n2292 GNDA.n2254 3.4105
R27212 GNDA.n2300 GNDA.n2254 3.4105
R27213 GNDA.n2291 GNDA.n2254 3.4105
R27214 GNDA.n2302 GNDA.n2254 3.4105
R27215 GNDA.n2290 GNDA.n2254 3.4105
R27216 GNDA.n2304 GNDA.n2254 3.4105
R27217 GNDA.n2289 GNDA.n2254 3.4105
R27218 GNDA.n2306 GNDA.n2254 3.4105
R27219 GNDA.n2288 GNDA.n2254 3.4105
R27220 GNDA.n2308 GNDA.n2254 3.4105
R27221 GNDA.n2287 GNDA.n2254 3.4105
R27222 GNDA.n2310 GNDA.n2254 3.4105
R27223 GNDA.n2286 GNDA.n2254 3.4105
R27224 GNDA.n2312 GNDA.n2254 3.4105
R27225 GNDA.n2285 GNDA.n2254 3.4105
R27226 GNDA.n2314 GNDA.n2254 3.4105
R27227 GNDA.n2284 GNDA.n2254 3.4105
R27228 GNDA.n2316 GNDA.n2254 3.4105
R27229 GNDA.n2283 GNDA.n2254 3.4105
R27230 GNDA.n2318 GNDA.n2254 3.4105
R27231 GNDA.n2282 GNDA.n2254 3.4105
R27232 GNDA.n2320 GNDA.n2254 3.4105
R27233 GNDA.n2281 GNDA.n2254 3.4105
R27234 GNDA.n2322 GNDA.n2254 3.4105
R27235 GNDA.n2280 GNDA.n2254 3.4105
R27236 GNDA.n2324 GNDA.n2254 3.4105
R27237 GNDA.n2649 GNDA.n2254 3.4105
R27238 GNDA.n2651 GNDA.n2254 3.4105
R27239 GNDA.n2653 GNDA.n2270 3.4105
R27240 GNDA.n2294 GNDA.n2270 3.4105
R27241 GNDA.n2296 GNDA.n2270 3.4105
R27242 GNDA.n2293 GNDA.n2270 3.4105
R27243 GNDA.n2298 GNDA.n2270 3.4105
R27244 GNDA.n2292 GNDA.n2270 3.4105
R27245 GNDA.n2300 GNDA.n2270 3.4105
R27246 GNDA.n2291 GNDA.n2270 3.4105
R27247 GNDA.n2302 GNDA.n2270 3.4105
R27248 GNDA.n2290 GNDA.n2270 3.4105
R27249 GNDA.n2304 GNDA.n2270 3.4105
R27250 GNDA.n2289 GNDA.n2270 3.4105
R27251 GNDA.n2306 GNDA.n2270 3.4105
R27252 GNDA.n2288 GNDA.n2270 3.4105
R27253 GNDA.n2308 GNDA.n2270 3.4105
R27254 GNDA.n2287 GNDA.n2270 3.4105
R27255 GNDA.n2310 GNDA.n2270 3.4105
R27256 GNDA.n2286 GNDA.n2270 3.4105
R27257 GNDA.n2312 GNDA.n2270 3.4105
R27258 GNDA.n2285 GNDA.n2270 3.4105
R27259 GNDA.n2314 GNDA.n2270 3.4105
R27260 GNDA.n2284 GNDA.n2270 3.4105
R27261 GNDA.n2316 GNDA.n2270 3.4105
R27262 GNDA.n2283 GNDA.n2270 3.4105
R27263 GNDA.n2318 GNDA.n2270 3.4105
R27264 GNDA.n2282 GNDA.n2270 3.4105
R27265 GNDA.n2320 GNDA.n2270 3.4105
R27266 GNDA.n2281 GNDA.n2270 3.4105
R27267 GNDA.n2322 GNDA.n2270 3.4105
R27268 GNDA.n2280 GNDA.n2270 3.4105
R27269 GNDA.n2324 GNDA.n2270 3.4105
R27270 GNDA.n2649 GNDA.n2270 3.4105
R27271 GNDA.n2651 GNDA.n2270 3.4105
R27272 GNDA.n2653 GNDA.n2253 3.4105
R27273 GNDA.n2294 GNDA.n2253 3.4105
R27274 GNDA.n2296 GNDA.n2253 3.4105
R27275 GNDA.n2293 GNDA.n2253 3.4105
R27276 GNDA.n2298 GNDA.n2253 3.4105
R27277 GNDA.n2292 GNDA.n2253 3.4105
R27278 GNDA.n2300 GNDA.n2253 3.4105
R27279 GNDA.n2291 GNDA.n2253 3.4105
R27280 GNDA.n2302 GNDA.n2253 3.4105
R27281 GNDA.n2290 GNDA.n2253 3.4105
R27282 GNDA.n2304 GNDA.n2253 3.4105
R27283 GNDA.n2289 GNDA.n2253 3.4105
R27284 GNDA.n2306 GNDA.n2253 3.4105
R27285 GNDA.n2288 GNDA.n2253 3.4105
R27286 GNDA.n2308 GNDA.n2253 3.4105
R27287 GNDA.n2287 GNDA.n2253 3.4105
R27288 GNDA.n2310 GNDA.n2253 3.4105
R27289 GNDA.n2286 GNDA.n2253 3.4105
R27290 GNDA.n2312 GNDA.n2253 3.4105
R27291 GNDA.n2285 GNDA.n2253 3.4105
R27292 GNDA.n2314 GNDA.n2253 3.4105
R27293 GNDA.n2284 GNDA.n2253 3.4105
R27294 GNDA.n2316 GNDA.n2253 3.4105
R27295 GNDA.n2283 GNDA.n2253 3.4105
R27296 GNDA.n2318 GNDA.n2253 3.4105
R27297 GNDA.n2282 GNDA.n2253 3.4105
R27298 GNDA.n2320 GNDA.n2253 3.4105
R27299 GNDA.n2281 GNDA.n2253 3.4105
R27300 GNDA.n2322 GNDA.n2253 3.4105
R27301 GNDA.n2280 GNDA.n2253 3.4105
R27302 GNDA.n2324 GNDA.n2253 3.4105
R27303 GNDA.n2649 GNDA.n2253 3.4105
R27304 GNDA.n2651 GNDA.n2253 3.4105
R27305 GNDA.n2653 GNDA.n2271 3.4105
R27306 GNDA.n2294 GNDA.n2271 3.4105
R27307 GNDA.n2296 GNDA.n2271 3.4105
R27308 GNDA.n2293 GNDA.n2271 3.4105
R27309 GNDA.n2298 GNDA.n2271 3.4105
R27310 GNDA.n2292 GNDA.n2271 3.4105
R27311 GNDA.n2300 GNDA.n2271 3.4105
R27312 GNDA.n2291 GNDA.n2271 3.4105
R27313 GNDA.n2302 GNDA.n2271 3.4105
R27314 GNDA.n2290 GNDA.n2271 3.4105
R27315 GNDA.n2304 GNDA.n2271 3.4105
R27316 GNDA.n2289 GNDA.n2271 3.4105
R27317 GNDA.n2306 GNDA.n2271 3.4105
R27318 GNDA.n2288 GNDA.n2271 3.4105
R27319 GNDA.n2308 GNDA.n2271 3.4105
R27320 GNDA.n2287 GNDA.n2271 3.4105
R27321 GNDA.n2310 GNDA.n2271 3.4105
R27322 GNDA.n2286 GNDA.n2271 3.4105
R27323 GNDA.n2312 GNDA.n2271 3.4105
R27324 GNDA.n2285 GNDA.n2271 3.4105
R27325 GNDA.n2314 GNDA.n2271 3.4105
R27326 GNDA.n2284 GNDA.n2271 3.4105
R27327 GNDA.n2316 GNDA.n2271 3.4105
R27328 GNDA.n2283 GNDA.n2271 3.4105
R27329 GNDA.n2318 GNDA.n2271 3.4105
R27330 GNDA.n2282 GNDA.n2271 3.4105
R27331 GNDA.n2320 GNDA.n2271 3.4105
R27332 GNDA.n2281 GNDA.n2271 3.4105
R27333 GNDA.n2322 GNDA.n2271 3.4105
R27334 GNDA.n2280 GNDA.n2271 3.4105
R27335 GNDA.n2324 GNDA.n2271 3.4105
R27336 GNDA.n2649 GNDA.n2271 3.4105
R27337 GNDA.n2651 GNDA.n2271 3.4105
R27338 GNDA.n2653 GNDA.n2252 3.4105
R27339 GNDA.n2294 GNDA.n2252 3.4105
R27340 GNDA.n2296 GNDA.n2252 3.4105
R27341 GNDA.n2293 GNDA.n2252 3.4105
R27342 GNDA.n2298 GNDA.n2252 3.4105
R27343 GNDA.n2292 GNDA.n2252 3.4105
R27344 GNDA.n2300 GNDA.n2252 3.4105
R27345 GNDA.n2291 GNDA.n2252 3.4105
R27346 GNDA.n2302 GNDA.n2252 3.4105
R27347 GNDA.n2290 GNDA.n2252 3.4105
R27348 GNDA.n2304 GNDA.n2252 3.4105
R27349 GNDA.n2289 GNDA.n2252 3.4105
R27350 GNDA.n2306 GNDA.n2252 3.4105
R27351 GNDA.n2288 GNDA.n2252 3.4105
R27352 GNDA.n2308 GNDA.n2252 3.4105
R27353 GNDA.n2287 GNDA.n2252 3.4105
R27354 GNDA.n2310 GNDA.n2252 3.4105
R27355 GNDA.n2286 GNDA.n2252 3.4105
R27356 GNDA.n2312 GNDA.n2252 3.4105
R27357 GNDA.n2285 GNDA.n2252 3.4105
R27358 GNDA.n2314 GNDA.n2252 3.4105
R27359 GNDA.n2284 GNDA.n2252 3.4105
R27360 GNDA.n2316 GNDA.n2252 3.4105
R27361 GNDA.n2283 GNDA.n2252 3.4105
R27362 GNDA.n2318 GNDA.n2252 3.4105
R27363 GNDA.n2282 GNDA.n2252 3.4105
R27364 GNDA.n2320 GNDA.n2252 3.4105
R27365 GNDA.n2281 GNDA.n2252 3.4105
R27366 GNDA.n2322 GNDA.n2252 3.4105
R27367 GNDA.n2280 GNDA.n2252 3.4105
R27368 GNDA.n2324 GNDA.n2252 3.4105
R27369 GNDA.n2649 GNDA.n2252 3.4105
R27370 GNDA.n2651 GNDA.n2252 3.4105
R27371 GNDA.n2653 GNDA.n2272 3.4105
R27372 GNDA.n2294 GNDA.n2272 3.4105
R27373 GNDA.n2296 GNDA.n2272 3.4105
R27374 GNDA.n2293 GNDA.n2272 3.4105
R27375 GNDA.n2298 GNDA.n2272 3.4105
R27376 GNDA.n2292 GNDA.n2272 3.4105
R27377 GNDA.n2300 GNDA.n2272 3.4105
R27378 GNDA.n2291 GNDA.n2272 3.4105
R27379 GNDA.n2302 GNDA.n2272 3.4105
R27380 GNDA.n2290 GNDA.n2272 3.4105
R27381 GNDA.n2304 GNDA.n2272 3.4105
R27382 GNDA.n2289 GNDA.n2272 3.4105
R27383 GNDA.n2306 GNDA.n2272 3.4105
R27384 GNDA.n2288 GNDA.n2272 3.4105
R27385 GNDA.n2308 GNDA.n2272 3.4105
R27386 GNDA.n2287 GNDA.n2272 3.4105
R27387 GNDA.n2310 GNDA.n2272 3.4105
R27388 GNDA.n2286 GNDA.n2272 3.4105
R27389 GNDA.n2312 GNDA.n2272 3.4105
R27390 GNDA.n2285 GNDA.n2272 3.4105
R27391 GNDA.n2314 GNDA.n2272 3.4105
R27392 GNDA.n2284 GNDA.n2272 3.4105
R27393 GNDA.n2316 GNDA.n2272 3.4105
R27394 GNDA.n2283 GNDA.n2272 3.4105
R27395 GNDA.n2318 GNDA.n2272 3.4105
R27396 GNDA.n2282 GNDA.n2272 3.4105
R27397 GNDA.n2320 GNDA.n2272 3.4105
R27398 GNDA.n2281 GNDA.n2272 3.4105
R27399 GNDA.n2322 GNDA.n2272 3.4105
R27400 GNDA.n2280 GNDA.n2272 3.4105
R27401 GNDA.n2324 GNDA.n2272 3.4105
R27402 GNDA.n2649 GNDA.n2272 3.4105
R27403 GNDA.n2651 GNDA.n2272 3.4105
R27404 GNDA.n2653 GNDA.n2251 3.4105
R27405 GNDA.n2294 GNDA.n2251 3.4105
R27406 GNDA.n2296 GNDA.n2251 3.4105
R27407 GNDA.n2293 GNDA.n2251 3.4105
R27408 GNDA.n2298 GNDA.n2251 3.4105
R27409 GNDA.n2292 GNDA.n2251 3.4105
R27410 GNDA.n2300 GNDA.n2251 3.4105
R27411 GNDA.n2291 GNDA.n2251 3.4105
R27412 GNDA.n2302 GNDA.n2251 3.4105
R27413 GNDA.n2290 GNDA.n2251 3.4105
R27414 GNDA.n2304 GNDA.n2251 3.4105
R27415 GNDA.n2289 GNDA.n2251 3.4105
R27416 GNDA.n2306 GNDA.n2251 3.4105
R27417 GNDA.n2288 GNDA.n2251 3.4105
R27418 GNDA.n2308 GNDA.n2251 3.4105
R27419 GNDA.n2287 GNDA.n2251 3.4105
R27420 GNDA.n2310 GNDA.n2251 3.4105
R27421 GNDA.n2286 GNDA.n2251 3.4105
R27422 GNDA.n2312 GNDA.n2251 3.4105
R27423 GNDA.n2285 GNDA.n2251 3.4105
R27424 GNDA.n2314 GNDA.n2251 3.4105
R27425 GNDA.n2284 GNDA.n2251 3.4105
R27426 GNDA.n2316 GNDA.n2251 3.4105
R27427 GNDA.n2283 GNDA.n2251 3.4105
R27428 GNDA.n2318 GNDA.n2251 3.4105
R27429 GNDA.n2282 GNDA.n2251 3.4105
R27430 GNDA.n2320 GNDA.n2251 3.4105
R27431 GNDA.n2281 GNDA.n2251 3.4105
R27432 GNDA.n2322 GNDA.n2251 3.4105
R27433 GNDA.n2280 GNDA.n2251 3.4105
R27434 GNDA.n2324 GNDA.n2251 3.4105
R27435 GNDA.n2649 GNDA.n2251 3.4105
R27436 GNDA.n2651 GNDA.n2251 3.4105
R27437 GNDA.n2653 GNDA.n2273 3.4105
R27438 GNDA.n2294 GNDA.n2273 3.4105
R27439 GNDA.n2296 GNDA.n2273 3.4105
R27440 GNDA.n2293 GNDA.n2273 3.4105
R27441 GNDA.n2298 GNDA.n2273 3.4105
R27442 GNDA.n2292 GNDA.n2273 3.4105
R27443 GNDA.n2300 GNDA.n2273 3.4105
R27444 GNDA.n2291 GNDA.n2273 3.4105
R27445 GNDA.n2302 GNDA.n2273 3.4105
R27446 GNDA.n2290 GNDA.n2273 3.4105
R27447 GNDA.n2304 GNDA.n2273 3.4105
R27448 GNDA.n2289 GNDA.n2273 3.4105
R27449 GNDA.n2306 GNDA.n2273 3.4105
R27450 GNDA.n2288 GNDA.n2273 3.4105
R27451 GNDA.n2308 GNDA.n2273 3.4105
R27452 GNDA.n2287 GNDA.n2273 3.4105
R27453 GNDA.n2310 GNDA.n2273 3.4105
R27454 GNDA.n2286 GNDA.n2273 3.4105
R27455 GNDA.n2312 GNDA.n2273 3.4105
R27456 GNDA.n2285 GNDA.n2273 3.4105
R27457 GNDA.n2314 GNDA.n2273 3.4105
R27458 GNDA.n2284 GNDA.n2273 3.4105
R27459 GNDA.n2316 GNDA.n2273 3.4105
R27460 GNDA.n2283 GNDA.n2273 3.4105
R27461 GNDA.n2318 GNDA.n2273 3.4105
R27462 GNDA.n2282 GNDA.n2273 3.4105
R27463 GNDA.n2320 GNDA.n2273 3.4105
R27464 GNDA.n2281 GNDA.n2273 3.4105
R27465 GNDA.n2322 GNDA.n2273 3.4105
R27466 GNDA.n2280 GNDA.n2273 3.4105
R27467 GNDA.n2324 GNDA.n2273 3.4105
R27468 GNDA.n2649 GNDA.n2273 3.4105
R27469 GNDA.n2651 GNDA.n2273 3.4105
R27470 GNDA.n2653 GNDA.n2250 3.4105
R27471 GNDA.n2294 GNDA.n2250 3.4105
R27472 GNDA.n2296 GNDA.n2250 3.4105
R27473 GNDA.n2293 GNDA.n2250 3.4105
R27474 GNDA.n2298 GNDA.n2250 3.4105
R27475 GNDA.n2292 GNDA.n2250 3.4105
R27476 GNDA.n2300 GNDA.n2250 3.4105
R27477 GNDA.n2291 GNDA.n2250 3.4105
R27478 GNDA.n2302 GNDA.n2250 3.4105
R27479 GNDA.n2290 GNDA.n2250 3.4105
R27480 GNDA.n2304 GNDA.n2250 3.4105
R27481 GNDA.n2289 GNDA.n2250 3.4105
R27482 GNDA.n2306 GNDA.n2250 3.4105
R27483 GNDA.n2288 GNDA.n2250 3.4105
R27484 GNDA.n2308 GNDA.n2250 3.4105
R27485 GNDA.n2287 GNDA.n2250 3.4105
R27486 GNDA.n2310 GNDA.n2250 3.4105
R27487 GNDA.n2286 GNDA.n2250 3.4105
R27488 GNDA.n2312 GNDA.n2250 3.4105
R27489 GNDA.n2285 GNDA.n2250 3.4105
R27490 GNDA.n2314 GNDA.n2250 3.4105
R27491 GNDA.n2284 GNDA.n2250 3.4105
R27492 GNDA.n2316 GNDA.n2250 3.4105
R27493 GNDA.n2283 GNDA.n2250 3.4105
R27494 GNDA.n2318 GNDA.n2250 3.4105
R27495 GNDA.n2282 GNDA.n2250 3.4105
R27496 GNDA.n2320 GNDA.n2250 3.4105
R27497 GNDA.n2281 GNDA.n2250 3.4105
R27498 GNDA.n2322 GNDA.n2250 3.4105
R27499 GNDA.n2280 GNDA.n2250 3.4105
R27500 GNDA.n2324 GNDA.n2250 3.4105
R27501 GNDA.n2649 GNDA.n2250 3.4105
R27502 GNDA.n2651 GNDA.n2250 3.4105
R27503 GNDA.n2653 GNDA.n2274 3.4105
R27504 GNDA.n2294 GNDA.n2274 3.4105
R27505 GNDA.n2296 GNDA.n2274 3.4105
R27506 GNDA.n2293 GNDA.n2274 3.4105
R27507 GNDA.n2298 GNDA.n2274 3.4105
R27508 GNDA.n2292 GNDA.n2274 3.4105
R27509 GNDA.n2300 GNDA.n2274 3.4105
R27510 GNDA.n2291 GNDA.n2274 3.4105
R27511 GNDA.n2302 GNDA.n2274 3.4105
R27512 GNDA.n2290 GNDA.n2274 3.4105
R27513 GNDA.n2304 GNDA.n2274 3.4105
R27514 GNDA.n2289 GNDA.n2274 3.4105
R27515 GNDA.n2306 GNDA.n2274 3.4105
R27516 GNDA.n2288 GNDA.n2274 3.4105
R27517 GNDA.n2308 GNDA.n2274 3.4105
R27518 GNDA.n2287 GNDA.n2274 3.4105
R27519 GNDA.n2310 GNDA.n2274 3.4105
R27520 GNDA.n2286 GNDA.n2274 3.4105
R27521 GNDA.n2312 GNDA.n2274 3.4105
R27522 GNDA.n2285 GNDA.n2274 3.4105
R27523 GNDA.n2314 GNDA.n2274 3.4105
R27524 GNDA.n2284 GNDA.n2274 3.4105
R27525 GNDA.n2316 GNDA.n2274 3.4105
R27526 GNDA.n2283 GNDA.n2274 3.4105
R27527 GNDA.n2318 GNDA.n2274 3.4105
R27528 GNDA.n2282 GNDA.n2274 3.4105
R27529 GNDA.n2320 GNDA.n2274 3.4105
R27530 GNDA.n2281 GNDA.n2274 3.4105
R27531 GNDA.n2322 GNDA.n2274 3.4105
R27532 GNDA.n2280 GNDA.n2274 3.4105
R27533 GNDA.n2324 GNDA.n2274 3.4105
R27534 GNDA.n2649 GNDA.n2274 3.4105
R27535 GNDA.n2651 GNDA.n2274 3.4105
R27536 GNDA.n2653 GNDA.n2249 3.4105
R27537 GNDA.n2294 GNDA.n2249 3.4105
R27538 GNDA.n2296 GNDA.n2249 3.4105
R27539 GNDA.n2293 GNDA.n2249 3.4105
R27540 GNDA.n2298 GNDA.n2249 3.4105
R27541 GNDA.n2292 GNDA.n2249 3.4105
R27542 GNDA.n2300 GNDA.n2249 3.4105
R27543 GNDA.n2291 GNDA.n2249 3.4105
R27544 GNDA.n2302 GNDA.n2249 3.4105
R27545 GNDA.n2290 GNDA.n2249 3.4105
R27546 GNDA.n2304 GNDA.n2249 3.4105
R27547 GNDA.n2289 GNDA.n2249 3.4105
R27548 GNDA.n2306 GNDA.n2249 3.4105
R27549 GNDA.n2288 GNDA.n2249 3.4105
R27550 GNDA.n2308 GNDA.n2249 3.4105
R27551 GNDA.n2287 GNDA.n2249 3.4105
R27552 GNDA.n2310 GNDA.n2249 3.4105
R27553 GNDA.n2286 GNDA.n2249 3.4105
R27554 GNDA.n2312 GNDA.n2249 3.4105
R27555 GNDA.n2285 GNDA.n2249 3.4105
R27556 GNDA.n2314 GNDA.n2249 3.4105
R27557 GNDA.n2284 GNDA.n2249 3.4105
R27558 GNDA.n2316 GNDA.n2249 3.4105
R27559 GNDA.n2283 GNDA.n2249 3.4105
R27560 GNDA.n2318 GNDA.n2249 3.4105
R27561 GNDA.n2282 GNDA.n2249 3.4105
R27562 GNDA.n2320 GNDA.n2249 3.4105
R27563 GNDA.n2281 GNDA.n2249 3.4105
R27564 GNDA.n2322 GNDA.n2249 3.4105
R27565 GNDA.n2280 GNDA.n2249 3.4105
R27566 GNDA.n2324 GNDA.n2249 3.4105
R27567 GNDA.n2649 GNDA.n2249 3.4105
R27568 GNDA.n2651 GNDA.n2249 3.4105
R27569 GNDA.n2653 GNDA.n2275 3.4105
R27570 GNDA.n2294 GNDA.n2275 3.4105
R27571 GNDA.n2296 GNDA.n2275 3.4105
R27572 GNDA.n2293 GNDA.n2275 3.4105
R27573 GNDA.n2298 GNDA.n2275 3.4105
R27574 GNDA.n2292 GNDA.n2275 3.4105
R27575 GNDA.n2300 GNDA.n2275 3.4105
R27576 GNDA.n2291 GNDA.n2275 3.4105
R27577 GNDA.n2302 GNDA.n2275 3.4105
R27578 GNDA.n2290 GNDA.n2275 3.4105
R27579 GNDA.n2304 GNDA.n2275 3.4105
R27580 GNDA.n2289 GNDA.n2275 3.4105
R27581 GNDA.n2306 GNDA.n2275 3.4105
R27582 GNDA.n2288 GNDA.n2275 3.4105
R27583 GNDA.n2308 GNDA.n2275 3.4105
R27584 GNDA.n2287 GNDA.n2275 3.4105
R27585 GNDA.n2310 GNDA.n2275 3.4105
R27586 GNDA.n2286 GNDA.n2275 3.4105
R27587 GNDA.n2312 GNDA.n2275 3.4105
R27588 GNDA.n2285 GNDA.n2275 3.4105
R27589 GNDA.n2314 GNDA.n2275 3.4105
R27590 GNDA.n2284 GNDA.n2275 3.4105
R27591 GNDA.n2316 GNDA.n2275 3.4105
R27592 GNDA.n2283 GNDA.n2275 3.4105
R27593 GNDA.n2318 GNDA.n2275 3.4105
R27594 GNDA.n2282 GNDA.n2275 3.4105
R27595 GNDA.n2320 GNDA.n2275 3.4105
R27596 GNDA.n2281 GNDA.n2275 3.4105
R27597 GNDA.n2322 GNDA.n2275 3.4105
R27598 GNDA.n2280 GNDA.n2275 3.4105
R27599 GNDA.n2324 GNDA.n2275 3.4105
R27600 GNDA.n2649 GNDA.n2275 3.4105
R27601 GNDA.n2651 GNDA.n2275 3.4105
R27602 GNDA.n2653 GNDA.n2248 3.4105
R27603 GNDA.n2294 GNDA.n2248 3.4105
R27604 GNDA.n2296 GNDA.n2248 3.4105
R27605 GNDA.n2293 GNDA.n2248 3.4105
R27606 GNDA.n2298 GNDA.n2248 3.4105
R27607 GNDA.n2292 GNDA.n2248 3.4105
R27608 GNDA.n2300 GNDA.n2248 3.4105
R27609 GNDA.n2291 GNDA.n2248 3.4105
R27610 GNDA.n2302 GNDA.n2248 3.4105
R27611 GNDA.n2290 GNDA.n2248 3.4105
R27612 GNDA.n2304 GNDA.n2248 3.4105
R27613 GNDA.n2289 GNDA.n2248 3.4105
R27614 GNDA.n2306 GNDA.n2248 3.4105
R27615 GNDA.n2288 GNDA.n2248 3.4105
R27616 GNDA.n2308 GNDA.n2248 3.4105
R27617 GNDA.n2287 GNDA.n2248 3.4105
R27618 GNDA.n2310 GNDA.n2248 3.4105
R27619 GNDA.n2286 GNDA.n2248 3.4105
R27620 GNDA.n2312 GNDA.n2248 3.4105
R27621 GNDA.n2285 GNDA.n2248 3.4105
R27622 GNDA.n2314 GNDA.n2248 3.4105
R27623 GNDA.n2284 GNDA.n2248 3.4105
R27624 GNDA.n2316 GNDA.n2248 3.4105
R27625 GNDA.n2283 GNDA.n2248 3.4105
R27626 GNDA.n2318 GNDA.n2248 3.4105
R27627 GNDA.n2282 GNDA.n2248 3.4105
R27628 GNDA.n2320 GNDA.n2248 3.4105
R27629 GNDA.n2281 GNDA.n2248 3.4105
R27630 GNDA.n2322 GNDA.n2248 3.4105
R27631 GNDA.n2280 GNDA.n2248 3.4105
R27632 GNDA.n2324 GNDA.n2248 3.4105
R27633 GNDA.n2649 GNDA.n2248 3.4105
R27634 GNDA.n2651 GNDA.n2248 3.4105
R27635 GNDA.n2653 GNDA.n2276 3.4105
R27636 GNDA.n2294 GNDA.n2276 3.4105
R27637 GNDA.n2296 GNDA.n2276 3.4105
R27638 GNDA.n2293 GNDA.n2276 3.4105
R27639 GNDA.n2298 GNDA.n2276 3.4105
R27640 GNDA.n2292 GNDA.n2276 3.4105
R27641 GNDA.n2300 GNDA.n2276 3.4105
R27642 GNDA.n2291 GNDA.n2276 3.4105
R27643 GNDA.n2302 GNDA.n2276 3.4105
R27644 GNDA.n2290 GNDA.n2276 3.4105
R27645 GNDA.n2304 GNDA.n2276 3.4105
R27646 GNDA.n2289 GNDA.n2276 3.4105
R27647 GNDA.n2306 GNDA.n2276 3.4105
R27648 GNDA.n2288 GNDA.n2276 3.4105
R27649 GNDA.n2308 GNDA.n2276 3.4105
R27650 GNDA.n2287 GNDA.n2276 3.4105
R27651 GNDA.n2310 GNDA.n2276 3.4105
R27652 GNDA.n2286 GNDA.n2276 3.4105
R27653 GNDA.n2312 GNDA.n2276 3.4105
R27654 GNDA.n2285 GNDA.n2276 3.4105
R27655 GNDA.n2314 GNDA.n2276 3.4105
R27656 GNDA.n2284 GNDA.n2276 3.4105
R27657 GNDA.n2316 GNDA.n2276 3.4105
R27658 GNDA.n2283 GNDA.n2276 3.4105
R27659 GNDA.n2318 GNDA.n2276 3.4105
R27660 GNDA.n2282 GNDA.n2276 3.4105
R27661 GNDA.n2320 GNDA.n2276 3.4105
R27662 GNDA.n2281 GNDA.n2276 3.4105
R27663 GNDA.n2322 GNDA.n2276 3.4105
R27664 GNDA.n2280 GNDA.n2276 3.4105
R27665 GNDA.n2324 GNDA.n2276 3.4105
R27666 GNDA.n2649 GNDA.n2276 3.4105
R27667 GNDA.n2651 GNDA.n2276 3.4105
R27668 GNDA.n2653 GNDA.n2247 3.4105
R27669 GNDA.n2294 GNDA.n2247 3.4105
R27670 GNDA.n2296 GNDA.n2247 3.4105
R27671 GNDA.n2293 GNDA.n2247 3.4105
R27672 GNDA.n2298 GNDA.n2247 3.4105
R27673 GNDA.n2292 GNDA.n2247 3.4105
R27674 GNDA.n2300 GNDA.n2247 3.4105
R27675 GNDA.n2291 GNDA.n2247 3.4105
R27676 GNDA.n2302 GNDA.n2247 3.4105
R27677 GNDA.n2290 GNDA.n2247 3.4105
R27678 GNDA.n2304 GNDA.n2247 3.4105
R27679 GNDA.n2289 GNDA.n2247 3.4105
R27680 GNDA.n2306 GNDA.n2247 3.4105
R27681 GNDA.n2288 GNDA.n2247 3.4105
R27682 GNDA.n2308 GNDA.n2247 3.4105
R27683 GNDA.n2287 GNDA.n2247 3.4105
R27684 GNDA.n2310 GNDA.n2247 3.4105
R27685 GNDA.n2286 GNDA.n2247 3.4105
R27686 GNDA.n2312 GNDA.n2247 3.4105
R27687 GNDA.n2285 GNDA.n2247 3.4105
R27688 GNDA.n2314 GNDA.n2247 3.4105
R27689 GNDA.n2284 GNDA.n2247 3.4105
R27690 GNDA.n2316 GNDA.n2247 3.4105
R27691 GNDA.n2283 GNDA.n2247 3.4105
R27692 GNDA.n2318 GNDA.n2247 3.4105
R27693 GNDA.n2282 GNDA.n2247 3.4105
R27694 GNDA.n2320 GNDA.n2247 3.4105
R27695 GNDA.n2281 GNDA.n2247 3.4105
R27696 GNDA.n2322 GNDA.n2247 3.4105
R27697 GNDA.n2280 GNDA.n2247 3.4105
R27698 GNDA.n2324 GNDA.n2247 3.4105
R27699 GNDA.n2649 GNDA.n2247 3.4105
R27700 GNDA.n2651 GNDA.n2247 3.4105
R27701 GNDA.n2653 GNDA.n2277 3.4105
R27702 GNDA.n2294 GNDA.n2277 3.4105
R27703 GNDA.n2296 GNDA.n2277 3.4105
R27704 GNDA.n2293 GNDA.n2277 3.4105
R27705 GNDA.n2298 GNDA.n2277 3.4105
R27706 GNDA.n2292 GNDA.n2277 3.4105
R27707 GNDA.n2300 GNDA.n2277 3.4105
R27708 GNDA.n2291 GNDA.n2277 3.4105
R27709 GNDA.n2302 GNDA.n2277 3.4105
R27710 GNDA.n2290 GNDA.n2277 3.4105
R27711 GNDA.n2304 GNDA.n2277 3.4105
R27712 GNDA.n2289 GNDA.n2277 3.4105
R27713 GNDA.n2306 GNDA.n2277 3.4105
R27714 GNDA.n2288 GNDA.n2277 3.4105
R27715 GNDA.n2308 GNDA.n2277 3.4105
R27716 GNDA.n2287 GNDA.n2277 3.4105
R27717 GNDA.n2310 GNDA.n2277 3.4105
R27718 GNDA.n2286 GNDA.n2277 3.4105
R27719 GNDA.n2312 GNDA.n2277 3.4105
R27720 GNDA.n2285 GNDA.n2277 3.4105
R27721 GNDA.n2314 GNDA.n2277 3.4105
R27722 GNDA.n2284 GNDA.n2277 3.4105
R27723 GNDA.n2316 GNDA.n2277 3.4105
R27724 GNDA.n2283 GNDA.n2277 3.4105
R27725 GNDA.n2318 GNDA.n2277 3.4105
R27726 GNDA.n2282 GNDA.n2277 3.4105
R27727 GNDA.n2320 GNDA.n2277 3.4105
R27728 GNDA.n2281 GNDA.n2277 3.4105
R27729 GNDA.n2322 GNDA.n2277 3.4105
R27730 GNDA.n2280 GNDA.n2277 3.4105
R27731 GNDA.n2324 GNDA.n2277 3.4105
R27732 GNDA.n2649 GNDA.n2277 3.4105
R27733 GNDA.n2651 GNDA.n2277 3.4105
R27734 GNDA.n2653 GNDA.n2246 3.4105
R27735 GNDA.n2294 GNDA.n2246 3.4105
R27736 GNDA.n2296 GNDA.n2246 3.4105
R27737 GNDA.n2293 GNDA.n2246 3.4105
R27738 GNDA.n2298 GNDA.n2246 3.4105
R27739 GNDA.n2292 GNDA.n2246 3.4105
R27740 GNDA.n2300 GNDA.n2246 3.4105
R27741 GNDA.n2291 GNDA.n2246 3.4105
R27742 GNDA.n2302 GNDA.n2246 3.4105
R27743 GNDA.n2290 GNDA.n2246 3.4105
R27744 GNDA.n2304 GNDA.n2246 3.4105
R27745 GNDA.n2289 GNDA.n2246 3.4105
R27746 GNDA.n2306 GNDA.n2246 3.4105
R27747 GNDA.n2288 GNDA.n2246 3.4105
R27748 GNDA.n2308 GNDA.n2246 3.4105
R27749 GNDA.n2287 GNDA.n2246 3.4105
R27750 GNDA.n2310 GNDA.n2246 3.4105
R27751 GNDA.n2286 GNDA.n2246 3.4105
R27752 GNDA.n2312 GNDA.n2246 3.4105
R27753 GNDA.n2285 GNDA.n2246 3.4105
R27754 GNDA.n2314 GNDA.n2246 3.4105
R27755 GNDA.n2284 GNDA.n2246 3.4105
R27756 GNDA.n2316 GNDA.n2246 3.4105
R27757 GNDA.n2283 GNDA.n2246 3.4105
R27758 GNDA.n2318 GNDA.n2246 3.4105
R27759 GNDA.n2282 GNDA.n2246 3.4105
R27760 GNDA.n2320 GNDA.n2246 3.4105
R27761 GNDA.n2281 GNDA.n2246 3.4105
R27762 GNDA.n2322 GNDA.n2246 3.4105
R27763 GNDA.n2280 GNDA.n2246 3.4105
R27764 GNDA.n2324 GNDA.n2246 3.4105
R27765 GNDA.n2649 GNDA.n2246 3.4105
R27766 GNDA.n2651 GNDA.n2246 3.4105
R27767 GNDA.n2653 GNDA.n2278 3.4105
R27768 GNDA.n2294 GNDA.n2278 3.4105
R27769 GNDA.n2296 GNDA.n2278 3.4105
R27770 GNDA.n2293 GNDA.n2278 3.4105
R27771 GNDA.n2298 GNDA.n2278 3.4105
R27772 GNDA.n2292 GNDA.n2278 3.4105
R27773 GNDA.n2300 GNDA.n2278 3.4105
R27774 GNDA.n2291 GNDA.n2278 3.4105
R27775 GNDA.n2302 GNDA.n2278 3.4105
R27776 GNDA.n2290 GNDA.n2278 3.4105
R27777 GNDA.n2304 GNDA.n2278 3.4105
R27778 GNDA.n2289 GNDA.n2278 3.4105
R27779 GNDA.n2306 GNDA.n2278 3.4105
R27780 GNDA.n2288 GNDA.n2278 3.4105
R27781 GNDA.n2308 GNDA.n2278 3.4105
R27782 GNDA.n2287 GNDA.n2278 3.4105
R27783 GNDA.n2310 GNDA.n2278 3.4105
R27784 GNDA.n2286 GNDA.n2278 3.4105
R27785 GNDA.n2312 GNDA.n2278 3.4105
R27786 GNDA.n2285 GNDA.n2278 3.4105
R27787 GNDA.n2314 GNDA.n2278 3.4105
R27788 GNDA.n2284 GNDA.n2278 3.4105
R27789 GNDA.n2316 GNDA.n2278 3.4105
R27790 GNDA.n2283 GNDA.n2278 3.4105
R27791 GNDA.n2318 GNDA.n2278 3.4105
R27792 GNDA.n2282 GNDA.n2278 3.4105
R27793 GNDA.n2320 GNDA.n2278 3.4105
R27794 GNDA.n2281 GNDA.n2278 3.4105
R27795 GNDA.n2322 GNDA.n2278 3.4105
R27796 GNDA.n2280 GNDA.n2278 3.4105
R27797 GNDA.n2324 GNDA.n2278 3.4105
R27798 GNDA.n2649 GNDA.n2278 3.4105
R27799 GNDA.n2651 GNDA.n2278 3.4105
R27800 GNDA.n2653 GNDA.n2245 3.4105
R27801 GNDA.n2294 GNDA.n2245 3.4105
R27802 GNDA.n2296 GNDA.n2245 3.4105
R27803 GNDA.n2293 GNDA.n2245 3.4105
R27804 GNDA.n2298 GNDA.n2245 3.4105
R27805 GNDA.n2292 GNDA.n2245 3.4105
R27806 GNDA.n2300 GNDA.n2245 3.4105
R27807 GNDA.n2291 GNDA.n2245 3.4105
R27808 GNDA.n2302 GNDA.n2245 3.4105
R27809 GNDA.n2290 GNDA.n2245 3.4105
R27810 GNDA.n2304 GNDA.n2245 3.4105
R27811 GNDA.n2289 GNDA.n2245 3.4105
R27812 GNDA.n2306 GNDA.n2245 3.4105
R27813 GNDA.n2288 GNDA.n2245 3.4105
R27814 GNDA.n2308 GNDA.n2245 3.4105
R27815 GNDA.n2287 GNDA.n2245 3.4105
R27816 GNDA.n2310 GNDA.n2245 3.4105
R27817 GNDA.n2286 GNDA.n2245 3.4105
R27818 GNDA.n2312 GNDA.n2245 3.4105
R27819 GNDA.n2285 GNDA.n2245 3.4105
R27820 GNDA.n2314 GNDA.n2245 3.4105
R27821 GNDA.n2284 GNDA.n2245 3.4105
R27822 GNDA.n2316 GNDA.n2245 3.4105
R27823 GNDA.n2283 GNDA.n2245 3.4105
R27824 GNDA.n2318 GNDA.n2245 3.4105
R27825 GNDA.n2282 GNDA.n2245 3.4105
R27826 GNDA.n2320 GNDA.n2245 3.4105
R27827 GNDA.n2281 GNDA.n2245 3.4105
R27828 GNDA.n2322 GNDA.n2245 3.4105
R27829 GNDA.n2280 GNDA.n2245 3.4105
R27830 GNDA.n2324 GNDA.n2245 3.4105
R27831 GNDA.n2649 GNDA.n2245 3.4105
R27832 GNDA.n2651 GNDA.n2245 3.4105
R27833 GNDA.n2653 GNDA.n2652 3.4105
R27834 GNDA.n2652 GNDA.n2294 3.4105
R27835 GNDA.n2652 GNDA.n2296 3.4105
R27836 GNDA.n2652 GNDA.n2293 3.4105
R27837 GNDA.n2652 GNDA.n2298 3.4105
R27838 GNDA.n2652 GNDA.n2292 3.4105
R27839 GNDA.n2652 GNDA.n2300 3.4105
R27840 GNDA.n2652 GNDA.n2291 3.4105
R27841 GNDA.n2652 GNDA.n2302 3.4105
R27842 GNDA.n2652 GNDA.n2290 3.4105
R27843 GNDA.n2652 GNDA.n2304 3.4105
R27844 GNDA.n2652 GNDA.n2289 3.4105
R27845 GNDA.n2652 GNDA.n2306 3.4105
R27846 GNDA.n2652 GNDA.n2288 3.4105
R27847 GNDA.n2652 GNDA.n2308 3.4105
R27848 GNDA.n2652 GNDA.n2287 3.4105
R27849 GNDA.n2652 GNDA.n2310 3.4105
R27850 GNDA.n2652 GNDA.n2286 3.4105
R27851 GNDA.n2652 GNDA.n2312 3.4105
R27852 GNDA.n2652 GNDA.n2285 3.4105
R27853 GNDA.n2652 GNDA.n2314 3.4105
R27854 GNDA.n2652 GNDA.n2284 3.4105
R27855 GNDA.n2652 GNDA.n2316 3.4105
R27856 GNDA.n2652 GNDA.n2283 3.4105
R27857 GNDA.n2652 GNDA.n2318 3.4105
R27858 GNDA.n2652 GNDA.n2282 3.4105
R27859 GNDA.n2652 GNDA.n2320 3.4105
R27860 GNDA.n2652 GNDA.n2281 3.4105
R27861 GNDA.n2652 GNDA.n2322 3.4105
R27862 GNDA.n2652 GNDA.n2280 3.4105
R27863 GNDA.n2652 GNDA.n2324 3.4105
R27864 GNDA.n2652 GNDA.n2651 3.4105
R27865 GNDA.n2408 GNDA.n2359 3.4105
R27866 GNDA.n2408 GNDA.n2376 3.4105
R27867 GNDA.n2614 GNDA.n2408 3.4105
R27868 GNDA.n2566 GNDA.n2361 3.4105
R27869 GNDA.n2566 GNDA.n2358 3.4105
R27870 GNDA.n2566 GNDA.n2362 3.4105
R27871 GNDA.n2566 GNDA.n2357 3.4105
R27872 GNDA.n2566 GNDA.n2363 3.4105
R27873 GNDA.n2566 GNDA.n2356 3.4105
R27874 GNDA.n2566 GNDA.n2364 3.4105
R27875 GNDA.n2566 GNDA.n2355 3.4105
R27876 GNDA.n2566 GNDA.n2365 3.4105
R27877 GNDA.n2566 GNDA.n2354 3.4105
R27878 GNDA.n2566 GNDA.n2366 3.4105
R27879 GNDA.n2566 GNDA.n2353 3.4105
R27880 GNDA.n2566 GNDA.n2367 3.4105
R27881 GNDA.n2566 GNDA.n2352 3.4105
R27882 GNDA.n2566 GNDA.n2368 3.4105
R27883 GNDA.n2566 GNDA.n2351 3.4105
R27884 GNDA.n2566 GNDA.n2369 3.4105
R27885 GNDA.n2566 GNDA.n2350 3.4105
R27886 GNDA.n2566 GNDA.n2370 3.4105
R27887 GNDA.n2566 GNDA.n2349 3.4105
R27888 GNDA.n2566 GNDA.n2371 3.4105
R27889 GNDA.n2566 GNDA.n2348 3.4105
R27890 GNDA.n2566 GNDA.n2372 3.4105
R27891 GNDA.n2566 GNDA.n2347 3.4105
R27892 GNDA.n2566 GNDA.n2373 3.4105
R27893 GNDA.n2566 GNDA.n2346 3.4105
R27894 GNDA.n2566 GNDA.n2374 3.4105
R27895 GNDA.n2566 GNDA.n2345 3.4105
R27896 GNDA.n2566 GNDA.n2375 3.4105
R27897 GNDA.n2566 GNDA.n2376 3.4105
R27898 GNDA.n2614 GNDA.n2566 3.4105
R27899 GNDA.n2392 GNDA.n2360 3.4105
R27900 GNDA.n2392 GNDA.n2359 3.4105
R27901 GNDA.n2392 GNDA.n2361 3.4105
R27902 GNDA.n2392 GNDA.n2358 3.4105
R27903 GNDA.n2392 GNDA.n2362 3.4105
R27904 GNDA.n2392 GNDA.n2357 3.4105
R27905 GNDA.n2392 GNDA.n2363 3.4105
R27906 GNDA.n2392 GNDA.n2356 3.4105
R27907 GNDA.n2392 GNDA.n2364 3.4105
R27908 GNDA.n2392 GNDA.n2355 3.4105
R27909 GNDA.n2392 GNDA.n2365 3.4105
R27910 GNDA.n2392 GNDA.n2354 3.4105
R27911 GNDA.n2392 GNDA.n2366 3.4105
R27912 GNDA.n2392 GNDA.n2353 3.4105
R27913 GNDA.n2392 GNDA.n2367 3.4105
R27914 GNDA.n2392 GNDA.n2352 3.4105
R27915 GNDA.n2392 GNDA.n2368 3.4105
R27916 GNDA.n2392 GNDA.n2351 3.4105
R27917 GNDA.n2392 GNDA.n2369 3.4105
R27918 GNDA.n2392 GNDA.n2350 3.4105
R27919 GNDA.n2392 GNDA.n2370 3.4105
R27920 GNDA.n2392 GNDA.n2349 3.4105
R27921 GNDA.n2392 GNDA.n2371 3.4105
R27922 GNDA.n2392 GNDA.n2348 3.4105
R27923 GNDA.n2392 GNDA.n2372 3.4105
R27924 GNDA.n2392 GNDA.n2347 3.4105
R27925 GNDA.n2392 GNDA.n2373 3.4105
R27926 GNDA.n2392 GNDA.n2346 3.4105
R27927 GNDA.n2392 GNDA.n2374 3.4105
R27928 GNDA.n2392 GNDA.n2345 3.4105
R27929 GNDA.n2392 GNDA.n2375 3.4105
R27930 GNDA.n2392 GNDA.n2376 3.4105
R27931 GNDA.n2614 GNDA.n2392 3.4105
R27932 GNDA.n2568 GNDA.n2360 3.4105
R27933 GNDA.n2568 GNDA.n2359 3.4105
R27934 GNDA.n2568 GNDA.n2361 3.4105
R27935 GNDA.n2568 GNDA.n2358 3.4105
R27936 GNDA.n2568 GNDA.n2362 3.4105
R27937 GNDA.n2568 GNDA.n2357 3.4105
R27938 GNDA.n2568 GNDA.n2363 3.4105
R27939 GNDA.n2568 GNDA.n2356 3.4105
R27940 GNDA.n2568 GNDA.n2364 3.4105
R27941 GNDA.n2568 GNDA.n2355 3.4105
R27942 GNDA.n2568 GNDA.n2365 3.4105
R27943 GNDA.n2568 GNDA.n2354 3.4105
R27944 GNDA.n2568 GNDA.n2366 3.4105
R27945 GNDA.n2568 GNDA.n2353 3.4105
R27946 GNDA.n2568 GNDA.n2367 3.4105
R27947 GNDA.n2568 GNDA.n2352 3.4105
R27948 GNDA.n2568 GNDA.n2368 3.4105
R27949 GNDA.n2568 GNDA.n2351 3.4105
R27950 GNDA.n2568 GNDA.n2369 3.4105
R27951 GNDA.n2568 GNDA.n2350 3.4105
R27952 GNDA.n2568 GNDA.n2370 3.4105
R27953 GNDA.n2568 GNDA.n2349 3.4105
R27954 GNDA.n2568 GNDA.n2371 3.4105
R27955 GNDA.n2568 GNDA.n2348 3.4105
R27956 GNDA.n2568 GNDA.n2372 3.4105
R27957 GNDA.n2568 GNDA.n2347 3.4105
R27958 GNDA.n2568 GNDA.n2373 3.4105
R27959 GNDA.n2568 GNDA.n2346 3.4105
R27960 GNDA.n2568 GNDA.n2374 3.4105
R27961 GNDA.n2568 GNDA.n2345 3.4105
R27962 GNDA.n2568 GNDA.n2375 3.4105
R27963 GNDA.n2568 GNDA.n2376 3.4105
R27964 GNDA.n2614 GNDA.n2568 3.4105
R27965 GNDA.n2391 GNDA.n2360 3.4105
R27966 GNDA.n2391 GNDA.n2359 3.4105
R27967 GNDA.n2391 GNDA.n2361 3.4105
R27968 GNDA.n2391 GNDA.n2358 3.4105
R27969 GNDA.n2391 GNDA.n2362 3.4105
R27970 GNDA.n2391 GNDA.n2357 3.4105
R27971 GNDA.n2391 GNDA.n2363 3.4105
R27972 GNDA.n2391 GNDA.n2356 3.4105
R27973 GNDA.n2391 GNDA.n2364 3.4105
R27974 GNDA.n2391 GNDA.n2355 3.4105
R27975 GNDA.n2391 GNDA.n2365 3.4105
R27976 GNDA.n2391 GNDA.n2354 3.4105
R27977 GNDA.n2391 GNDA.n2366 3.4105
R27978 GNDA.n2391 GNDA.n2353 3.4105
R27979 GNDA.n2391 GNDA.n2367 3.4105
R27980 GNDA.n2391 GNDA.n2352 3.4105
R27981 GNDA.n2391 GNDA.n2368 3.4105
R27982 GNDA.n2391 GNDA.n2351 3.4105
R27983 GNDA.n2391 GNDA.n2369 3.4105
R27984 GNDA.n2391 GNDA.n2350 3.4105
R27985 GNDA.n2391 GNDA.n2370 3.4105
R27986 GNDA.n2391 GNDA.n2349 3.4105
R27987 GNDA.n2391 GNDA.n2371 3.4105
R27988 GNDA.n2391 GNDA.n2348 3.4105
R27989 GNDA.n2391 GNDA.n2372 3.4105
R27990 GNDA.n2391 GNDA.n2347 3.4105
R27991 GNDA.n2391 GNDA.n2373 3.4105
R27992 GNDA.n2391 GNDA.n2346 3.4105
R27993 GNDA.n2391 GNDA.n2374 3.4105
R27994 GNDA.n2391 GNDA.n2345 3.4105
R27995 GNDA.n2391 GNDA.n2375 3.4105
R27996 GNDA.n2391 GNDA.n2376 3.4105
R27997 GNDA.n2614 GNDA.n2391 3.4105
R27998 GNDA.n2570 GNDA.n2360 3.4105
R27999 GNDA.n2570 GNDA.n2359 3.4105
R28000 GNDA.n2570 GNDA.n2361 3.4105
R28001 GNDA.n2570 GNDA.n2358 3.4105
R28002 GNDA.n2570 GNDA.n2362 3.4105
R28003 GNDA.n2570 GNDA.n2357 3.4105
R28004 GNDA.n2570 GNDA.n2363 3.4105
R28005 GNDA.n2570 GNDA.n2356 3.4105
R28006 GNDA.n2570 GNDA.n2364 3.4105
R28007 GNDA.n2570 GNDA.n2355 3.4105
R28008 GNDA.n2570 GNDA.n2365 3.4105
R28009 GNDA.n2570 GNDA.n2354 3.4105
R28010 GNDA.n2570 GNDA.n2366 3.4105
R28011 GNDA.n2570 GNDA.n2353 3.4105
R28012 GNDA.n2570 GNDA.n2367 3.4105
R28013 GNDA.n2570 GNDA.n2352 3.4105
R28014 GNDA.n2570 GNDA.n2368 3.4105
R28015 GNDA.n2570 GNDA.n2351 3.4105
R28016 GNDA.n2570 GNDA.n2369 3.4105
R28017 GNDA.n2570 GNDA.n2350 3.4105
R28018 GNDA.n2570 GNDA.n2370 3.4105
R28019 GNDA.n2570 GNDA.n2349 3.4105
R28020 GNDA.n2570 GNDA.n2371 3.4105
R28021 GNDA.n2570 GNDA.n2348 3.4105
R28022 GNDA.n2570 GNDA.n2372 3.4105
R28023 GNDA.n2570 GNDA.n2347 3.4105
R28024 GNDA.n2570 GNDA.n2373 3.4105
R28025 GNDA.n2570 GNDA.n2346 3.4105
R28026 GNDA.n2570 GNDA.n2374 3.4105
R28027 GNDA.n2570 GNDA.n2345 3.4105
R28028 GNDA.n2570 GNDA.n2375 3.4105
R28029 GNDA.n2570 GNDA.n2376 3.4105
R28030 GNDA.n2614 GNDA.n2570 3.4105
R28031 GNDA.n2390 GNDA.n2360 3.4105
R28032 GNDA.n2390 GNDA.n2359 3.4105
R28033 GNDA.n2390 GNDA.n2361 3.4105
R28034 GNDA.n2390 GNDA.n2358 3.4105
R28035 GNDA.n2390 GNDA.n2362 3.4105
R28036 GNDA.n2390 GNDA.n2357 3.4105
R28037 GNDA.n2390 GNDA.n2363 3.4105
R28038 GNDA.n2390 GNDA.n2356 3.4105
R28039 GNDA.n2390 GNDA.n2364 3.4105
R28040 GNDA.n2390 GNDA.n2355 3.4105
R28041 GNDA.n2390 GNDA.n2365 3.4105
R28042 GNDA.n2390 GNDA.n2354 3.4105
R28043 GNDA.n2390 GNDA.n2366 3.4105
R28044 GNDA.n2390 GNDA.n2353 3.4105
R28045 GNDA.n2390 GNDA.n2367 3.4105
R28046 GNDA.n2390 GNDA.n2352 3.4105
R28047 GNDA.n2390 GNDA.n2368 3.4105
R28048 GNDA.n2390 GNDA.n2351 3.4105
R28049 GNDA.n2390 GNDA.n2369 3.4105
R28050 GNDA.n2390 GNDA.n2350 3.4105
R28051 GNDA.n2390 GNDA.n2370 3.4105
R28052 GNDA.n2390 GNDA.n2349 3.4105
R28053 GNDA.n2390 GNDA.n2371 3.4105
R28054 GNDA.n2390 GNDA.n2348 3.4105
R28055 GNDA.n2390 GNDA.n2372 3.4105
R28056 GNDA.n2390 GNDA.n2347 3.4105
R28057 GNDA.n2390 GNDA.n2373 3.4105
R28058 GNDA.n2390 GNDA.n2346 3.4105
R28059 GNDA.n2390 GNDA.n2374 3.4105
R28060 GNDA.n2390 GNDA.n2345 3.4105
R28061 GNDA.n2390 GNDA.n2375 3.4105
R28062 GNDA.n2390 GNDA.n2376 3.4105
R28063 GNDA.n2614 GNDA.n2390 3.4105
R28064 GNDA.n2572 GNDA.n2360 3.4105
R28065 GNDA.n2572 GNDA.n2359 3.4105
R28066 GNDA.n2572 GNDA.n2361 3.4105
R28067 GNDA.n2572 GNDA.n2358 3.4105
R28068 GNDA.n2572 GNDA.n2362 3.4105
R28069 GNDA.n2572 GNDA.n2357 3.4105
R28070 GNDA.n2572 GNDA.n2363 3.4105
R28071 GNDA.n2572 GNDA.n2356 3.4105
R28072 GNDA.n2572 GNDA.n2364 3.4105
R28073 GNDA.n2572 GNDA.n2355 3.4105
R28074 GNDA.n2572 GNDA.n2365 3.4105
R28075 GNDA.n2572 GNDA.n2354 3.4105
R28076 GNDA.n2572 GNDA.n2366 3.4105
R28077 GNDA.n2572 GNDA.n2353 3.4105
R28078 GNDA.n2572 GNDA.n2367 3.4105
R28079 GNDA.n2572 GNDA.n2352 3.4105
R28080 GNDA.n2572 GNDA.n2368 3.4105
R28081 GNDA.n2572 GNDA.n2351 3.4105
R28082 GNDA.n2572 GNDA.n2369 3.4105
R28083 GNDA.n2572 GNDA.n2350 3.4105
R28084 GNDA.n2572 GNDA.n2370 3.4105
R28085 GNDA.n2572 GNDA.n2349 3.4105
R28086 GNDA.n2572 GNDA.n2371 3.4105
R28087 GNDA.n2572 GNDA.n2348 3.4105
R28088 GNDA.n2572 GNDA.n2372 3.4105
R28089 GNDA.n2572 GNDA.n2347 3.4105
R28090 GNDA.n2572 GNDA.n2373 3.4105
R28091 GNDA.n2572 GNDA.n2346 3.4105
R28092 GNDA.n2572 GNDA.n2374 3.4105
R28093 GNDA.n2572 GNDA.n2345 3.4105
R28094 GNDA.n2572 GNDA.n2375 3.4105
R28095 GNDA.n2572 GNDA.n2376 3.4105
R28096 GNDA.n2614 GNDA.n2572 3.4105
R28097 GNDA.n2389 GNDA.n2360 3.4105
R28098 GNDA.n2389 GNDA.n2359 3.4105
R28099 GNDA.n2389 GNDA.n2361 3.4105
R28100 GNDA.n2389 GNDA.n2358 3.4105
R28101 GNDA.n2389 GNDA.n2362 3.4105
R28102 GNDA.n2389 GNDA.n2357 3.4105
R28103 GNDA.n2389 GNDA.n2363 3.4105
R28104 GNDA.n2389 GNDA.n2356 3.4105
R28105 GNDA.n2389 GNDA.n2364 3.4105
R28106 GNDA.n2389 GNDA.n2355 3.4105
R28107 GNDA.n2389 GNDA.n2365 3.4105
R28108 GNDA.n2389 GNDA.n2354 3.4105
R28109 GNDA.n2389 GNDA.n2366 3.4105
R28110 GNDA.n2389 GNDA.n2353 3.4105
R28111 GNDA.n2389 GNDA.n2367 3.4105
R28112 GNDA.n2389 GNDA.n2352 3.4105
R28113 GNDA.n2389 GNDA.n2368 3.4105
R28114 GNDA.n2389 GNDA.n2351 3.4105
R28115 GNDA.n2389 GNDA.n2369 3.4105
R28116 GNDA.n2389 GNDA.n2350 3.4105
R28117 GNDA.n2389 GNDA.n2370 3.4105
R28118 GNDA.n2389 GNDA.n2349 3.4105
R28119 GNDA.n2389 GNDA.n2371 3.4105
R28120 GNDA.n2389 GNDA.n2348 3.4105
R28121 GNDA.n2389 GNDA.n2372 3.4105
R28122 GNDA.n2389 GNDA.n2347 3.4105
R28123 GNDA.n2389 GNDA.n2373 3.4105
R28124 GNDA.n2389 GNDA.n2346 3.4105
R28125 GNDA.n2389 GNDA.n2374 3.4105
R28126 GNDA.n2389 GNDA.n2345 3.4105
R28127 GNDA.n2389 GNDA.n2375 3.4105
R28128 GNDA.n2389 GNDA.n2376 3.4105
R28129 GNDA.n2614 GNDA.n2389 3.4105
R28130 GNDA.n2574 GNDA.n2360 3.4105
R28131 GNDA.n2574 GNDA.n2359 3.4105
R28132 GNDA.n2574 GNDA.n2361 3.4105
R28133 GNDA.n2574 GNDA.n2358 3.4105
R28134 GNDA.n2574 GNDA.n2362 3.4105
R28135 GNDA.n2574 GNDA.n2357 3.4105
R28136 GNDA.n2574 GNDA.n2363 3.4105
R28137 GNDA.n2574 GNDA.n2356 3.4105
R28138 GNDA.n2574 GNDA.n2364 3.4105
R28139 GNDA.n2574 GNDA.n2355 3.4105
R28140 GNDA.n2574 GNDA.n2365 3.4105
R28141 GNDA.n2574 GNDA.n2354 3.4105
R28142 GNDA.n2574 GNDA.n2366 3.4105
R28143 GNDA.n2574 GNDA.n2353 3.4105
R28144 GNDA.n2574 GNDA.n2367 3.4105
R28145 GNDA.n2574 GNDA.n2352 3.4105
R28146 GNDA.n2574 GNDA.n2368 3.4105
R28147 GNDA.n2574 GNDA.n2351 3.4105
R28148 GNDA.n2574 GNDA.n2369 3.4105
R28149 GNDA.n2574 GNDA.n2350 3.4105
R28150 GNDA.n2574 GNDA.n2370 3.4105
R28151 GNDA.n2574 GNDA.n2349 3.4105
R28152 GNDA.n2574 GNDA.n2371 3.4105
R28153 GNDA.n2574 GNDA.n2348 3.4105
R28154 GNDA.n2574 GNDA.n2372 3.4105
R28155 GNDA.n2574 GNDA.n2347 3.4105
R28156 GNDA.n2574 GNDA.n2373 3.4105
R28157 GNDA.n2574 GNDA.n2346 3.4105
R28158 GNDA.n2574 GNDA.n2374 3.4105
R28159 GNDA.n2574 GNDA.n2345 3.4105
R28160 GNDA.n2574 GNDA.n2375 3.4105
R28161 GNDA.n2574 GNDA.n2376 3.4105
R28162 GNDA.n2614 GNDA.n2574 3.4105
R28163 GNDA.n2388 GNDA.n2360 3.4105
R28164 GNDA.n2388 GNDA.n2359 3.4105
R28165 GNDA.n2388 GNDA.n2361 3.4105
R28166 GNDA.n2388 GNDA.n2358 3.4105
R28167 GNDA.n2388 GNDA.n2362 3.4105
R28168 GNDA.n2388 GNDA.n2357 3.4105
R28169 GNDA.n2388 GNDA.n2363 3.4105
R28170 GNDA.n2388 GNDA.n2356 3.4105
R28171 GNDA.n2388 GNDA.n2364 3.4105
R28172 GNDA.n2388 GNDA.n2355 3.4105
R28173 GNDA.n2388 GNDA.n2365 3.4105
R28174 GNDA.n2388 GNDA.n2354 3.4105
R28175 GNDA.n2388 GNDA.n2366 3.4105
R28176 GNDA.n2388 GNDA.n2353 3.4105
R28177 GNDA.n2388 GNDA.n2367 3.4105
R28178 GNDA.n2388 GNDA.n2352 3.4105
R28179 GNDA.n2388 GNDA.n2368 3.4105
R28180 GNDA.n2388 GNDA.n2351 3.4105
R28181 GNDA.n2388 GNDA.n2369 3.4105
R28182 GNDA.n2388 GNDA.n2350 3.4105
R28183 GNDA.n2388 GNDA.n2370 3.4105
R28184 GNDA.n2388 GNDA.n2349 3.4105
R28185 GNDA.n2388 GNDA.n2371 3.4105
R28186 GNDA.n2388 GNDA.n2348 3.4105
R28187 GNDA.n2388 GNDA.n2372 3.4105
R28188 GNDA.n2388 GNDA.n2347 3.4105
R28189 GNDA.n2388 GNDA.n2373 3.4105
R28190 GNDA.n2388 GNDA.n2346 3.4105
R28191 GNDA.n2388 GNDA.n2374 3.4105
R28192 GNDA.n2388 GNDA.n2345 3.4105
R28193 GNDA.n2388 GNDA.n2375 3.4105
R28194 GNDA.n2388 GNDA.n2376 3.4105
R28195 GNDA.n2614 GNDA.n2388 3.4105
R28196 GNDA.n2576 GNDA.n2360 3.4105
R28197 GNDA.n2576 GNDA.n2359 3.4105
R28198 GNDA.n2576 GNDA.n2361 3.4105
R28199 GNDA.n2576 GNDA.n2358 3.4105
R28200 GNDA.n2576 GNDA.n2362 3.4105
R28201 GNDA.n2576 GNDA.n2357 3.4105
R28202 GNDA.n2576 GNDA.n2363 3.4105
R28203 GNDA.n2576 GNDA.n2356 3.4105
R28204 GNDA.n2576 GNDA.n2364 3.4105
R28205 GNDA.n2576 GNDA.n2355 3.4105
R28206 GNDA.n2576 GNDA.n2365 3.4105
R28207 GNDA.n2576 GNDA.n2354 3.4105
R28208 GNDA.n2576 GNDA.n2366 3.4105
R28209 GNDA.n2576 GNDA.n2353 3.4105
R28210 GNDA.n2576 GNDA.n2367 3.4105
R28211 GNDA.n2576 GNDA.n2352 3.4105
R28212 GNDA.n2576 GNDA.n2368 3.4105
R28213 GNDA.n2576 GNDA.n2351 3.4105
R28214 GNDA.n2576 GNDA.n2369 3.4105
R28215 GNDA.n2576 GNDA.n2350 3.4105
R28216 GNDA.n2576 GNDA.n2370 3.4105
R28217 GNDA.n2576 GNDA.n2349 3.4105
R28218 GNDA.n2576 GNDA.n2371 3.4105
R28219 GNDA.n2576 GNDA.n2348 3.4105
R28220 GNDA.n2576 GNDA.n2372 3.4105
R28221 GNDA.n2576 GNDA.n2347 3.4105
R28222 GNDA.n2576 GNDA.n2373 3.4105
R28223 GNDA.n2576 GNDA.n2346 3.4105
R28224 GNDA.n2576 GNDA.n2374 3.4105
R28225 GNDA.n2576 GNDA.n2345 3.4105
R28226 GNDA.n2576 GNDA.n2375 3.4105
R28227 GNDA.n2576 GNDA.n2376 3.4105
R28228 GNDA.n2614 GNDA.n2576 3.4105
R28229 GNDA.n2387 GNDA.n2360 3.4105
R28230 GNDA.n2387 GNDA.n2359 3.4105
R28231 GNDA.n2387 GNDA.n2361 3.4105
R28232 GNDA.n2387 GNDA.n2358 3.4105
R28233 GNDA.n2387 GNDA.n2362 3.4105
R28234 GNDA.n2387 GNDA.n2357 3.4105
R28235 GNDA.n2387 GNDA.n2363 3.4105
R28236 GNDA.n2387 GNDA.n2356 3.4105
R28237 GNDA.n2387 GNDA.n2364 3.4105
R28238 GNDA.n2387 GNDA.n2355 3.4105
R28239 GNDA.n2387 GNDA.n2365 3.4105
R28240 GNDA.n2387 GNDA.n2354 3.4105
R28241 GNDA.n2387 GNDA.n2366 3.4105
R28242 GNDA.n2387 GNDA.n2353 3.4105
R28243 GNDA.n2387 GNDA.n2367 3.4105
R28244 GNDA.n2387 GNDA.n2352 3.4105
R28245 GNDA.n2387 GNDA.n2368 3.4105
R28246 GNDA.n2387 GNDA.n2351 3.4105
R28247 GNDA.n2387 GNDA.n2369 3.4105
R28248 GNDA.n2387 GNDA.n2350 3.4105
R28249 GNDA.n2387 GNDA.n2370 3.4105
R28250 GNDA.n2387 GNDA.n2349 3.4105
R28251 GNDA.n2387 GNDA.n2371 3.4105
R28252 GNDA.n2387 GNDA.n2348 3.4105
R28253 GNDA.n2387 GNDA.n2372 3.4105
R28254 GNDA.n2387 GNDA.n2347 3.4105
R28255 GNDA.n2387 GNDA.n2373 3.4105
R28256 GNDA.n2387 GNDA.n2346 3.4105
R28257 GNDA.n2387 GNDA.n2374 3.4105
R28258 GNDA.n2387 GNDA.n2345 3.4105
R28259 GNDA.n2387 GNDA.n2375 3.4105
R28260 GNDA.n2387 GNDA.n2376 3.4105
R28261 GNDA.n2614 GNDA.n2387 3.4105
R28262 GNDA.n2578 GNDA.n2360 3.4105
R28263 GNDA.n2578 GNDA.n2359 3.4105
R28264 GNDA.n2578 GNDA.n2361 3.4105
R28265 GNDA.n2578 GNDA.n2358 3.4105
R28266 GNDA.n2578 GNDA.n2362 3.4105
R28267 GNDA.n2578 GNDA.n2357 3.4105
R28268 GNDA.n2578 GNDA.n2363 3.4105
R28269 GNDA.n2578 GNDA.n2356 3.4105
R28270 GNDA.n2578 GNDA.n2364 3.4105
R28271 GNDA.n2578 GNDA.n2355 3.4105
R28272 GNDA.n2578 GNDA.n2365 3.4105
R28273 GNDA.n2578 GNDA.n2354 3.4105
R28274 GNDA.n2578 GNDA.n2366 3.4105
R28275 GNDA.n2578 GNDA.n2353 3.4105
R28276 GNDA.n2578 GNDA.n2367 3.4105
R28277 GNDA.n2578 GNDA.n2352 3.4105
R28278 GNDA.n2578 GNDA.n2368 3.4105
R28279 GNDA.n2578 GNDA.n2351 3.4105
R28280 GNDA.n2578 GNDA.n2369 3.4105
R28281 GNDA.n2578 GNDA.n2350 3.4105
R28282 GNDA.n2578 GNDA.n2370 3.4105
R28283 GNDA.n2578 GNDA.n2349 3.4105
R28284 GNDA.n2578 GNDA.n2371 3.4105
R28285 GNDA.n2578 GNDA.n2348 3.4105
R28286 GNDA.n2578 GNDA.n2372 3.4105
R28287 GNDA.n2578 GNDA.n2347 3.4105
R28288 GNDA.n2578 GNDA.n2373 3.4105
R28289 GNDA.n2578 GNDA.n2346 3.4105
R28290 GNDA.n2578 GNDA.n2374 3.4105
R28291 GNDA.n2578 GNDA.n2345 3.4105
R28292 GNDA.n2578 GNDA.n2375 3.4105
R28293 GNDA.n2578 GNDA.n2376 3.4105
R28294 GNDA.n2614 GNDA.n2578 3.4105
R28295 GNDA.n2386 GNDA.n2360 3.4105
R28296 GNDA.n2386 GNDA.n2359 3.4105
R28297 GNDA.n2386 GNDA.n2361 3.4105
R28298 GNDA.n2386 GNDA.n2358 3.4105
R28299 GNDA.n2386 GNDA.n2362 3.4105
R28300 GNDA.n2386 GNDA.n2357 3.4105
R28301 GNDA.n2386 GNDA.n2363 3.4105
R28302 GNDA.n2386 GNDA.n2356 3.4105
R28303 GNDA.n2386 GNDA.n2364 3.4105
R28304 GNDA.n2386 GNDA.n2355 3.4105
R28305 GNDA.n2386 GNDA.n2365 3.4105
R28306 GNDA.n2386 GNDA.n2354 3.4105
R28307 GNDA.n2386 GNDA.n2366 3.4105
R28308 GNDA.n2386 GNDA.n2353 3.4105
R28309 GNDA.n2386 GNDA.n2367 3.4105
R28310 GNDA.n2386 GNDA.n2352 3.4105
R28311 GNDA.n2386 GNDA.n2368 3.4105
R28312 GNDA.n2386 GNDA.n2351 3.4105
R28313 GNDA.n2386 GNDA.n2369 3.4105
R28314 GNDA.n2386 GNDA.n2350 3.4105
R28315 GNDA.n2386 GNDA.n2370 3.4105
R28316 GNDA.n2386 GNDA.n2349 3.4105
R28317 GNDA.n2386 GNDA.n2371 3.4105
R28318 GNDA.n2386 GNDA.n2348 3.4105
R28319 GNDA.n2386 GNDA.n2372 3.4105
R28320 GNDA.n2386 GNDA.n2347 3.4105
R28321 GNDA.n2386 GNDA.n2373 3.4105
R28322 GNDA.n2386 GNDA.n2346 3.4105
R28323 GNDA.n2386 GNDA.n2374 3.4105
R28324 GNDA.n2386 GNDA.n2345 3.4105
R28325 GNDA.n2386 GNDA.n2375 3.4105
R28326 GNDA.n2386 GNDA.n2376 3.4105
R28327 GNDA.n2614 GNDA.n2386 3.4105
R28328 GNDA.n2580 GNDA.n2360 3.4105
R28329 GNDA.n2580 GNDA.n2359 3.4105
R28330 GNDA.n2580 GNDA.n2361 3.4105
R28331 GNDA.n2580 GNDA.n2358 3.4105
R28332 GNDA.n2580 GNDA.n2362 3.4105
R28333 GNDA.n2580 GNDA.n2357 3.4105
R28334 GNDA.n2580 GNDA.n2363 3.4105
R28335 GNDA.n2580 GNDA.n2356 3.4105
R28336 GNDA.n2580 GNDA.n2364 3.4105
R28337 GNDA.n2580 GNDA.n2355 3.4105
R28338 GNDA.n2580 GNDA.n2365 3.4105
R28339 GNDA.n2580 GNDA.n2354 3.4105
R28340 GNDA.n2580 GNDA.n2366 3.4105
R28341 GNDA.n2580 GNDA.n2353 3.4105
R28342 GNDA.n2580 GNDA.n2367 3.4105
R28343 GNDA.n2580 GNDA.n2352 3.4105
R28344 GNDA.n2580 GNDA.n2368 3.4105
R28345 GNDA.n2580 GNDA.n2351 3.4105
R28346 GNDA.n2580 GNDA.n2369 3.4105
R28347 GNDA.n2580 GNDA.n2350 3.4105
R28348 GNDA.n2580 GNDA.n2370 3.4105
R28349 GNDA.n2580 GNDA.n2349 3.4105
R28350 GNDA.n2580 GNDA.n2371 3.4105
R28351 GNDA.n2580 GNDA.n2348 3.4105
R28352 GNDA.n2580 GNDA.n2372 3.4105
R28353 GNDA.n2580 GNDA.n2347 3.4105
R28354 GNDA.n2580 GNDA.n2373 3.4105
R28355 GNDA.n2580 GNDA.n2346 3.4105
R28356 GNDA.n2580 GNDA.n2374 3.4105
R28357 GNDA.n2580 GNDA.n2345 3.4105
R28358 GNDA.n2580 GNDA.n2375 3.4105
R28359 GNDA.n2580 GNDA.n2376 3.4105
R28360 GNDA.n2614 GNDA.n2580 3.4105
R28361 GNDA.n2385 GNDA.n2360 3.4105
R28362 GNDA.n2385 GNDA.n2359 3.4105
R28363 GNDA.n2385 GNDA.n2361 3.4105
R28364 GNDA.n2385 GNDA.n2358 3.4105
R28365 GNDA.n2385 GNDA.n2362 3.4105
R28366 GNDA.n2385 GNDA.n2357 3.4105
R28367 GNDA.n2385 GNDA.n2363 3.4105
R28368 GNDA.n2385 GNDA.n2356 3.4105
R28369 GNDA.n2385 GNDA.n2364 3.4105
R28370 GNDA.n2385 GNDA.n2355 3.4105
R28371 GNDA.n2385 GNDA.n2365 3.4105
R28372 GNDA.n2385 GNDA.n2354 3.4105
R28373 GNDA.n2385 GNDA.n2366 3.4105
R28374 GNDA.n2385 GNDA.n2353 3.4105
R28375 GNDA.n2385 GNDA.n2367 3.4105
R28376 GNDA.n2385 GNDA.n2352 3.4105
R28377 GNDA.n2385 GNDA.n2368 3.4105
R28378 GNDA.n2385 GNDA.n2351 3.4105
R28379 GNDA.n2385 GNDA.n2369 3.4105
R28380 GNDA.n2385 GNDA.n2350 3.4105
R28381 GNDA.n2385 GNDA.n2370 3.4105
R28382 GNDA.n2385 GNDA.n2349 3.4105
R28383 GNDA.n2385 GNDA.n2371 3.4105
R28384 GNDA.n2385 GNDA.n2348 3.4105
R28385 GNDA.n2385 GNDA.n2372 3.4105
R28386 GNDA.n2385 GNDA.n2347 3.4105
R28387 GNDA.n2385 GNDA.n2373 3.4105
R28388 GNDA.n2385 GNDA.n2346 3.4105
R28389 GNDA.n2385 GNDA.n2374 3.4105
R28390 GNDA.n2385 GNDA.n2345 3.4105
R28391 GNDA.n2385 GNDA.n2375 3.4105
R28392 GNDA.n2385 GNDA.n2376 3.4105
R28393 GNDA.n2614 GNDA.n2385 3.4105
R28394 GNDA.n2582 GNDA.n2360 3.4105
R28395 GNDA.n2582 GNDA.n2359 3.4105
R28396 GNDA.n2582 GNDA.n2361 3.4105
R28397 GNDA.n2582 GNDA.n2358 3.4105
R28398 GNDA.n2582 GNDA.n2362 3.4105
R28399 GNDA.n2582 GNDA.n2357 3.4105
R28400 GNDA.n2582 GNDA.n2363 3.4105
R28401 GNDA.n2582 GNDA.n2356 3.4105
R28402 GNDA.n2582 GNDA.n2364 3.4105
R28403 GNDA.n2582 GNDA.n2355 3.4105
R28404 GNDA.n2582 GNDA.n2365 3.4105
R28405 GNDA.n2582 GNDA.n2354 3.4105
R28406 GNDA.n2582 GNDA.n2366 3.4105
R28407 GNDA.n2582 GNDA.n2353 3.4105
R28408 GNDA.n2582 GNDA.n2367 3.4105
R28409 GNDA.n2582 GNDA.n2352 3.4105
R28410 GNDA.n2582 GNDA.n2368 3.4105
R28411 GNDA.n2582 GNDA.n2351 3.4105
R28412 GNDA.n2582 GNDA.n2369 3.4105
R28413 GNDA.n2582 GNDA.n2350 3.4105
R28414 GNDA.n2582 GNDA.n2370 3.4105
R28415 GNDA.n2582 GNDA.n2349 3.4105
R28416 GNDA.n2582 GNDA.n2371 3.4105
R28417 GNDA.n2582 GNDA.n2348 3.4105
R28418 GNDA.n2582 GNDA.n2372 3.4105
R28419 GNDA.n2582 GNDA.n2347 3.4105
R28420 GNDA.n2582 GNDA.n2373 3.4105
R28421 GNDA.n2582 GNDA.n2346 3.4105
R28422 GNDA.n2582 GNDA.n2374 3.4105
R28423 GNDA.n2582 GNDA.n2345 3.4105
R28424 GNDA.n2582 GNDA.n2375 3.4105
R28425 GNDA.n2582 GNDA.n2376 3.4105
R28426 GNDA.n2614 GNDA.n2582 3.4105
R28427 GNDA.n2384 GNDA.n2360 3.4105
R28428 GNDA.n2384 GNDA.n2359 3.4105
R28429 GNDA.n2384 GNDA.n2361 3.4105
R28430 GNDA.n2384 GNDA.n2358 3.4105
R28431 GNDA.n2384 GNDA.n2362 3.4105
R28432 GNDA.n2384 GNDA.n2357 3.4105
R28433 GNDA.n2384 GNDA.n2363 3.4105
R28434 GNDA.n2384 GNDA.n2356 3.4105
R28435 GNDA.n2384 GNDA.n2364 3.4105
R28436 GNDA.n2384 GNDA.n2355 3.4105
R28437 GNDA.n2384 GNDA.n2365 3.4105
R28438 GNDA.n2384 GNDA.n2354 3.4105
R28439 GNDA.n2384 GNDA.n2366 3.4105
R28440 GNDA.n2384 GNDA.n2353 3.4105
R28441 GNDA.n2384 GNDA.n2367 3.4105
R28442 GNDA.n2384 GNDA.n2352 3.4105
R28443 GNDA.n2384 GNDA.n2368 3.4105
R28444 GNDA.n2384 GNDA.n2351 3.4105
R28445 GNDA.n2384 GNDA.n2369 3.4105
R28446 GNDA.n2384 GNDA.n2350 3.4105
R28447 GNDA.n2384 GNDA.n2370 3.4105
R28448 GNDA.n2384 GNDA.n2349 3.4105
R28449 GNDA.n2384 GNDA.n2371 3.4105
R28450 GNDA.n2384 GNDA.n2348 3.4105
R28451 GNDA.n2384 GNDA.n2372 3.4105
R28452 GNDA.n2384 GNDA.n2347 3.4105
R28453 GNDA.n2384 GNDA.n2373 3.4105
R28454 GNDA.n2384 GNDA.n2346 3.4105
R28455 GNDA.n2384 GNDA.n2374 3.4105
R28456 GNDA.n2384 GNDA.n2345 3.4105
R28457 GNDA.n2384 GNDA.n2375 3.4105
R28458 GNDA.n2384 GNDA.n2376 3.4105
R28459 GNDA.n2614 GNDA.n2384 3.4105
R28460 GNDA.n2584 GNDA.n2360 3.4105
R28461 GNDA.n2584 GNDA.n2359 3.4105
R28462 GNDA.n2584 GNDA.n2361 3.4105
R28463 GNDA.n2584 GNDA.n2358 3.4105
R28464 GNDA.n2584 GNDA.n2362 3.4105
R28465 GNDA.n2584 GNDA.n2357 3.4105
R28466 GNDA.n2584 GNDA.n2363 3.4105
R28467 GNDA.n2584 GNDA.n2356 3.4105
R28468 GNDA.n2584 GNDA.n2364 3.4105
R28469 GNDA.n2584 GNDA.n2355 3.4105
R28470 GNDA.n2584 GNDA.n2365 3.4105
R28471 GNDA.n2584 GNDA.n2354 3.4105
R28472 GNDA.n2584 GNDA.n2366 3.4105
R28473 GNDA.n2584 GNDA.n2353 3.4105
R28474 GNDA.n2584 GNDA.n2367 3.4105
R28475 GNDA.n2584 GNDA.n2352 3.4105
R28476 GNDA.n2584 GNDA.n2368 3.4105
R28477 GNDA.n2584 GNDA.n2351 3.4105
R28478 GNDA.n2584 GNDA.n2369 3.4105
R28479 GNDA.n2584 GNDA.n2350 3.4105
R28480 GNDA.n2584 GNDA.n2370 3.4105
R28481 GNDA.n2584 GNDA.n2349 3.4105
R28482 GNDA.n2584 GNDA.n2371 3.4105
R28483 GNDA.n2584 GNDA.n2348 3.4105
R28484 GNDA.n2584 GNDA.n2372 3.4105
R28485 GNDA.n2584 GNDA.n2347 3.4105
R28486 GNDA.n2584 GNDA.n2373 3.4105
R28487 GNDA.n2584 GNDA.n2346 3.4105
R28488 GNDA.n2584 GNDA.n2374 3.4105
R28489 GNDA.n2584 GNDA.n2345 3.4105
R28490 GNDA.n2584 GNDA.n2375 3.4105
R28491 GNDA.n2584 GNDA.n2376 3.4105
R28492 GNDA.n2614 GNDA.n2584 3.4105
R28493 GNDA.n2383 GNDA.n2360 3.4105
R28494 GNDA.n2383 GNDA.n2359 3.4105
R28495 GNDA.n2383 GNDA.n2361 3.4105
R28496 GNDA.n2383 GNDA.n2358 3.4105
R28497 GNDA.n2383 GNDA.n2362 3.4105
R28498 GNDA.n2383 GNDA.n2357 3.4105
R28499 GNDA.n2383 GNDA.n2363 3.4105
R28500 GNDA.n2383 GNDA.n2356 3.4105
R28501 GNDA.n2383 GNDA.n2364 3.4105
R28502 GNDA.n2383 GNDA.n2355 3.4105
R28503 GNDA.n2383 GNDA.n2365 3.4105
R28504 GNDA.n2383 GNDA.n2354 3.4105
R28505 GNDA.n2383 GNDA.n2366 3.4105
R28506 GNDA.n2383 GNDA.n2353 3.4105
R28507 GNDA.n2383 GNDA.n2367 3.4105
R28508 GNDA.n2383 GNDA.n2352 3.4105
R28509 GNDA.n2383 GNDA.n2368 3.4105
R28510 GNDA.n2383 GNDA.n2351 3.4105
R28511 GNDA.n2383 GNDA.n2369 3.4105
R28512 GNDA.n2383 GNDA.n2350 3.4105
R28513 GNDA.n2383 GNDA.n2370 3.4105
R28514 GNDA.n2383 GNDA.n2349 3.4105
R28515 GNDA.n2383 GNDA.n2371 3.4105
R28516 GNDA.n2383 GNDA.n2348 3.4105
R28517 GNDA.n2383 GNDA.n2372 3.4105
R28518 GNDA.n2383 GNDA.n2347 3.4105
R28519 GNDA.n2383 GNDA.n2373 3.4105
R28520 GNDA.n2383 GNDA.n2346 3.4105
R28521 GNDA.n2383 GNDA.n2374 3.4105
R28522 GNDA.n2383 GNDA.n2345 3.4105
R28523 GNDA.n2383 GNDA.n2375 3.4105
R28524 GNDA.n2383 GNDA.n2376 3.4105
R28525 GNDA.n2614 GNDA.n2383 3.4105
R28526 GNDA.n2586 GNDA.n2360 3.4105
R28527 GNDA.n2586 GNDA.n2359 3.4105
R28528 GNDA.n2586 GNDA.n2361 3.4105
R28529 GNDA.n2586 GNDA.n2358 3.4105
R28530 GNDA.n2586 GNDA.n2362 3.4105
R28531 GNDA.n2586 GNDA.n2357 3.4105
R28532 GNDA.n2586 GNDA.n2363 3.4105
R28533 GNDA.n2586 GNDA.n2356 3.4105
R28534 GNDA.n2586 GNDA.n2364 3.4105
R28535 GNDA.n2586 GNDA.n2355 3.4105
R28536 GNDA.n2586 GNDA.n2365 3.4105
R28537 GNDA.n2586 GNDA.n2354 3.4105
R28538 GNDA.n2586 GNDA.n2366 3.4105
R28539 GNDA.n2586 GNDA.n2353 3.4105
R28540 GNDA.n2586 GNDA.n2367 3.4105
R28541 GNDA.n2586 GNDA.n2352 3.4105
R28542 GNDA.n2586 GNDA.n2368 3.4105
R28543 GNDA.n2586 GNDA.n2351 3.4105
R28544 GNDA.n2586 GNDA.n2369 3.4105
R28545 GNDA.n2586 GNDA.n2350 3.4105
R28546 GNDA.n2586 GNDA.n2370 3.4105
R28547 GNDA.n2586 GNDA.n2349 3.4105
R28548 GNDA.n2586 GNDA.n2371 3.4105
R28549 GNDA.n2586 GNDA.n2348 3.4105
R28550 GNDA.n2586 GNDA.n2372 3.4105
R28551 GNDA.n2586 GNDA.n2347 3.4105
R28552 GNDA.n2586 GNDA.n2373 3.4105
R28553 GNDA.n2586 GNDA.n2346 3.4105
R28554 GNDA.n2586 GNDA.n2374 3.4105
R28555 GNDA.n2586 GNDA.n2345 3.4105
R28556 GNDA.n2586 GNDA.n2375 3.4105
R28557 GNDA.n2586 GNDA.n2376 3.4105
R28558 GNDA.n2614 GNDA.n2586 3.4105
R28559 GNDA.n2382 GNDA.n2360 3.4105
R28560 GNDA.n2382 GNDA.n2359 3.4105
R28561 GNDA.n2382 GNDA.n2361 3.4105
R28562 GNDA.n2382 GNDA.n2358 3.4105
R28563 GNDA.n2382 GNDA.n2362 3.4105
R28564 GNDA.n2382 GNDA.n2357 3.4105
R28565 GNDA.n2382 GNDA.n2363 3.4105
R28566 GNDA.n2382 GNDA.n2356 3.4105
R28567 GNDA.n2382 GNDA.n2364 3.4105
R28568 GNDA.n2382 GNDA.n2355 3.4105
R28569 GNDA.n2382 GNDA.n2365 3.4105
R28570 GNDA.n2382 GNDA.n2354 3.4105
R28571 GNDA.n2382 GNDA.n2366 3.4105
R28572 GNDA.n2382 GNDA.n2353 3.4105
R28573 GNDA.n2382 GNDA.n2367 3.4105
R28574 GNDA.n2382 GNDA.n2352 3.4105
R28575 GNDA.n2382 GNDA.n2368 3.4105
R28576 GNDA.n2382 GNDA.n2351 3.4105
R28577 GNDA.n2382 GNDA.n2369 3.4105
R28578 GNDA.n2382 GNDA.n2350 3.4105
R28579 GNDA.n2382 GNDA.n2370 3.4105
R28580 GNDA.n2382 GNDA.n2349 3.4105
R28581 GNDA.n2382 GNDA.n2371 3.4105
R28582 GNDA.n2382 GNDA.n2348 3.4105
R28583 GNDA.n2382 GNDA.n2372 3.4105
R28584 GNDA.n2382 GNDA.n2347 3.4105
R28585 GNDA.n2382 GNDA.n2373 3.4105
R28586 GNDA.n2382 GNDA.n2346 3.4105
R28587 GNDA.n2382 GNDA.n2374 3.4105
R28588 GNDA.n2382 GNDA.n2345 3.4105
R28589 GNDA.n2382 GNDA.n2375 3.4105
R28590 GNDA.n2382 GNDA.n2376 3.4105
R28591 GNDA.n2614 GNDA.n2382 3.4105
R28592 GNDA.n2588 GNDA.n2360 3.4105
R28593 GNDA.n2588 GNDA.n2359 3.4105
R28594 GNDA.n2588 GNDA.n2361 3.4105
R28595 GNDA.n2588 GNDA.n2358 3.4105
R28596 GNDA.n2588 GNDA.n2362 3.4105
R28597 GNDA.n2588 GNDA.n2357 3.4105
R28598 GNDA.n2588 GNDA.n2363 3.4105
R28599 GNDA.n2588 GNDA.n2356 3.4105
R28600 GNDA.n2588 GNDA.n2364 3.4105
R28601 GNDA.n2588 GNDA.n2355 3.4105
R28602 GNDA.n2588 GNDA.n2365 3.4105
R28603 GNDA.n2588 GNDA.n2354 3.4105
R28604 GNDA.n2588 GNDA.n2366 3.4105
R28605 GNDA.n2588 GNDA.n2353 3.4105
R28606 GNDA.n2588 GNDA.n2367 3.4105
R28607 GNDA.n2588 GNDA.n2352 3.4105
R28608 GNDA.n2588 GNDA.n2368 3.4105
R28609 GNDA.n2588 GNDA.n2351 3.4105
R28610 GNDA.n2588 GNDA.n2369 3.4105
R28611 GNDA.n2588 GNDA.n2350 3.4105
R28612 GNDA.n2588 GNDA.n2370 3.4105
R28613 GNDA.n2588 GNDA.n2349 3.4105
R28614 GNDA.n2588 GNDA.n2371 3.4105
R28615 GNDA.n2588 GNDA.n2348 3.4105
R28616 GNDA.n2588 GNDA.n2372 3.4105
R28617 GNDA.n2588 GNDA.n2347 3.4105
R28618 GNDA.n2588 GNDA.n2373 3.4105
R28619 GNDA.n2588 GNDA.n2346 3.4105
R28620 GNDA.n2588 GNDA.n2374 3.4105
R28621 GNDA.n2588 GNDA.n2345 3.4105
R28622 GNDA.n2588 GNDA.n2375 3.4105
R28623 GNDA.n2588 GNDA.n2376 3.4105
R28624 GNDA.n2614 GNDA.n2588 3.4105
R28625 GNDA.n2381 GNDA.n2360 3.4105
R28626 GNDA.n2381 GNDA.n2359 3.4105
R28627 GNDA.n2381 GNDA.n2361 3.4105
R28628 GNDA.n2381 GNDA.n2358 3.4105
R28629 GNDA.n2381 GNDA.n2362 3.4105
R28630 GNDA.n2381 GNDA.n2357 3.4105
R28631 GNDA.n2381 GNDA.n2363 3.4105
R28632 GNDA.n2381 GNDA.n2356 3.4105
R28633 GNDA.n2381 GNDA.n2364 3.4105
R28634 GNDA.n2381 GNDA.n2355 3.4105
R28635 GNDA.n2381 GNDA.n2365 3.4105
R28636 GNDA.n2381 GNDA.n2354 3.4105
R28637 GNDA.n2381 GNDA.n2366 3.4105
R28638 GNDA.n2381 GNDA.n2353 3.4105
R28639 GNDA.n2381 GNDA.n2367 3.4105
R28640 GNDA.n2381 GNDA.n2352 3.4105
R28641 GNDA.n2381 GNDA.n2368 3.4105
R28642 GNDA.n2381 GNDA.n2351 3.4105
R28643 GNDA.n2381 GNDA.n2369 3.4105
R28644 GNDA.n2381 GNDA.n2350 3.4105
R28645 GNDA.n2381 GNDA.n2370 3.4105
R28646 GNDA.n2381 GNDA.n2349 3.4105
R28647 GNDA.n2381 GNDA.n2371 3.4105
R28648 GNDA.n2381 GNDA.n2348 3.4105
R28649 GNDA.n2381 GNDA.n2372 3.4105
R28650 GNDA.n2381 GNDA.n2347 3.4105
R28651 GNDA.n2381 GNDA.n2373 3.4105
R28652 GNDA.n2381 GNDA.n2346 3.4105
R28653 GNDA.n2381 GNDA.n2374 3.4105
R28654 GNDA.n2381 GNDA.n2345 3.4105
R28655 GNDA.n2381 GNDA.n2375 3.4105
R28656 GNDA.n2381 GNDA.n2376 3.4105
R28657 GNDA.n2614 GNDA.n2381 3.4105
R28658 GNDA.n2590 GNDA.n2360 3.4105
R28659 GNDA.n2590 GNDA.n2359 3.4105
R28660 GNDA.n2590 GNDA.n2361 3.4105
R28661 GNDA.n2590 GNDA.n2358 3.4105
R28662 GNDA.n2590 GNDA.n2362 3.4105
R28663 GNDA.n2590 GNDA.n2357 3.4105
R28664 GNDA.n2590 GNDA.n2363 3.4105
R28665 GNDA.n2590 GNDA.n2356 3.4105
R28666 GNDA.n2590 GNDA.n2364 3.4105
R28667 GNDA.n2590 GNDA.n2355 3.4105
R28668 GNDA.n2590 GNDA.n2365 3.4105
R28669 GNDA.n2590 GNDA.n2354 3.4105
R28670 GNDA.n2590 GNDA.n2366 3.4105
R28671 GNDA.n2590 GNDA.n2353 3.4105
R28672 GNDA.n2590 GNDA.n2367 3.4105
R28673 GNDA.n2590 GNDA.n2352 3.4105
R28674 GNDA.n2590 GNDA.n2368 3.4105
R28675 GNDA.n2590 GNDA.n2351 3.4105
R28676 GNDA.n2590 GNDA.n2369 3.4105
R28677 GNDA.n2590 GNDA.n2350 3.4105
R28678 GNDA.n2590 GNDA.n2370 3.4105
R28679 GNDA.n2590 GNDA.n2349 3.4105
R28680 GNDA.n2590 GNDA.n2371 3.4105
R28681 GNDA.n2590 GNDA.n2348 3.4105
R28682 GNDA.n2590 GNDA.n2372 3.4105
R28683 GNDA.n2590 GNDA.n2347 3.4105
R28684 GNDA.n2590 GNDA.n2373 3.4105
R28685 GNDA.n2590 GNDA.n2346 3.4105
R28686 GNDA.n2590 GNDA.n2374 3.4105
R28687 GNDA.n2590 GNDA.n2345 3.4105
R28688 GNDA.n2590 GNDA.n2375 3.4105
R28689 GNDA.n2590 GNDA.n2376 3.4105
R28690 GNDA.n2614 GNDA.n2590 3.4105
R28691 GNDA.n2380 GNDA.n2360 3.4105
R28692 GNDA.n2380 GNDA.n2359 3.4105
R28693 GNDA.n2380 GNDA.n2361 3.4105
R28694 GNDA.n2380 GNDA.n2358 3.4105
R28695 GNDA.n2380 GNDA.n2362 3.4105
R28696 GNDA.n2380 GNDA.n2357 3.4105
R28697 GNDA.n2380 GNDA.n2363 3.4105
R28698 GNDA.n2380 GNDA.n2356 3.4105
R28699 GNDA.n2380 GNDA.n2364 3.4105
R28700 GNDA.n2380 GNDA.n2355 3.4105
R28701 GNDA.n2380 GNDA.n2365 3.4105
R28702 GNDA.n2380 GNDA.n2354 3.4105
R28703 GNDA.n2380 GNDA.n2366 3.4105
R28704 GNDA.n2380 GNDA.n2353 3.4105
R28705 GNDA.n2380 GNDA.n2367 3.4105
R28706 GNDA.n2380 GNDA.n2352 3.4105
R28707 GNDA.n2380 GNDA.n2368 3.4105
R28708 GNDA.n2380 GNDA.n2351 3.4105
R28709 GNDA.n2380 GNDA.n2369 3.4105
R28710 GNDA.n2380 GNDA.n2350 3.4105
R28711 GNDA.n2380 GNDA.n2370 3.4105
R28712 GNDA.n2380 GNDA.n2349 3.4105
R28713 GNDA.n2380 GNDA.n2371 3.4105
R28714 GNDA.n2380 GNDA.n2348 3.4105
R28715 GNDA.n2380 GNDA.n2372 3.4105
R28716 GNDA.n2380 GNDA.n2347 3.4105
R28717 GNDA.n2380 GNDA.n2373 3.4105
R28718 GNDA.n2380 GNDA.n2346 3.4105
R28719 GNDA.n2380 GNDA.n2374 3.4105
R28720 GNDA.n2380 GNDA.n2345 3.4105
R28721 GNDA.n2380 GNDA.n2375 3.4105
R28722 GNDA.n2380 GNDA.n2376 3.4105
R28723 GNDA.n2614 GNDA.n2380 3.4105
R28724 GNDA.n2592 GNDA.n2360 3.4105
R28725 GNDA.n2592 GNDA.n2359 3.4105
R28726 GNDA.n2592 GNDA.n2361 3.4105
R28727 GNDA.n2592 GNDA.n2358 3.4105
R28728 GNDA.n2592 GNDA.n2362 3.4105
R28729 GNDA.n2592 GNDA.n2357 3.4105
R28730 GNDA.n2592 GNDA.n2363 3.4105
R28731 GNDA.n2592 GNDA.n2356 3.4105
R28732 GNDA.n2592 GNDA.n2364 3.4105
R28733 GNDA.n2592 GNDA.n2355 3.4105
R28734 GNDA.n2592 GNDA.n2365 3.4105
R28735 GNDA.n2592 GNDA.n2354 3.4105
R28736 GNDA.n2592 GNDA.n2366 3.4105
R28737 GNDA.n2592 GNDA.n2353 3.4105
R28738 GNDA.n2592 GNDA.n2367 3.4105
R28739 GNDA.n2592 GNDA.n2352 3.4105
R28740 GNDA.n2592 GNDA.n2368 3.4105
R28741 GNDA.n2592 GNDA.n2351 3.4105
R28742 GNDA.n2592 GNDA.n2369 3.4105
R28743 GNDA.n2592 GNDA.n2350 3.4105
R28744 GNDA.n2592 GNDA.n2370 3.4105
R28745 GNDA.n2592 GNDA.n2349 3.4105
R28746 GNDA.n2592 GNDA.n2371 3.4105
R28747 GNDA.n2592 GNDA.n2348 3.4105
R28748 GNDA.n2592 GNDA.n2372 3.4105
R28749 GNDA.n2592 GNDA.n2347 3.4105
R28750 GNDA.n2592 GNDA.n2373 3.4105
R28751 GNDA.n2592 GNDA.n2346 3.4105
R28752 GNDA.n2592 GNDA.n2374 3.4105
R28753 GNDA.n2592 GNDA.n2345 3.4105
R28754 GNDA.n2592 GNDA.n2375 3.4105
R28755 GNDA.n2592 GNDA.n2376 3.4105
R28756 GNDA.n2614 GNDA.n2592 3.4105
R28757 GNDA.n2379 GNDA.n2360 3.4105
R28758 GNDA.n2379 GNDA.n2359 3.4105
R28759 GNDA.n2379 GNDA.n2361 3.4105
R28760 GNDA.n2379 GNDA.n2358 3.4105
R28761 GNDA.n2379 GNDA.n2362 3.4105
R28762 GNDA.n2379 GNDA.n2357 3.4105
R28763 GNDA.n2379 GNDA.n2363 3.4105
R28764 GNDA.n2379 GNDA.n2356 3.4105
R28765 GNDA.n2379 GNDA.n2364 3.4105
R28766 GNDA.n2379 GNDA.n2355 3.4105
R28767 GNDA.n2379 GNDA.n2365 3.4105
R28768 GNDA.n2379 GNDA.n2354 3.4105
R28769 GNDA.n2379 GNDA.n2366 3.4105
R28770 GNDA.n2379 GNDA.n2353 3.4105
R28771 GNDA.n2379 GNDA.n2367 3.4105
R28772 GNDA.n2379 GNDA.n2352 3.4105
R28773 GNDA.n2379 GNDA.n2368 3.4105
R28774 GNDA.n2379 GNDA.n2351 3.4105
R28775 GNDA.n2379 GNDA.n2369 3.4105
R28776 GNDA.n2379 GNDA.n2350 3.4105
R28777 GNDA.n2379 GNDA.n2370 3.4105
R28778 GNDA.n2379 GNDA.n2349 3.4105
R28779 GNDA.n2379 GNDA.n2371 3.4105
R28780 GNDA.n2379 GNDA.n2348 3.4105
R28781 GNDA.n2379 GNDA.n2372 3.4105
R28782 GNDA.n2379 GNDA.n2347 3.4105
R28783 GNDA.n2379 GNDA.n2373 3.4105
R28784 GNDA.n2379 GNDA.n2346 3.4105
R28785 GNDA.n2379 GNDA.n2374 3.4105
R28786 GNDA.n2379 GNDA.n2345 3.4105
R28787 GNDA.n2379 GNDA.n2375 3.4105
R28788 GNDA.n2379 GNDA.n2376 3.4105
R28789 GNDA.n2614 GNDA.n2379 3.4105
R28790 GNDA.n2594 GNDA.n2360 3.4105
R28791 GNDA.n2594 GNDA.n2359 3.4105
R28792 GNDA.n2594 GNDA.n2361 3.4105
R28793 GNDA.n2594 GNDA.n2358 3.4105
R28794 GNDA.n2594 GNDA.n2362 3.4105
R28795 GNDA.n2594 GNDA.n2357 3.4105
R28796 GNDA.n2594 GNDA.n2363 3.4105
R28797 GNDA.n2594 GNDA.n2356 3.4105
R28798 GNDA.n2594 GNDA.n2364 3.4105
R28799 GNDA.n2594 GNDA.n2355 3.4105
R28800 GNDA.n2594 GNDA.n2365 3.4105
R28801 GNDA.n2594 GNDA.n2354 3.4105
R28802 GNDA.n2594 GNDA.n2366 3.4105
R28803 GNDA.n2594 GNDA.n2353 3.4105
R28804 GNDA.n2594 GNDA.n2367 3.4105
R28805 GNDA.n2594 GNDA.n2352 3.4105
R28806 GNDA.n2594 GNDA.n2368 3.4105
R28807 GNDA.n2594 GNDA.n2351 3.4105
R28808 GNDA.n2594 GNDA.n2369 3.4105
R28809 GNDA.n2594 GNDA.n2350 3.4105
R28810 GNDA.n2594 GNDA.n2370 3.4105
R28811 GNDA.n2594 GNDA.n2349 3.4105
R28812 GNDA.n2594 GNDA.n2371 3.4105
R28813 GNDA.n2594 GNDA.n2348 3.4105
R28814 GNDA.n2594 GNDA.n2372 3.4105
R28815 GNDA.n2594 GNDA.n2347 3.4105
R28816 GNDA.n2594 GNDA.n2373 3.4105
R28817 GNDA.n2594 GNDA.n2346 3.4105
R28818 GNDA.n2594 GNDA.n2374 3.4105
R28819 GNDA.n2594 GNDA.n2345 3.4105
R28820 GNDA.n2594 GNDA.n2375 3.4105
R28821 GNDA.n2594 GNDA.n2376 3.4105
R28822 GNDA.n2614 GNDA.n2594 3.4105
R28823 GNDA.n2378 GNDA.n2360 3.4105
R28824 GNDA.n2378 GNDA.n2359 3.4105
R28825 GNDA.n2378 GNDA.n2361 3.4105
R28826 GNDA.n2378 GNDA.n2358 3.4105
R28827 GNDA.n2378 GNDA.n2362 3.4105
R28828 GNDA.n2378 GNDA.n2357 3.4105
R28829 GNDA.n2378 GNDA.n2363 3.4105
R28830 GNDA.n2378 GNDA.n2356 3.4105
R28831 GNDA.n2378 GNDA.n2364 3.4105
R28832 GNDA.n2378 GNDA.n2355 3.4105
R28833 GNDA.n2378 GNDA.n2365 3.4105
R28834 GNDA.n2378 GNDA.n2354 3.4105
R28835 GNDA.n2378 GNDA.n2366 3.4105
R28836 GNDA.n2378 GNDA.n2353 3.4105
R28837 GNDA.n2378 GNDA.n2367 3.4105
R28838 GNDA.n2378 GNDA.n2352 3.4105
R28839 GNDA.n2378 GNDA.n2368 3.4105
R28840 GNDA.n2378 GNDA.n2351 3.4105
R28841 GNDA.n2378 GNDA.n2369 3.4105
R28842 GNDA.n2378 GNDA.n2350 3.4105
R28843 GNDA.n2378 GNDA.n2370 3.4105
R28844 GNDA.n2378 GNDA.n2349 3.4105
R28845 GNDA.n2378 GNDA.n2371 3.4105
R28846 GNDA.n2378 GNDA.n2348 3.4105
R28847 GNDA.n2378 GNDA.n2372 3.4105
R28848 GNDA.n2378 GNDA.n2347 3.4105
R28849 GNDA.n2378 GNDA.n2373 3.4105
R28850 GNDA.n2378 GNDA.n2346 3.4105
R28851 GNDA.n2378 GNDA.n2374 3.4105
R28852 GNDA.n2378 GNDA.n2345 3.4105
R28853 GNDA.n2378 GNDA.n2375 3.4105
R28854 GNDA.n2378 GNDA.n2376 3.4105
R28855 GNDA.n2614 GNDA.n2378 3.4105
R28856 GNDA.n2613 GNDA.n2360 3.4105
R28857 GNDA.n2613 GNDA.n2359 3.4105
R28858 GNDA.n2613 GNDA.n2361 3.4105
R28859 GNDA.n2613 GNDA.n2358 3.4105
R28860 GNDA.n2613 GNDA.n2362 3.4105
R28861 GNDA.n2613 GNDA.n2357 3.4105
R28862 GNDA.n2613 GNDA.n2363 3.4105
R28863 GNDA.n2613 GNDA.n2356 3.4105
R28864 GNDA.n2613 GNDA.n2364 3.4105
R28865 GNDA.n2613 GNDA.n2355 3.4105
R28866 GNDA.n2613 GNDA.n2365 3.4105
R28867 GNDA.n2613 GNDA.n2354 3.4105
R28868 GNDA.n2613 GNDA.n2366 3.4105
R28869 GNDA.n2613 GNDA.n2353 3.4105
R28870 GNDA.n2613 GNDA.n2367 3.4105
R28871 GNDA.n2613 GNDA.n2352 3.4105
R28872 GNDA.n2613 GNDA.n2368 3.4105
R28873 GNDA.n2613 GNDA.n2351 3.4105
R28874 GNDA.n2613 GNDA.n2369 3.4105
R28875 GNDA.n2613 GNDA.n2350 3.4105
R28876 GNDA.n2613 GNDA.n2370 3.4105
R28877 GNDA.n2613 GNDA.n2349 3.4105
R28878 GNDA.n2613 GNDA.n2371 3.4105
R28879 GNDA.n2613 GNDA.n2348 3.4105
R28880 GNDA.n2613 GNDA.n2372 3.4105
R28881 GNDA.n2613 GNDA.n2347 3.4105
R28882 GNDA.n2613 GNDA.n2373 3.4105
R28883 GNDA.n2613 GNDA.n2346 3.4105
R28884 GNDA.n2613 GNDA.n2374 3.4105
R28885 GNDA.n2613 GNDA.n2345 3.4105
R28886 GNDA.n2613 GNDA.n2375 3.4105
R28887 GNDA.n2613 GNDA.n2376 3.4105
R28888 GNDA.n2614 GNDA.n2613 3.4105
R28889 GNDA.n2377 GNDA.n2360 3.4105
R28890 GNDA.n2377 GNDA.n2359 3.4105
R28891 GNDA.n2377 GNDA.n2361 3.4105
R28892 GNDA.n2377 GNDA.n2358 3.4105
R28893 GNDA.n2377 GNDA.n2362 3.4105
R28894 GNDA.n2377 GNDA.n2357 3.4105
R28895 GNDA.n2377 GNDA.n2363 3.4105
R28896 GNDA.n2377 GNDA.n2356 3.4105
R28897 GNDA.n2377 GNDA.n2364 3.4105
R28898 GNDA.n2377 GNDA.n2355 3.4105
R28899 GNDA.n2377 GNDA.n2365 3.4105
R28900 GNDA.n2377 GNDA.n2354 3.4105
R28901 GNDA.n2377 GNDA.n2366 3.4105
R28902 GNDA.n2377 GNDA.n2353 3.4105
R28903 GNDA.n2377 GNDA.n2367 3.4105
R28904 GNDA.n2377 GNDA.n2352 3.4105
R28905 GNDA.n2377 GNDA.n2368 3.4105
R28906 GNDA.n2377 GNDA.n2351 3.4105
R28907 GNDA.n2377 GNDA.n2369 3.4105
R28908 GNDA.n2377 GNDA.n2350 3.4105
R28909 GNDA.n2377 GNDA.n2370 3.4105
R28910 GNDA.n2377 GNDA.n2349 3.4105
R28911 GNDA.n2377 GNDA.n2371 3.4105
R28912 GNDA.n2377 GNDA.n2348 3.4105
R28913 GNDA.n2377 GNDA.n2372 3.4105
R28914 GNDA.n2377 GNDA.n2347 3.4105
R28915 GNDA.n2377 GNDA.n2373 3.4105
R28916 GNDA.n2377 GNDA.n2346 3.4105
R28917 GNDA.n2377 GNDA.n2374 3.4105
R28918 GNDA.n2377 GNDA.n2345 3.4105
R28919 GNDA.n2377 GNDA.n2375 3.4105
R28920 GNDA.n2377 GNDA.n2376 3.4105
R28921 GNDA.n2614 GNDA.n2377 3.4105
R28922 GNDA.n2615 GNDA.n2360 3.4105
R28923 GNDA.n2615 GNDA.n2359 3.4105
R28924 GNDA.n2615 GNDA.n2361 3.4105
R28925 GNDA.n2615 GNDA.n2358 3.4105
R28926 GNDA.n2615 GNDA.n2362 3.4105
R28927 GNDA.n2615 GNDA.n2357 3.4105
R28928 GNDA.n2615 GNDA.n2363 3.4105
R28929 GNDA.n2615 GNDA.n2356 3.4105
R28930 GNDA.n2615 GNDA.n2364 3.4105
R28931 GNDA.n2615 GNDA.n2355 3.4105
R28932 GNDA.n2615 GNDA.n2365 3.4105
R28933 GNDA.n2615 GNDA.n2354 3.4105
R28934 GNDA.n2615 GNDA.n2366 3.4105
R28935 GNDA.n2615 GNDA.n2353 3.4105
R28936 GNDA.n2615 GNDA.n2367 3.4105
R28937 GNDA.n2615 GNDA.n2352 3.4105
R28938 GNDA.n2615 GNDA.n2368 3.4105
R28939 GNDA.n2615 GNDA.n2351 3.4105
R28940 GNDA.n2615 GNDA.n2369 3.4105
R28941 GNDA.n2615 GNDA.n2350 3.4105
R28942 GNDA.n2615 GNDA.n2370 3.4105
R28943 GNDA.n2615 GNDA.n2349 3.4105
R28944 GNDA.n2615 GNDA.n2371 3.4105
R28945 GNDA.n2615 GNDA.n2348 3.4105
R28946 GNDA.n2615 GNDA.n2372 3.4105
R28947 GNDA.n2615 GNDA.n2347 3.4105
R28948 GNDA.n2615 GNDA.n2373 3.4105
R28949 GNDA.n2615 GNDA.n2346 3.4105
R28950 GNDA.n2615 GNDA.n2374 3.4105
R28951 GNDA.n2615 GNDA.n2345 3.4105
R28952 GNDA.n2615 GNDA.n2375 3.4105
R28953 GNDA.n2615 GNDA.n2344 3.4105
R28954 GNDA.n2615 GNDA.n2376 3.4105
R28955 GNDA.n2615 GNDA.n2614 3.4105
R28956 GNDA.n5403 GNDA.n5402 3.08383
R28957 GNDA.n637 GNDA.n636 3.08383
R28958 GNDA.n5324 GNDA.n763 3.04346
R28959 GNDA.n5016 GNDA.n5015 3.00528
R28960 GNDA.n5350 GNDA.n5349 3.00528
R28961 GNDA.n4910 GNDA.n4906 2.69842
R28962 GNDA.n5276 GNDA.n5275 2.6629
R28963 GNDA.n5081 GNDA.n872 2.6629
R28964 GNDA.n5223 GNDA.n815 2.6629
R28965 GNDA.n4721 GNDA.n4720 2.6629
R28966 GNDA.n4633 GNDA.n1259 2.6629
R28967 GNDA.n1783 GNDA.n1782 2.6629
R28968 GNDA.n4818 GNDA.n4817 2.6629
R28969 GNDA.n1233 GNDA.n1232 2.6629
R28970 GNDA.n4544 GNDA.n4543 2.6629
R28971 GNDA.n4451 GNDA.n1653 2.6629
R28972 GNDA.n4850 GNDA.n1151 2.6629
R28973 GNDA.n1510 GNDA.n1398 2.6629
R28974 GNDA.n5029 GNDA.n941 2.6629
R28975 GNDA.n5187 GNDA.n5186 2.6629
R28976 GNDA.n4445 GNDA.n4444 2.6629
R28977 GNDA.n5542 GNDA.n5541 2.57991
R28978 GNDA.n578 GNDA.n577 2.57939
R28979 GNDA.n355 GNDA.n353 2.54738
R28980 GNDA.n268 GNDA.n267 2.54738
R28981 GNDA.n181 GNDA.n180 2.54738
R28982 GNDA.n451 GNDA.n450 2.54738
R28983 GNDA.n444 GNDA.n443 2.54738
R28984 GNDA.n617 GNDA.n27 2.46404
R28985 GNDA.n614 GNDA.n612 2.46404
R28986 GNDA.n5276 GNDA.n5223 2.4581
R28987 GNDA.n5334 GNDA.n5333 2.4581
R28988 GNDA.n5187 GNDA.n872 2.4581
R28989 GNDA.n5136 GNDA.n815 2.4581
R28990 GNDA.n4721 GNDA.n1233 2.4581
R28991 GNDA.n4634 GNDA.n4633 2.4581
R28992 GNDA.n1782 GNDA.n1259 2.4581
R28993 GNDA.n1821 GNDA.n1820 2.4581
R28994 GNDA.n1232 GNDA.n1214 2.4581
R28995 GNDA.n4544 GNDA.n1398 2.4581
R28996 GNDA.n4452 GNDA.n4451 2.4581
R28997 GNDA.n1510 GNDA.n1509 2.4581
R28998 GNDA.n5186 GNDA.n882 2.4581
R28999 GNDA.n4445 GNDA.n1653 2.4581
R29000 GNDA.n4353 GNDA.n4352 2.4581
R29001 GNDA.n4886 GNDA.n4885 2.41717
R29002 GNDA.n977 GNDA.n976 2.39683
R29003 GNDA.n1067 GNDA.n1066 2.30736
R29004 GNDA.n2075 GNDA.n2074 2.30736
R29005 GNDA.n4113 GNDA.n3686 2.30736
R29006 GNDA.n4092 GNDA.n4091 2.30736
R29007 GNDA.n4011 GNDA.n4010 2.30736
R29008 GNDA.n3930 GNDA.n3929 2.30736
R29009 GNDA.n4234 GNDA.n4233 2.30736
R29010 GNDA.n3849 GNDA.n3848 2.30736
R29011 GNDA.n3768 GNDA.n3767 2.30736
R29012 GNDA.n3560 GNDA.n3552 2.30736
R29013 GNDA.n4239 GNDA.n1999 2.30736
R29014 GNDA.n3455 GNDA.n3454 2.30736
R29015 GNDA.n3366 GNDA.n3365 2.30736
R29016 GNDA.n3283 GNDA.n3282 2.30736
R29017 GNDA.n3207 GNDA.n3206 2.30736
R29018 GNDA.n3104 GNDA.n3103 2.30736
R29019 GNDA.n3049 GNDA.n3048 2.30736
R29020 GNDA.n2973 GNDA.n2972 2.30736
R29021 GNDA.n2870 GNDA.n2869 2.30736
R29022 GNDA.n2815 GNDA.n2814 2.30736
R29023 GNDA.n2737 GNDA.n2736 2.30736
R29024 GNDA.n5597 GNDA.n5596 2.30736
R29025 GNDA.n572 GNDA.n571 2.30736
R29026 GNDA.n316 GNDA.n315 2.30736
R29027 GNDA.n262 GNDA.n261 2.30736
R29028 GNDA.n143 GNDA.n142 2.30736
R29029 GNDA.n506 GNDA.n505 2.30736
R29030 GNDA.n409 GNDA.n404 2.30736
R29031 GNDA.n2203 GNDA.n2202 2.29914
R29032 GNDA.n3625 GNDA.n3624 2.29914
R29033 GNDA.n2208 GNDA.n2207 2.29914
R29034 GNDA.n3620 GNDA.n3619 2.29878
R29035 GNDA.n4901 GNDA.n4900 2.29738
R29036 GNDA.n2217 GNDA.n2213 2.26187
R29037 GNDA.n3633 GNDA.n3629 2.26187
R29038 GNDA.n5066 GNDA.n5065 2.26187
R29039 GNDA.n5321 GNDA.n5320 2.26187
R29040 GNDA.n4167 GNDA.n3641 2.26187
R29041 GNDA.n3398 GNDA.n3394 2.26187
R29042 GNDA.n5445 GNDA.n5444 2.26187
R29043 GNDA.n5414 GNDA.n690 2.26187
R29044 GNDA.n2191 GNDA.n693 2.26187
R29045 GNDA.n2194 GNDA.n2189 2.26187
R29046 GNDA.n3614 GNDA.n3610 2.26187
R29047 GNDA.n4905 GNDA.n950 2.26187
R29048 GNDA.n4909 GNDA.n4908 2.26187
R29049 GNDA.n4908 GNDA.n947 2.26187
R29050 GNDA.n2214 GNDA.n2212 2.26187
R29051 GNDA.n2214 GNDA.n2213 2.26187
R29052 GNDA.n3630 GNDA.n3628 2.26187
R29053 GNDA.n3630 GNDA.n3629 2.26187
R29054 GNDA.n5322 GNDA.n5321 2.26187
R29055 GNDA.n5048 GNDA.n5047 2.26187
R29056 GNDA.n4177 GNDA.n3512 2.26187
R29057 GNDA.n4173 GNDA.n3597 2.26187
R29058 GNDA.n4169 GNDA.n3602 2.26187
R29059 GNDA.n4161 GNDA.n3644 2.26187
R29060 GNDA.n4157 GNDA.n3649 2.26187
R29061 GNDA.n4153 GNDA.n3654 2.26187
R29062 GNDA.n4149 GNDA.n3659 2.26187
R29063 GNDA.n3395 GNDA.n3394 2.26187
R29064 GNDA.n2683 GNDA.n2682 2.26187
R29065 GNDA.n2195 GNDA.n2194 2.26187
R29066 GNDA.n5428 GNDA.n5427 2.26187
R29067 GNDA.n5485 GNDA.n664 2.26187
R29068 GNDA.n686 GNDA.n685 2.26187
R29069 GNDA.n5486 GNDA.n5485 2.26187
R29070 GNDA.n28 GNDA.n26 2.26187
R29071 GNDA.n5529 GNDA.n29 2.26187
R29072 GNDA.n5530 GNDA.n5529 2.26187
R29073 GNDA.n373 GNDA.n372 2.26187
R29074 GNDA.n4902 GNDA.n949 2.26187
R29075 GNDA.n4186 GNDA.n4185 2.25831
R29076 GNDA.n4187 GNDA.n4186 2.24241
R29077 GNDA.n3510 GNDA.n3509 2.24241
R29078 GNDA.n3292 GNDA.n3291 2.24241
R29079 GNDA.n3293 GNDA.n3290 2.24241
R29080 GNDA.n2218 GNDA.n2212 2.24063
R29081 GNDA.n3634 GNDA.n3628 2.24063
R29082 GNDA.n3635 GNDA.n3608 2.24063
R29083 GNDA.n3627 GNDA.n3607 2.24063
R29084 GNDA.n5065 GNDA.n5064 2.24063
R29085 GNDA.n5047 GNDA.n767 2.24063
R29086 GNDA.n5050 GNDA.n5049 2.24063
R29087 GNDA.n5320 GNDA.n5319 2.24063
R29088 GNDA.n4891 GNDA.n4890 2.24063
R29089 GNDA.n4889 GNDA.n4888 2.24063
R29090 GNDA.n4178 GNDA.n4177 2.24063
R29091 GNDA.n3595 GNDA.n3513 2.24063
R29092 GNDA.n4174 GNDA.n4173 2.24063
R29093 GNDA.n3600 GNDA.n3598 2.24063
R29094 GNDA.n4170 GNDA.n4169 2.24063
R29095 GNDA.n3605 GNDA.n3603 2.24063
R29096 GNDA.n4162 GNDA.n4161 2.24063
R29097 GNDA.n3647 GNDA.n3645 2.24063
R29098 GNDA.n4158 GNDA.n4157 2.24063
R29099 GNDA.n3652 GNDA.n3650 2.24063
R29100 GNDA.n4154 GNDA.n4153 2.24063
R29101 GNDA.n3657 GNDA.n3655 2.24063
R29102 GNDA.n4150 GNDA.n4149 2.24063
R29103 GNDA.n4148 GNDA.n3660 2.24063
R29104 GNDA.n4165 GNDA.n3641 2.24063
R29105 GNDA.n4166 GNDA.n3642 2.24063
R29106 GNDA.n3399 GNDA.n3393 2.24063
R29107 GNDA.n2682 GNDA.n2240 2.24063
R29108 GNDA.n2681 GNDA.n2679 2.24063
R29109 GNDA.n2825 GNDA.n2238 2.24063
R29110 GNDA.n2239 GNDA.n2237 2.24063
R29111 GNDA.n2822 GNDA.n2821 2.24063
R29112 GNDA.n2912 GNDA.n2235 2.24063
R29113 GNDA.n2236 GNDA.n2234 2.24063
R29114 GNDA.n2909 GNDA.n2908 2.24063
R29115 GNDA.n2916 GNDA.n2231 2.24063
R29116 GNDA.n2233 GNDA.n2232 2.24063
R29117 GNDA.n2917 GNDA.n2186 2.24063
R29118 GNDA.n3059 GNDA.n2154 2.24063
R29119 GNDA.n2155 GNDA.n2153 2.24063
R29120 GNDA.n3056 GNDA.n3055 2.24063
R29121 GNDA.n3146 GNDA.n2151 2.24063
R29122 GNDA.n2152 GNDA.n2150 2.24063
R29123 GNDA.n3143 GNDA.n3142 2.24063
R29124 GNDA.n3150 GNDA.n2116 2.24063
R29125 GNDA.n2149 GNDA.n2148 2.24063
R29126 GNDA.n3151 GNDA.n2147 2.24063
R29127 GNDA.n3294 GNDA.n3289 2.24063
R29128 GNDA.n3309 GNDA.n2029 2.24063
R29129 GNDA.n2031 GNDA.n2030 2.24063
R29130 GNDA.n3310 GNDA.n2028 2.24063
R29131 GNDA.n2224 GNDA.n2156 2.24063
R29132 GNDA.n2228 GNDA.n2227 2.24063
R29133 GNDA.n2222 GNDA.n2209 2.24063
R29134 GNDA.n2211 GNDA.n2210 2.24063
R29135 GNDA.n2223 GNDA.n2188 2.24063
R29136 GNDA.n5431 GNDA.n5422 2.24063
R29137 GNDA.n5432 GNDA.n5418 2.24063
R29138 GNDA.n5433 GNDA.n655 2.24063
R29139 GNDA.n5437 GNDA.n5436 2.24063
R29140 GNDA.n5443 GNDA.n679 2.24063
R29141 GNDA.n5416 GNDA.n5415 2.24063
R29142 GNDA.n2192 GNDA.n696 2.24063
R29143 GNDA.n2198 GNDA.n2189 2.24063
R29144 GNDA.n685 GNDA.n682 2.24063
R29145 GNDA.n684 GNDA.n681 2.24063
R29146 GNDA.n5489 GNDA.n5484 2.24063
R29147 GNDA.n5490 GNDA.n664 2.24063
R29148 GNDA.n5494 GNDA.n657 2.24063
R29149 GNDA.n659 GNDA.n658 2.24063
R29150 GNDA.n5495 GNDA.n656 2.24063
R29151 GNDA.n5499 GNDA.n652 2.24063
R29152 GNDA.n654 GNDA.n653 2.24063
R29153 GNDA.n5500 GNDA.n651 2.24063
R29154 GNDA.n3615 GNDA.n3614 2.24063
R29155 GNDA.n3611 GNDA.n3609 2.24063
R29156 GNDA.n5503 GNDA.n5502 2.24063
R29157 GNDA.n650 GNDA.n648 2.24063
R29158 GNDA.n5533 GNDA.n5528 2.24063
R29159 GNDA.n5534 GNDA.n29 2.24063
R29160 GNDA.n5539 GNDA.n27 2.24063
R29161 GNDA.n5540 GNDA.n26 2.24063
R29162 GNDA.n445 GNDA.n373 2.24063
R29163 GNDA.n375 GNDA.n371 2.24063
R29164 GNDA.n449 GNDA.n368 2.24063
R29165 GNDA.n370 GNDA.n369 2.24063
R29166 GNDA.n450 GNDA.n97 2.24063
R29167 GNDA.n364 GNDA.n183 2.24063
R29168 GNDA.n365 GNDA.n182 2.24063
R29169 GNDA.n366 GNDA.n181 2.24063
R29170 GNDA.n360 GNDA.n270 2.24063
R29171 GNDA.n361 GNDA.n269 2.24063
R29172 GNDA.n362 GNDA.n268 2.24063
R29173 GNDA.n354 GNDA.n25 2.24063
R29174 GNDA.n357 GNDA.n356 2.24063
R29175 GNDA.n358 GNDA.n355 2.24063
R29176 GNDA.n606 GNDA.n600 2.24063
R29177 GNDA.n602 GNDA.n601 2.24063
R29178 GNDA.n607 GNDA.n580 2.24063
R29179 GNDA.n612 GNDA.n43 2.24063
R29180 GNDA.n44 GNDA.n42 2.24063
R29181 GNDA.n4906 GNDA.n949 2.24063
R29182 GNDA.n3637 GNDA.n3636 2.24063
R29183 GNDA.n5150 GNDA.n5051 2.24063
R29184 GNDA.n5149 GNDA.n5148 2.24063
R29185 GNDA.n5323 GNDA.n764 2.24063
R29186 GNDA.n4892 GNDA.n1108 2.24063
R29187 GNDA.n3395 GNDA.n1972 2.24063
R29188 GNDA.n2226 GNDA.n2225 2.24063
R29189 GNDA.n5427 GNDA.n5426 2.24063
R29190 GNDA.n5435 GNDA.n5434 2.24063
R29191 GNDA.n5446 GNDA.n5445 2.24063
R29192 GNDA.n5448 GNDA.n5447 2.24063
R29193 GNDA.n5442 GNDA.n690 2.24063
R29194 GNDA.n5441 GNDA.n5440 2.24063
R29195 GNDA.n5413 GNDA.n693 2.24063
R29196 GNDA.n5412 GNDA.n5411 2.24063
R29197 GNDA.n2197 GNDA.n2196 2.24063
R29198 GNDA.n5501 GNDA.n647 2.24063
R29199 GNDA.n5536 GNDA.n5535 2.24063
R29200 GNDA.n609 GNDA.n608 2.24063
R29201 GNDA.n4901 GNDA.n950 2.24063
R29202 GNDA.n4910 GNDA.n4909 2.24063
R29203 GNDA.n4912 GNDA.n4911 2.24063
R29204 GNDA.n5063 GNDA.n5054 2.22018
R29205 GNDA.n5147 GNDA.n5067 2.22018
R29206 GNDA.n4885 GNDA.n1109 2.22018
R29207 GNDA.n5410 GNDA.n700 2.22018
R29208 GNDA.n5459 GNDA.n663 2.22018
R29209 GNDA.n5453 GNDA.n5452 2.22018
R29210 GNDA.n5507 GNDA.n5506 2.22018
R29211 GNDA.n599 GNDA.n589 2.22018
R29212 GNDA.n5527 GNDA.n34 2.22018
R29213 GNDA.n1513 GNDA.n1398 2.18124
R29214 GNDA.n4597 GNDA.n1233 2.18124
R29215 GNDA.n5188 GNDA.n5187 2.18124
R29216 GNDA.n1934 GNDA.n1653 2.18124
R29217 GNDA.n1379 GNDA.n1259 2.18124
R29218 GNDA.n5223 GNDA.n816 2.18124
R29219 GNDA.n4893 GNDA.n4892 2.16717
R29220 GNDA.n5335 GNDA.n5334 2.1509
R29221 GNDA.n5137 GNDA.n5136 2.1509
R29222 GNDA.n4652 GNDA.n4634 2.1509
R29223 GNDA.n1820 GNDA.n1819 2.1509
R29224 GNDA.n4752 GNDA.n1214 2.1509
R29225 GNDA.n4478 GNDA.n4452 2.1509
R29226 GNDA.n1509 GNDA.n1508 2.1509
R29227 GNDA.n888 GNDA.n882 2.1509
R29228 GNDA.n4379 GNDA.n4353 2.1509
R29229 GNDA.n5275 GNDA.n5274 2.13383
R29230 GNDA.n5082 GNDA.n5081 2.13383
R29231 GNDA.n4720 GNDA.n1234 2.13383
R29232 GNDA.n1471 GNDA.n1151 2.13383
R29233 GNDA.n1783 GNDA.n1781 2.13383
R29234 GNDA.n4817 GNDA.n1192 2.13383
R29235 GNDA.n4543 GNDA.n1632 2.13383
R29236 GNDA.n5002 GNDA.n941 2.13383
R29237 GNDA.n4444 GNDA.n1936 2.13383
R29238 GNDA.n3304 GNDA.n3302 2.09414
R29239 GNDA.n4182 GNDA.n1970 2.09414
R29240 GNDA.n4278 GNDA.n4277 2.09414
R29241 GNDA.n3300 GNDA.n3298 2.09414
R29242 GNDA.n4547 GNDA.n1398 2.08643
R29243 GNDA.n1233 GNDA.n847 2.08643
R29244 GNDA.n5187 GNDA.n881 2.08643
R29245 GNDA.n4448 GNDA.n1653 2.08643
R29246 GNDA.n4630 GNDA.n1259 2.08643
R29247 GNDA.n5223 GNDA.n5222 2.08643
R29248 GNDA.n5306 GNDA.n769 2.04803
R29249 GNDA.n5311 GNDA.n5308 2.04803
R29250 GNDA.n5161 GNDA.n5160 2.04803
R29251 GNDA.n5275 GNDA.n809 1.9461
R29252 GNDA.n5081 GNDA.n739 1.9461
R29253 GNDA.n4720 GNDA.n4719 1.9461
R29254 GNDA.n1784 GNDA.n1783 1.9461
R29255 GNDA.n4817 GNDA.n4816 1.9461
R29256 GNDA.n4543 GNDA.n4542 1.9461
R29257 GNDA.n1474 GNDA.n1151 1.9461
R29258 GNDA.n5005 GNDA.n941 1.9461
R29259 GNDA.n4444 GNDA.n4443 1.9461
R29260 GNDA.n2202 GNDA.n2200 1.93383
R29261 GNDA.n3624 GNDA.n3622 1.93383
R29262 GNDA.n3619 GNDA.n3617 1.93383
R29263 GNDA.n2207 GNDA.n2205 1.93383
R29264 GNDA.n2225 GNDA.n2223 1.82342
R29265 GNDA.n3640 GNDA.n3639 1.82342
R29266 GNDA.n5319 GNDA.n5318 1.71925
R29267 GNDA.n2492 GNDA.n2490 1.70567
R29268 GNDA.n2492 GNDA.n2489 1.70567
R29269 GNDA.n2492 GNDA.n2488 1.70567
R29270 GNDA.n2492 GNDA.n2487 1.70567
R29271 GNDA.n2492 GNDA.n2486 1.70567
R29272 GNDA.n2492 GNDA.n2485 1.70567
R29273 GNDA.n2492 GNDA.n2484 1.70567
R29274 GNDA.n2492 GNDA.n2483 1.70567
R29275 GNDA.n2492 GNDA.n2482 1.70567
R29276 GNDA.n2492 GNDA.n2481 1.70567
R29277 GNDA.n2492 GNDA.n2480 1.70567
R29278 GNDA.n2492 GNDA.n2479 1.70567
R29279 GNDA.n2492 GNDA.n2478 1.70567
R29280 GNDA.n2492 GNDA.n2477 1.70567
R29281 GNDA.n2492 GNDA.n2476 1.70567
R29282 GNDA.n2492 GNDA.n2475 1.70567
R29283 GNDA.n2491 GNDA.n954 1.70567
R29284 GNDA.n2539 GNDA.n2473 1.70567
R29285 GNDA.n2473 GNDA.n2472 1.70567
R29286 GNDA.n2473 GNDA.n2471 1.70567
R29287 GNDA.n2473 GNDA.n2470 1.70567
R29288 GNDA.n2473 GNDA.n2469 1.70567
R29289 GNDA.n2473 GNDA.n2468 1.70567
R29290 GNDA.n2473 GNDA.n2467 1.70567
R29291 GNDA.n2473 GNDA.n2466 1.70567
R29292 GNDA.n2473 GNDA.n2465 1.70567
R29293 GNDA.n2473 GNDA.n2464 1.70567
R29294 GNDA.n2473 GNDA.n2463 1.70567
R29295 GNDA.n2473 GNDA.n2462 1.70567
R29296 GNDA.n2473 GNDA.n2461 1.70567
R29297 GNDA.n2473 GNDA.n2460 1.70567
R29298 GNDA.n2473 GNDA.n2459 1.70567
R29299 GNDA.n2473 GNDA.n2458 1.70567
R29300 GNDA.n2493 GNDA.n2474 1.70567
R29301 GNDA.n2494 GNDA.n954 1.70567
R29302 GNDA.n2496 GNDA.n2474 1.70567
R29303 GNDA.n2497 GNDA.n954 1.70567
R29304 GNDA.n2499 GNDA.n2474 1.70567
R29305 GNDA.n2500 GNDA.n954 1.70567
R29306 GNDA.n2502 GNDA.n2474 1.70567
R29307 GNDA.n2503 GNDA.n954 1.70567
R29308 GNDA.n2505 GNDA.n2474 1.70567
R29309 GNDA.n2506 GNDA.n954 1.70567
R29310 GNDA.n2508 GNDA.n2474 1.70567
R29311 GNDA.n2509 GNDA.n954 1.70567
R29312 GNDA.n2511 GNDA.n2474 1.70567
R29313 GNDA.n2512 GNDA.n954 1.70567
R29314 GNDA.n2514 GNDA.n2474 1.70567
R29315 GNDA.n2515 GNDA.n954 1.70567
R29316 GNDA.n2517 GNDA.n2474 1.70567
R29317 GNDA.n2518 GNDA.n954 1.70567
R29318 GNDA.n2520 GNDA.n2474 1.70567
R29319 GNDA.n2521 GNDA.n954 1.70567
R29320 GNDA.n2523 GNDA.n2474 1.70567
R29321 GNDA.n2524 GNDA.n954 1.70567
R29322 GNDA.n2526 GNDA.n2474 1.70567
R29323 GNDA.n2527 GNDA.n954 1.70567
R29324 GNDA.n2529 GNDA.n2474 1.70567
R29325 GNDA.n2530 GNDA.n954 1.70567
R29326 GNDA.n2532 GNDA.n2474 1.70567
R29327 GNDA.n2533 GNDA.n954 1.70567
R29328 GNDA.n2535 GNDA.n2474 1.70567
R29329 GNDA.n2536 GNDA.n954 1.70567
R29330 GNDA.n2538 GNDA.n2474 1.70567
R29331 GNDA.n2541 GNDA.n954 1.70567
R29332 GNDA.n2544 GNDA.n2425 1.70567
R29333 GNDA.n2474 GNDA.n2409 1.70567
R29334 GNDA.n2650 GNDA.n2262 1.70567
R29335 GNDA.n2650 GNDA.n2631 1.70567
R29336 GNDA.n2650 GNDA.n2630 1.70567
R29337 GNDA.n2650 GNDA.n2629 1.70567
R29338 GNDA.n2650 GNDA.n2628 1.70567
R29339 GNDA.n2650 GNDA.n2627 1.70567
R29340 GNDA.n2650 GNDA.n2626 1.70567
R29341 GNDA.n2650 GNDA.n2625 1.70567
R29342 GNDA.n2650 GNDA.n2624 1.70567
R29343 GNDA.n2650 GNDA.n2623 1.70567
R29344 GNDA.n2650 GNDA.n2622 1.70567
R29345 GNDA.n2650 GNDA.n2621 1.70567
R29346 GNDA.n2650 GNDA.n2620 1.70567
R29347 GNDA.n2650 GNDA.n2619 1.70567
R29348 GNDA.n2650 GNDA.n2618 1.70567
R29349 GNDA.n2650 GNDA.n2617 1.70567
R29350 GNDA.n2295 GNDA.n2261 1.70567
R29351 GNDA.n2297 GNDA.n2261 1.70567
R29352 GNDA.n2299 GNDA.n2261 1.70567
R29353 GNDA.n2301 GNDA.n2261 1.70567
R29354 GNDA.n2303 GNDA.n2261 1.70567
R29355 GNDA.n2305 GNDA.n2261 1.70567
R29356 GNDA.n2307 GNDA.n2261 1.70567
R29357 GNDA.n2309 GNDA.n2261 1.70567
R29358 GNDA.n2311 GNDA.n2261 1.70567
R29359 GNDA.n2313 GNDA.n2261 1.70567
R29360 GNDA.n2315 GNDA.n2261 1.70567
R29361 GNDA.n2317 GNDA.n2261 1.70567
R29362 GNDA.n2319 GNDA.n2261 1.70567
R29363 GNDA.n2321 GNDA.n2261 1.70567
R29364 GNDA.n2323 GNDA.n2261 1.70567
R29365 GNDA.n2616 GNDA.n2342 1.70567
R29366 GNDA.n2648 GNDA.n2632 1.70567
R29367 GNDA.n2342 GNDA.n2341 1.70567
R29368 GNDA.n2648 GNDA.n2633 1.70567
R29369 GNDA.n2342 GNDA.n2340 1.70567
R29370 GNDA.n2648 GNDA.n2634 1.70567
R29371 GNDA.n2342 GNDA.n2339 1.70567
R29372 GNDA.n2648 GNDA.n2635 1.70567
R29373 GNDA.n2342 GNDA.n2338 1.70567
R29374 GNDA.n2648 GNDA.n2636 1.70567
R29375 GNDA.n2342 GNDA.n2337 1.70567
R29376 GNDA.n2648 GNDA.n2637 1.70567
R29377 GNDA.n2342 GNDA.n2336 1.70567
R29378 GNDA.n2648 GNDA.n2638 1.70567
R29379 GNDA.n2342 GNDA.n2335 1.70567
R29380 GNDA.n2648 GNDA.n2639 1.70567
R29381 GNDA.n2342 GNDA.n2334 1.70567
R29382 GNDA.n2648 GNDA.n2640 1.70567
R29383 GNDA.n2342 GNDA.n2333 1.70567
R29384 GNDA.n2648 GNDA.n2641 1.70567
R29385 GNDA.n2342 GNDA.n2332 1.70567
R29386 GNDA.n2648 GNDA.n2642 1.70567
R29387 GNDA.n2342 GNDA.n2331 1.70567
R29388 GNDA.n2648 GNDA.n2643 1.70567
R29389 GNDA.n2342 GNDA.n2330 1.70567
R29390 GNDA.n2648 GNDA.n2644 1.70567
R29391 GNDA.n2342 GNDA.n2329 1.70567
R29392 GNDA.n2648 GNDA.n2645 1.70567
R29393 GNDA.n2342 GNDA.n2328 1.70567
R29394 GNDA.n2648 GNDA.n2646 1.70567
R29395 GNDA.n2342 GNDA.n2327 1.70567
R29396 GNDA.n2648 GNDA.n2647 1.70567
R29397 GNDA.n2342 GNDA.n2326 1.70567
R29398 GNDA.n2648 GNDA.n2279 1.70567
R29399 GNDA.n2652 GNDA.n2325 1.70567
R29400 GNDA.n2561 GNDA.n2360 1.70567
R29401 GNDA.n2562 GNDA.n2560 1.70567
R29402 GNDA.n2562 GNDA.n2559 1.70567
R29403 GNDA.n2562 GNDA.n2558 1.70567
R29404 GNDA.n2562 GNDA.n2557 1.70567
R29405 GNDA.n2562 GNDA.n2556 1.70567
R29406 GNDA.n2562 GNDA.n2555 1.70567
R29407 GNDA.n2562 GNDA.n2554 1.70567
R29408 GNDA.n2562 GNDA.n2553 1.70567
R29409 GNDA.n2562 GNDA.n2552 1.70567
R29410 GNDA.n2562 GNDA.n2551 1.70567
R29411 GNDA.n2562 GNDA.n2550 1.70567
R29412 GNDA.n2562 GNDA.n2549 1.70567
R29413 GNDA.n2562 GNDA.n2548 1.70567
R29414 GNDA.n2562 GNDA.n2547 1.70567
R29415 GNDA.n2562 GNDA.n2546 1.70567
R29416 GNDA.n2562 GNDA.n2545 1.70567
R29417 GNDA.n2563 GNDA.n2562 1.70567
R29418 GNDA.n2408 GNDA.n2407 1.70567
R29419 GNDA.n2408 GNDA.n2406 1.70567
R29420 GNDA.n2408 GNDA.n2405 1.70567
R29421 GNDA.n2408 GNDA.n2404 1.70567
R29422 GNDA.n2408 GNDA.n2403 1.70567
R29423 GNDA.n2408 GNDA.n2402 1.70567
R29424 GNDA.n2408 GNDA.n2401 1.70567
R29425 GNDA.n2408 GNDA.n2400 1.70567
R29426 GNDA.n2408 GNDA.n2399 1.70567
R29427 GNDA.n2408 GNDA.n2398 1.70567
R29428 GNDA.n2408 GNDA.n2397 1.70567
R29429 GNDA.n2408 GNDA.n2396 1.70567
R29430 GNDA.n2408 GNDA.n2395 1.70567
R29431 GNDA.n2408 GNDA.n2394 1.70567
R29432 GNDA.n2408 GNDA.n2393 1.70567
R29433 GNDA.n2566 GNDA.n2565 1.70567
R29434 GNDA.n2610 GNDA.n2595 1.70567
R29435 GNDA.n2564 GNDA.n2344 1.70567
R29436 GNDA.n2610 GNDA.n2596 1.70567
R29437 GNDA.n2567 GNDA.n2344 1.70567
R29438 GNDA.n2610 GNDA.n2597 1.70567
R29439 GNDA.n2569 GNDA.n2344 1.70567
R29440 GNDA.n2610 GNDA.n2598 1.70567
R29441 GNDA.n2571 GNDA.n2344 1.70567
R29442 GNDA.n2610 GNDA.n2599 1.70567
R29443 GNDA.n2573 GNDA.n2344 1.70567
R29444 GNDA.n2610 GNDA.n2600 1.70567
R29445 GNDA.n2575 GNDA.n2344 1.70567
R29446 GNDA.n2610 GNDA.n2601 1.70567
R29447 GNDA.n2577 GNDA.n2344 1.70567
R29448 GNDA.n2610 GNDA.n2602 1.70567
R29449 GNDA.n2579 GNDA.n2344 1.70567
R29450 GNDA.n2610 GNDA.n2603 1.70567
R29451 GNDA.n2581 GNDA.n2344 1.70567
R29452 GNDA.n2610 GNDA.n2604 1.70567
R29453 GNDA.n2583 GNDA.n2344 1.70567
R29454 GNDA.n2610 GNDA.n2605 1.70567
R29455 GNDA.n2585 GNDA.n2344 1.70567
R29456 GNDA.n2610 GNDA.n2606 1.70567
R29457 GNDA.n2587 GNDA.n2344 1.70567
R29458 GNDA.n2610 GNDA.n2607 1.70567
R29459 GNDA.n2589 GNDA.n2344 1.70567
R29460 GNDA.n2610 GNDA.n2608 1.70567
R29461 GNDA.n2591 GNDA.n2344 1.70567
R29462 GNDA.n2610 GNDA.n2609 1.70567
R29463 GNDA.n2593 GNDA.n2344 1.70567
R29464 GNDA.n2611 GNDA.n2610 1.70567
R29465 GNDA.n2612 GNDA.n2344 1.70567
R29466 GNDA.n2610 GNDA.n2343 1.70567
R29467 GNDA.n2817 GNDA.n2750 1.69433
R29468 GNDA.n2817 GNDA.n2747 1.69433
R29469 GNDA.n2817 GNDA.n2744 1.69433
R29470 GNDA.n2879 GNDA.n2161 1.69433
R29471 GNDA.n2888 GNDA.n2161 1.69433
R29472 GNDA.n2897 GNDA.n2161 1.69433
R29473 GNDA.n2975 GNDA.n2171 1.69433
R29474 GNDA.n2975 GNDA.n2168 1.69433
R29475 GNDA.n2975 GNDA.n2165 1.69433
R29476 GNDA.n3051 GNDA.n2984 1.69433
R29477 GNDA.n3051 GNDA.n2981 1.69433
R29478 GNDA.n3051 GNDA.n2978 1.69433
R29479 GNDA.n3113 GNDA.n2122 1.69433
R29480 GNDA.n3122 GNDA.n2122 1.69433
R29481 GNDA.n3131 GNDA.n2122 1.69433
R29482 GNDA.n3209 GNDA.n2132 1.69433
R29483 GNDA.n3209 GNDA.n2129 1.69433
R29484 GNDA.n3209 GNDA.n2126 1.69433
R29485 GNDA.n3285 GNDA.n3218 1.69433
R29486 GNDA.n3285 GNDA.n3215 1.69433
R29487 GNDA.n3285 GNDA.n3212 1.69433
R29488 GNDA.n3368 GNDA.n2013 1.69433
R29489 GNDA.n3368 GNDA.n2010 1.69433
R29490 GNDA.n3368 GNDA.n2007 1.69433
R29491 GNDA.n3457 GNDA.n3378 1.69433
R29492 GNDA.n3457 GNDA.n3375 1.69433
R29493 GNDA.n3457 GNDA.n3372 1.69433
R29494 GNDA.n2084 GNDA.n2003 1.69433
R29495 GNDA.n2093 GNDA.n2003 1.69433
R29496 GNDA.n2102 GNDA.n2003 1.69433
R29497 GNDA.n4237 GNDA.n3470 1.69433
R29498 GNDA.n4237 GNDA.n3466 1.69433
R29499 GNDA.n4237 GNDA.n3461 1.69433
R29500 GNDA.n3549 GNDA.n3486 1.69433
R29501 GNDA.n3538 GNDA.n3486 1.69433
R29502 GNDA.n3525 GNDA.n3486 1.69433
R29503 GNDA.n3770 GNDA.n3699 1.69433
R29504 GNDA.n3770 GNDA.n3696 1.69433
R29505 GNDA.n3770 GNDA.n3693 1.69433
R29506 GNDA.n3851 GNDA.n3780 1.69433
R29507 GNDA.n3851 GNDA.n3777 1.69433
R29508 GNDA.n3851 GNDA.n3774 1.69433
R29509 GNDA.n4236 GNDA.n3483 1.69433
R29510 GNDA.n4236 GNDA.n3480 1.69433
R29511 GNDA.n4236 GNDA.n3477 1.69433
R29512 GNDA.n3932 GNDA.n3861 1.69433
R29513 GNDA.n3932 GNDA.n3858 1.69433
R29514 GNDA.n3932 GNDA.n3855 1.69433
R29515 GNDA.n4013 GNDA.n3942 1.69433
R29516 GNDA.n4013 GNDA.n3939 1.69433
R29517 GNDA.n4013 GNDA.n3936 1.69433
R29518 GNDA.n4094 GNDA.n4023 1.69433
R29519 GNDA.n4094 GNDA.n4020 1.69433
R29520 GNDA.n4094 GNDA.n4017 1.69433
R29521 GNDA.n4111 GNDA.n4107 1.69433
R29522 GNDA.n4111 GNDA.n4103 1.69433
R29523 GNDA.n4111 GNDA.n4098 1.69433
R29524 GNDA.n508 GNDA.n81 1.69433
R29525 GNDA.n508 GNDA.n78 1.69433
R29526 GNDA.n508 GNDA.n75 1.69433
R29527 GNDA.n152 GNDA.n84 1.69433
R29528 GNDA.n161 GNDA.n84 1.69433
R29529 GNDA.n170 GNDA.n84 1.69433
R29530 GNDA.n264 GNDA.n197 1.69433
R29531 GNDA.n264 GNDA.n194 1.69433
R29532 GNDA.n264 GNDA.n191 1.69433
R29533 GNDA.n325 GNDA.n0 1.69433
R29534 GNDA.n334 GNDA.n0 1.69433
R29535 GNDA.n343 GNDA.n0 1.69433
R29536 GNDA.n574 GNDA.n57 1.69433
R29537 GNDA.n574 GNDA.n54 1.69433
R29538 GNDA.n574 GNDA.n51 1.69433
R29539 GNDA.n5599 GNDA.n10 1.69433
R29540 GNDA.n5599 GNDA.n7 1.69433
R29541 GNDA.n5599 GNDA.n4 1.69433
R29542 GNDA.n4897 GNDA.n964 1.69433
R29543 GNDA.n4897 GNDA.n961 1.69433
R29544 GNDA.n4897 GNDA.n958 1.69433
R29545 GNDA.n4896 GNDA.n1039 1.69433
R29546 GNDA.n4896 GNDA.n1036 1.69433
R29547 GNDA.n4896 GNDA.n1033 1.69433
R29548 GNDA.n2741 GNDA.n2664 1.69337
R29549 GNDA.n2741 GNDA.n2663 1.69337
R29550 GNDA.n2741 GNDA.n2661 1.69337
R29551 GNDA.n2741 GNDA.n2660 1.69337
R29552 GNDA.n2741 GNDA.n2658 1.69337
R29553 GNDA.n2741 GNDA.n2657 1.69337
R29554 GNDA.n2741 GNDA.n2655 1.69337
R29555 GNDA.n2741 GNDA.n2654 1.69337
R29556 GNDA.n509 GNDA.n70 1.69337
R29557 GNDA.n509 GNDA.n69 1.69337
R29558 GNDA.n509 GNDA.n67 1.69337
R29559 GNDA.n509 GNDA.n66 1.69337
R29560 GNDA.n509 GNDA.n64 1.69337
R29561 GNDA.n509 GNDA.n63 1.69337
R29562 GNDA.n509 GNDA.n61 1.69337
R29563 GNDA.n509 GNDA.n60 1.69337
R29564 GNDA.n2817 GNDA.n2752 1.6924
R29565 GNDA.n2817 GNDA.n2751 1.6924
R29566 GNDA.n2817 GNDA.n2749 1.6924
R29567 GNDA.n2817 GNDA.n2748 1.6924
R29568 GNDA.n2817 GNDA.n2746 1.6924
R29569 GNDA.n2817 GNDA.n2745 1.6924
R29570 GNDA.n2817 GNDA.n2743 1.6924
R29571 GNDA.n2817 GNDA.n2742 1.6924
R29572 GNDA.n2873 GNDA.n2161 1.6924
R29573 GNDA.n2876 GNDA.n2161 1.6924
R29574 GNDA.n2882 GNDA.n2161 1.6924
R29575 GNDA.n2885 GNDA.n2161 1.6924
R29576 GNDA.n2891 GNDA.n2161 1.6924
R29577 GNDA.n2894 GNDA.n2161 1.6924
R29578 GNDA.n2900 GNDA.n2161 1.6924
R29579 GNDA.n2903 GNDA.n2161 1.6924
R29580 GNDA.n2975 GNDA.n2173 1.6924
R29581 GNDA.n2975 GNDA.n2172 1.6924
R29582 GNDA.n2975 GNDA.n2170 1.6924
R29583 GNDA.n2975 GNDA.n2169 1.6924
R29584 GNDA.n2975 GNDA.n2167 1.6924
R29585 GNDA.n2975 GNDA.n2166 1.6924
R29586 GNDA.n2975 GNDA.n2164 1.6924
R29587 GNDA.n2975 GNDA.n2163 1.6924
R29588 GNDA.n3051 GNDA.n2986 1.6924
R29589 GNDA.n3051 GNDA.n2985 1.6924
R29590 GNDA.n3051 GNDA.n2983 1.6924
R29591 GNDA.n3051 GNDA.n2982 1.6924
R29592 GNDA.n3051 GNDA.n2980 1.6924
R29593 GNDA.n3051 GNDA.n2979 1.6924
R29594 GNDA.n3051 GNDA.n2977 1.6924
R29595 GNDA.n3051 GNDA.n2976 1.6924
R29596 GNDA.n3107 GNDA.n2122 1.6924
R29597 GNDA.n3110 GNDA.n2122 1.6924
R29598 GNDA.n3116 GNDA.n2122 1.6924
R29599 GNDA.n3119 GNDA.n2122 1.6924
R29600 GNDA.n3125 GNDA.n2122 1.6924
R29601 GNDA.n3128 GNDA.n2122 1.6924
R29602 GNDA.n3134 GNDA.n2122 1.6924
R29603 GNDA.n3137 GNDA.n2122 1.6924
R29604 GNDA.n3209 GNDA.n2134 1.6924
R29605 GNDA.n3209 GNDA.n2133 1.6924
R29606 GNDA.n3209 GNDA.n2131 1.6924
R29607 GNDA.n3209 GNDA.n2130 1.6924
R29608 GNDA.n3209 GNDA.n2128 1.6924
R29609 GNDA.n3209 GNDA.n2127 1.6924
R29610 GNDA.n3209 GNDA.n2125 1.6924
R29611 GNDA.n3209 GNDA.n2124 1.6924
R29612 GNDA.n3285 GNDA.n3220 1.6924
R29613 GNDA.n3285 GNDA.n3219 1.6924
R29614 GNDA.n3285 GNDA.n3217 1.6924
R29615 GNDA.n3285 GNDA.n3216 1.6924
R29616 GNDA.n3285 GNDA.n3214 1.6924
R29617 GNDA.n3285 GNDA.n3213 1.6924
R29618 GNDA.n3285 GNDA.n3211 1.6924
R29619 GNDA.n3285 GNDA.n3210 1.6924
R29620 GNDA.n3368 GNDA.n2015 1.6924
R29621 GNDA.n3368 GNDA.n2014 1.6924
R29622 GNDA.n3368 GNDA.n2012 1.6924
R29623 GNDA.n3368 GNDA.n2011 1.6924
R29624 GNDA.n3368 GNDA.n2009 1.6924
R29625 GNDA.n3368 GNDA.n2008 1.6924
R29626 GNDA.n3368 GNDA.n2006 1.6924
R29627 GNDA.n3368 GNDA.n2005 1.6924
R29628 GNDA.n3457 GNDA.n3380 1.6924
R29629 GNDA.n3457 GNDA.n3379 1.6924
R29630 GNDA.n3457 GNDA.n3377 1.6924
R29631 GNDA.n3457 GNDA.n3376 1.6924
R29632 GNDA.n3457 GNDA.n3374 1.6924
R29633 GNDA.n3457 GNDA.n3373 1.6924
R29634 GNDA.n3457 GNDA.n3371 1.6924
R29635 GNDA.n3457 GNDA.n3370 1.6924
R29636 GNDA.n2078 GNDA.n2003 1.6924
R29637 GNDA.n2081 GNDA.n2003 1.6924
R29638 GNDA.n2087 GNDA.n2003 1.6924
R29639 GNDA.n2090 GNDA.n2003 1.6924
R29640 GNDA.n2096 GNDA.n2003 1.6924
R29641 GNDA.n2099 GNDA.n2003 1.6924
R29642 GNDA.n2105 GNDA.n2003 1.6924
R29643 GNDA.n2108 GNDA.n2003 1.6924
R29644 GNDA.n4237 GNDA.n3473 1.6924
R29645 GNDA.n4237 GNDA.n3472 1.6924
R29646 GNDA.n4237 GNDA.n3469 1.6924
R29647 GNDA.n4237 GNDA.n3467 1.6924
R29648 GNDA.n4237 GNDA.n3464 1.6924
R29649 GNDA.n4237 GNDA.n3463 1.6924
R29650 GNDA.n4237 GNDA.n3460 1.6924
R29651 GNDA.n4237 GNDA.n3458 1.6924
R29652 GNDA.n3557 GNDA.n3486 1.6924
R29653 GNDA.n3554 GNDA.n3486 1.6924
R29654 GNDA.n3546 GNDA.n3486 1.6924
R29655 GNDA.n3541 GNDA.n3486 1.6924
R29656 GNDA.n3533 GNDA.n3486 1.6924
R29657 GNDA.n3530 GNDA.n3486 1.6924
R29658 GNDA.n3522 GNDA.n3486 1.6924
R29659 GNDA.n3517 GNDA.n3486 1.6924
R29660 GNDA.n3770 GNDA.n3701 1.6924
R29661 GNDA.n3770 GNDA.n3700 1.6924
R29662 GNDA.n3770 GNDA.n3698 1.6924
R29663 GNDA.n3770 GNDA.n3697 1.6924
R29664 GNDA.n3770 GNDA.n3695 1.6924
R29665 GNDA.n3770 GNDA.n3694 1.6924
R29666 GNDA.n3770 GNDA.n3692 1.6924
R29667 GNDA.n3770 GNDA.n3691 1.6924
R29668 GNDA.n3851 GNDA.n3782 1.6924
R29669 GNDA.n3851 GNDA.n3781 1.6924
R29670 GNDA.n3851 GNDA.n3779 1.6924
R29671 GNDA.n3851 GNDA.n3778 1.6924
R29672 GNDA.n3851 GNDA.n3776 1.6924
R29673 GNDA.n3851 GNDA.n3775 1.6924
R29674 GNDA.n3851 GNDA.n3773 1.6924
R29675 GNDA.n3851 GNDA.n3772 1.6924
R29676 GNDA.n4236 GNDA.n3485 1.6924
R29677 GNDA.n4236 GNDA.n3484 1.6924
R29678 GNDA.n4236 GNDA.n3482 1.6924
R29679 GNDA.n4236 GNDA.n3481 1.6924
R29680 GNDA.n4236 GNDA.n3479 1.6924
R29681 GNDA.n4236 GNDA.n3478 1.6924
R29682 GNDA.n4236 GNDA.n3476 1.6924
R29683 GNDA.n4236 GNDA.n3475 1.6924
R29684 GNDA.n3932 GNDA.n3863 1.6924
R29685 GNDA.n3932 GNDA.n3862 1.6924
R29686 GNDA.n3932 GNDA.n3860 1.6924
R29687 GNDA.n3932 GNDA.n3859 1.6924
R29688 GNDA.n3932 GNDA.n3857 1.6924
R29689 GNDA.n3932 GNDA.n3856 1.6924
R29690 GNDA.n3932 GNDA.n3854 1.6924
R29691 GNDA.n3932 GNDA.n3853 1.6924
R29692 GNDA.n4013 GNDA.n3944 1.6924
R29693 GNDA.n4013 GNDA.n3943 1.6924
R29694 GNDA.n4013 GNDA.n3941 1.6924
R29695 GNDA.n4013 GNDA.n3940 1.6924
R29696 GNDA.n4013 GNDA.n3938 1.6924
R29697 GNDA.n4013 GNDA.n3937 1.6924
R29698 GNDA.n4013 GNDA.n3935 1.6924
R29699 GNDA.n4013 GNDA.n3934 1.6924
R29700 GNDA.n4094 GNDA.n4025 1.6924
R29701 GNDA.n4094 GNDA.n4024 1.6924
R29702 GNDA.n4094 GNDA.n4022 1.6924
R29703 GNDA.n4094 GNDA.n4021 1.6924
R29704 GNDA.n4094 GNDA.n4019 1.6924
R29705 GNDA.n4094 GNDA.n4018 1.6924
R29706 GNDA.n4094 GNDA.n4016 1.6924
R29707 GNDA.n4094 GNDA.n4015 1.6924
R29708 GNDA.n4111 GNDA.n4110 1.6924
R29709 GNDA.n4111 GNDA.n4109 1.6924
R29710 GNDA.n4111 GNDA.n4106 1.6924
R29711 GNDA.n4111 GNDA.n4104 1.6924
R29712 GNDA.n4111 GNDA.n4101 1.6924
R29713 GNDA.n4111 GNDA.n4100 1.6924
R29714 GNDA.n4111 GNDA.n4097 1.6924
R29715 GNDA.n4111 GNDA.n4095 1.6924
R29716 GNDA.n508 GNDA.n83 1.6924
R29717 GNDA.n508 GNDA.n82 1.6924
R29718 GNDA.n508 GNDA.n80 1.6924
R29719 GNDA.n508 GNDA.n79 1.6924
R29720 GNDA.n508 GNDA.n77 1.6924
R29721 GNDA.n508 GNDA.n76 1.6924
R29722 GNDA.n508 GNDA.n74 1.6924
R29723 GNDA.n508 GNDA.n73 1.6924
R29724 GNDA.n146 GNDA.n84 1.6924
R29725 GNDA.n149 GNDA.n84 1.6924
R29726 GNDA.n155 GNDA.n84 1.6924
R29727 GNDA.n158 GNDA.n84 1.6924
R29728 GNDA.n164 GNDA.n84 1.6924
R29729 GNDA.n167 GNDA.n84 1.6924
R29730 GNDA.n173 GNDA.n84 1.6924
R29731 GNDA.n176 GNDA.n84 1.6924
R29732 GNDA.n264 GNDA.n199 1.6924
R29733 GNDA.n264 GNDA.n198 1.6924
R29734 GNDA.n264 GNDA.n196 1.6924
R29735 GNDA.n264 GNDA.n195 1.6924
R29736 GNDA.n264 GNDA.n193 1.6924
R29737 GNDA.n264 GNDA.n192 1.6924
R29738 GNDA.n264 GNDA.n190 1.6924
R29739 GNDA.n264 GNDA.n189 1.6924
R29740 GNDA.n319 GNDA.n0 1.6924
R29741 GNDA.n322 GNDA.n0 1.6924
R29742 GNDA.n328 GNDA.n0 1.6924
R29743 GNDA.n331 GNDA.n0 1.6924
R29744 GNDA.n337 GNDA.n0 1.6924
R29745 GNDA.n340 GNDA.n0 1.6924
R29746 GNDA.n346 GNDA.n0 1.6924
R29747 GNDA.n349 GNDA.n0 1.6924
R29748 GNDA.n574 GNDA.n59 1.6924
R29749 GNDA.n574 GNDA.n58 1.6924
R29750 GNDA.n574 GNDA.n56 1.6924
R29751 GNDA.n574 GNDA.n55 1.6924
R29752 GNDA.n574 GNDA.n53 1.6924
R29753 GNDA.n574 GNDA.n52 1.6924
R29754 GNDA.n574 GNDA.n50 1.6924
R29755 GNDA.n574 GNDA.n49 1.6924
R29756 GNDA.n5599 GNDA.n12 1.6924
R29757 GNDA.n5599 GNDA.n11 1.6924
R29758 GNDA.n5599 GNDA.n9 1.6924
R29759 GNDA.n5599 GNDA.n8 1.6924
R29760 GNDA.n5599 GNDA.n6 1.6924
R29761 GNDA.n5599 GNDA.n5 1.6924
R29762 GNDA.n5599 GNDA.n3 1.6924
R29763 GNDA.n5599 GNDA.n2 1.6924
R29764 GNDA.n4897 GNDA.n1029 1.6924
R29765 GNDA.n4897 GNDA.n965 1.6924
R29766 GNDA.n4897 GNDA.n963 1.6924
R29767 GNDA.n4897 GNDA.n962 1.6924
R29768 GNDA.n4897 GNDA.n960 1.6924
R29769 GNDA.n4897 GNDA.n959 1.6924
R29770 GNDA.n4897 GNDA.n957 1.6924
R29771 GNDA.n4897 GNDA.n956 1.6924
R29772 GNDA.n4896 GNDA.n1041 1.6924
R29773 GNDA.n4896 GNDA.n1040 1.6924
R29774 GNDA.n4896 GNDA.n1038 1.6924
R29775 GNDA.n4896 GNDA.n1037 1.6924
R29776 GNDA.n4896 GNDA.n1035 1.6924
R29777 GNDA.n4896 GNDA.n1034 1.6924
R29778 GNDA.n4896 GNDA.n1032 1.6924
R29779 GNDA.n4896 GNDA.n1031 1.6924
R29780 GNDA.n2741 GNDA.n2740 1.6924
R29781 GNDA.n2741 GNDA.n2662 1.6924
R29782 GNDA.n2741 GNDA.n2659 1.6924
R29783 GNDA.n2741 GNDA.n2656 1.6924
R29784 GNDA.n509 GNDA.n71 1.6924
R29785 GNDA.n509 GNDA.n68 1.6924
R29786 GNDA.n509 GNDA.n65 1.6924
R29787 GNDA.n509 GNDA.n62 1.6924
R29788 GNDA.n5422 GNDA.n5421 1.65675
R29789 GNDA.n5426 GNDA.n5425 1.65675
R29790 GNDA.n588 GNDA.n583 1.56997
R29791 GNDA.n33 GNDA.n32 1.56997
R29792 GNDA.n5332 GNDA.n5331 1.47392
R29793 GNDA.n4852 GNDA.n4851 1.47392
R29794 GNDA.n1829 GNDA.n1705 1.47392
R29795 GNDA.n4825 GNDA.n1188 1.47392
R29796 GNDA.n5031 GNDA.n5030 1.47392
R29797 GNDA.n4342 GNDA.n1957 1.47392
R29798 GNDA.n5470 GNDA.n665 1.44719
R29799 GNDA.n5483 GNDA.n5482 1.44719
R29800 GNDA.n587 GNDA.n585 1.26092
R29801 GNDA.n4274 GNDA.n4273 1.24761
R29802 GNDA.n2113 GNDA.n2112 1.24759
R29803 GNDA_2 GNDA.n5599 1.24042
R29804 GNDA.n5440 GNDA.n5439 1.13592
R29805 GNDA.n5497 GNDA.n655 1.13592
R29806 GNDA.n3638 GNDA.n3625 1.09425
R29807 GNDA.n2209 GNDA.n2208 1.09425
R29808 GNDA.n3636 GNDA.n3634 1.07342
R29809 GNDA.n2219 GNDA.n2218 1.06821
R29810 GNDA.n682 GNDA.n665 1.063
R29811 GNDA.n5484 GNDA.n5483 1.063
R29812 GNDA.n4922 GNDA.n4912 1.05258
R29813 GNDA.n5415 GNDA.n5413 0.984875
R29814 GNDA.n5501 GNDA.n5500 0.984875
R29815 GNDA.n619 GNDA.n617 0.975928
R29816 GNDA.n615 GNDA.n614 0.975928
R29817 GNDA.n5294 GNDA.n5293 0.8197
R29818 GNDA.n5280 GNDA.n810 0.8197
R29819 GNDA.n5287 GNDA.n5281 0.8197
R29820 GNDA.n5286 GNDA.n5283 0.8197
R29821 GNDA.n5300 GNDA.n779 0.8197
R29822 GNDA.n789 GNDA.n786 0.8197
R29823 GNDA.n791 GNDA.n790 0.8197
R29824 GNDA.n5335 GNDA.n756 0.8197
R29825 GNDA.n5365 GNDA.n5364 0.8197
R29826 GNDA.n5351 GNDA.n740 0.8197
R29827 GNDA.n5358 GNDA.n5352 0.8197
R29828 GNDA.n5357 GNDA.n5354 0.8197
R29829 GNDA.n5371 GNDA.n718 0.8197
R29830 GNDA.n5076 GNDA.n5073 0.8197
R29831 GNDA.n5079 GNDA.n5078 0.8197
R29832 GNDA.n5137 GNDA.n5080 0.8197
R29833 GNDA.n4718 GNDA.n1236 0.8197
R29834 GNDA.n4715 GNDA.n4714 0.8197
R29835 GNDA.n4711 GNDA.n1239 0.8197
R29836 GNDA.n4710 GNDA.n1240 0.8197
R29837 GNDA.n4644 GNDA.n4641 0.8197
R29838 GNDA.n4645 GNDA.n4635 0.8197
R29839 GNDA.n4649 GNDA.n4648 0.8197
R29840 GNDA.n4653 GNDA.n4652 0.8197
R29841 GNDA.n1809 GNDA.n1808 0.8197
R29842 GNDA.n1805 GNDA.n1804 0.8197
R29843 GNDA.n1801 GNDA.n1785 0.8197
R29844 GNDA.n1800 GNDA.n1797 0.8197
R29845 GNDA.n1793 GNDA.n1790 0.8197
R29846 GNDA.n1787 GNDA.n1709 0.8197
R29847 GNDA.n1816 GNDA.n1815 0.8197
R29848 GNDA.n1819 GNDA.n1708 0.8197
R29849 GNDA.n4813 GNDA.n1193 0.8197
R29850 GNDA.n4812 GNDA.n1195 0.8197
R29851 GNDA.n4746 GNDA.n4728 0.8197
R29852 GNDA.n4745 GNDA.n4743 0.8197
R29853 GNDA.n4739 GNDA.n4738 0.8197
R29854 GNDA.n4735 GNDA.n4731 0.8197
R29855 GNDA.n4734 GNDA.n1215 0.8197
R29856 GNDA.n4753 GNDA.n4752 0.8197
R29857 GNDA.n4539 GNDA.n1633 0.8197
R29858 GNDA.n4538 GNDA.n1634 0.8197
R29859 GNDA.n4457 GNDA.n4454 0.8197
R29860 GNDA.n4460 GNDA.n4459 0.8197
R29861 GNDA.n4470 GNDA.n4467 0.8197
R29862 GNDA.n4471 GNDA.n4453 0.8197
R29863 GNDA.n4475 GNDA.n4474 0.8197
R29864 GNDA.n4479 GNDA.n4478 0.8197
R29865 GNDA.n1498 GNDA.n1497 0.8197
R29866 GNDA.n1495 GNDA.n1494 0.8197
R29867 GNDA.n1491 GNDA.n1475 0.8197
R29868 GNDA.n1490 GNDA.n1487 0.8197
R29869 GNDA.n1483 GNDA.n1480 0.8197
R29870 GNDA.n1477 GNDA.n1401 0.8197
R29871 GNDA.n1505 GNDA.n1504 0.8197
R29872 GNDA.n1508 GNDA.n1400 0.8197
R29873 GNDA.n5007 GNDA.n5006 0.8197
R29874 GNDA.n5013 GNDA.n4929 0.8197
R29875 GNDA.n5012 GNDA.n4930 0.8197
R29876 GNDA.n4936 GNDA.n4935 0.8197
R29877 GNDA.n5172 GNDA.n5171 0.8197
R29878 GNDA.n892 GNDA.n891 0.8197
R29879 GNDA.n5180 GNDA.n887 0.8197
R29880 GNDA.n5179 GNDA.n888 0.8197
R29881 GNDA.n4440 GNDA.n1937 0.8197
R29882 GNDA.n4439 GNDA.n1938 0.8197
R29883 GNDA.n4358 GNDA.n4355 0.8197
R29884 GNDA.n4361 GNDA.n4360 0.8197
R29885 GNDA.n4371 GNDA.n4368 0.8197
R29886 GNDA.n4372 GNDA.n4354 0.8197
R29887 GNDA.n4376 GNDA.n4375 0.8197
R29888 GNDA.n4380 GNDA.n4379 0.8197
R29889 GNDA.n4151 GNDA.n4147 0.776542
R29890 GNDA.n4155 GNDA.n3656 0.776542
R29891 GNDA.n4159 GNDA.n3651 0.776542
R29892 GNDA.n4163 GNDA.n3646 0.776542
R29893 GNDA.n4171 GNDA.n3604 0.776542
R29894 GNDA.n4175 GNDA.n3599 0.776542
R29895 GNDA.n4179 GNDA.n3594 0.776542
R29896 GNDA.n5151 GNDA.n5150 0.776542
R29897 GNDA.n3400 GNDA.n3399 0.776542
R29898 GNDA.n3311 GNDA.n3310 0.776542
R29899 GNDA.n3142 GNDA.n3141 0.776542
R29900 GNDA.n3055 GNDA.n3054 0.776542
R29901 GNDA.n2918 GNDA.n2917 0.776542
R29902 GNDA.n2908 GNDA.n2907 0.776542
R29903 GNDA.n2821 GNDA.n2820 0.776542
R29904 GNDA.n2686 GNDA.n2685 0.776542
R29905 GNDA.n3152 GNDA.n3151 0.776542
R29906 GNDA.n4189 GNDA.n4188 0.77295
R29907 GNDA.n3289 GNDA.n3288 0.77295
R29908 GNDA.n4897 GNDA.n954 0.723198
R29909 GNDA.n3625 GNDA.n3620 0.688
R29910 GNDA.n2208 GNDA.n2203 0.688
R29911 GNDA.n5318 GNDA.n767 0.65675
R29912 GNDA.n2741 GNDA.n2653 0.655048
R29913 GNDA.n5541 GNDA.n5540 0.578165
R29914 GNDA.n611 GNDA.n578 0.576795
R29915 GNDA.n578 GNDA.n45 0.568015
R29916 GNDA.n5541 GNDA.n25 0.567378
R29917 GNDA.n5282 GNDA_2 0.5637
R29918 GNDA.n5353 GNDA_2 0.5637
R29919 GNDA_2 GNDA.n4636 0.5637
R29920 GNDA_2 GNDA.n1786 0.5637
R29921 GNDA.n4742 GNDA_2 0.5637
R29922 GNDA.n4464 GNDA_2 0.5637
R29923 GNDA_2 GNDA.n1476 0.5637
R29924 GNDA.n4933 GNDA_2 0.5637
R29925 GNDA.n4365 GNDA_2 0.5637
R29926 GNDA.n5405 GNDA.n5403 0.5005
R29927 GNDA.n5402 GNDA.n5399 0.5005
R29928 GNDA.n639 GNDA.n637 0.5005
R29929 GNDA.n636 GNDA.n633 0.5005
R29930 GNDA.n5020 GNDA.n745 0.458833
R29931 GNDA.n600 GNDA.n599 0.427583
R29932 GNDA.n5528 GNDA.n5527 0.427583
R29933 GNDA.n3620 GNDA.n3615 0.40675
R29934 GNDA.n2203 GNDA.n2198 0.40675
R29935 GNDA.n5535 GNDA.n5534 0.40675
R29936 GNDA.n608 GNDA.n607 0.40675
R29937 GNDA.n5446 GNDA.n688 0.359875
R29938 GNDA.n5491 GNDA.n5490 0.359875
R29939 GNDA.n5345 GNDA.n5344 0.34425
R29940 GNDA.n4274 GNDA.n1973 0.324972
R29941 GNDA.n3292 GNDA.n2113 0.32313
R29942 GNDA.n2562 GNDA.n2544 0.286759
R29943 GNDA.n4178 GNDA.n4176 0.28175
R29944 GNDA.n4174 GNDA.n4172 0.28175
R29945 GNDA.n4162 GNDA.n4160 0.28175
R29946 GNDA.n4158 GNDA.n4156 0.28175
R29947 GNDA.n4154 GNDA.n4152 0.28175
R29948 GNDA.n2823 GNDA.n2240 0.28175
R29949 GNDA.n2910 GNDA.n2825 0.28175
R29950 GNDA.n2914 GNDA.n2912 0.28175
R29951 GNDA.n3144 GNDA.n3059 0.28175
R29952 GNDA.n447 GNDA.n445 0.28175
R29953 GNDA.n368 GNDA.n367 0.28175
R29954 GNDA.n364 GNDA.n363 0.28175
R29955 GNDA.n360 GNDA.n359 0.28175
R29956 GNDA.n3296 GNDA.n2116 0.271333
R29957 GNDA.n5301 GNDA_2 0.2565
R29958 GNDA.n5372 GNDA_2 0.2565
R29959 GNDA.n4639 GNDA_2 0.2565
R29960 GNDA.n1794 GNDA_2 0.2565
R29961 GNDA.n4730 GNDA_2 0.2565
R29962 GNDA_2 GNDA.n4463 0.2565
R29963 GNDA.n1484 GNDA_2 0.2565
R29964 GNDA_2 GNDA.n4932 0.2565
R29965 GNDA_2 GNDA.n4364 0.2565
R29966 GNDA.n2650 GNDA.n2615 0.230359
R29967 GNDA.n5411 GNDA.n5410 0.229667
R29968 GNDA.n5492 GNDA.n663 0.229667
R29969 GNDA.n5453 GNDA.n5448 0.229667
R29970 GNDA.n5483 GNDA.n665 0.229667
R29971 GNDA.n5506 GNDA.n5505 0.229667
R29972 GNDA.n4924 GNDA.n4922 0.229667
R29973 GNDA.n5434 GNDA.n5432 0.214042
R29974 GNDA.n5443 GNDA.n5442 0.214042
R29975 GNDA.n5496 GNDA.n5495 0.214042
R29976 GNDA.n4275 GNDA.n1972 0.198417
R29977 GNDA.n3148 GNDA.n3146 0.198417
R29978 GNDA.n3307 GNDA.n3305 0.198417
R29979 GNDA.n5064 GNDA.n5063 0.188
R29980 GNDA.n5148 GNDA.n5147 0.188
R29981 GNDA.n4183 GNDA.n4180 0.188
R29982 GNDA.n5345 GNDA.n745 0.15675
R29983 GNDA.n5021 GNDA.n5020 0.151542
R29984 GNDA.n5343 GNDA.n5342 0.151542
R29985 GNDA.n5324 GNDA.n5323 0.147453
R29986 GNDA.n2034 GNDA.n2033 0.146333
R29987 GNDA.n2035 GNDA.n2034 0.146333
R29988 GNDA.n2036 GNDA.n2035 0.146333
R29989 GNDA.n2040 GNDA.n2039 0.146333
R29990 GNDA.n2041 GNDA.n2040 0.146333
R29991 GNDA.n2042 GNDA.n2041 0.146333
R29992 GNDA.n2046 GNDA.n2045 0.146333
R29993 GNDA.n2047 GNDA.n2046 0.146333
R29994 GNDA.n2048 GNDA.n2047 0.146333
R29995 GNDA.n2052 GNDA.n2051 0.146333
R29996 GNDA.n2053 GNDA.n2052 0.146333
R29997 GNDA.n2054 GNDA.n2053 0.146333
R29998 GNDA.n4145 GNDA.n4144 0.146333
R29999 GNDA.n4144 GNDA.n3665 0.146333
R30000 GNDA.n4140 GNDA.n3665 0.146333
R30001 GNDA.n4134 GNDA.n3670 0.146333
R30002 GNDA.n4134 GNDA.n4133 0.146333
R30003 GNDA.n4133 GNDA.n4132 0.146333
R30004 GNDA.n4127 GNDA.n4126 0.146333
R30005 GNDA.n4126 GNDA.n3680 0.146333
R30006 GNDA.n4122 GNDA.n3680 0.146333
R30007 GNDA.n4116 GNDA.n3685 0.146333
R30008 GNDA.n4116 GNDA.n4115 0.146333
R30009 GNDA.n4115 GNDA.n4114 0.146333
R30010 GNDA.n4050 GNDA.n4045 0.146333
R30011 GNDA.n4054 GNDA.n4045 0.146333
R30012 GNDA.n4055 GNDA.n4054 0.146333
R30013 GNDA.n4063 GNDA.n4062 0.146333
R30014 GNDA.n4066 GNDA.n4063 0.146333
R30015 GNDA.n4066 GNDA.n4037 0.146333
R30016 GNDA.n4074 GNDA.n4033 0.146333
R30017 GNDA.n4078 GNDA.n4033 0.146333
R30018 GNDA.n4079 GNDA.n4078 0.146333
R30019 GNDA.n4087 GNDA.n4086 0.146333
R30020 GNDA.n4090 GNDA.n4087 0.146333
R30021 GNDA.n4090 GNDA.n4027 0.146333
R30022 GNDA.n3969 GNDA.n3964 0.146333
R30023 GNDA.n3973 GNDA.n3964 0.146333
R30024 GNDA.n3974 GNDA.n3973 0.146333
R30025 GNDA.n3982 GNDA.n3981 0.146333
R30026 GNDA.n3985 GNDA.n3982 0.146333
R30027 GNDA.n3985 GNDA.n3956 0.146333
R30028 GNDA.n3993 GNDA.n3952 0.146333
R30029 GNDA.n3997 GNDA.n3952 0.146333
R30030 GNDA.n3998 GNDA.n3997 0.146333
R30031 GNDA.n4006 GNDA.n4005 0.146333
R30032 GNDA.n4009 GNDA.n4006 0.146333
R30033 GNDA.n4009 GNDA.n3946 0.146333
R30034 GNDA.n3888 GNDA.n3883 0.146333
R30035 GNDA.n3892 GNDA.n3883 0.146333
R30036 GNDA.n3893 GNDA.n3892 0.146333
R30037 GNDA.n3901 GNDA.n3900 0.146333
R30038 GNDA.n3904 GNDA.n3901 0.146333
R30039 GNDA.n3904 GNDA.n3875 0.146333
R30040 GNDA.n3912 GNDA.n3871 0.146333
R30041 GNDA.n3916 GNDA.n3871 0.146333
R30042 GNDA.n3917 GNDA.n3916 0.146333
R30043 GNDA.n3925 GNDA.n3924 0.146333
R30044 GNDA.n3928 GNDA.n3925 0.146333
R30045 GNDA.n3928 GNDA.n3865 0.146333
R30046 GNDA.n4192 GNDA.n3506 0.146333
R30047 GNDA.n4196 GNDA.n3506 0.146333
R30048 GNDA.n4197 GNDA.n4196 0.146333
R30049 GNDA.n4205 GNDA.n4204 0.146333
R30050 GNDA.n4208 GNDA.n4205 0.146333
R30051 GNDA.n4208 GNDA.n3498 0.146333
R30052 GNDA.n4216 GNDA.n3494 0.146333
R30053 GNDA.n4220 GNDA.n3494 0.146333
R30054 GNDA.n4221 GNDA.n4220 0.146333
R30055 GNDA.n4229 GNDA.n4228 0.146333
R30056 GNDA.n4232 GNDA.n4229 0.146333
R30057 GNDA.n4232 GNDA.n3488 0.146333
R30058 GNDA.n3807 GNDA.n3802 0.146333
R30059 GNDA.n3811 GNDA.n3802 0.146333
R30060 GNDA.n3812 GNDA.n3811 0.146333
R30061 GNDA.n3820 GNDA.n3819 0.146333
R30062 GNDA.n3823 GNDA.n3820 0.146333
R30063 GNDA.n3823 GNDA.n3794 0.146333
R30064 GNDA.n3831 GNDA.n3790 0.146333
R30065 GNDA.n3835 GNDA.n3790 0.146333
R30066 GNDA.n3836 GNDA.n3835 0.146333
R30067 GNDA.n3844 GNDA.n3843 0.146333
R30068 GNDA.n3847 GNDA.n3844 0.146333
R30069 GNDA.n3847 GNDA.n3784 0.146333
R30070 GNDA.n3726 GNDA.n3721 0.146333
R30071 GNDA.n3730 GNDA.n3721 0.146333
R30072 GNDA.n3731 GNDA.n3730 0.146333
R30073 GNDA.n3739 GNDA.n3738 0.146333
R30074 GNDA.n3742 GNDA.n3739 0.146333
R30075 GNDA.n3742 GNDA.n3713 0.146333
R30076 GNDA.n3750 GNDA.n3709 0.146333
R30077 GNDA.n3754 GNDA.n3709 0.146333
R30078 GNDA.n3755 GNDA.n3754 0.146333
R30079 GNDA.n3763 GNDA.n3762 0.146333
R30080 GNDA.n3766 GNDA.n3763 0.146333
R30081 GNDA.n3766 GNDA.n3703 0.146333
R30082 GNDA.n3592 GNDA.n3591 0.146333
R30083 GNDA.n3591 GNDA.n3519 0.146333
R30084 GNDA.n3587 GNDA.n3519 0.146333
R30085 GNDA.n3581 GNDA.n3527 0.146333
R30086 GNDA.n3581 GNDA.n3580 0.146333
R30087 GNDA.n3580 GNDA.n3579 0.146333
R30088 GNDA.n3574 GNDA.n3573 0.146333
R30089 GNDA.n3573 GNDA.n3543 0.146333
R30090 GNDA.n3569 GNDA.n3543 0.146333
R30091 GNDA.n3563 GNDA.n3551 0.146333
R30092 GNDA.n3563 GNDA.n3562 0.146333
R30093 GNDA.n3562 GNDA.n3561 0.146333
R30094 GNDA.n4271 GNDA.n4270 0.146333
R30095 GNDA.n4270 GNDA.n1978 0.146333
R30096 GNDA.n4266 GNDA.n1978 0.146333
R30097 GNDA.n4260 GNDA.n1983 0.146333
R30098 GNDA.n4260 GNDA.n4259 0.146333
R30099 GNDA.n4259 GNDA.n4258 0.146333
R30100 GNDA.n4253 GNDA.n4252 0.146333
R30101 GNDA.n4252 GNDA.n1993 0.146333
R30102 GNDA.n4248 GNDA.n1993 0.146333
R30103 GNDA.n4242 GNDA.n1998 0.146333
R30104 GNDA.n4242 GNDA.n4241 0.146333
R30105 GNDA.n4241 GNDA.n4240 0.146333
R30106 GNDA.n1065 GNDA.n1061 0.146333
R30107 GNDA.n1069 GNDA.n1061 0.146333
R30108 GNDA.n1070 GNDA.n1069 0.146333
R30109 GNDA.n1078 GNDA.n1077 0.146333
R30110 GNDA.n1081 GNDA.n1078 0.146333
R30111 GNDA.n1081 GNDA.n1053 0.146333
R30112 GNDA.n1089 GNDA.n1049 0.146333
R30113 GNDA.n1093 GNDA.n1049 0.146333
R30114 GNDA.n1094 GNDA.n1093 0.146333
R30115 GNDA.n1102 GNDA.n1101 0.146333
R30116 GNDA.n1105 GNDA.n1102 0.146333
R30117 GNDA.n1105 GNDA.n1043 0.146333
R30118 GNDA.n3403 GNDA.n3392 0.146333
R30119 GNDA.n3409 GNDA.n3392 0.146333
R30120 GNDA.n3410 GNDA.n3409 0.146333
R30121 GNDA.n3420 GNDA.n3419 0.146333
R30122 GNDA.n3423 GNDA.n3420 0.146333
R30123 GNDA.n3423 GNDA.n3388 0.146333
R30124 GNDA.n3433 GNDA.n3386 0.146333
R30125 GNDA.n3439 GNDA.n3386 0.146333
R30126 GNDA.n3440 GNDA.n3439 0.146333
R30127 GNDA.n3450 GNDA.n3449 0.146333
R30128 GNDA.n3453 GNDA.n3450 0.146333
R30129 GNDA.n3453 GNDA.n3382 0.146333
R30130 GNDA.n3314 GNDA.n2027 0.146333
R30131 GNDA.n3320 GNDA.n2027 0.146333
R30132 GNDA.n3321 GNDA.n3320 0.146333
R30133 GNDA.n3331 GNDA.n3330 0.146333
R30134 GNDA.n3334 GNDA.n3331 0.146333
R30135 GNDA.n3334 GNDA.n2023 0.146333
R30136 GNDA.n3344 GNDA.n2021 0.146333
R30137 GNDA.n3350 GNDA.n2021 0.146333
R30138 GNDA.n3351 GNDA.n3350 0.146333
R30139 GNDA.n3361 GNDA.n3360 0.146333
R30140 GNDA.n3364 GNDA.n3361 0.146333
R30141 GNDA.n3364 GNDA.n2017 0.146333
R30142 GNDA.n3232 GNDA.n2120 0.146333
R30143 GNDA.n3237 GNDA.n3232 0.146333
R30144 GNDA.n3238 GNDA.n3237 0.146333
R30145 GNDA.n3248 GNDA.n3247 0.146333
R30146 GNDA.n3251 GNDA.n3248 0.146333
R30147 GNDA.n3251 GNDA.n3228 0.146333
R30148 GNDA.n3261 GNDA.n3226 0.146333
R30149 GNDA.n3267 GNDA.n3226 0.146333
R30150 GNDA.n3268 GNDA.n3267 0.146333
R30151 GNDA.n3278 GNDA.n3277 0.146333
R30152 GNDA.n3281 GNDA.n3278 0.146333
R30153 GNDA.n3281 GNDA.n3222 0.146333
R30154 GNDA.n3155 GNDA.n2146 0.146333
R30155 GNDA.n3161 GNDA.n2146 0.146333
R30156 GNDA.n3162 GNDA.n3161 0.146333
R30157 GNDA.n3172 GNDA.n3171 0.146333
R30158 GNDA.n3175 GNDA.n3172 0.146333
R30159 GNDA.n3175 GNDA.n2142 0.146333
R30160 GNDA.n3185 GNDA.n2140 0.146333
R30161 GNDA.n3191 GNDA.n2140 0.146333
R30162 GNDA.n3192 GNDA.n3191 0.146333
R30163 GNDA.n3202 GNDA.n3201 0.146333
R30164 GNDA.n3205 GNDA.n3202 0.146333
R30165 GNDA.n3205 GNDA.n2136 0.146333
R30166 GNDA.n3063 GNDA.n3062 0.146333
R30167 GNDA.n3064 GNDA.n3063 0.146333
R30168 GNDA.n3065 GNDA.n3064 0.146333
R30169 GNDA.n3069 GNDA.n3068 0.146333
R30170 GNDA.n3070 GNDA.n3069 0.146333
R30171 GNDA.n3071 GNDA.n3070 0.146333
R30172 GNDA.n3075 GNDA.n3074 0.146333
R30173 GNDA.n3076 GNDA.n3075 0.146333
R30174 GNDA.n3077 GNDA.n3076 0.146333
R30175 GNDA.n3081 GNDA.n3080 0.146333
R30176 GNDA.n3082 GNDA.n3081 0.146333
R30177 GNDA.n3083 GNDA.n3082 0.146333
R30178 GNDA.n2998 GNDA.n2159 0.146333
R30179 GNDA.n3003 GNDA.n2998 0.146333
R30180 GNDA.n3004 GNDA.n3003 0.146333
R30181 GNDA.n3014 GNDA.n3013 0.146333
R30182 GNDA.n3017 GNDA.n3014 0.146333
R30183 GNDA.n3017 GNDA.n2994 0.146333
R30184 GNDA.n3027 GNDA.n2992 0.146333
R30185 GNDA.n3033 GNDA.n2992 0.146333
R30186 GNDA.n3034 GNDA.n3033 0.146333
R30187 GNDA.n3044 GNDA.n3043 0.146333
R30188 GNDA.n3047 GNDA.n3044 0.146333
R30189 GNDA.n3047 GNDA.n2988 0.146333
R30190 GNDA.n2921 GNDA.n2185 0.146333
R30191 GNDA.n2927 GNDA.n2185 0.146333
R30192 GNDA.n2928 GNDA.n2927 0.146333
R30193 GNDA.n2938 GNDA.n2937 0.146333
R30194 GNDA.n2941 GNDA.n2938 0.146333
R30195 GNDA.n2941 GNDA.n2181 0.146333
R30196 GNDA.n2951 GNDA.n2179 0.146333
R30197 GNDA.n2957 GNDA.n2179 0.146333
R30198 GNDA.n2958 GNDA.n2957 0.146333
R30199 GNDA.n2968 GNDA.n2967 0.146333
R30200 GNDA.n2971 GNDA.n2968 0.146333
R30201 GNDA.n2971 GNDA.n2175 0.146333
R30202 GNDA.n2829 GNDA.n2828 0.146333
R30203 GNDA.n2830 GNDA.n2829 0.146333
R30204 GNDA.n2831 GNDA.n2830 0.146333
R30205 GNDA.n2835 GNDA.n2834 0.146333
R30206 GNDA.n2836 GNDA.n2835 0.146333
R30207 GNDA.n2837 GNDA.n2836 0.146333
R30208 GNDA.n2841 GNDA.n2840 0.146333
R30209 GNDA.n2842 GNDA.n2841 0.146333
R30210 GNDA.n2843 GNDA.n2842 0.146333
R30211 GNDA.n2847 GNDA.n2846 0.146333
R30212 GNDA.n2848 GNDA.n2847 0.146333
R30213 GNDA.n2849 GNDA.n2848 0.146333
R30214 GNDA.n2764 GNDA.n2243 0.146333
R30215 GNDA.n2769 GNDA.n2764 0.146333
R30216 GNDA.n2770 GNDA.n2769 0.146333
R30217 GNDA.n2780 GNDA.n2779 0.146333
R30218 GNDA.n2783 GNDA.n2780 0.146333
R30219 GNDA.n2783 GNDA.n2760 0.146333
R30220 GNDA.n2793 GNDA.n2758 0.146333
R30221 GNDA.n2799 GNDA.n2758 0.146333
R30222 GNDA.n2800 GNDA.n2799 0.146333
R30223 GNDA.n2810 GNDA.n2809 0.146333
R30224 GNDA.n2813 GNDA.n2810 0.146333
R30225 GNDA.n2813 GNDA.n2754 0.146333
R30226 GNDA.n2691 GNDA.n2688 0.146333
R30227 GNDA.n2694 GNDA.n2691 0.146333
R30228 GNDA.n2694 GNDA.n2676 0.146333
R30229 GNDA.n2704 GNDA.n2674 0.146333
R30230 GNDA.n2708 GNDA.n2674 0.146333
R30231 GNDA.n2711 GNDA.n2708 0.146333
R30232 GNDA.n2721 GNDA.n2718 0.146333
R30233 GNDA.n2724 GNDA.n2721 0.146333
R30234 GNDA.n2724 GNDA.n2670 0.146333
R30235 GNDA.n2733 GNDA.n2667 0.146333
R30236 GNDA.n2738 GNDA.n2667 0.146333
R30237 GNDA.n2738 GNDA.n2668 0.146333
R30238 GNDA.n5545 GNDA.n24 0.146333
R30239 GNDA.n5551 GNDA.n24 0.146333
R30240 GNDA.n5552 GNDA.n5551 0.146333
R30241 GNDA.n5562 GNDA.n5561 0.146333
R30242 GNDA.n5565 GNDA.n5562 0.146333
R30243 GNDA.n5565 GNDA.n20 0.146333
R30244 GNDA.n5575 GNDA.n18 0.146333
R30245 GNDA.n5581 GNDA.n18 0.146333
R30246 GNDA.n5582 GNDA.n5581 0.146333
R30247 GNDA.n5592 GNDA.n5591 0.146333
R30248 GNDA.n5595 GNDA.n5592 0.146333
R30249 GNDA.n5595 GNDA.n14 0.146333
R30250 GNDA.n521 GNDA.n47 0.146333
R30251 GNDA.n526 GNDA.n521 0.146333
R30252 GNDA.n527 GNDA.n526 0.146333
R30253 GNDA.n537 GNDA.n536 0.146333
R30254 GNDA.n540 GNDA.n537 0.146333
R30255 GNDA.n540 GNDA.n517 0.146333
R30256 GNDA.n550 GNDA.n515 0.146333
R30257 GNDA.n556 GNDA.n515 0.146333
R30258 GNDA.n557 GNDA.n556 0.146333
R30259 GNDA.n567 GNDA.n566 0.146333
R30260 GNDA.n570 GNDA.n567 0.146333
R30261 GNDA.n570 GNDA.n511 0.146333
R30262 GNDA.n275 GNDA.n274 0.146333
R30263 GNDA.n276 GNDA.n275 0.146333
R30264 GNDA.n277 GNDA.n276 0.146333
R30265 GNDA.n281 GNDA.n280 0.146333
R30266 GNDA.n282 GNDA.n281 0.146333
R30267 GNDA.n283 GNDA.n282 0.146333
R30268 GNDA.n287 GNDA.n286 0.146333
R30269 GNDA.n288 GNDA.n287 0.146333
R30270 GNDA.n289 GNDA.n288 0.146333
R30271 GNDA.n293 GNDA.n292 0.146333
R30272 GNDA.n294 GNDA.n293 0.146333
R30273 GNDA.n295 GNDA.n294 0.146333
R30274 GNDA.n211 GNDA.n187 0.146333
R30275 GNDA.n216 GNDA.n211 0.146333
R30276 GNDA.n217 GNDA.n216 0.146333
R30277 GNDA.n227 GNDA.n226 0.146333
R30278 GNDA.n230 GNDA.n227 0.146333
R30279 GNDA.n230 GNDA.n207 0.146333
R30280 GNDA.n240 GNDA.n205 0.146333
R30281 GNDA.n246 GNDA.n205 0.146333
R30282 GNDA.n247 GNDA.n246 0.146333
R30283 GNDA.n257 GNDA.n256 0.146333
R30284 GNDA.n260 GNDA.n257 0.146333
R30285 GNDA.n260 GNDA.n201 0.146333
R30286 GNDA.n102 GNDA.n101 0.146333
R30287 GNDA.n103 GNDA.n102 0.146333
R30288 GNDA.n104 GNDA.n103 0.146333
R30289 GNDA.n108 GNDA.n107 0.146333
R30290 GNDA.n109 GNDA.n108 0.146333
R30291 GNDA.n110 GNDA.n109 0.146333
R30292 GNDA.n114 GNDA.n113 0.146333
R30293 GNDA.n115 GNDA.n114 0.146333
R30294 GNDA.n116 GNDA.n115 0.146333
R30295 GNDA.n120 GNDA.n119 0.146333
R30296 GNDA.n121 GNDA.n120 0.146333
R30297 GNDA.n122 GNDA.n121 0.146333
R30298 GNDA.n454 GNDA.n96 0.146333
R30299 GNDA.n460 GNDA.n96 0.146333
R30300 GNDA.n461 GNDA.n460 0.146333
R30301 GNDA.n471 GNDA.n470 0.146333
R30302 GNDA.n474 GNDA.n471 0.146333
R30303 GNDA.n474 GNDA.n92 0.146333
R30304 GNDA.n484 GNDA.n90 0.146333
R30305 GNDA.n490 GNDA.n90 0.146333
R30306 GNDA.n491 GNDA.n490 0.146333
R30307 GNDA.n501 GNDA.n500 0.146333
R30308 GNDA.n504 GNDA.n501 0.146333
R30309 GNDA.n504 GNDA.n86 0.146333
R30310 GNDA.n441 GNDA.n440 0.146333
R30311 GNDA.n440 GNDA.n379 0.146333
R30312 GNDA.n436 GNDA.n379 0.146333
R30313 GNDA.n430 GNDA.n385 0.146333
R30314 GNDA.n430 GNDA.n429 0.146333
R30315 GNDA.n429 GNDA.n428 0.146333
R30316 GNDA.n423 GNDA.n422 0.146333
R30317 GNDA.n422 GNDA.n397 0.146333
R30318 GNDA.n418 GNDA.n397 0.146333
R30319 GNDA.n412 GNDA.n403 0.146333
R30320 GNDA.n412 GNDA.n411 0.146333
R30321 GNDA.n411 GNDA.n410 0.146333
R30322 GNDA.n984 GNDA.n976 0.146333
R30323 GNDA.n985 GNDA.n984 0.146333
R30324 GNDA.n995 GNDA.n994 0.146333
R30325 GNDA.n996 GNDA.n995 0.146333
R30326 GNDA.n996 GNDA.n972 0.146333
R30327 GNDA.n1006 GNDA.n970 0.146333
R30328 GNDA.n1014 GNDA.n970 0.146333
R30329 GNDA.n1015 GNDA.n1014 0.146333
R30330 GNDA.n1025 GNDA.n1024 0.146333
R30331 GNDA.n1026 GNDA.n1025 0.146333
R30332 GNDA.n1026 GNDA.n951 0.146333
R30333 GNDA.n980 GNDA.n979 0.146333
R30334 GNDA.n983 GNDA.n980 0.146333
R30335 GNDA.n983 GNDA.n975 0.146333
R30336 GNDA.n993 GNDA.n973 0.146333
R30337 GNDA.n999 GNDA.n973 0.146333
R30338 GNDA.n1000 GNDA.n999 0.146333
R30339 GNDA.n1010 GNDA.n1009 0.146333
R30340 GNDA.n1013 GNDA.n1010 0.146333
R30341 GNDA.n1013 GNDA.n969 0.146333
R30342 GNDA.n1023 GNDA.n967 0.146333
R30343 GNDA.n1027 GNDA.n967 0.146333
R30344 GNDA.n1027 GNDA.n952 0.146333
R30345 GNDA.n2111 GNDA.n2033 0.135917
R30346 GNDA.n2037 GNDA.n2036 0.135917
R30347 GNDA.n2039 GNDA.n2038 0.135917
R30348 GNDA.n2043 GNDA.n2042 0.135917
R30349 GNDA.n2045 GNDA.n2044 0.135917
R30350 GNDA.n2049 GNDA.n2048 0.135917
R30351 GNDA.n2051 GNDA.n2050 0.135917
R30352 GNDA.n4146 GNDA.n4145 0.135917
R30353 GNDA.n4140 GNDA.n4139 0.135917
R30354 GNDA.n4138 GNDA.n3670 0.135917
R30355 GNDA.n4132 GNDA.n3675 0.135917
R30356 GNDA.n4128 GNDA.n4127 0.135917
R30357 GNDA.n4122 GNDA.n4121 0.135917
R30358 GNDA.n4120 GNDA.n3685 0.135917
R30359 GNDA.n4050 GNDA.n4048 0.135917
R30360 GNDA.n4058 GNDA.n4055 0.135917
R30361 GNDA.n4062 GNDA.n4041 0.135917
R30362 GNDA.n4070 GNDA.n4037 0.135917
R30363 GNDA.n4074 GNDA.n4071 0.135917
R30364 GNDA.n4082 GNDA.n4079 0.135917
R30365 GNDA.n4086 GNDA.n4029 0.135917
R30366 GNDA.n3969 GNDA.n3967 0.135917
R30367 GNDA.n3977 GNDA.n3974 0.135917
R30368 GNDA.n3981 GNDA.n3960 0.135917
R30369 GNDA.n3989 GNDA.n3956 0.135917
R30370 GNDA.n3993 GNDA.n3990 0.135917
R30371 GNDA.n4001 GNDA.n3998 0.135917
R30372 GNDA.n4005 GNDA.n3948 0.135917
R30373 GNDA.n3888 GNDA.n3886 0.135917
R30374 GNDA.n3896 GNDA.n3893 0.135917
R30375 GNDA.n3900 GNDA.n3879 0.135917
R30376 GNDA.n3908 GNDA.n3875 0.135917
R30377 GNDA.n3912 GNDA.n3909 0.135917
R30378 GNDA.n3920 GNDA.n3917 0.135917
R30379 GNDA.n3924 GNDA.n3867 0.135917
R30380 GNDA.n4192 GNDA.n4190 0.135917
R30381 GNDA.n4200 GNDA.n4197 0.135917
R30382 GNDA.n4204 GNDA.n3502 0.135917
R30383 GNDA.n4212 GNDA.n3498 0.135917
R30384 GNDA.n4216 GNDA.n4213 0.135917
R30385 GNDA.n4224 GNDA.n4221 0.135917
R30386 GNDA.n4228 GNDA.n3490 0.135917
R30387 GNDA.n3807 GNDA.n3805 0.135917
R30388 GNDA.n3815 GNDA.n3812 0.135917
R30389 GNDA.n3819 GNDA.n3798 0.135917
R30390 GNDA.n3827 GNDA.n3794 0.135917
R30391 GNDA.n3831 GNDA.n3828 0.135917
R30392 GNDA.n3839 GNDA.n3836 0.135917
R30393 GNDA.n3843 GNDA.n3786 0.135917
R30394 GNDA.n3726 GNDA.n3724 0.135917
R30395 GNDA.n3734 GNDA.n3731 0.135917
R30396 GNDA.n3738 GNDA.n3717 0.135917
R30397 GNDA.n3746 GNDA.n3713 0.135917
R30398 GNDA.n3750 GNDA.n3747 0.135917
R30399 GNDA.n3758 GNDA.n3755 0.135917
R30400 GNDA.n3762 GNDA.n3705 0.135917
R30401 GNDA.n3593 GNDA.n3592 0.135917
R30402 GNDA.n3587 GNDA.n3586 0.135917
R30403 GNDA.n3585 GNDA.n3527 0.135917
R30404 GNDA.n3579 GNDA.n3535 0.135917
R30405 GNDA.n3575 GNDA.n3574 0.135917
R30406 GNDA.n3569 GNDA.n3568 0.135917
R30407 GNDA.n3567 GNDA.n3551 0.135917
R30408 GNDA.n4272 GNDA.n4271 0.135917
R30409 GNDA.n4266 GNDA.n4265 0.135917
R30410 GNDA.n4264 GNDA.n1983 0.135917
R30411 GNDA.n4258 GNDA.n1988 0.135917
R30412 GNDA.n4254 GNDA.n4253 0.135917
R30413 GNDA.n4248 GNDA.n4247 0.135917
R30414 GNDA.n4246 GNDA.n1998 0.135917
R30415 GNDA.n1073 GNDA.n1070 0.135917
R30416 GNDA.n1077 GNDA.n1057 0.135917
R30417 GNDA.n1085 GNDA.n1053 0.135917
R30418 GNDA.n1089 GNDA.n1086 0.135917
R30419 GNDA.n1097 GNDA.n1094 0.135917
R30420 GNDA.n1101 GNDA.n1045 0.135917
R30421 GNDA.n4894 GNDA.n1043 0.135917
R30422 GNDA.n3403 GNDA.n3401 0.135917
R30423 GNDA.n3413 GNDA.n3410 0.135917
R30424 GNDA.n3419 GNDA.n3390 0.135917
R30425 GNDA.n3429 GNDA.n3388 0.135917
R30426 GNDA.n3433 GNDA.n3430 0.135917
R30427 GNDA.n3443 GNDA.n3440 0.135917
R30428 GNDA.n3449 GNDA.n3384 0.135917
R30429 GNDA.n3314 GNDA.n3312 0.135917
R30430 GNDA.n3324 GNDA.n3321 0.135917
R30431 GNDA.n3330 GNDA.n2025 0.135917
R30432 GNDA.n3340 GNDA.n2023 0.135917
R30433 GNDA.n3344 GNDA.n3341 0.135917
R30434 GNDA.n3354 GNDA.n3351 0.135917
R30435 GNDA.n3360 GNDA.n2019 0.135917
R30436 GNDA.n3287 GNDA.n2120 0.135917
R30437 GNDA.n3241 GNDA.n3238 0.135917
R30438 GNDA.n3247 GNDA.n3230 0.135917
R30439 GNDA.n3257 GNDA.n3228 0.135917
R30440 GNDA.n3261 GNDA.n3258 0.135917
R30441 GNDA.n3271 GNDA.n3268 0.135917
R30442 GNDA.n3277 GNDA.n3224 0.135917
R30443 GNDA.n3155 GNDA.n3153 0.135917
R30444 GNDA.n3165 GNDA.n3162 0.135917
R30445 GNDA.n3171 GNDA.n2144 0.135917
R30446 GNDA.n3181 GNDA.n2142 0.135917
R30447 GNDA.n3185 GNDA.n3182 0.135917
R30448 GNDA.n3195 GNDA.n3192 0.135917
R30449 GNDA.n3201 GNDA.n2138 0.135917
R30450 GNDA.n3140 GNDA.n3062 0.135917
R30451 GNDA.n3066 GNDA.n3065 0.135917
R30452 GNDA.n3068 GNDA.n3067 0.135917
R30453 GNDA.n3072 GNDA.n3071 0.135917
R30454 GNDA.n3074 GNDA.n3073 0.135917
R30455 GNDA.n3078 GNDA.n3077 0.135917
R30456 GNDA.n3080 GNDA.n3079 0.135917
R30457 GNDA.n3053 GNDA.n2159 0.135917
R30458 GNDA.n3007 GNDA.n3004 0.135917
R30459 GNDA.n3013 GNDA.n2996 0.135917
R30460 GNDA.n3023 GNDA.n2994 0.135917
R30461 GNDA.n3027 GNDA.n3024 0.135917
R30462 GNDA.n3037 GNDA.n3034 0.135917
R30463 GNDA.n3043 GNDA.n2990 0.135917
R30464 GNDA.n2921 GNDA.n2919 0.135917
R30465 GNDA.n2931 GNDA.n2928 0.135917
R30466 GNDA.n2937 GNDA.n2183 0.135917
R30467 GNDA.n2947 GNDA.n2181 0.135917
R30468 GNDA.n2951 GNDA.n2948 0.135917
R30469 GNDA.n2961 GNDA.n2958 0.135917
R30470 GNDA.n2967 GNDA.n2177 0.135917
R30471 GNDA.n2906 GNDA.n2828 0.135917
R30472 GNDA.n2832 GNDA.n2831 0.135917
R30473 GNDA.n2834 GNDA.n2833 0.135917
R30474 GNDA.n2838 GNDA.n2837 0.135917
R30475 GNDA.n2840 GNDA.n2839 0.135917
R30476 GNDA.n2844 GNDA.n2843 0.135917
R30477 GNDA.n2846 GNDA.n2845 0.135917
R30478 GNDA.n2819 GNDA.n2243 0.135917
R30479 GNDA.n2773 GNDA.n2770 0.135917
R30480 GNDA.n2779 GNDA.n2762 0.135917
R30481 GNDA.n2789 GNDA.n2760 0.135917
R30482 GNDA.n2793 GNDA.n2790 0.135917
R30483 GNDA.n2803 GNDA.n2800 0.135917
R30484 GNDA.n2809 GNDA.n2756 0.135917
R30485 GNDA.n2688 GNDA.n2678 0.135917
R30486 GNDA.n2698 GNDA.n2676 0.135917
R30487 GNDA.n2704 GNDA.n2701 0.135917
R30488 GNDA.n2714 GNDA.n2711 0.135917
R30489 GNDA.n2718 GNDA.n2672 0.135917
R30490 GNDA.n2728 GNDA.n2670 0.135917
R30491 GNDA.n2733 GNDA.n2731 0.135917
R30492 GNDA.n5545 GNDA.n5543 0.135917
R30493 GNDA.n5555 GNDA.n5552 0.135917
R30494 GNDA.n5561 GNDA.n22 0.135917
R30495 GNDA.n5571 GNDA.n20 0.135917
R30496 GNDA.n5575 GNDA.n5572 0.135917
R30497 GNDA.n5585 GNDA.n5582 0.135917
R30498 GNDA.n5591 GNDA.n16 0.135917
R30499 GNDA.n576 GNDA.n47 0.135917
R30500 GNDA.n530 GNDA.n527 0.135917
R30501 GNDA.n536 GNDA.n519 0.135917
R30502 GNDA.n546 GNDA.n517 0.135917
R30503 GNDA.n550 GNDA.n547 0.135917
R30504 GNDA.n560 GNDA.n557 0.135917
R30505 GNDA.n566 GNDA.n513 0.135917
R30506 GNDA.n352 GNDA.n274 0.135917
R30507 GNDA.n278 GNDA.n277 0.135917
R30508 GNDA.n280 GNDA.n279 0.135917
R30509 GNDA.n284 GNDA.n283 0.135917
R30510 GNDA.n286 GNDA.n285 0.135917
R30511 GNDA.n290 GNDA.n289 0.135917
R30512 GNDA.n292 GNDA.n291 0.135917
R30513 GNDA.n266 GNDA.n187 0.135917
R30514 GNDA.n220 GNDA.n217 0.135917
R30515 GNDA.n226 GNDA.n209 0.135917
R30516 GNDA.n236 GNDA.n207 0.135917
R30517 GNDA.n240 GNDA.n237 0.135917
R30518 GNDA.n250 GNDA.n247 0.135917
R30519 GNDA.n256 GNDA.n203 0.135917
R30520 GNDA.n179 GNDA.n101 0.135917
R30521 GNDA.n105 GNDA.n104 0.135917
R30522 GNDA.n107 GNDA.n106 0.135917
R30523 GNDA.n111 GNDA.n110 0.135917
R30524 GNDA.n113 GNDA.n112 0.135917
R30525 GNDA.n117 GNDA.n116 0.135917
R30526 GNDA.n119 GNDA.n118 0.135917
R30527 GNDA.n454 GNDA.n452 0.135917
R30528 GNDA.n464 GNDA.n461 0.135917
R30529 GNDA.n470 GNDA.n94 0.135917
R30530 GNDA.n480 GNDA.n92 0.135917
R30531 GNDA.n484 GNDA.n481 0.135917
R30532 GNDA.n494 GNDA.n491 0.135917
R30533 GNDA.n500 GNDA.n88 0.135917
R30534 GNDA.n442 GNDA.n441 0.135917
R30535 GNDA.n436 GNDA.n435 0.135917
R30536 GNDA.n434 GNDA.n385 0.135917
R30537 GNDA.n428 GNDA.n391 0.135917
R30538 GNDA.n424 GNDA.n423 0.135917
R30539 GNDA.n418 GNDA.n417 0.135917
R30540 GNDA.n416 GNDA.n403 0.135917
R30541 GNDA.n986 GNDA.n985 0.135917
R30542 GNDA.n994 GNDA.n974 0.135917
R30543 GNDA.n1004 GNDA.n972 0.135917
R30544 GNDA.n1006 GNDA.n1005 0.135917
R30545 GNDA.n1016 GNDA.n1015 0.135917
R30546 GNDA.n1024 GNDA.n968 0.135917
R30547 GNDA.n4900 GNDA.n951 0.135917
R30548 GNDA.n989 GNDA.n975 0.135917
R30549 GNDA.n993 GNDA.n990 0.135917
R30550 GNDA.n1003 GNDA.n1000 0.135917
R30551 GNDA.n1009 GNDA.n971 0.135917
R30552 GNDA.n1019 GNDA.n969 0.135917
R30553 GNDA.n1023 GNDA.n1020 0.135917
R30554 GNDA.n4899 GNDA.n952 0.135917
R30555 GNDA.n4897 GNDA.n4896 0.135331
R30556 GNDA.n4275 GNDA.n4274 0.125674
R30557 GNDA.n3305 GNDA.n2113 0.125568
R30558 GNDA.n2038 GNDA.n2037 0.1255
R30559 GNDA.n2044 GNDA.n2043 0.1255
R30560 GNDA.n2050 GNDA.n2049 0.1255
R30561 GNDA.n4139 GNDA.n4138 0.1255
R30562 GNDA.n4128 GNDA.n3675 0.1255
R30563 GNDA.n4121 GNDA.n4120 0.1255
R30564 GNDA.n4058 GNDA.n4041 0.1255
R30565 GNDA.n4071 GNDA.n4070 0.1255
R30566 GNDA.n4082 GNDA.n4029 0.1255
R30567 GNDA.n3977 GNDA.n3960 0.1255
R30568 GNDA.n3990 GNDA.n3989 0.1255
R30569 GNDA.n4001 GNDA.n3948 0.1255
R30570 GNDA.n3896 GNDA.n3879 0.1255
R30571 GNDA.n3909 GNDA.n3908 0.1255
R30572 GNDA.n3920 GNDA.n3867 0.1255
R30573 GNDA.n4200 GNDA.n3502 0.1255
R30574 GNDA.n4213 GNDA.n4212 0.1255
R30575 GNDA.n4224 GNDA.n3490 0.1255
R30576 GNDA.n3815 GNDA.n3798 0.1255
R30577 GNDA.n3828 GNDA.n3827 0.1255
R30578 GNDA.n3839 GNDA.n3786 0.1255
R30579 GNDA.n3734 GNDA.n3717 0.1255
R30580 GNDA.n3747 GNDA.n3746 0.1255
R30581 GNDA.n3758 GNDA.n3705 0.1255
R30582 GNDA.n3586 GNDA.n3585 0.1255
R30583 GNDA.n3575 GNDA.n3535 0.1255
R30584 GNDA.n3568 GNDA.n3567 0.1255
R30585 GNDA.n4265 GNDA.n4264 0.1255
R30586 GNDA.n4254 GNDA.n1988 0.1255
R30587 GNDA.n4247 GNDA.n4246 0.1255
R30588 GNDA.n5146 GNDA.n5068 0.1255
R30589 GNDA.n5062 GNDA.n5055 0.1255
R30590 GNDA.n1073 GNDA.n1057 0.1255
R30591 GNDA.n1086 GNDA.n1085 0.1255
R30592 GNDA.n1097 GNDA.n1045 0.1255
R30593 GNDA.n4884 GNDA.n1110 0.1255
R30594 GNDA.n4170 GNDA.n4168 0.1255
R30595 GNDA.n3413 GNDA.n3390 0.1255
R30596 GNDA.n3430 GNDA.n3429 0.1255
R30597 GNDA.n3443 GNDA.n3384 0.1255
R30598 GNDA.n3324 GNDA.n2025 0.1255
R30599 GNDA.n3341 GNDA.n3340 0.1255
R30600 GNDA.n3354 GNDA.n2019 0.1255
R30601 GNDA.n3241 GNDA.n3230 0.1255
R30602 GNDA.n3258 GNDA.n3257 0.1255
R30603 GNDA.n3271 GNDA.n3224 0.1255
R30604 GNDA.n3165 GNDA.n2144 0.1255
R30605 GNDA.n3182 GNDA.n3181 0.1255
R30606 GNDA.n3195 GNDA.n2138 0.1255
R30607 GNDA.n3067 GNDA.n3066 0.1255
R30608 GNDA.n3073 GNDA.n3072 0.1255
R30609 GNDA.n3079 GNDA.n3078 0.1255
R30610 GNDA.n3007 GNDA.n2996 0.1255
R30611 GNDA.n3024 GNDA.n3023 0.1255
R30612 GNDA.n3037 GNDA.n2990 0.1255
R30613 GNDA.n2931 GNDA.n2183 0.1255
R30614 GNDA.n2948 GNDA.n2947 0.1255
R30615 GNDA.n2961 GNDA.n2177 0.1255
R30616 GNDA.n2833 GNDA.n2832 0.1255
R30617 GNDA.n2839 GNDA.n2838 0.1255
R30618 GNDA.n2845 GNDA.n2844 0.1255
R30619 GNDA.n2773 GNDA.n2762 0.1255
R30620 GNDA.n2790 GNDA.n2789 0.1255
R30621 GNDA.n2803 GNDA.n2756 0.1255
R30622 GNDA.n2701 GNDA.n2698 0.1255
R30623 GNDA.n2714 GNDA.n2672 0.1255
R30624 GNDA.n2731 GNDA.n2728 0.1255
R30625 GNDA.n3057 GNDA.n2156 0.1255
R30626 GNDA.n5409 GNDA.n701 0.1255
R30627 GNDA.n5461 GNDA.n5460 0.1255
R30628 GNDA.n5454 GNDA.n678 0.1255
R30629 GNDA.n645 GNDA.n631 0.1255
R30630 GNDA.n5526 GNDA.n35 0.1255
R30631 GNDA.n598 GNDA.n597 0.1255
R30632 GNDA.n5555 GNDA.n22 0.1255
R30633 GNDA.n5572 GNDA.n5571 0.1255
R30634 GNDA.n5585 GNDA.n16 0.1255
R30635 GNDA.n530 GNDA.n519 0.1255
R30636 GNDA.n547 GNDA.n546 0.1255
R30637 GNDA.n560 GNDA.n513 0.1255
R30638 GNDA.n279 GNDA.n278 0.1255
R30639 GNDA.n285 GNDA.n284 0.1255
R30640 GNDA.n291 GNDA.n290 0.1255
R30641 GNDA.n220 GNDA.n209 0.1255
R30642 GNDA.n237 GNDA.n236 0.1255
R30643 GNDA.n250 GNDA.n203 0.1255
R30644 GNDA.n106 GNDA.n105 0.1255
R30645 GNDA.n112 GNDA.n111 0.1255
R30646 GNDA.n118 GNDA.n117 0.1255
R30647 GNDA.n464 GNDA.n94 0.1255
R30648 GNDA.n481 GNDA.n480 0.1255
R30649 GNDA.n494 GNDA.n88 0.1255
R30650 GNDA.n435 GNDA.n434 0.1255
R30651 GNDA.n424 GNDA.n391 0.1255
R30652 GNDA.n417 GNDA.n416 0.1255
R30653 GNDA.n986 GNDA.n974 0.1255
R30654 GNDA.n1005 GNDA.n1004 0.1255
R30655 GNDA.n1016 GNDA.n968 0.1255
R30656 GNDA.n990 GNDA.n989 0.1255
R30657 GNDA.n1003 GNDA.n971 0.1255
R30658 GNDA.n1020 GNDA.n1019 0.1255
R30659 GNDA.n5470 GNDA.n5469 0.123287
R30660 GNDA.n5482 GNDA.n5481 0.12293
R30661 GNDA.n2196 GNDA.n2192 0.0994583
R30662 GNDA.n5504 GNDA.n649 0.0994583
R30663 GNDA.n4187 GNDA.n4183 0.09425
R30664 GNDA.n3296 GNDA.n3295 0.09425
R30665 GNDA.n3457 GNDA.n3368 0.08275
R30666 GNDA.n2614 GNDA 0.0817953
R30667 GNDA.n2055 GNDA.n2032 0.0734167
R30668 GNDA.n2056 GNDA.n2055 0.0734167
R30669 GNDA.n2057 GNDA.n2056 0.0734167
R30670 GNDA.n2061 GNDA.n2060 0.0734167
R30671 GNDA.n2062 GNDA.n2061 0.0734167
R30672 GNDA.n2063 GNDA.n2062 0.0734167
R30673 GNDA.n2067 GNDA.n2066 0.0734167
R30674 GNDA.n2068 GNDA.n2067 0.0734167
R30675 GNDA.n2069 GNDA.n2068 0.0734167
R30676 GNDA.n2073 GNDA.n2072 0.0734167
R30677 GNDA.n2074 GNDA.n2073 0.0734167
R30678 GNDA.n4143 GNDA.n3661 0.0734167
R30679 GNDA.n4143 GNDA.n4142 0.0734167
R30680 GNDA.n4142 GNDA.n4141 0.0734167
R30681 GNDA.n4136 GNDA.n4135 0.0734167
R30682 GNDA.n4135 GNDA.n3671 0.0734167
R30683 GNDA.n4131 GNDA.n3671 0.0734167
R30684 GNDA.n4125 GNDA.n3676 0.0734167
R30685 GNDA.n4125 GNDA.n4124 0.0734167
R30686 GNDA.n4124 GNDA.n4123 0.0734167
R30687 GNDA.n4118 GNDA.n4117 0.0734167
R30688 GNDA.n4117 GNDA.n3686 0.0734167
R30689 GNDA.n4052 GNDA.n4051 0.0734167
R30690 GNDA.n4053 GNDA.n4052 0.0734167
R30691 GNDA.n4053 GNDA.n4044 0.0734167
R30692 GNDA.n4061 GNDA.n4040 0.0734167
R30693 GNDA.n4067 GNDA.n4040 0.0734167
R30694 GNDA.n4068 GNDA.n4067 0.0734167
R30695 GNDA.n4076 GNDA.n4075 0.0734167
R30696 GNDA.n4077 GNDA.n4076 0.0734167
R30697 GNDA.n4077 GNDA.n4032 0.0734167
R30698 GNDA.n4085 GNDA.n4028 0.0734167
R30699 GNDA.n4091 GNDA.n4028 0.0734167
R30700 GNDA.n3971 GNDA.n3970 0.0734167
R30701 GNDA.n3972 GNDA.n3971 0.0734167
R30702 GNDA.n3972 GNDA.n3963 0.0734167
R30703 GNDA.n3980 GNDA.n3959 0.0734167
R30704 GNDA.n3986 GNDA.n3959 0.0734167
R30705 GNDA.n3987 GNDA.n3986 0.0734167
R30706 GNDA.n3995 GNDA.n3994 0.0734167
R30707 GNDA.n3996 GNDA.n3995 0.0734167
R30708 GNDA.n3996 GNDA.n3951 0.0734167
R30709 GNDA.n4004 GNDA.n3947 0.0734167
R30710 GNDA.n4010 GNDA.n3947 0.0734167
R30711 GNDA.n3890 GNDA.n3889 0.0734167
R30712 GNDA.n3891 GNDA.n3890 0.0734167
R30713 GNDA.n3891 GNDA.n3882 0.0734167
R30714 GNDA.n3899 GNDA.n3878 0.0734167
R30715 GNDA.n3905 GNDA.n3878 0.0734167
R30716 GNDA.n3906 GNDA.n3905 0.0734167
R30717 GNDA.n3914 GNDA.n3913 0.0734167
R30718 GNDA.n3915 GNDA.n3914 0.0734167
R30719 GNDA.n3915 GNDA.n3870 0.0734167
R30720 GNDA.n3923 GNDA.n3866 0.0734167
R30721 GNDA.n3929 GNDA.n3866 0.0734167
R30722 GNDA.n4194 GNDA.n4193 0.0734167
R30723 GNDA.n4195 GNDA.n4194 0.0734167
R30724 GNDA.n4195 GNDA.n3505 0.0734167
R30725 GNDA.n4203 GNDA.n3501 0.0734167
R30726 GNDA.n4209 GNDA.n3501 0.0734167
R30727 GNDA.n4210 GNDA.n4209 0.0734167
R30728 GNDA.n4218 GNDA.n4217 0.0734167
R30729 GNDA.n4219 GNDA.n4218 0.0734167
R30730 GNDA.n4219 GNDA.n3493 0.0734167
R30731 GNDA.n4227 GNDA.n3489 0.0734167
R30732 GNDA.n4233 GNDA.n3489 0.0734167
R30733 GNDA.n3809 GNDA.n3808 0.0734167
R30734 GNDA.n3810 GNDA.n3809 0.0734167
R30735 GNDA.n3810 GNDA.n3801 0.0734167
R30736 GNDA.n3818 GNDA.n3797 0.0734167
R30737 GNDA.n3824 GNDA.n3797 0.0734167
R30738 GNDA.n3825 GNDA.n3824 0.0734167
R30739 GNDA.n3833 GNDA.n3832 0.0734167
R30740 GNDA.n3834 GNDA.n3833 0.0734167
R30741 GNDA.n3834 GNDA.n3789 0.0734167
R30742 GNDA.n3842 GNDA.n3785 0.0734167
R30743 GNDA.n3848 GNDA.n3785 0.0734167
R30744 GNDA.n3728 GNDA.n3727 0.0734167
R30745 GNDA.n3729 GNDA.n3728 0.0734167
R30746 GNDA.n3729 GNDA.n3720 0.0734167
R30747 GNDA.n3737 GNDA.n3716 0.0734167
R30748 GNDA.n3743 GNDA.n3716 0.0734167
R30749 GNDA.n3744 GNDA.n3743 0.0734167
R30750 GNDA.n3752 GNDA.n3751 0.0734167
R30751 GNDA.n3753 GNDA.n3752 0.0734167
R30752 GNDA.n3753 GNDA.n3708 0.0734167
R30753 GNDA.n3761 GNDA.n3704 0.0734167
R30754 GNDA.n3767 GNDA.n3704 0.0734167
R30755 GNDA.n3590 GNDA.n3514 0.0734167
R30756 GNDA.n3590 GNDA.n3589 0.0734167
R30757 GNDA.n3589 GNDA.n3588 0.0734167
R30758 GNDA.n3583 GNDA.n3582 0.0734167
R30759 GNDA.n3582 GNDA.n3528 0.0734167
R30760 GNDA.n3578 GNDA.n3528 0.0734167
R30761 GNDA.n3572 GNDA.n3536 0.0734167
R30762 GNDA.n3572 GNDA.n3571 0.0734167
R30763 GNDA.n3571 GNDA.n3570 0.0734167
R30764 GNDA.n3565 GNDA.n3564 0.0734167
R30765 GNDA.n3564 GNDA.n3552 0.0734167
R30766 GNDA.n4269 GNDA.n1974 0.0734167
R30767 GNDA.n4269 GNDA.n4268 0.0734167
R30768 GNDA.n4268 GNDA.n4267 0.0734167
R30769 GNDA.n4262 GNDA.n4261 0.0734167
R30770 GNDA.n4261 GNDA.n1984 0.0734167
R30771 GNDA.n4257 GNDA.n1984 0.0734167
R30772 GNDA.n4251 GNDA.n1989 0.0734167
R30773 GNDA.n4251 GNDA.n4250 0.0734167
R30774 GNDA.n4250 GNDA.n4249 0.0734167
R30775 GNDA.n4244 GNDA.n4243 0.0734167
R30776 GNDA.n4243 GNDA.n1999 0.0734167
R30777 GNDA.n1068 GNDA.n1067 0.0734167
R30778 GNDA.n1068 GNDA.n1060 0.0734167
R30779 GNDA.n1076 GNDA.n1056 0.0734167
R30780 GNDA.n1082 GNDA.n1056 0.0734167
R30781 GNDA.n1083 GNDA.n1082 0.0734167
R30782 GNDA.n1091 GNDA.n1090 0.0734167
R30783 GNDA.n1092 GNDA.n1091 0.0734167
R30784 GNDA.n1092 GNDA.n1048 0.0734167
R30785 GNDA.n1100 GNDA.n1044 0.0734167
R30786 GNDA.n1106 GNDA.n1044 0.0734167
R30787 GNDA.n1107 GNDA.n1106 0.0734167
R30788 GNDA.n4165 GNDA.n4164 0.0734167
R30789 GNDA.n3405 GNDA.n3404 0.0734167
R30790 GNDA.n3406 GNDA.n3405 0.0734167
R30791 GNDA.n3406 GNDA.n3391 0.0734167
R30792 GNDA.n3416 GNDA.n3389 0.0734167
R30793 GNDA.n3424 GNDA.n3389 0.0734167
R30794 GNDA.n3425 GNDA.n3424 0.0734167
R30795 GNDA.n3435 GNDA.n3434 0.0734167
R30796 GNDA.n3436 GNDA.n3435 0.0734167
R30797 GNDA.n3436 GNDA.n3385 0.0734167
R30798 GNDA.n3446 GNDA.n3383 0.0734167
R30799 GNDA.n3454 GNDA.n3383 0.0734167
R30800 GNDA.n3316 GNDA.n3315 0.0734167
R30801 GNDA.n3317 GNDA.n3316 0.0734167
R30802 GNDA.n3317 GNDA.n2026 0.0734167
R30803 GNDA.n3327 GNDA.n2024 0.0734167
R30804 GNDA.n3335 GNDA.n2024 0.0734167
R30805 GNDA.n3336 GNDA.n3335 0.0734167
R30806 GNDA.n3346 GNDA.n3345 0.0734167
R30807 GNDA.n3347 GNDA.n3346 0.0734167
R30808 GNDA.n3347 GNDA.n2020 0.0734167
R30809 GNDA.n3357 GNDA.n2018 0.0734167
R30810 GNDA.n3365 GNDA.n2018 0.0734167
R30811 GNDA.n3233 GNDA.n2119 0.0734167
R30812 GNDA.n3234 GNDA.n3233 0.0734167
R30813 GNDA.n3234 GNDA.n3231 0.0734167
R30814 GNDA.n3244 GNDA.n3229 0.0734167
R30815 GNDA.n3252 GNDA.n3229 0.0734167
R30816 GNDA.n3253 GNDA.n3252 0.0734167
R30817 GNDA.n3263 GNDA.n3262 0.0734167
R30818 GNDA.n3264 GNDA.n3263 0.0734167
R30819 GNDA.n3264 GNDA.n3225 0.0734167
R30820 GNDA.n3274 GNDA.n3223 0.0734167
R30821 GNDA.n3282 GNDA.n3223 0.0734167
R30822 GNDA.n3157 GNDA.n3156 0.0734167
R30823 GNDA.n3158 GNDA.n3157 0.0734167
R30824 GNDA.n3158 GNDA.n2145 0.0734167
R30825 GNDA.n3168 GNDA.n2143 0.0734167
R30826 GNDA.n3176 GNDA.n2143 0.0734167
R30827 GNDA.n3177 GNDA.n3176 0.0734167
R30828 GNDA.n3187 GNDA.n3186 0.0734167
R30829 GNDA.n3188 GNDA.n3187 0.0734167
R30830 GNDA.n3188 GNDA.n2139 0.0734167
R30831 GNDA.n3198 GNDA.n2137 0.0734167
R30832 GNDA.n3206 GNDA.n2137 0.0734167
R30833 GNDA.n3084 GNDA.n3061 0.0734167
R30834 GNDA.n3085 GNDA.n3084 0.0734167
R30835 GNDA.n3086 GNDA.n3085 0.0734167
R30836 GNDA.n3090 GNDA.n3089 0.0734167
R30837 GNDA.n3091 GNDA.n3090 0.0734167
R30838 GNDA.n3092 GNDA.n3091 0.0734167
R30839 GNDA.n3096 GNDA.n3095 0.0734167
R30840 GNDA.n3097 GNDA.n3096 0.0734167
R30841 GNDA.n3098 GNDA.n3097 0.0734167
R30842 GNDA.n3102 GNDA.n3101 0.0734167
R30843 GNDA.n3103 GNDA.n3102 0.0734167
R30844 GNDA.n2999 GNDA.n2158 0.0734167
R30845 GNDA.n3000 GNDA.n2999 0.0734167
R30846 GNDA.n3000 GNDA.n2997 0.0734167
R30847 GNDA.n3010 GNDA.n2995 0.0734167
R30848 GNDA.n3018 GNDA.n2995 0.0734167
R30849 GNDA.n3019 GNDA.n3018 0.0734167
R30850 GNDA.n3029 GNDA.n3028 0.0734167
R30851 GNDA.n3030 GNDA.n3029 0.0734167
R30852 GNDA.n3030 GNDA.n2991 0.0734167
R30853 GNDA.n3040 GNDA.n2989 0.0734167
R30854 GNDA.n3048 GNDA.n2989 0.0734167
R30855 GNDA.n2923 GNDA.n2922 0.0734167
R30856 GNDA.n2924 GNDA.n2923 0.0734167
R30857 GNDA.n2924 GNDA.n2184 0.0734167
R30858 GNDA.n2934 GNDA.n2182 0.0734167
R30859 GNDA.n2942 GNDA.n2182 0.0734167
R30860 GNDA.n2943 GNDA.n2942 0.0734167
R30861 GNDA.n2953 GNDA.n2952 0.0734167
R30862 GNDA.n2954 GNDA.n2953 0.0734167
R30863 GNDA.n2954 GNDA.n2178 0.0734167
R30864 GNDA.n2964 GNDA.n2176 0.0734167
R30865 GNDA.n2972 GNDA.n2176 0.0734167
R30866 GNDA.n2850 GNDA.n2827 0.0734167
R30867 GNDA.n2851 GNDA.n2850 0.0734167
R30868 GNDA.n2852 GNDA.n2851 0.0734167
R30869 GNDA.n2856 GNDA.n2855 0.0734167
R30870 GNDA.n2857 GNDA.n2856 0.0734167
R30871 GNDA.n2858 GNDA.n2857 0.0734167
R30872 GNDA.n2862 GNDA.n2861 0.0734167
R30873 GNDA.n2863 GNDA.n2862 0.0734167
R30874 GNDA.n2864 GNDA.n2863 0.0734167
R30875 GNDA.n2868 GNDA.n2867 0.0734167
R30876 GNDA.n2869 GNDA.n2868 0.0734167
R30877 GNDA.n2765 GNDA.n2242 0.0734167
R30878 GNDA.n2766 GNDA.n2765 0.0734167
R30879 GNDA.n2766 GNDA.n2763 0.0734167
R30880 GNDA.n2776 GNDA.n2761 0.0734167
R30881 GNDA.n2784 GNDA.n2761 0.0734167
R30882 GNDA.n2785 GNDA.n2784 0.0734167
R30883 GNDA.n2795 GNDA.n2794 0.0734167
R30884 GNDA.n2796 GNDA.n2795 0.0734167
R30885 GNDA.n2796 GNDA.n2757 0.0734167
R30886 GNDA.n2806 GNDA.n2755 0.0734167
R30887 GNDA.n2814 GNDA.n2755 0.0734167
R30888 GNDA.n2687 GNDA.n2677 0.0734167
R30889 GNDA.n2695 GNDA.n2677 0.0734167
R30890 GNDA.n2696 GNDA.n2695 0.0734167
R30891 GNDA.n2706 GNDA.n2705 0.0734167
R30892 GNDA.n2707 GNDA.n2706 0.0734167
R30893 GNDA.n2707 GNDA.n2673 0.0734167
R30894 GNDA.n2717 GNDA.n2671 0.0734167
R30895 GNDA.n2725 GNDA.n2671 0.0734167
R30896 GNDA.n2726 GNDA.n2725 0.0734167
R30897 GNDA.n2735 GNDA.n2734 0.0734167
R30898 GNDA.n2737 GNDA.n2735 0.0734167
R30899 GNDA.n2231 GNDA.n2230 0.0734167
R30900 GNDA.n5547 GNDA.n5546 0.0734167
R30901 GNDA.n5548 GNDA.n5547 0.0734167
R30902 GNDA.n5548 GNDA.n23 0.0734167
R30903 GNDA.n5558 GNDA.n21 0.0734167
R30904 GNDA.n5566 GNDA.n21 0.0734167
R30905 GNDA.n5567 GNDA.n5566 0.0734167
R30906 GNDA.n5577 GNDA.n5576 0.0734167
R30907 GNDA.n5578 GNDA.n5577 0.0734167
R30908 GNDA.n5578 GNDA.n17 0.0734167
R30909 GNDA.n5588 GNDA.n15 0.0734167
R30910 GNDA.n5596 GNDA.n15 0.0734167
R30911 GNDA.n522 GNDA.n46 0.0734167
R30912 GNDA.n523 GNDA.n522 0.0734167
R30913 GNDA.n523 GNDA.n520 0.0734167
R30914 GNDA.n533 GNDA.n518 0.0734167
R30915 GNDA.n541 GNDA.n518 0.0734167
R30916 GNDA.n542 GNDA.n541 0.0734167
R30917 GNDA.n552 GNDA.n551 0.0734167
R30918 GNDA.n553 GNDA.n552 0.0734167
R30919 GNDA.n553 GNDA.n514 0.0734167
R30920 GNDA.n563 GNDA.n512 0.0734167
R30921 GNDA.n571 GNDA.n512 0.0734167
R30922 GNDA.n296 GNDA.n273 0.0734167
R30923 GNDA.n297 GNDA.n296 0.0734167
R30924 GNDA.n298 GNDA.n297 0.0734167
R30925 GNDA.n302 GNDA.n301 0.0734167
R30926 GNDA.n303 GNDA.n302 0.0734167
R30927 GNDA.n304 GNDA.n303 0.0734167
R30928 GNDA.n308 GNDA.n307 0.0734167
R30929 GNDA.n309 GNDA.n308 0.0734167
R30930 GNDA.n310 GNDA.n309 0.0734167
R30931 GNDA.n314 GNDA.n313 0.0734167
R30932 GNDA.n315 GNDA.n314 0.0734167
R30933 GNDA.n212 GNDA.n186 0.0734167
R30934 GNDA.n213 GNDA.n212 0.0734167
R30935 GNDA.n213 GNDA.n210 0.0734167
R30936 GNDA.n223 GNDA.n208 0.0734167
R30937 GNDA.n231 GNDA.n208 0.0734167
R30938 GNDA.n232 GNDA.n231 0.0734167
R30939 GNDA.n242 GNDA.n241 0.0734167
R30940 GNDA.n243 GNDA.n242 0.0734167
R30941 GNDA.n243 GNDA.n204 0.0734167
R30942 GNDA.n253 GNDA.n202 0.0734167
R30943 GNDA.n261 GNDA.n202 0.0734167
R30944 GNDA.n123 GNDA.n100 0.0734167
R30945 GNDA.n124 GNDA.n123 0.0734167
R30946 GNDA.n125 GNDA.n124 0.0734167
R30947 GNDA.n129 GNDA.n128 0.0734167
R30948 GNDA.n130 GNDA.n129 0.0734167
R30949 GNDA.n131 GNDA.n130 0.0734167
R30950 GNDA.n135 GNDA.n134 0.0734167
R30951 GNDA.n136 GNDA.n135 0.0734167
R30952 GNDA.n137 GNDA.n136 0.0734167
R30953 GNDA.n141 GNDA.n140 0.0734167
R30954 GNDA.n142 GNDA.n141 0.0734167
R30955 GNDA.n456 GNDA.n455 0.0734167
R30956 GNDA.n457 GNDA.n456 0.0734167
R30957 GNDA.n457 GNDA.n95 0.0734167
R30958 GNDA.n467 GNDA.n93 0.0734167
R30959 GNDA.n475 GNDA.n93 0.0734167
R30960 GNDA.n476 GNDA.n475 0.0734167
R30961 GNDA.n486 GNDA.n485 0.0734167
R30962 GNDA.n487 GNDA.n486 0.0734167
R30963 GNDA.n487 GNDA.n89 0.0734167
R30964 GNDA.n497 GNDA.n87 0.0734167
R30965 GNDA.n505 GNDA.n87 0.0734167
R30966 GNDA.n439 GNDA.n376 0.0734167
R30967 GNDA.n439 GNDA.n438 0.0734167
R30968 GNDA.n438 GNDA.n437 0.0734167
R30969 GNDA.n432 GNDA.n431 0.0734167
R30970 GNDA.n431 GNDA.n386 0.0734167
R30971 GNDA.n427 GNDA.n386 0.0734167
R30972 GNDA.n421 GNDA.n392 0.0734167
R30973 GNDA.n421 GNDA.n420 0.0734167
R30974 GNDA.n420 GNDA.n419 0.0734167
R30975 GNDA.n414 GNDA.n413 0.0734167
R30976 GNDA.n413 GNDA.n404 0.0734167
R30977 GNDA.n2112 GNDA.n2032 0.0682083
R30978 GNDA.n2058 GNDA.n2057 0.0682083
R30979 GNDA.n2060 GNDA.n2059 0.0682083
R30980 GNDA.n2064 GNDA.n2063 0.0682083
R30981 GNDA.n2066 GNDA.n2065 0.0682083
R30982 GNDA.n2070 GNDA.n2069 0.0682083
R30983 GNDA.n2072 GNDA.n2071 0.0682083
R30984 GNDA.n4147 GNDA.n3661 0.0682083
R30985 GNDA.n4141 GNDA.n3666 0.0682083
R30986 GNDA.n4137 GNDA.n4136 0.0682083
R30987 GNDA.n4131 GNDA.n4130 0.0682083
R30988 GNDA.n4129 GNDA.n3676 0.0682083
R30989 GNDA.n4123 GNDA.n3681 0.0682083
R30990 GNDA.n4119 GNDA.n4118 0.0682083
R30991 GNDA.n4051 GNDA.n3656 0.0682083
R30992 GNDA.n4059 GNDA.n4044 0.0682083
R30993 GNDA.n4061 GNDA.n4060 0.0682083
R30994 GNDA.n4069 GNDA.n4068 0.0682083
R30995 GNDA.n4075 GNDA.n4036 0.0682083
R30996 GNDA.n4083 GNDA.n4032 0.0682083
R30997 GNDA.n4085 GNDA.n4084 0.0682083
R30998 GNDA.n3970 GNDA.n3651 0.0682083
R30999 GNDA.n3978 GNDA.n3963 0.0682083
R31000 GNDA.n3980 GNDA.n3979 0.0682083
R31001 GNDA.n3988 GNDA.n3987 0.0682083
R31002 GNDA.n3994 GNDA.n3955 0.0682083
R31003 GNDA.n4002 GNDA.n3951 0.0682083
R31004 GNDA.n4004 GNDA.n4003 0.0682083
R31005 GNDA.n3889 GNDA.n3646 0.0682083
R31006 GNDA.n3897 GNDA.n3882 0.0682083
R31007 GNDA.n3899 GNDA.n3898 0.0682083
R31008 GNDA.n3907 GNDA.n3906 0.0682083
R31009 GNDA.n3913 GNDA.n3874 0.0682083
R31010 GNDA.n3921 GNDA.n3870 0.0682083
R31011 GNDA.n3923 GNDA.n3922 0.0682083
R31012 GNDA.n4193 GNDA.n4189 0.0682083
R31013 GNDA.n4201 GNDA.n3505 0.0682083
R31014 GNDA.n4203 GNDA.n4202 0.0682083
R31015 GNDA.n4211 GNDA.n4210 0.0682083
R31016 GNDA.n4217 GNDA.n3497 0.0682083
R31017 GNDA.n4225 GNDA.n3493 0.0682083
R31018 GNDA.n4227 GNDA.n4226 0.0682083
R31019 GNDA.n3808 GNDA.n3604 0.0682083
R31020 GNDA.n3816 GNDA.n3801 0.0682083
R31021 GNDA.n3818 GNDA.n3817 0.0682083
R31022 GNDA.n3826 GNDA.n3825 0.0682083
R31023 GNDA.n3832 GNDA.n3793 0.0682083
R31024 GNDA.n3840 GNDA.n3789 0.0682083
R31025 GNDA.n3842 GNDA.n3841 0.0682083
R31026 GNDA.n3727 GNDA.n3599 0.0682083
R31027 GNDA.n3735 GNDA.n3720 0.0682083
R31028 GNDA.n3737 GNDA.n3736 0.0682083
R31029 GNDA.n3745 GNDA.n3744 0.0682083
R31030 GNDA.n3751 GNDA.n3712 0.0682083
R31031 GNDA.n3759 GNDA.n3708 0.0682083
R31032 GNDA.n3761 GNDA.n3760 0.0682083
R31033 GNDA.n3594 GNDA.n3514 0.0682083
R31034 GNDA.n3588 GNDA.n3520 0.0682083
R31035 GNDA.n3584 GNDA.n3583 0.0682083
R31036 GNDA.n3578 GNDA.n3577 0.0682083
R31037 GNDA.n3576 GNDA.n3536 0.0682083
R31038 GNDA.n3570 GNDA.n3544 0.0682083
R31039 GNDA.n3566 GNDA.n3565 0.0682083
R31040 GNDA.n4273 GNDA.n1974 0.0682083
R31041 GNDA.n4267 GNDA.n1979 0.0682083
R31042 GNDA.n4263 GNDA.n4262 0.0682083
R31043 GNDA.n4257 GNDA.n4256 0.0682083
R31044 GNDA.n4255 GNDA.n1989 0.0682083
R31045 GNDA.n4249 GNDA.n1994 0.0682083
R31046 GNDA.n4245 GNDA.n4244 0.0682083
R31047 GNDA.n1074 GNDA.n1060 0.0682083
R31048 GNDA.n1076 GNDA.n1075 0.0682083
R31049 GNDA.n1084 GNDA.n1083 0.0682083
R31050 GNDA.n1090 GNDA.n1052 0.0682083
R31051 GNDA.n1098 GNDA.n1048 0.0682083
R31052 GNDA.n1100 GNDA.n1099 0.0682083
R31053 GNDA.n4893 GNDA.n1107 0.0682083
R31054 GNDA.n3404 GNDA.n3400 0.0682083
R31055 GNDA.n3414 GNDA.n3391 0.0682083
R31056 GNDA.n3416 GNDA.n3415 0.0682083
R31057 GNDA.n3426 GNDA.n3425 0.0682083
R31058 GNDA.n3434 GNDA.n3387 0.0682083
R31059 GNDA.n3444 GNDA.n3385 0.0682083
R31060 GNDA.n3446 GNDA.n3445 0.0682083
R31061 GNDA.n3315 GNDA.n3311 0.0682083
R31062 GNDA.n3325 GNDA.n2026 0.0682083
R31063 GNDA.n3327 GNDA.n3326 0.0682083
R31064 GNDA.n3337 GNDA.n3336 0.0682083
R31065 GNDA.n3345 GNDA.n2022 0.0682083
R31066 GNDA.n3355 GNDA.n2020 0.0682083
R31067 GNDA.n3357 GNDA.n3356 0.0682083
R31068 GNDA.n3288 GNDA.n2119 0.0682083
R31069 GNDA.n3242 GNDA.n3231 0.0682083
R31070 GNDA.n3244 GNDA.n3243 0.0682083
R31071 GNDA.n3254 GNDA.n3253 0.0682083
R31072 GNDA.n3262 GNDA.n3227 0.0682083
R31073 GNDA.n3272 GNDA.n3225 0.0682083
R31074 GNDA.n3274 GNDA.n3273 0.0682083
R31075 GNDA.n3156 GNDA.n3152 0.0682083
R31076 GNDA.n3166 GNDA.n2145 0.0682083
R31077 GNDA.n3168 GNDA.n3167 0.0682083
R31078 GNDA.n3178 GNDA.n3177 0.0682083
R31079 GNDA.n3186 GNDA.n2141 0.0682083
R31080 GNDA.n3196 GNDA.n2139 0.0682083
R31081 GNDA.n3198 GNDA.n3197 0.0682083
R31082 GNDA.n3141 GNDA.n3061 0.0682083
R31083 GNDA.n3087 GNDA.n3086 0.0682083
R31084 GNDA.n3089 GNDA.n3088 0.0682083
R31085 GNDA.n3093 GNDA.n3092 0.0682083
R31086 GNDA.n3095 GNDA.n3094 0.0682083
R31087 GNDA.n3099 GNDA.n3098 0.0682083
R31088 GNDA.n3101 GNDA.n3100 0.0682083
R31089 GNDA.n3054 GNDA.n2158 0.0682083
R31090 GNDA.n3008 GNDA.n2997 0.0682083
R31091 GNDA.n3010 GNDA.n3009 0.0682083
R31092 GNDA.n3020 GNDA.n3019 0.0682083
R31093 GNDA.n3028 GNDA.n2993 0.0682083
R31094 GNDA.n3038 GNDA.n2991 0.0682083
R31095 GNDA.n3040 GNDA.n3039 0.0682083
R31096 GNDA.n2922 GNDA.n2918 0.0682083
R31097 GNDA.n2932 GNDA.n2184 0.0682083
R31098 GNDA.n2934 GNDA.n2933 0.0682083
R31099 GNDA.n2944 GNDA.n2943 0.0682083
R31100 GNDA.n2952 GNDA.n2180 0.0682083
R31101 GNDA.n2962 GNDA.n2178 0.0682083
R31102 GNDA.n2964 GNDA.n2963 0.0682083
R31103 GNDA.n2907 GNDA.n2827 0.0682083
R31104 GNDA.n2853 GNDA.n2852 0.0682083
R31105 GNDA.n2855 GNDA.n2854 0.0682083
R31106 GNDA.n2859 GNDA.n2858 0.0682083
R31107 GNDA.n2861 GNDA.n2860 0.0682083
R31108 GNDA.n2865 GNDA.n2864 0.0682083
R31109 GNDA.n2867 GNDA.n2866 0.0682083
R31110 GNDA.n2820 GNDA.n2242 0.0682083
R31111 GNDA.n2774 GNDA.n2763 0.0682083
R31112 GNDA.n2776 GNDA.n2775 0.0682083
R31113 GNDA.n2786 GNDA.n2785 0.0682083
R31114 GNDA.n2794 GNDA.n2759 0.0682083
R31115 GNDA.n2804 GNDA.n2757 0.0682083
R31116 GNDA.n2806 GNDA.n2805 0.0682083
R31117 GNDA.n2687 GNDA.n2686 0.0682083
R31118 GNDA.n2697 GNDA.n2696 0.0682083
R31119 GNDA.n2705 GNDA.n2675 0.0682083
R31120 GNDA.n2715 GNDA.n2673 0.0682083
R31121 GNDA.n2717 GNDA.n2716 0.0682083
R31122 GNDA.n2727 GNDA.n2726 0.0682083
R31123 GNDA.n2734 GNDA.n2669 0.0682083
R31124 GNDA.n5546 GNDA.n5542 0.0682083
R31125 GNDA.n5556 GNDA.n23 0.0682083
R31126 GNDA.n5558 GNDA.n5557 0.0682083
R31127 GNDA.n5568 GNDA.n5567 0.0682083
R31128 GNDA.n5576 GNDA.n19 0.0682083
R31129 GNDA.n5586 GNDA.n17 0.0682083
R31130 GNDA.n5588 GNDA.n5587 0.0682083
R31131 GNDA.n577 GNDA.n46 0.0682083
R31132 GNDA.n531 GNDA.n520 0.0682083
R31133 GNDA.n533 GNDA.n532 0.0682083
R31134 GNDA.n543 GNDA.n542 0.0682083
R31135 GNDA.n551 GNDA.n516 0.0682083
R31136 GNDA.n561 GNDA.n514 0.0682083
R31137 GNDA.n563 GNDA.n562 0.0682083
R31138 GNDA.n353 GNDA.n273 0.0682083
R31139 GNDA.n299 GNDA.n298 0.0682083
R31140 GNDA.n301 GNDA.n300 0.0682083
R31141 GNDA.n305 GNDA.n304 0.0682083
R31142 GNDA.n307 GNDA.n306 0.0682083
R31143 GNDA.n311 GNDA.n310 0.0682083
R31144 GNDA.n313 GNDA.n312 0.0682083
R31145 GNDA.n267 GNDA.n186 0.0682083
R31146 GNDA.n221 GNDA.n210 0.0682083
R31147 GNDA.n223 GNDA.n222 0.0682083
R31148 GNDA.n233 GNDA.n232 0.0682083
R31149 GNDA.n241 GNDA.n206 0.0682083
R31150 GNDA.n251 GNDA.n204 0.0682083
R31151 GNDA.n253 GNDA.n252 0.0682083
R31152 GNDA.n180 GNDA.n100 0.0682083
R31153 GNDA.n126 GNDA.n125 0.0682083
R31154 GNDA.n128 GNDA.n127 0.0682083
R31155 GNDA.n132 GNDA.n131 0.0682083
R31156 GNDA.n134 GNDA.n133 0.0682083
R31157 GNDA.n138 GNDA.n137 0.0682083
R31158 GNDA.n140 GNDA.n139 0.0682083
R31159 GNDA.n455 GNDA.n451 0.0682083
R31160 GNDA.n465 GNDA.n95 0.0682083
R31161 GNDA.n467 GNDA.n466 0.0682083
R31162 GNDA.n477 GNDA.n476 0.0682083
R31163 GNDA.n485 GNDA.n91 0.0682083
R31164 GNDA.n495 GNDA.n89 0.0682083
R31165 GNDA.n497 GNDA.n496 0.0682083
R31166 GNDA.n443 GNDA.n376 0.0682083
R31167 GNDA.n437 GNDA.n380 0.0682083
R31168 GNDA.n433 GNDA.n432 0.0682083
R31169 GNDA.n427 GNDA.n426 0.0682083
R31170 GNDA.n425 GNDA.n392 0.0682083
R31171 GNDA.n419 GNDA.n398 0.0682083
R31172 GNDA.n415 GNDA.n414 0.0682083
R31173 GNDA.n1066 GNDA.n1065 0.0672139
R31174 GNDA.n2075 GNDA.n2054 0.0672139
R31175 GNDA.n4114 GNDA.n4113 0.0672139
R31176 GNDA.n4092 GNDA.n4027 0.0672139
R31177 GNDA.n4011 GNDA.n3946 0.0672139
R31178 GNDA.n3930 GNDA.n3865 0.0672139
R31179 GNDA.n4234 GNDA.n3488 0.0672139
R31180 GNDA.n3849 GNDA.n3784 0.0672139
R31181 GNDA.n3768 GNDA.n3703 0.0672139
R31182 GNDA.n3561 GNDA.n3560 0.0672139
R31183 GNDA.n4240 GNDA.n4239 0.0672139
R31184 GNDA.n3455 GNDA.n3382 0.0672139
R31185 GNDA.n3366 GNDA.n2017 0.0672139
R31186 GNDA.n3283 GNDA.n3222 0.0672139
R31187 GNDA.n3207 GNDA.n2136 0.0672139
R31188 GNDA.n3104 GNDA.n3083 0.0672139
R31189 GNDA.n3049 GNDA.n2988 0.0672139
R31190 GNDA.n2973 GNDA.n2175 0.0672139
R31191 GNDA.n2870 GNDA.n2849 0.0672139
R31192 GNDA.n2815 GNDA.n2754 0.0672139
R31193 GNDA.n2736 GNDA.n2668 0.0672139
R31194 GNDA.n5597 GNDA.n14 0.0672139
R31195 GNDA.n572 GNDA.n511 0.0672139
R31196 GNDA.n316 GNDA.n295 0.0672139
R31197 GNDA.n262 GNDA.n201 0.0672139
R31198 GNDA.n143 GNDA.n122 0.0672139
R31199 GNDA.n506 GNDA.n86 0.0672139
R31200 GNDA.n410 GNDA.n409 0.0672139
R31201 GNDA.n979 GNDA.n977 0.0667303
R31202 GNDA.n2059 GNDA.n2058 0.063
R31203 GNDA.n2065 GNDA.n2064 0.063
R31204 GNDA.n2071 GNDA.n2070 0.063
R31205 GNDA.n4137 GNDA.n3666 0.063
R31206 GNDA.n4130 GNDA.n4129 0.063
R31207 GNDA.n4119 GNDA.n3681 0.063
R31208 GNDA.n4060 GNDA.n4059 0.063
R31209 GNDA.n4069 GNDA.n4036 0.063
R31210 GNDA.n4084 GNDA.n4083 0.063
R31211 GNDA.n3979 GNDA.n3978 0.063
R31212 GNDA.n3988 GNDA.n3955 0.063
R31213 GNDA.n4003 GNDA.n4002 0.063
R31214 GNDA.n3898 GNDA.n3897 0.063
R31215 GNDA.n3907 GNDA.n3874 0.063
R31216 GNDA.n3922 GNDA.n3921 0.063
R31217 GNDA.n4202 GNDA.n4201 0.063
R31218 GNDA.n4211 GNDA.n3497 0.063
R31219 GNDA.n4226 GNDA.n4225 0.063
R31220 GNDA.n3817 GNDA.n3816 0.063
R31221 GNDA.n3826 GNDA.n3793 0.063
R31222 GNDA.n3841 GNDA.n3840 0.063
R31223 GNDA.n3736 GNDA.n3735 0.063
R31224 GNDA.n3745 GNDA.n3712 0.063
R31225 GNDA.n3760 GNDA.n3759 0.063
R31226 GNDA.n3584 GNDA.n3520 0.063
R31227 GNDA.n3577 GNDA.n3576 0.063
R31228 GNDA.n3566 GNDA.n3544 0.063
R31229 GNDA.n4263 GNDA.n1979 0.063
R31230 GNDA.n4256 GNDA.n4255 0.063
R31231 GNDA.n4245 GNDA.n1994 0.063
R31232 GNDA.n1075 GNDA.n1074 0.063
R31233 GNDA.n1084 GNDA.n1052 0.063
R31234 GNDA.n1099 GNDA.n1098 0.063
R31235 GNDA.n3415 GNDA.n3414 0.063
R31236 GNDA.n3426 GNDA.n3387 0.063
R31237 GNDA.n3445 GNDA.n3444 0.063
R31238 GNDA.n3326 GNDA.n3325 0.063
R31239 GNDA.n3337 GNDA.n2022 0.063
R31240 GNDA.n3356 GNDA.n3355 0.063
R31241 GNDA.n3243 GNDA.n3242 0.063
R31242 GNDA.n3254 GNDA.n3227 0.063
R31243 GNDA.n3273 GNDA.n3272 0.063
R31244 GNDA.n3167 GNDA.n3166 0.063
R31245 GNDA.n3178 GNDA.n2141 0.063
R31246 GNDA.n3197 GNDA.n3196 0.063
R31247 GNDA.n3088 GNDA.n3087 0.063
R31248 GNDA.n3094 GNDA.n3093 0.063
R31249 GNDA.n3100 GNDA.n3099 0.063
R31250 GNDA.n3009 GNDA.n3008 0.063
R31251 GNDA.n3020 GNDA.n2993 0.063
R31252 GNDA.n3039 GNDA.n3038 0.063
R31253 GNDA.n2933 GNDA.n2932 0.063
R31254 GNDA.n2944 GNDA.n2180 0.063
R31255 GNDA.n2963 GNDA.n2962 0.063
R31256 GNDA.n2854 GNDA.n2853 0.063
R31257 GNDA.n2860 GNDA.n2859 0.063
R31258 GNDA.n2866 GNDA.n2865 0.063
R31259 GNDA.n2775 GNDA.n2774 0.063
R31260 GNDA.n2786 GNDA.n2759 0.063
R31261 GNDA.n2805 GNDA.n2804 0.063
R31262 GNDA.n2697 GNDA.n2675 0.063
R31263 GNDA.n2716 GNDA.n2715 0.063
R31264 GNDA.n2727 GNDA.n2669 0.063
R31265 GNDA.n599 GNDA.n588 0.063
R31266 GNDA.n5527 GNDA.n33 0.063
R31267 GNDA.n5557 GNDA.n5556 0.063
R31268 GNDA.n5568 GNDA.n19 0.063
R31269 GNDA.n5587 GNDA.n5586 0.063
R31270 GNDA.n532 GNDA.n531 0.063
R31271 GNDA.n543 GNDA.n516 0.063
R31272 GNDA.n562 GNDA.n561 0.063
R31273 GNDA.n300 GNDA.n299 0.063
R31274 GNDA.n306 GNDA.n305 0.063
R31275 GNDA.n312 GNDA.n311 0.063
R31276 GNDA.n222 GNDA.n221 0.063
R31277 GNDA.n233 GNDA.n206 0.063
R31278 GNDA.n252 GNDA.n251 0.063
R31279 GNDA.n127 GNDA.n126 0.063
R31280 GNDA.n133 GNDA.n132 0.063
R31281 GNDA.n139 GNDA.n138 0.063
R31282 GNDA.n466 GNDA.n465 0.063
R31283 GNDA.n477 GNDA.n91 0.063
R31284 GNDA.n496 GNDA.n495 0.063
R31285 GNDA.n433 GNDA.n380 0.063
R31286 GNDA.n426 GNDA.n425 0.063
R31287 GNDA.n415 GNDA.n398 0.063
R31288 GNDA.n5021 GNDA.n4924 0.063
R31289 GNDA.n5344 GNDA.n5343 0.063
R31290 GNDA.n5068 GNDA.n5067 0.0626438
R31291 GNDA.n5055 GNDA.n5054 0.0626438
R31292 GNDA.n1110 GNDA.n1109 0.0626438
R31293 GNDA.n701 GNDA.n700 0.0626438
R31294 GNDA.n5460 GNDA.n5459 0.0626438
R31295 GNDA.n5452 GNDA.n678 0.0626438
R31296 GNDA.n5507 GNDA.n631 0.0626438
R31297 GNDA.n35 GNDA.n34 0.0626438
R31298 GNDA.n597 GNDA.n589 0.0626438
R31299 GNDA.n588 GNDA.n587 0.0577917
R31300 GNDA.n585 GNDA.n33 0.0577917
R31301 GNDA.n2107 GNDA.n2106 0.0553333
R31302 GNDA.n2098 GNDA.n2097 0.0553333
R31303 GNDA.n2089 GNDA.n2088 0.0553333
R31304 GNDA.n2080 GNDA.n2079 0.0553333
R31305 GNDA.n4096 GNDA.n3664 0.0553333
R31306 GNDA.n3673 GNDA.n3672 0.0553333
R31307 GNDA.n4105 GNDA.n3679 0.0553333
R31308 GNDA.n3688 GNDA.n3687 0.0553333
R31309 GNDA.n4047 GNDA.n4046 0.0553333
R31310 GNDA.n4065 GNDA.n4064 0.0553333
R31311 GNDA.n4035 GNDA.n4034 0.0553333
R31312 GNDA.n4089 GNDA.n4088 0.0553333
R31313 GNDA.n3966 GNDA.n3965 0.0553333
R31314 GNDA.n3984 GNDA.n3983 0.0553333
R31315 GNDA.n3954 GNDA.n3953 0.0553333
R31316 GNDA.n4008 GNDA.n4007 0.0553333
R31317 GNDA.n3885 GNDA.n3884 0.0553333
R31318 GNDA.n3903 GNDA.n3902 0.0553333
R31319 GNDA.n3873 GNDA.n3872 0.0553333
R31320 GNDA.n3927 GNDA.n3926 0.0553333
R31321 GNDA.n3508 GNDA.n3507 0.0553333
R31322 GNDA.n4207 GNDA.n4206 0.0553333
R31323 GNDA.n3496 GNDA.n3495 0.0553333
R31324 GNDA.n4231 GNDA.n4230 0.0553333
R31325 GNDA.n3804 GNDA.n3803 0.0553333
R31326 GNDA.n3822 GNDA.n3821 0.0553333
R31327 GNDA.n3792 GNDA.n3791 0.0553333
R31328 GNDA.n3846 GNDA.n3845 0.0553333
R31329 GNDA.n3723 GNDA.n3722 0.0553333
R31330 GNDA.n3741 GNDA.n3740 0.0553333
R31331 GNDA.n3711 GNDA.n3710 0.0553333
R31332 GNDA.n3765 GNDA.n3764 0.0553333
R31333 GNDA.n3521 GNDA.n3518 0.0553333
R31334 GNDA.n3532 GNDA.n3531 0.0553333
R31335 GNDA.n3545 GNDA.n3542 0.0553333
R31336 GNDA.n3556 GNDA.n3555 0.0553333
R31337 GNDA.n3459 GNDA.n1977 0.0553333
R31338 GNDA.n1986 GNDA.n1985 0.0553333
R31339 GNDA.n3468 GNDA.n1992 0.0553333
R31340 GNDA.n2001 GNDA.n2000 0.0553333
R31341 GNDA.n1063 GNDA.n1062 0.0553333
R31342 GNDA.n1080 GNDA.n1079 0.0553333
R31343 GNDA.n1051 GNDA.n1050 0.0553333
R31344 GNDA.n1104 GNDA.n1103 0.0553333
R31345 GNDA.n3408 GNDA.n3407 0.0553333
R31346 GNDA.n3422 GNDA.n3421 0.0553333
R31347 GNDA.n3438 GNDA.n3437 0.0553333
R31348 GNDA.n3452 GNDA.n3451 0.0553333
R31349 GNDA.n3319 GNDA.n3318 0.0553333
R31350 GNDA.n3333 GNDA.n3332 0.0553333
R31351 GNDA.n3349 GNDA.n3348 0.0553333
R31352 GNDA.n3363 GNDA.n3362 0.0553333
R31353 GNDA.n3236 GNDA.n3235 0.0553333
R31354 GNDA.n3250 GNDA.n3249 0.0553333
R31355 GNDA.n3266 GNDA.n3265 0.0553333
R31356 GNDA.n3280 GNDA.n3279 0.0553333
R31357 GNDA.n3160 GNDA.n3159 0.0553333
R31358 GNDA.n3174 GNDA.n3173 0.0553333
R31359 GNDA.n3190 GNDA.n3189 0.0553333
R31360 GNDA.n3204 GNDA.n3203 0.0553333
R31361 GNDA.n3136 GNDA.n3135 0.0553333
R31362 GNDA.n3127 GNDA.n3126 0.0553333
R31363 GNDA.n3118 GNDA.n3117 0.0553333
R31364 GNDA.n3109 GNDA.n3108 0.0553333
R31365 GNDA.n3002 GNDA.n3001 0.0553333
R31366 GNDA.n3016 GNDA.n3015 0.0553333
R31367 GNDA.n3032 GNDA.n3031 0.0553333
R31368 GNDA.n3046 GNDA.n3045 0.0553333
R31369 GNDA.n2926 GNDA.n2925 0.0553333
R31370 GNDA.n2940 GNDA.n2939 0.0553333
R31371 GNDA.n2956 GNDA.n2955 0.0553333
R31372 GNDA.n2970 GNDA.n2969 0.0553333
R31373 GNDA.n2902 GNDA.n2901 0.0553333
R31374 GNDA.n2893 GNDA.n2892 0.0553333
R31375 GNDA.n2884 GNDA.n2883 0.0553333
R31376 GNDA.n2875 GNDA.n2874 0.0553333
R31377 GNDA.n2768 GNDA.n2767 0.0553333
R31378 GNDA.n2782 GNDA.n2781 0.0553333
R31379 GNDA.n2798 GNDA.n2797 0.0553333
R31380 GNDA.n2812 GNDA.n2811 0.0553333
R31381 GNDA.n2690 GNDA.n2689 0.0553333
R31382 GNDA.n2693 GNDA.n2692 0.0553333
R31383 GNDA.n2703 GNDA.n2702 0.0553333
R31384 GNDA.n2710 GNDA.n2709 0.0553333
R31385 GNDA.n2720 GNDA.n2719 0.0553333
R31386 GNDA.n2723 GNDA.n2722 0.0553333
R31387 GNDA.n2732 GNDA.n2665 0.0553333
R31388 GNDA.n2739 GNDA.n2666 0.0553333
R31389 GNDA.n5550 GNDA.n5549 0.0553333
R31390 GNDA.n5564 GNDA.n5563 0.0553333
R31391 GNDA.n5580 GNDA.n5579 0.0553333
R31392 GNDA.n5594 GNDA.n5593 0.0553333
R31393 GNDA.n525 GNDA.n524 0.0553333
R31394 GNDA.n539 GNDA.n538 0.0553333
R31395 GNDA.n555 GNDA.n554 0.0553333
R31396 GNDA.n569 GNDA.n568 0.0553333
R31397 GNDA.n348 GNDA.n347 0.0553333
R31398 GNDA.n339 GNDA.n338 0.0553333
R31399 GNDA.n330 GNDA.n329 0.0553333
R31400 GNDA.n321 GNDA.n320 0.0553333
R31401 GNDA.n215 GNDA.n214 0.0553333
R31402 GNDA.n229 GNDA.n228 0.0553333
R31403 GNDA.n245 GNDA.n244 0.0553333
R31404 GNDA.n259 GNDA.n258 0.0553333
R31405 GNDA.n175 GNDA.n174 0.0553333
R31406 GNDA.n166 GNDA.n165 0.0553333
R31407 GNDA.n157 GNDA.n156 0.0553333
R31408 GNDA.n148 GNDA.n147 0.0553333
R31409 GNDA.n459 GNDA.n458 0.0553333
R31410 GNDA.n473 GNDA.n472 0.0553333
R31411 GNDA.n489 GNDA.n488 0.0553333
R31412 GNDA.n503 GNDA.n502 0.0553333
R31413 GNDA.n378 GNDA.n377 0.0553333
R31414 GNDA.n382 GNDA.n381 0.0553333
R31415 GNDA.n388 GNDA.n387 0.0553333
R31416 GNDA.n390 GNDA.n389 0.0553333
R31417 GNDA.n396 GNDA.n395 0.0553333
R31418 GNDA.n400 GNDA.n399 0.0553333
R31419 GNDA.n406 GNDA.n405 0.0553333
R31420 GNDA.n408 GNDA.n407 0.0553333
R31421 GNDA.n982 GNDA.n981 0.0553333
R31422 GNDA.n998 GNDA.n997 0.0553333
R31423 GNDA.n1012 GNDA.n1011 0.0553333
R31424 GNDA.n1028 GNDA.n966 0.0553333
R31425 GNDA.n5301 GNDA_2 0.0517
R31426 GNDA.n5372 GNDA_2 0.0517
R31427 GNDA_2 GNDA.n4639 0.0517
R31428 GNDA.n1794 GNDA_2 0.0517
R31429 GNDA_2 GNDA.n4730 0.0517
R31430 GNDA.n4463 GNDA_2 0.0517
R31431 GNDA.n1484 GNDA_2 0.0517
R31432 GNDA.n4932 GNDA_2 0.0517
R31433 GNDA.n4364 GNDA_2 0.0517
R31434 GNDA.n2110 GNDA.n2109 0.0514167
R31435 GNDA.n2104 GNDA.n2103 0.0514167
R31436 GNDA.n2101 GNDA.n2100 0.0514167
R31437 GNDA.n2095 GNDA.n2094 0.0514167
R31438 GNDA.n2092 GNDA.n2091 0.0514167
R31439 GNDA.n2086 GNDA.n2085 0.0514167
R31440 GNDA.n2083 GNDA.n2082 0.0514167
R31441 GNDA.n2077 GNDA.n2076 0.0514167
R31442 GNDA.n3663 GNDA.n3662 0.0514167
R31443 GNDA.n3668 GNDA.n3667 0.0514167
R31444 GNDA.n4099 GNDA.n3669 0.0514167
R31445 GNDA.n4102 GNDA.n3674 0.0514167
R31446 GNDA.n3678 GNDA.n3677 0.0514167
R31447 GNDA.n3683 GNDA.n3682 0.0514167
R31448 GNDA.n4108 GNDA.n3684 0.0514167
R31449 GNDA.n4112 GNDA.n3689 0.0514167
R31450 GNDA.n4049 GNDA.n4014 0.0514167
R31451 GNDA.n4057 GNDA.n4056 0.0514167
R31452 GNDA.n4043 GNDA.n4042 0.0514167
R31453 GNDA.n4039 GNDA.n4038 0.0514167
R31454 GNDA.n4073 GNDA.n4072 0.0514167
R31455 GNDA.n4081 GNDA.n4080 0.0514167
R31456 GNDA.n4031 GNDA.n4030 0.0514167
R31457 GNDA.n4093 GNDA.n4026 0.0514167
R31458 GNDA.n3968 GNDA.n3933 0.0514167
R31459 GNDA.n3976 GNDA.n3975 0.0514167
R31460 GNDA.n3962 GNDA.n3961 0.0514167
R31461 GNDA.n3958 GNDA.n3957 0.0514167
R31462 GNDA.n3992 GNDA.n3991 0.0514167
R31463 GNDA.n4000 GNDA.n3999 0.0514167
R31464 GNDA.n3950 GNDA.n3949 0.0514167
R31465 GNDA.n4012 GNDA.n3945 0.0514167
R31466 GNDA.n3887 GNDA.n3852 0.0514167
R31467 GNDA.n3895 GNDA.n3894 0.0514167
R31468 GNDA.n3881 GNDA.n3880 0.0514167
R31469 GNDA.n3877 GNDA.n3876 0.0514167
R31470 GNDA.n3911 GNDA.n3910 0.0514167
R31471 GNDA.n3919 GNDA.n3918 0.0514167
R31472 GNDA.n3869 GNDA.n3868 0.0514167
R31473 GNDA.n3931 GNDA.n3864 0.0514167
R31474 GNDA.n4191 GNDA.n3474 0.0514167
R31475 GNDA.n4199 GNDA.n4198 0.0514167
R31476 GNDA.n3504 GNDA.n3503 0.0514167
R31477 GNDA.n3500 GNDA.n3499 0.0514167
R31478 GNDA.n4215 GNDA.n4214 0.0514167
R31479 GNDA.n4223 GNDA.n4222 0.0514167
R31480 GNDA.n3492 GNDA.n3491 0.0514167
R31481 GNDA.n4235 GNDA.n3487 0.0514167
R31482 GNDA.n3806 GNDA.n3771 0.0514167
R31483 GNDA.n3814 GNDA.n3813 0.0514167
R31484 GNDA.n3800 GNDA.n3799 0.0514167
R31485 GNDA.n3796 GNDA.n3795 0.0514167
R31486 GNDA.n3830 GNDA.n3829 0.0514167
R31487 GNDA.n3838 GNDA.n3837 0.0514167
R31488 GNDA.n3788 GNDA.n3787 0.0514167
R31489 GNDA.n3850 GNDA.n3783 0.0514167
R31490 GNDA.n3725 GNDA.n3690 0.0514167
R31491 GNDA.n3733 GNDA.n3732 0.0514167
R31492 GNDA.n3719 GNDA.n3718 0.0514167
R31493 GNDA.n3715 GNDA.n3714 0.0514167
R31494 GNDA.n3749 GNDA.n3748 0.0514167
R31495 GNDA.n3757 GNDA.n3756 0.0514167
R31496 GNDA.n3707 GNDA.n3706 0.0514167
R31497 GNDA.n3769 GNDA.n3702 0.0514167
R31498 GNDA.n3516 GNDA.n3515 0.0514167
R31499 GNDA.n3524 GNDA.n3523 0.0514167
R31500 GNDA.n3529 GNDA.n3526 0.0514167
R31501 GNDA.n3537 GNDA.n3534 0.0514167
R31502 GNDA.n3540 GNDA.n3539 0.0514167
R31503 GNDA.n3548 GNDA.n3547 0.0514167
R31504 GNDA.n3553 GNDA.n3550 0.0514167
R31505 GNDA.n3559 GNDA.n3558 0.0514167
R31506 GNDA.n1976 GNDA.n1975 0.0514167
R31507 GNDA.n1981 GNDA.n1980 0.0514167
R31508 GNDA.n3462 GNDA.n1982 0.0514167
R31509 GNDA.n3465 GNDA.n1987 0.0514167
R31510 GNDA.n1991 GNDA.n1990 0.0514167
R31511 GNDA.n1996 GNDA.n1995 0.0514167
R31512 GNDA.n3471 GNDA.n1997 0.0514167
R31513 GNDA.n4238 GNDA.n2002 0.0514167
R31514 GNDA.n1064 GNDA.n1030 0.0514167
R31515 GNDA.n1072 GNDA.n1071 0.0514167
R31516 GNDA.n1059 GNDA.n1058 0.0514167
R31517 GNDA.n1055 GNDA.n1054 0.0514167
R31518 GNDA.n1088 GNDA.n1087 0.0514167
R31519 GNDA.n1096 GNDA.n1095 0.0514167
R31520 GNDA.n1047 GNDA.n1046 0.0514167
R31521 GNDA.n4895 GNDA.n1042 0.0514167
R31522 GNDA.n3402 GNDA.n3369 0.0514167
R31523 GNDA.n3412 GNDA.n3411 0.0514167
R31524 GNDA.n3418 GNDA.n3417 0.0514167
R31525 GNDA.n3428 GNDA.n3427 0.0514167
R31526 GNDA.n3432 GNDA.n3431 0.0514167
R31527 GNDA.n3442 GNDA.n3441 0.0514167
R31528 GNDA.n3448 GNDA.n3447 0.0514167
R31529 GNDA.n3456 GNDA.n3381 0.0514167
R31530 GNDA.n3313 GNDA.n2004 0.0514167
R31531 GNDA.n3323 GNDA.n3322 0.0514167
R31532 GNDA.n3329 GNDA.n3328 0.0514167
R31533 GNDA.n3339 GNDA.n3338 0.0514167
R31534 GNDA.n3343 GNDA.n3342 0.0514167
R31535 GNDA.n3353 GNDA.n3352 0.0514167
R31536 GNDA.n3359 GNDA.n3358 0.0514167
R31537 GNDA.n3367 GNDA.n2016 0.0514167
R31538 GNDA.n3286 GNDA.n2121 0.0514167
R31539 GNDA.n3240 GNDA.n3239 0.0514167
R31540 GNDA.n3246 GNDA.n3245 0.0514167
R31541 GNDA.n3256 GNDA.n3255 0.0514167
R31542 GNDA.n3260 GNDA.n3259 0.0514167
R31543 GNDA.n3270 GNDA.n3269 0.0514167
R31544 GNDA.n3276 GNDA.n3275 0.0514167
R31545 GNDA.n3284 GNDA.n3221 0.0514167
R31546 GNDA.n3154 GNDA.n2123 0.0514167
R31547 GNDA.n3164 GNDA.n3163 0.0514167
R31548 GNDA.n3170 GNDA.n3169 0.0514167
R31549 GNDA.n3180 GNDA.n3179 0.0514167
R31550 GNDA.n3184 GNDA.n3183 0.0514167
R31551 GNDA.n3194 GNDA.n3193 0.0514167
R31552 GNDA.n3200 GNDA.n3199 0.0514167
R31553 GNDA.n3208 GNDA.n2135 0.0514167
R31554 GNDA.n3139 GNDA.n3138 0.0514167
R31555 GNDA.n3133 GNDA.n3132 0.0514167
R31556 GNDA.n3130 GNDA.n3129 0.0514167
R31557 GNDA.n3124 GNDA.n3123 0.0514167
R31558 GNDA.n3121 GNDA.n3120 0.0514167
R31559 GNDA.n3115 GNDA.n3114 0.0514167
R31560 GNDA.n3112 GNDA.n3111 0.0514167
R31561 GNDA.n3106 GNDA.n3105 0.0514167
R31562 GNDA.n3052 GNDA.n2160 0.0514167
R31563 GNDA.n3006 GNDA.n3005 0.0514167
R31564 GNDA.n3012 GNDA.n3011 0.0514167
R31565 GNDA.n3022 GNDA.n3021 0.0514167
R31566 GNDA.n3026 GNDA.n3025 0.0514167
R31567 GNDA.n3036 GNDA.n3035 0.0514167
R31568 GNDA.n3042 GNDA.n3041 0.0514167
R31569 GNDA.n3050 GNDA.n2987 0.0514167
R31570 GNDA.n2920 GNDA.n2162 0.0514167
R31571 GNDA.n2930 GNDA.n2929 0.0514167
R31572 GNDA.n2936 GNDA.n2935 0.0514167
R31573 GNDA.n2946 GNDA.n2945 0.0514167
R31574 GNDA.n2950 GNDA.n2949 0.0514167
R31575 GNDA.n2960 GNDA.n2959 0.0514167
R31576 GNDA.n2966 GNDA.n2965 0.0514167
R31577 GNDA.n2974 GNDA.n2174 0.0514167
R31578 GNDA.n2905 GNDA.n2904 0.0514167
R31579 GNDA.n2899 GNDA.n2898 0.0514167
R31580 GNDA.n2896 GNDA.n2895 0.0514167
R31581 GNDA.n2890 GNDA.n2889 0.0514167
R31582 GNDA.n2887 GNDA.n2886 0.0514167
R31583 GNDA.n2881 GNDA.n2880 0.0514167
R31584 GNDA.n2878 GNDA.n2877 0.0514167
R31585 GNDA.n2872 GNDA.n2871 0.0514167
R31586 GNDA.n2818 GNDA.n2244 0.0514167
R31587 GNDA.n2772 GNDA.n2771 0.0514167
R31588 GNDA.n2778 GNDA.n2777 0.0514167
R31589 GNDA.n2788 GNDA.n2787 0.0514167
R31590 GNDA.n2792 GNDA.n2791 0.0514167
R31591 GNDA.n2802 GNDA.n2801 0.0514167
R31592 GNDA.n2808 GNDA.n2807 0.0514167
R31593 GNDA.n2816 GNDA.n2753 0.0514167
R31594 GNDA.n5544 GNDA.n1 0.0514167
R31595 GNDA.n5554 GNDA.n5553 0.0514167
R31596 GNDA.n5560 GNDA.n5559 0.0514167
R31597 GNDA.n5570 GNDA.n5569 0.0514167
R31598 GNDA.n5574 GNDA.n5573 0.0514167
R31599 GNDA.n5584 GNDA.n5583 0.0514167
R31600 GNDA.n5590 GNDA.n5589 0.0514167
R31601 GNDA.n5598 GNDA.n13 0.0514167
R31602 GNDA.n575 GNDA.n48 0.0514167
R31603 GNDA.n529 GNDA.n528 0.0514167
R31604 GNDA.n535 GNDA.n534 0.0514167
R31605 GNDA.n545 GNDA.n544 0.0514167
R31606 GNDA.n549 GNDA.n548 0.0514167
R31607 GNDA.n559 GNDA.n558 0.0514167
R31608 GNDA.n565 GNDA.n564 0.0514167
R31609 GNDA.n573 GNDA.n510 0.0514167
R31610 GNDA.n351 GNDA.n350 0.0514167
R31611 GNDA.n345 GNDA.n344 0.0514167
R31612 GNDA.n342 GNDA.n341 0.0514167
R31613 GNDA.n336 GNDA.n335 0.0514167
R31614 GNDA.n333 GNDA.n332 0.0514167
R31615 GNDA.n327 GNDA.n326 0.0514167
R31616 GNDA.n324 GNDA.n323 0.0514167
R31617 GNDA.n318 GNDA.n317 0.0514167
R31618 GNDA.n265 GNDA.n188 0.0514167
R31619 GNDA.n219 GNDA.n218 0.0514167
R31620 GNDA.n225 GNDA.n224 0.0514167
R31621 GNDA.n235 GNDA.n234 0.0514167
R31622 GNDA.n239 GNDA.n238 0.0514167
R31623 GNDA.n249 GNDA.n248 0.0514167
R31624 GNDA.n255 GNDA.n254 0.0514167
R31625 GNDA.n263 GNDA.n200 0.0514167
R31626 GNDA.n178 GNDA.n177 0.0514167
R31627 GNDA.n172 GNDA.n171 0.0514167
R31628 GNDA.n169 GNDA.n168 0.0514167
R31629 GNDA.n163 GNDA.n162 0.0514167
R31630 GNDA.n160 GNDA.n159 0.0514167
R31631 GNDA.n154 GNDA.n153 0.0514167
R31632 GNDA.n151 GNDA.n150 0.0514167
R31633 GNDA.n145 GNDA.n144 0.0514167
R31634 GNDA.n453 GNDA.n72 0.0514167
R31635 GNDA.n463 GNDA.n462 0.0514167
R31636 GNDA.n469 GNDA.n468 0.0514167
R31637 GNDA.n479 GNDA.n478 0.0514167
R31638 GNDA.n483 GNDA.n482 0.0514167
R31639 GNDA.n493 GNDA.n492 0.0514167
R31640 GNDA.n499 GNDA.n498 0.0514167
R31641 GNDA.n507 GNDA.n85 0.0514167
R31642 GNDA.n978 GNDA.n955 0.0514167
R31643 GNDA.n988 GNDA.n987 0.0514167
R31644 GNDA.n992 GNDA.n991 0.0514167
R31645 GNDA.n1002 GNDA.n1001 0.0514167
R31646 GNDA.n1008 GNDA.n1007 0.0514167
R31647 GNDA.n1018 GNDA.n1017 0.0514167
R31648 GNDA.n1022 GNDA.n1021 0.0514167
R31649 GNDA.n4898 GNDA.n953 0.0514167
R31650 GNDA.n2700 GNDA.n2699 0.0475
R31651 GNDA.n2713 GNDA.n2712 0.0475
R31652 GNDA.n2730 GNDA.n2729 0.0475
R31653 GNDA.n384 GNDA.n383 0.0475
R31654 GNDA.n394 GNDA.n393 0.0475
R31655 GNDA.n402 GNDA.n401 0.0475
R31656 GNDA.n3615 GNDA.n3609 0.0421667
R31657 GNDA.n3627 GNDA.n3608 0.0421667
R31658 GNDA.n5049 GNDA.n767 0.0421667
R31659 GNDA.n4890 GNDA.n4889 0.0421667
R31660 GNDA.n4187 GNDA.n3510 0.0421667
R31661 GNDA.n4178 GNDA.n3595 0.0421667
R31662 GNDA.n4174 GNDA.n3600 0.0421667
R31663 GNDA.n4170 GNDA.n3605 0.0421667
R31664 GNDA.n4166 GNDA.n4165 0.0421667
R31665 GNDA.n4162 GNDA.n3647 0.0421667
R31666 GNDA.n4158 GNDA.n3652 0.0421667
R31667 GNDA.n4154 GNDA.n3657 0.0421667
R31668 GNDA.n4150 GNDA.n4148 0.0421667
R31669 GNDA.n2681 GNDA.n2240 0.0421667
R31670 GNDA.n2825 GNDA.n2237 0.0421667
R31671 GNDA.n2912 GNDA.n2234 0.0421667
R31672 GNDA.n2232 GNDA.n2231 0.0421667
R31673 GNDA.n2227 GNDA.n2156 0.0421667
R31674 GNDA.n3059 GNDA.n2153 0.0421667
R31675 GNDA.n3146 GNDA.n2150 0.0421667
R31676 GNDA.n2148 GNDA.n2116 0.0421667
R31677 GNDA.n3293 GNDA.n3292 0.0421667
R31678 GNDA.n2030 GNDA.n2029 0.0421667
R31679 GNDA.n2210 GNDA.n2209 0.0421667
R31680 GNDA.n5436 GNDA.n655 0.0421667
R31681 GNDA.n653 GNDA.n652 0.0421667
R31682 GNDA.n658 GNDA.n657 0.0421667
R31683 GNDA.n684 GNDA.n682 0.0421667
R31684 GNDA.n5503 GNDA.n650 0.0421667
R31685 GNDA.n601 GNDA.n600 0.0421667
R31686 GNDA.n445 GNDA.n371 0.0421667
R31687 GNDA.n369 GNDA.n368 0.0421667
R31688 GNDA.n365 GNDA.n364 0.0421667
R31689 GNDA.n361 GNDA.n360 0.0421667
R31690 GNDA.n357 GNDA.n25 0.0421667
R31691 GNDA.n612 GNDA.n42 0.0421667
R31692 GNDA.n2108 GNDA.n2107 0.028198
R31693 GNDA.n2105 GNDA.n2104 0.028198
R31694 GNDA.n2099 GNDA.n2098 0.028198
R31695 GNDA.n2096 GNDA.n2095 0.028198
R31696 GNDA.n2090 GNDA.n2089 0.028198
R31697 GNDA.n2087 GNDA.n2086 0.028198
R31698 GNDA.n2081 GNDA.n2080 0.028198
R31699 GNDA.n2078 GNDA.n2077 0.028198
R31700 GNDA.n4095 GNDA.n3664 0.028198
R31701 GNDA.n4097 GNDA.n3667 0.028198
R31702 GNDA.n4100 GNDA.n3672 0.028198
R31703 GNDA.n4101 GNDA.n3674 0.028198
R31704 GNDA.n4104 GNDA.n3679 0.028198
R31705 GNDA.n4106 GNDA.n3682 0.028198
R31706 GNDA.n4109 GNDA.n3687 0.028198
R31707 GNDA.n4110 GNDA.n3689 0.028198
R31708 GNDA.n4046 GNDA.n4015 0.028198
R31709 GNDA.n4056 GNDA.n4016 0.028198
R31710 GNDA.n4064 GNDA.n4018 0.028198
R31711 GNDA.n4038 GNDA.n4019 0.028198
R31712 GNDA.n4034 GNDA.n4021 0.028198
R31713 GNDA.n4080 GNDA.n4022 0.028198
R31714 GNDA.n4088 GNDA.n4024 0.028198
R31715 GNDA.n4026 GNDA.n4025 0.028198
R31716 GNDA.n3965 GNDA.n3934 0.028198
R31717 GNDA.n3975 GNDA.n3935 0.028198
R31718 GNDA.n3983 GNDA.n3937 0.028198
R31719 GNDA.n3957 GNDA.n3938 0.028198
R31720 GNDA.n3953 GNDA.n3940 0.028198
R31721 GNDA.n3999 GNDA.n3941 0.028198
R31722 GNDA.n4007 GNDA.n3943 0.028198
R31723 GNDA.n3945 GNDA.n3944 0.028198
R31724 GNDA.n3884 GNDA.n3853 0.028198
R31725 GNDA.n3894 GNDA.n3854 0.028198
R31726 GNDA.n3902 GNDA.n3856 0.028198
R31727 GNDA.n3876 GNDA.n3857 0.028198
R31728 GNDA.n3872 GNDA.n3859 0.028198
R31729 GNDA.n3918 GNDA.n3860 0.028198
R31730 GNDA.n3926 GNDA.n3862 0.028198
R31731 GNDA.n3864 GNDA.n3863 0.028198
R31732 GNDA.n3507 GNDA.n3475 0.028198
R31733 GNDA.n4198 GNDA.n3476 0.028198
R31734 GNDA.n4206 GNDA.n3478 0.028198
R31735 GNDA.n3499 GNDA.n3479 0.028198
R31736 GNDA.n3495 GNDA.n3481 0.028198
R31737 GNDA.n4222 GNDA.n3482 0.028198
R31738 GNDA.n4230 GNDA.n3484 0.028198
R31739 GNDA.n3487 GNDA.n3485 0.028198
R31740 GNDA.n3803 GNDA.n3772 0.028198
R31741 GNDA.n3813 GNDA.n3773 0.028198
R31742 GNDA.n3821 GNDA.n3775 0.028198
R31743 GNDA.n3795 GNDA.n3776 0.028198
R31744 GNDA.n3791 GNDA.n3778 0.028198
R31745 GNDA.n3837 GNDA.n3779 0.028198
R31746 GNDA.n3845 GNDA.n3781 0.028198
R31747 GNDA.n3783 GNDA.n3782 0.028198
R31748 GNDA.n3722 GNDA.n3691 0.028198
R31749 GNDA.n3732 GNDA.n3692 0.028198
R31750 GNDA.n3740 GNDA.n3694 0.028198
R31751 GNDA.n3714 GNDA.n3695 0.028198
R31752 GNDA.n3710 GNDA.n3697 0.028198
R31753 GNDA.n3756 GNDA.n3698 0.028198
R31754 GNDA.n3764 GNDA.n3700 0.028198
R31755 GNDA.n3702 GNDA.n3701 0.028198
R31756 GNDA.n3518 GNDA.n3517 0.028198
R31757 GNDA.n3523 GNDA.n3522 0.028198
R31758 GNDA.n3531 GNDA.n3530 0.028198
R31759 GNDA.n3534 GNDA.n3533 0.028198
R31760 GNDA.n3542 GNDA.n3541 0.028198
R31761 GNDA.n3547 GNDA.n3546 0.028198
R31762 GNDA.n3555 GNDA.n3554 0.028198
R31763 GNDA.n3558 GNDA.n3557 0.028198
R31764 GNDA.n3458 GNDA.n1977 0.028198
R31765 GNDA.n3460 GNDA.n1980 0.028198
R31766 GNDA.n3463 GNDA.n1985 0.028198
R31767 GNDA.n3464 GNDA.n1987 0.028198
R31768 GNDA.n3467 GNDA.n1992 0.028198
R31769 GNDA.n3469 GNDA.n1995 0.028198
R31770 GNDA.n3472 GNDA.n2000 0.028198
R31771 GNDA.n3473 GNDA.n2002 0.028198
R31772 GNDA.n1062 GNDA.n1031 0.028198
R31773 GNDA.n1071 GNDA.n1032 0.028198
R31774 GNDA.n1079 GNDA.n1034 0.028198
R31775 GNDA.n1054 GNDA.n1035 0.028198
R31776 GNDA.n1050 GNDA.n1037 0.028198
R31777 GNDA.n1095 GNDA.n1038 0.028198
R31778 GNDA.n1103 GNDA.n1040 0.028198
R31779 GNDA.n1042 GNDA.n1041 0.028198
R31780 GNDA.n3407 GNDA.n3370 0.028198
R31781 GNDA.n3411 GNDA.n3371 0.028198
R31782 GNDA.n3421 GNDA.n3373 0.028198
R31783 GNDA.n3427 GNDA.n3374 0.028198
R31784 GNDA.n3437 GNDA.n3376 0.028198
R31785 GNDA.n3441 GNDA.n3377 0.028198
R31786 GNDA.n3451 GNDA.n3379 0.028198
R31787 GNDA.n3381 GNDA.n3380 0.028198
R31788 GNDA.n3318 GNDA.n2005 0.028198
R31789 GNDA.n3322 GNDA.n2006 0.028198
R31790 GNDA.n3332 GNDA.n2008 0.028198
R31791 GNDA.n3338 GNDA.n2009 0.028198
R31792 GNDA.n3348 GNDA.n2011 0.028198
R31793 GNDA.n3352 GNDA.n2012 0.028198
R31794 GNDA.n3362 GNDA.n2014 0.028198
R31795 GNDA.n2016 GNDA.n2015 0.028198
R31796 GNDA.n3235 GNDA.n3210 0.028198
R31797 GNDA.n3239 GNDA.n3211 0.028198
R31798 GNDA.n3249 GNDA.n3213 0.028198
R31799 GNDA.n3255 GNDA.n3214 0.028198
R31800 GNDA.n3265 GNDA.n3216 0.028198
R31801 GNDA.n3269 GNDA.n3217 0.028198
R31802 GNDA.n3279 GNDA.n3219 0.028198
R31803 GNDA.n3221 GNDA.n3220 0.028198
R31804 GNDA.n3159 GNDA.n2124 0.028198
R31805 GNDA.n3163 GNDA.n2125 0.028198
R31806 GNDA.n3173 GNDA.n2127 0.028198
R31807 GNDA.n3179 GNDA.n2128 0.028198
R31808 GNDA.n3189 GNDA.n2130 0.028198
R31809 GNDA.n3193 GNDA.n2131 0.028198
R31810 GNDA.n3203 GNDA.n2133 0.028198
R31811 GNDA.n2135 GNDA.n2134 0.028198
R31812 GNDA.n3137 GNDA.n3136 0.028198
R31813 GNDA.n3134 GNDA.n3133 0.028198
R31814 GNDA.n3128 GNDA.n3127 0.028198
R31815 GNDA.n3125 GNDA.n3124 0.028198
R31816 GNDA.n3119 GNDA.n3118 0.028198
R31817 GNDA.n3116 GNDA.n3115 0.028198
R31818 GNDA.n3110 GNDA.n3109 0.028198
R31819 GNDA.n3107 GNDA.n3106 0.028198
R31820 GNDA.n3001 GNDA.n2976 0.028198
R31821 GNDA.n3005 GNDA.n2977 0.028198
R31822 GNDA.n3015 GNDA.n2979 0.028198
R31823 GNDA.n3021 GNDA.n2980 0.028198
R31824 GNDA.n3031 GNDA.n2982 0.028198
R31825 GNDA.n3035 GNDA.n2983 0.028198
R31826 GNDA.n3045 GNDA.n2985 0.028198
R31827 GNDA.n2987 GNDA.n2986 0.028198
R31828 GNDA.n2925 GNDA.n2163 0.028198
R31829 GNDA.n2929 GNDA.n2164 0.028198
R31830 GNDA.n2939 GNDA.n2166 0.028198
R31831 GNDA.n2945 GNDA.n2167 0.028198
R31832 GNDA.n2955 GNDA.n2169 0.028198
R31833 GNDA.n2959 GNDA.n2170 0.028198
R31834 GNDA.n2969 GNDA.n2172 0.028198
R31835 GNDA.n2174 GNDA.n2173 0.028198
R31836 GNDA.n2903 GNDA.n2902 0.028198
R31837 GNDA.n2900 GNDA.n2899 0.028198
R31838 GNDA.n2894 GNDA.n2893 0.028198
R31839 GNDA.n2891 GNDA.n2890 0.028198
R31840 GNDA.n2885 GNDA.n2884 0.028198
R31841 GNDA.n2882 GNDA.n2881 0.028198
R31842 GNDA.n2876 GNDA.n2875 0.028198
R31843 GNDA.n2873 GNDA.n2872 0.028198
R31844 GNDA.n2767 GNDA.n2742 0.028198
R31845 GNDA.n2771 GNDA.n2743 0.028198
R31846 GNDA.n2781 GNDA.n2745 0.028198
R31847 GNDA.n2787 GNDA.n2746 0.028198
R31848 GNDA.n2797 GNDA.n2748 0.028198
R31849 GNDA.n2801 GNDA.n2749 0.028198
R31850 GNDA.n2811 GNDA.n2751 0.028198
R31851 GNDA.n2753 GNDA.n2752 0.028198
R31852 GNDA.n2812 GNDA.n2752 0.028198
R31853 GNDA.n2808 GNDA.n2751 0.028198
R31854 GNDA.n2798 GNDA.n2749 0.028198
R31855 GNDA.n2792 GNDA.n2748 0.028198
R31856 GNDA.n2782 GNDA.n2746 0.028198
R31857 GNDA.n2778 GNDA.n2745 0.028198
R31858 GNDA.n2768 GNDA.n2743 0.028198
R31859 GNDA.n2742 GNDA.n2244 0.028198
R31860 GNDA.n2874 GNDA.n2873 0.028198
R31861 GNDA.n2877 GNDA.n2876 0.028198
R31862 GNDA.n2883 GNDA.n2882 0.028198
R31863 GNDA.n2886 GNDA.n2885 0.028198
R31864 GNDA.n2892 GNDA.n2891 0.028198
R31865 GNDA.n2895 GNDA.n2894 0.028198
R31866 GNDA.n2901 GNDA.n2900 0.028198
R31867 GNDA.n2904 GNDA.n2903 0.028198
R31868 GNDA.n2970 GNDA.n2173 0.028198
R31869 GNDA.n2966 GNDA.n2172 0.028198
R31870 GNDA.n2956 GNDA.n2170 0.028198
R31871 GNDA.n2950 GNDA.n2169 0.028198
R31872 GNDA.n2940 GNDA.n2167 0.028198
R31873 GNDA.n2936 GNDA.n2166 0.028198
R31874 GNDA.n2926 GNDA.n2164 0.028198
R31875 GNDA.n2920 GNDA.n2163 0.028198
R31876 GNDA.n3046 GNDA.n2986 0.028198
R31877 GNDA.n3042 GNDA.n2985 0.028198
R31878 GNDA.n3032 GNDA.n2983 0.028198
R31879 GNDA.n3026 GNDA.n2982 0.028198
R31880 GNDA.n3016 GNDA.n2980 0.028198
R31881 GNDA.n3012 GNDA.n2979 0.028198
R31882 GNDA.n3002 GNDA.n2977 0.028198
R31883 GNDA.n2976 GNDA.n2160 0.028198
R31884 GNDA.n3108 GNDA.n3107 0.028198
R31885 GNDA.n3111 GNDA.n3110 0.028198
R31886 GNDA.n3117 GNDA.n3116 0.028198
R31887 GNDA.n3120 GNDA.n3119 0.028198
R31888 GNDA.n3126 GNDA.n3125 0.028198
R31889 GNDA.n3129 GNDA.n3128 0.028198
R31890 GNDA.n3135 GNDA.n3134 0.028198
R31891 GNDA.n3138 GNDA.n3137 0.028198
R31892 GNDA.n3204 GNDA.n2134 0.028198
R31893 GNDA.n3200 GNDA.n2133 0.028198
R31894 GNDA.n3190 GNDA.n2131 0.028198
R31895 GNDA.n3184 GNDA.n2130 0.028198
R31896 GNDA.n3174 GNDA.n2128 0.028198
R31897 GNDA.n3170 GNDA.n2127 0.028198
R31898 GNDA.n3160 GNDA.n2125 0.028198
R31899 GNDA.n3154 GNDA.n2124 0.028198
R31900 GNDA.n3280 GNDA.n3220 0.028198
R31901 GNDA.n3276 GNDA.n3219 0.028198
R31902 GNDA.n3266 GNDA.n3217 0.028198
R31903 GNDA.n3260 GNDA.n3216 0.028198
R31904 GNDA.n3250 GNDA.n3214 0.028198
R31905 GNDA.n3246 GNDA.n3213 0.028198
R31906 GNDA.n3236 GNDA.n3211 0.028198
R31907 GNDA.n3210 GNDA.n2121 0.028198
R31908 GNDA.n3363 GNDA.n2015 0.028198
R31909 GNDA.n3359 GNDA.n2014 0.028198
R31910 GNDA.n3349 GNDA.n2012 0.028198
R31911 GNDA.n3343 GNDA.n2011 0.028198
R31912 GNDA.n3333 GNDA.n2009 0.028198
R31913 GNDA.n3329 GNDA.n2008 0.028198
R31914 GNDA.n3319 GNDA.n2006 0.028198
R31915 GNDA.n3313 GNDA.n2005 0.028198
R31916 GNDA.n3452 GNDA.n3380 0.028198
R31917 GNDA.n3448 GNDA.n3379 0.028198
R31918 GNDA.n3438 GNDA.n3377 0.028198
R31919 GNDA.n3432 GNDA.n3376 0.028198
R31920 GNDA.n3422 GNDA.n3374 0.028198
R31921 GNDA.n3418 GNDA.n3373 0.028198
R31922 GNDA.n3408 GNDA.n3371 0.028198
R31923 GNDA.n3402 GNDA.n3370 0.028198
R31924 GNDA.n2079 GNDA.n2078 0.028198
R31925 GNDA.n2082 GNDA.n2081 0.028198
R31926 GNDA.n2088 GNDA.n2087 0.028198
R31927 GNDA.n2091 GNDA.n2090 0.028198
R31928 GNDA.n2097 GNDA.n2096 0.028198
R31929 GNDA.n2100 GNDA.n2099 0.028198
R31930 GNDA.n2106 GNDA.n2105 0.028198
R31931 GNDA.n2109 GNDA.n2108 0.028198
R31932 GNDA.n3473 GNDA.n2001 0.028198
R31933 GNDA.n3472 GNDA.n3471 0.028198
R31934 GNDA.n3469 GNDA.n3468 0.028198
R31935 GNDA.n3467 GNDA.n1991 0.028198
R31936 GNDA.n3464 GNDA.n1986 0.028198
R31937 GNDA.n3463 GNDA.n3462 0.028198
R31938 GNDA.n3460 GNDA.n3459 0.028198
R31939 GNDA.n3458 GNDA.n1976 0.028198
R31940 GNDA.n3557 GNDA.n3556 0.028198
R31941 GNDA.n3554 GNDA.n3553 0.028198
R31942 GNDA.n3546 GNDA.n3545 0.028198
R31943 GNDA.n3541 GNDA.n3540 0.028198
R31944 GNDA.n3533 GNDA.n3532 0.028198
R31945 GNDA.n3530 GNDA.n3529 0.028198
R31946 GNDA.n3522 GNDA.n3521 0.028198
R31947 GNDA.n3517 GNDA.n3516 0.028198
R31948 GNDA.n3765 GNDA.n3701 0.028198
R31949 GNDA.n3707 GNDA.n3700 0.028198
R31950 GNDA.n3711 GNDA.n3698 0.028198
R31951 GNDA.n3749 GNDA.n3697 0.028198
R31952 GNDA.n3741 GNDA.n3695 0.028198
R31953 GNDA.n3719 GNDA.n3694 0.028198
R31954 GNDA.n3723 GNDA.n3692 0.028198
R31955 GNDA.n3725 GNDA.n3691 0.028198
R31956 GNDA.n3846 GNDA.n3782 0.028198
R31957 GNDA.n3788 GNDA.n3781 0.028198
R31958 GNDA.n3792 GNDA.n3779 0.028198
R31959 GNDA.n3830 GNDA.n3778 0.028198
R31960 GNDA.n3822 GNDA.n3776 0.028198
R31961 GNDA.n3800 GNDA.n3775 0.028198
R31962 GNDA.n3804 GNDA.n3773 0.028198
R31963 GNDA.n3806 GNDA.n3772 0.028198
R31964 GNDA.n4231 GNDA.n3485 0.028198
R31965 GNDA.n3492 GNDA.n3484 0.028198
R31966 GNDA.n3496 GNDA.n3482 0.028198
R31967 GNDA.n4215 GNDA.n3481 0.028198
R31968 GNDA.n4207 GNDA.n3479 0.028198
R31969 GNDA.n3504 GNDA.n3478 0.028198
R31970 GNDA.n3508 GNDA.n3476 0.028198
R31971 GNDA.n4191 GNDA.n3475 0.028198
R31972 GNDA.n3927 GNDA.n3863 0.028198
R31973 GNDA.n3869 GNDA.n3862 0.028198
R31974 GNDA.n3873 GNDA.n3860 0.028198
R31975 GNDA.n3911 GNDA.n3859 0.028198
R31976 GNDA.n3903 GNDA.n3857 0.028198
R31977 GNDA.n3881 GNDA.n3856 0.028198
R31978 GNDA.n3885 GNDA.n3854 0.028198
R31979 GNDA.n3887 GNDA.n3853 0.028198
R31980 GNDA.n4008 GNDA.n3944 0.028198
R31981 GNDA.n3950 GNDA.n3943 0.028198
R31982 GNDA.n3954 GNDA.n3941 0.028198
R31983 GNDA.n3992 GNDA.n3940 0.028198
R31984 GNDA.n3984 GNDA.n3938 0.028198
R31985 GNDA.n3962 GNDA.n3937 0.028198
R31986 GNDA.n3966 GNDA.n3935 0.028198
R31987 GNDA.n3968 GNDA.n3934 0.028198
R31988 GNDA.n4089 GNDA.n4025 0.028198
R31989 GNDA.n4031 GNDA.n4024 0.028198
R31990 GNDA.n4035 GNDA.n4022 0.028198
R31991 GNDA.n4073 GNDA.n4021 0.028198
R31992 GNDA.n4065 GNDA.n4019 0.028198
R31993 GNDA.n4043 GNDA.n4018 0.028198
R31994 GNDA.n4047 GNDA.n4016 0.028198
R31995 GNDA.n4049 GNDA.n4015 0.028198
R31996 GNDA.n4110 GNDA.n3688 0.028198
R31997 GNDA.n4109 GNDA.n4108 0.028198
R31998 GNDA.n4106 GNDA.n4105 0.028198
R31999 GNDA.n4104 GNDA.n3678 0.028198
R32000 GNDA.n4101 GNDA.n3673 0.028198
R32001 GNDA.n4100 GNDA.n4099 0.028198
R32002 GNDA.n4097 GNDA.n4096 0.028198
R32003 GNDA.n4095 GNDA.n3663 0.028198
R32004 GNDA.n5549 GNDA.n2 0.028198
R32005 GNDA.n5553 GNDA.n3 0.028198
R32006 GNDA.n5563 GNDA.n5 0.028198
R32007 GNDA.n5569 GNDA.n6 0.028198
R32008 GNDA.n5579 GNDA.n8 0.028198
R32009 GNDA.n5583 GNDA.n9 0.028198
R32010 GNDA.n5593 GNDA.n11 0.028198
R32011 GNDA.n13 GNDA.n12 0.028198
R32012 GNDA.n524 GNDA.n49 0.028198
R32013 GNDA.n528 GNDA.n50 0.028198
R32014 GNDA.n538 GNDA.n52 0.028198
R32015 GNDA.n544 GNDA.n53 0.028198
R32016 GNDA.n554 GNDA.n55 0.028198
R32017 GNDA.n558 GNDA.n56 0.028198
R32018 GNDA.n568 GNDA.n58 0.028198
R32019 GNDA.n510 GNDA.n59 0.028198
R32020 GNDA.n349 GNDA.n348 0.028198
R32021 GNDA.n346 GNDA.n345 0.028198
R32022 GNDA.n340 GNDA.n339 0.028198
R32023 GNDA.n337 GNDA.n336 0.028198
R32024 GNDA.n331 GNDA.n330 0.028198
R32025 GNDA.n328 GNDA.n327 0.028198
R32026 GNDA.n322 GNDA.n321 0.028198
R32027 GNDA.n319 GNDA.n318 0.028198
R32028 GNDA.n214 GNDA.n189 0.028198
R32029 GNDA.n218 GNDA.n190 0.028198
R32030 GNDA.n228 GNDA.n192 0.028198
R32031 GNDA.n234 GNDA.n193 0.028198
R32032 GNDA.n244 GNDA.n195 0.028198
R32033 GNDA.n248 GNDA.n196 0.028198
R32034 GNDA.n258 GNDA.n198 0.028198
R32035 GNDA.n200 GNDA.n199 0.028198
R32036 GNDA.n176 GNDA.n175 0.028198
R32037 GNDA.n173 GNDA.n172 0.028198
R32038 GNDA.n167 GNDA.n166 0.028198
R32039 GNDA.n164 GNDA.n163 0.028198
R32040 GNDA.n158 GNDA.n157 0.028198
R32041 GNDA.n155 GNDA.n154 0.028198
R32042 GNDA.n149 GNDA.n148 0.028198
R32043 GNDA.n146 GNDA.n145 0.028198
R32044 GNDA.n458 GNDA.n73 0.028198
R32045 GNDA.n462 GNDA.n74 0.028198
R32046 GNDA.n472 GNDA.n76 0.028198
R32047 GNDA.n478 GNDA.n77 0.028198
R32048 GNDA.n488 GNDA.n79 0.028198
R32049 GNDA.n492 GNDA.n80 0.028198
R32050 GNDA.n502 GNDA.n82 0.028198
R32051 GNDA.n85 GNDA.n83 0.028198
R32052 GNDA.n503 GNDA.n83 0.028198
R32053 GNDA.n499 GNDA.n82 0.028198
R32054 GNDA.n489 GNDA.n80 0.028198
R32055 GNDA.n483 GNDA.n79 0.028198
R32056 GNDA.n473 GNDA.n77 0.028198
R32057 GNDA.n469 GNDA.n76 0.028198
R32058 GNDA.n459 GNDA.n74 0.028198
R32059 GNDA.n453 GNDA.n73 0.028198
R32060 GNDA.n147 GNDA.n146 0.028198
R32061 GNDA.n150 GNDA.n149 0.028198
R32062 GNDA.n156 GNDA.n155 0.028198
R32063 GNDA.n159 GNDA.n158 0.028198
R32064 GNDA.n165 GNDA.n164 0.028198
R32065 GNDA.n168 GNDA.n167 0.028198
R32066 GNDA.n174 GNDA.n173 0.028198
R32067 GNDA.n177 GNDA.n176 0.028198
R32068 GNDA.n259 GNDA.n199 0.028198
R32069 GNDA.n255 GNDA.n198 0.028198
R32070 GNDA.n245 GNDA.n196 0.028198
R32071 GNDA.n239 GNDA.n195 0.028198
R32072 GNDA.n229 GNDA.n193 0.028198
R32073 GNDA.n225 GNDA.n192 0.028198
R32074 GNDA.n215 GNDA.n190 0.028198
R32075 GNDA.n189 GNDA.n188 0.028198
R32076 GNDA.n320 GNDA.n319 0.028198
R32077 GNDA.n323 GNDA.n322 0.028198
R32078 GNDA.n329 GNDA.n328 0.028198
R32079 GNDA.n332 GNDA.n331 0.028198
R32080 GNDA.n338 GNDA.n337 0.028198
R32081 GNDA.n341 GNDA.n340 0.028198
R32082 GNDA.n347 GNDA.n346 0.028198
R32083 GNDA.n350 GNDA.n349 0.028198
R32084 GNDA.n569 GNDA.n59 0.028198
R32085 GNDA.n565 GNDA.n58 0.028198
R32086 GNDA.n555 GNDA.n56 0.028198
R32087 GNDA.n549 GNDA.n55 0.028198
R32088 GNDA.n539 GNDA.n53 0.028198
R32089 GNDA.n535 GNDA.n52 0.028198
R32090 GNDA.n525 GNDA.n50 0.028198
R32091 GNDA.n49 GNDA.n48 0.028198
R32092 GNDA.n5594 GNDA.n12 0.028198
R32093 GNDA.n5590 GNDA.n11 0.028198
R32094 GNDA.n5580 GNDA.n9 0.028198
R32095 GNDA.n5574 GNDA.n8 0.028198
R32096 GNDA.n5564 GNDA.n6 0.028198
R32097 GNDA.n5560 GNDA.n5 0.028198
R32098 GNDA.n5550 GNDA.n3 0.028198
R32099 GNDA.n5544 GNDA.n2 0.028198
R32100 GNDA.n981 GNDA.n956 0.028198
R32101 GNDA.n987 GNDA.n957 0.028198
R32102 GNDA.n997 GNDA.n959 0.028198
R32103 GNDA.n1001 GNDA.n960 0.028198
R32104 GNDA.n1011 GNDA.n962 0.028198
R32105 GNDA.n1017 GNDA.n963 0.028198
R32106 GNDA.n966 GNDA.n965 0.028198
R32107 GNDA.n1029 GNDA.n953 0.028198
R32108 GNDA.n1029 GNDA.n1028 0.028198
R32109 GNDA.n1022 GNDA.n965 0.028198
R32110 GNDA.n1012 GNDA.n963 0.028198
R32111 GNDA.n1008 GNDA.n962 0.028198
R32112 GNDA.n998 GNDA.n960 0.028198
R32113 GNDA.n992 GNDA.n959 0.028198
R32114 GNDA.n982 GNDA.n957 0.028198
R32115 GNDA.n978 GNDA.n956 0.028198
R32116 GNDA.n1104 GNDA.n1041 0.028198
R32117 GNDA.n1047 GNDA.n1040 0.028198
R32118 GNDA.n1051 GNDA.n1038 0.028198
R32119 GNDA.n1088 GNDA.n1037 0.028198
R32120 GNDA.n1080 GNDA.n1035 0.028198
R32121 GNDA.n1059 GNDA.n1034 0.028198
R32122 GNDA.n1063 GNDA.n1032 0.028198
R32123 GNDA.n1064 GNDA.n1031 0.028198
R32124 GNDA.n2690 GNDA.n2656 0.028198
R32125 GNDA.n2702 GNDA.n2659 0.028198
R32126 GNDA.n2720 GNDA.n2662 0.028198
R32127 GNDA.n2740 GNDA.n2665 0.028198
R32128 GNDA.n2740 GNDA.n2739 0.028198
R32129 GNDA.n2723 GNDA.n2662 0.028198
R32130 GNDA.n2709 GNDA.n2659 0.028198
R32131 GNDA.n2693 GNDA.n2656 0.028198
R32132 GNDA.n378 GNDA.n62 0.028198
R32133 GNDA.n388 GNDA.n65 0.028198
R32134 GNDA.n396 GNDA.n68 0.028198
R32135 GNDA.n406 GNDA.n71 0.028198
R32136 GNDA.n407 GNDA.n71 0.028198
R32137 GNDA.n399 GNDA.n68 0.028198
R32138 GNDA.n389 GNDA.n65 0.028198
R32139 GNDA.n381 GNDA.n62 0.028198
R32140 GNDA.n2692 GNDA.n2657 0.0262697
R32141 GNDA.n2700 GNDA.n2658 0.0262697
R32142 GNDA.n2710 GNDA.n2660 0.0262697
R32143 GNDA.n2712 GNDA.n2661 0.0262697
R32144 GNDA.n2722 GNDA.n2663 0.0262697
R32145 GNDA.n2730 GNDA.n2664 0.0262697
R32146 GNDA.n2666 GNDA.n2654 0.0262697
R32147 GNDA.n2732 GNDA.n2664 0.0262697
R32148 GNDA.n2729 GNDA.n2663 0.0262697
R32149 GNDA.n2719 GNDA.n2661 0.0262697
R32150 GNDA.n2713 GNDA.n2660 0.0262697
R32151 GNDA.n2703 GNDA.n2658 0.0262697
R32152 GNDA.n2699 GNDA.n2657 0.0262697
R32153 GNDA.n2689 GNDA.n2655 0.0262697
R32154 GNDA.n382 GNDA.n63 0.0262697
R32155 GNDA.n384 GNDA.n64 0.0262697
R32156 GNDA.n390 GNDA.n66 0.0262697
R32157 GNDA.n394 GNDA.n67 0.0262697
R32158 GNDA.n400 GNDA.n69 0.0262697
R32159 GNDA.n402 GNDA.n70 0.0262697
R32160 GNDA.n408 GNDA.n60 0.0262697
R32161 GNDA.n405 GNDA.n70 0.0262697
R32162 GNDA.n401 GNDA.n69 0.0262697
R32163 GNDA.n395 GNDA.n67 0.0262697
R32164 GNDA.n393 GNDA.n66 0.0262697
R32165 GNDA.n387 GNDA.n64 0.0262697
R32166 GNDA.n383 GNDA.n63 0.0262697
R32167 GNDA.n377 GNDA.n61 0.0262697
R32168 GNDA.n2102 GNDA.n2101 0.0243392
R32169 GNDA.n2093 GNDA.n2092 0.0243392
R32170 GNDA.n2084 GNDA.n2083 0.0243392
R32171 GNDA.n4098 GNDA.n3669 0.0243392
R32172 GNDA.n4103 GNDA.n3677 0.0243392
R32173 GNDA.n4107 GNDA.n3684 0.0243392
R32174 GNDA.n4042 GNDA.n4017 0.0243392
R32175 GNDA.n4072 GNDA.n4020 0.0243392
R32176 GNDA.n4030 GNDA.n4023 0.0243392
R32177 GNDA.n3961 GNDA.n3936 0.0243392
R32178 GNDA.n3991 GNDA.n3939 0.0243392
R32179 GNDA.n3949 GNDA.n3942 0.0243392
R32180 GNDA.n3880 GNDA.n3855 0.0243392
R32181 GNDA.n3910 GNDA.n3858 0.0243392
R32182 GNDA.n3868 GNDA.n3861 0.0243392
R32183 GNDA.n3503 GNDA.n3477 0.0243392
R32184 GNDA.n4214 GNDA.n3480 0.0243392
R32185 GNDA.n3491 GNDA.n3483 0.0243392
R32186 GNDA.n3799 GNDA.n3774 0.0243392
R32187 GNDA.n3829 GNDA.n3777 0.0243392
R32188 GNDA.n3787 GNDA.n3780 0.0243392
R32189 GNDA.n3718 GNDA.n3693 0.0243392
R32190 GNDA.n3748 GNDA.n3696 0.0243392
R32191 GNDA.n3706 GNDA.n3699 0.0243392
R32192 GNDA.n3526 GNDA.n3525 0.0243392
R32193 GNDA.n3539 GNDA.n3538 0.0243392
R32194 GNDA.n3550 GNDA.n3549 0.0243392
R32195 GNDA.n3461 GNDA.n1982 0.0243392
R32196 GNDA.n3466 GNDA.n1990 0.0243392
R32197 GNDA.n3470 GNDA.n1997 0.0243392
R32198 GNDA.n1058 GNDA.n1033 0.0243392
R32199 GNDA.n1087 GNDA.n1036 0.0243392
R32200 GNDA.n1046 GNDA.n1039 0.0243392
R32201 GNDA.n3417 GNDA.n3372 0.0243392
R32202 GNDA.n3431 GNDA.n3375 0.0243392
R32203 GNDA.n3447 GNDA.n3378 0.0243392
R32204 GNDA.n3328 GNDA.n2007 0.0243392
R32205 GNDA.n3342 GNDA.n2010 0.0243392
R32206 GNDA.n3358 GNDA.n2013 0.0243392
R32207 GNDA.n3245 GNDA.n3212 0.0243392
R32208 GNDA.n3259 GNDA.n3215 0.0243392
R32209 GNDA.n3275 GNDA.n3218 0.0243392
R32210 GNDA.n3169 GNDA.n2126 0.0243392
R32211 GNDA.n3183 GNDA.n2129 0.0243392
R32212 GNDA.n3199 GNDA.n2132 0.0243392
R32213 GNDA.n3131 GNDA.n3130 0.0243392
R32214 GNDA.n3122 GNDA.n3121 0.0243392
R32215 GNDA.n3113 GNDA.n3112 0.0243392
R32216 GNDA.n3011 GNDA.n2978 0.0243392
R32217 GNDA.n3025 GNDA.n2981 0.0243392
R32218 GNDA.n3041 GNDA.n2984 0.0243392
R32219 GNDA.n2935 GNDA.n2165 0.0243392
R32220 GNDA.n2949 GNDA.n2168 0.0243392
R32221 GNDA.n2965 GNDA.n2171 0.0243392
R32222 GNDA.n2897 GNDA.n2896 0.0243392
R32223 GNDA.n2888 GNDA.n2887 0.0243392
R32224 GNDA.n2879 GNDA.n2878 0.0243392
R32225 GNDA.n2777 GNDA.n2744 0.0243392
R32226 GNDA.n2791 GNDA.n2747 0.0243392
R32227 GNDA.n2807 GNDA.n2750 0.0243392
R32228 GNDA.n2802 GNDA.n2750 0.0243392
R32229 GNDA.n2788 GNDA.n2747 0.0243392
R32230 GNDA.n2772 GNDA.n2744 0.0243392
R32231 GNDA.n2880 GNDA.n2879 0.0243392
R32232 GNDA.n2889 GNDA.n2888 0.0243392
R32233 GNDA.n2898 GNDA.n2897 0.0243392
R32234 GNDA.n2960 GNDA.n2171 0.0243392
R32235 GNDA.n2946 GNDA.n2168 0.0243392
R32236 GNDA.n2930 GNDA.n2165 0.0243392
R32237 GNDA.n3036 GNDA.n2984 0.0243392
R32238 GNDA.n3022 GNDA.n2981 0.0243392
R32239 GNDA.n3006 GNDA.n2978 0.0243392
R32240 GNDA.n3114 GNDA.n3113 0.0243392
R32241 GNDA.n3123 GNDA.n3122 0.0243392
R32242 GNDA.n3132 GNDA.n3131 0.0243392
R32243 GNDA.n3194 GNDA.n2132 0.0243392
R32244 GNDA.n3180 GNDA.n2129 0.0243392
R32245 GNDA.n3164 GNDA.n2126 0.0243392
R32246 GNDA.n3270 GNDA.n3218 0.0243392
R32247 GNDA.n3256 GNDA.n3215 0.0243392
R32248 GNDA.n3240 GNDA.n3212 0.0243392
R32249 GNDA.n3353 GNDA.n2013 0.0243392
R32250 GNDA.n3339 GNDA.n2010 0.0243392
R32251 GNDA.n3323 GNDA.n2007 0.0243392
R32252 GNDA.n3442 GNDA.n3378 0.0243392
R32253 GNDA.n3428 GNDA.n3375 0.0243392
R32254 GNDA.n3412 GNDA.n3372 0.0243392
R32255 GNDA.n2085 GNDA.n2084 0.0243392
R32256 GNDA.n2094 GNDA.n2093 0.0243392
R32257 GNDA.n2103 GNDA.n2102 0.0243392
R32258 GNDA.n3470 GNDA.n1996 0.0243392
R32259 GNDA.n3466 GNDA.n3465 0.0243392
R32260 GNDA.n3461 GNDA.n1981 0.0243392
R32261 GNDA.n3549 GNDA.n3548 0.0243392
R32262 GNDA.n3538 GNDA.n3537 0.0243392
R32263 GNDA.n3525 GNDA.n3524 0.0243392
R32264 GNDA.n3757 GNDA.n3699 0.0243392
R32265 GNDA.n3715 GNDA.n3696 0.0243392
R32266 GNDA.n3733 GNDA.n3693 0.0243392
R32267 GNDA.n3838 GNDA.n3780 0.0243392
R32268 GNDA.n3796 GNDA.n3777 0.0243392
R32269 GNDA.n3814 GNDA.n3774 0.0243392
R32270 GNDA.n4223 GNDA.n3483 0.0243392
R32271 GNDA.n3500 GNDA.n3480 0.0243392
R32272 GNDA.n4199 GNDA.n3477 0.0243392
R32273 GNDA.n3919 GNDA.n3861 0.0243392
R32274 GNDA.n3877 GNDA.n3858 0.0243392
R32275 GNDA.n3895 GNDA.n3855 0.0243392
R32276 GNDA.n4000 GNDA.n3942 0.0243392
R32277 GNDA.n3958 GNDA.n3939 0.0243392
R32278 GNDA.n3976 GNDA.n3936 0.0243392
R32279 GNDA.n4081 GNDA.n4023 0.0243392
R32280 GNDA.n4039 GNDA.n4020 0.0243392
R32281 GNDA.n4057 GNDA.n4017 0.0243392
R32282 GNDA.n4107 GNDA.n3683 0.0243392
R32283 GNDA.n4103 GNDA.n4102 0.0243392
R32284 GNDA.n4098 GNDA.n3668 0.0243392
R32285 GNDA.n5559 GNDA.n4 0.0243392
R32286 GNDA.n5573 GNDA.n7 0.0243392
R32287 GNDA.n5589 GNDA.n10 0.0243392
R32288 GNDA.n534 GNDA.n51 0.0243392
R32289 GNDA.n548 GNDA.n54 0.0243392
R32290 GNDA.n564 GNDA.n57 0.0243392
R32291 GNDA.n343 GNDA.n342 0.0243392
R32292 GNDA.n334 GNDA.n333 0.0243392
R32293 GNDA.n325 GNDA.n324 0.0243392
R32294 GNDA.n224 GNDA.n191 0.0243392
R32295 GNDA.n238 GNDA.n194 0.0243392
R32296 GNDA.n254 GNDA.n197 0.0243392
R32297 GNDA.n170 GNDA.n169 0.0243392
R32298 GNDA.n161 GNDA.n160 0.0243392
R32299 GNDA.n152 GNDA.n151 0.0243392
R32300 GNDA.n468 GNDA.n75 0.0243392
R32301 GNDA.n482 GNDA.n78 0.0243392
R32302 GNDA.n498 GNDA.n81 0.0243392
R32303 GNDA.n493 GNDA.n81 0.0243392
R32304 GNDA.n479 GNDA.n78 0.0243392
R32305 GNDA.n463 GNDA.n75 0.0243392
R32306 GNDA.n153 GNDA.n152 0.0243392
R32307 GNDA.n162 GNDA.n161 0.0243392
R32308 GNDA.n171 GNDA.n170 0.0243392
R32309 GNDA.n249 GNDA.n197 0.0243392
R32310 GNDA.n235 GNDA.n194 0.0243392
R32311 GNDA.n219 GNDA.n191 0.0243392
R32312 GNDA.n326 GNDA.n325 0.0243392
R32313 GNDA.n335 GNDA.n334 0.0243392
R32314 GNDA.n344 GNDA.n343 0.0243392
R32315 GNDA.n559 GNDA.n57 0.0243392
R32316 GNDA.n545 GNDA.n54 0.0243392
R32317 GNDA.n529 GNDA.n51 0.0243392
R32318 GNDA.n5584 GNDA.n10 0.0243392
R32319 GNDA.n5570 GNDA.n7 0.0243392
R32320 GNDA.n5554 GNDA.n4 0.0243392
R32321 GNDA.n991 GNDA.n958 0.0243392
R32322 GNDA.n1007 GNDA.n961 0.0243392
R32323 GNDA.n1021 GNDA.n964 0.0243392
R32324 GNDA.n1018 GNDA.n964 0.0243392
R32325 GNDA.n1002 GNDA.n961 0.0243392
R32326 GNDA.n988 GNDA.n958 0.0243392
R32327 GNDA.n1096 GNDA.n1039 0.0243392
R32328 GNDA.n1055 GNDA.n1036 0.0243392
R32329 GNDA.n1072 GNDA.n1033 0.0243392
R32330 GNDA.n2217 GNDA.n2216 0.0217373
R32331 GNDA.n2221 GNDA.n2211 0.0217373
R32332 GNDA.n2222 GNDA.n2221 0.0217373
R32333 GNDA.n2225 GNDA.n2224 0.0217373
R32334 GNDA.n2229 GNDA.n2228 0.0217373
R32335 GNDA.n2215 GNDA.n2212 0.0217373
R32336 GNDA.n2218 GNDA.n2217 0.0217373
R32337 GNDA.n4151 GNDA.n3660 0.0217373
R32338 GNDA.n4155 GNDA.n3655 0.0217373
R32339 GNDA.n4159 GNDA.n3650 0.0217373
R32340 GNDA.n4163 GNDA.n3645 0.0217373
R32341 GNDA.n4171 GNDA.n3603 0.0217373
R32342 GNDA.n4175 GNDA.n3598 0.0217373
R32343 GNDA.n4179 GNDA.n3513 0.0217373
R32344 GNDA.n3633 GNDA.n3632 0.0217373
R32345 GNDA.n3636 GNDA.n3635 0.0217373
R32346 GNDA.n3639 GNDA.n3607 0.0217373
R32347 GNDA.n3642 GNDA.n3606 0.0217373
R32348 GNDA.n3641 GNDA.n3606 0.0217373
R32349 GNDA.n3631 GNDA.n3628 0.0217373
R32350 GNDA.n3634 GNDA.n3633 0.0217373
R32351 GNDA.n3610 GNDA.n3609 0.0217373
R32352 GNDA.n3635 GNDA.n3626 0.0217373
R32353 GNDA.n3626 GNDA.n3607 0.0217373
R32354 GNDA.n5148 GNDA.n5066 0.0217373
R32355 GNDA.n5151 GNDA.n5050 0.0217373
R32356 GNDA.n5065 GNDA.n5052 0.0217373
R32357 GNDA.n5066 GNDA.n5053 0.0217373
R32358 GNDA.n5047 GNDA.n5046 0.0217373
R32359 GNDA.n5050 GNDA.n5046 0.0217373
R32360 GNDA.n4892 GNDA.n4891 0.0217373
R32361 GNDA.n4888 GNDA.n763 0.0217373
R32362 GNDA.n5320 GNDA.n765 0.0217373
R32363 GNDA.n5321 GNDA.n766 0.0217373
R32364 GNDA.n4891 GNDA.n4887 0.0217373
R32365 GNDA.n4888 GNDA.n4887 0.0217373
R32366 GNDA.n3393 GNDA.n1972 0.0217373
R32367 GNDA.n4167 GNDA.n4166 0.0217373
R32368 GNDA.n4177 GNDA.n3511 0.0217373
R32369 GNDA.n3513 GNDA.n3511 0.0217373
R32370 GNDA.n4173 GNDA.n3596 0.0217373
R32371 GNDA.n3598 GNDA.n3596 0.0217373
R32372 GNDA.n4169 GNDA.n3601 0.0217373
R32373 GNDA.n3603 GNDA.n3601 0.0217373
R32374 GNDA.n4161 GNDA.n3643 0.0217373
R32375 GNDA.n3645 GNDA.n3643 0.0217373
R32376 GNDA.n4157 GNDA.n3648 0.0217373
R32377 GNDA.n3650 GNDA.n3648 0.0217373
R32378 GNDA.n4153 GNDA.n3653 0.0217373
R32379 GNDA.n3655 GNDA.n3653 0.0217373
R32380 GNDA.n4149 GNDA.n3658 0.0217373
R32381 GNDA.n3660 GNDA.n3658 0.0217373
R32382 GNDA.n3642 GNDA.n3640 0.0217373
R32383 GNDA.n4168 GNDA.n4167 0.0217373
R32384 GNDA.n3398 GNDA.n3397 0.0217373
R32385 GNDA.n3396 GNDA.n3393 0.0217373
R32386 GNDA.n3399 GNDA.n3398 0.0217373
R32387 GNDA.n3308 GNDA.n2031 0.0217373
R32388 GNDA.n3309 GNDA.n3308 0.0217373
R32389 GNDA.n3149 GNDA.n2149 0.0217373
R32390 GNDA.n3150 GNDA.n3149 0.0217373
R32391 GNDA.n3060 GNDA.n2152 0.0217373
R32392 GNDA.n3060 GNDA.n2151 0.0217373
R32393 GNDA.n2157 GNDA.n2155 0.0217373
R32394 GNDA.n2157 GNDA.n2154 0.0217373
R32395 GNDA.n2915 GNDA.n2233 0.0217373
R32396 GNDA.n2916 GNDA.n2915 0.0217373
R32397 GNDA.n2826 GNDA.n2236 0.0217373
R32398 GNDA.n2826 GNDA.n2235 0.0217373
R32399 GNDA.n2241 GNDA.n2239 0.0217373
R32400 GNDA.n2241 GNDA.n2238 0.0217373
R32401 GNDA.n2685 GNDA.n2679 0.0217373
R32402 GNDA.n2822 GNDA.n2237 0.0217373
R32403 GNDA.n2909 GNDA.n2234 0.0217373
R32404 GNDA.n2232 GNDA.n2186 0.0217373
R32405 GNDA.n3056 GNDA.n2153 0.0217373
R32406 GNDA.n3143 GNDA.n2150 0.0217373
R32407 GNDA.n2148 GNDA.n2147 0.0217373
R32408 GNDA.n3294 GNDA.n3293 0.0217373
R32409 GNDA.n2030 GNDA.n2028 0.0217373
R32410 GNDA.n2682 GNDA.n2680 0.0217373
R32411 GNDA.n2680 GNDA.n2679 0.0217373
R32412 GNDA.n2824 GNDA.n2239 0.0217373
R32413 GNDA.n2821 GNDA.n2238 0.0217373
R32414 GNDA.n2823 GNDA.n2822 0.0217373
R32415 GNDA.n2911 GNDA.n2236 0.0217373
R32416 GNDA.n2908 GNDA.n2235 0.0217373
R32417 GNDA.n2910 GNDA.n2909 0.0217373
R32418 GNDA.n2913 GNDA.n2233 0.0217373
R32419 GNDA.n2917 GNDA.n2916 0.0217373
R32420 GNDA.n2914 GNDA.n2186 0.0217373
R32421 GNDA.n3058 GNDA.n2155 0.0217373
R32422 GNDA.n3055 GNDA.n2154 0.0217373
R32423 GNDA.n3057 GNDA.n3056 0.0217373
R32424 GNDA.n3145 GNDA.n2152 0.0217373
R32425 GNDA.n3142 GNDA.n2151 0.0217373
R32426 GNDA.n3144 GNDA.n3143 0.0217373
R32427 GNDA.n3147 GNDA.n2149 0.0217373
R32428 GNDA.n3151 GNDA.n3150 0.0217373
R32429 GNDA.n3148 GNDA.n2147 0.0217373
R32430 GNDA.n3295 GNDA.n3294 0.0217373
R32431 GNDA.n3306 GNDA.n2031 0.0217373
R32432 GNDA.n3310 GNDA.n3309 0.0217373
R32433 GNDA.n3307 GNDA.n2028 0.0217373
R32434 GNDA.n2224 GNDA.n2187 0.0217373
R32435 GNDA.n2228 GNDA.n2187 0.0217373
R32436 GNDA.n2210 GNDA.n2188 0.0217373
R32437 GNDA.n2219 GNDA.n2211 0.0217373
R32438 GNDA.n2223 GNDA.n2222 0.0217373
R32439 GNDA.n2220 GNDA.n2188 0.0217373
R32440 GNDA.n5411 GNDA.n696 0.0217373
R32441 GNDA.n5426 GNDA.n5418 0.0217373
R32442 GNDA.n5431 GNDA.n5430 0.0217373
R32443 GNDA.n5434 GNDA.n5433 0.0217373
R32444 GNDA.n5438 GNDA.n5437 0.0217373
R32445 GNDA.n5429 GNDA.n5418 0.0217373
R32446 GNDA.n5432 GNDA.n5431 0.0217373
R32447 GNDA.n5440 GNDA.n5416 0.0217373
R32448 GNDA.n653 GNDA.n651 0.0217373
R32449 GNDA.n5433 GNDA.n5417 0.0217373
R32450 GNDA.n5437 GNDA.n5417 0.0217373
R32451 GNDA.n658 GNDA.n656 0.0217373
R32452 GNDA.n5448 GNDA.n679 0.0217373
R32453 GNDA.n688 GNDA.n681 0.0217373
R32454 GNDA.n5444 GNDA.n680 0.0217373
R32455 GNDA.n5414 GNDA.n691 0.0217373
R32456 GNDA.n2191 GNDA.n694 0.0217373
R32457 GNDA.n2193 GNDA.n2189 0.0217373
R32458 GNDA.n689 GNDA.n679 0.0217373
R32459 GNDA.n5444 GNDA.n5443 0.0217373
R32460 GNDA.n5416 GNDA.n692 0.0217373
R32461 GNDA.n5415 GNDA.n5414 0.0217373
R32462 GNDA.n696 GNDA.n695 0.0217373
R32463 GNDA.n2192 GNDA.n2191 0.0217373
R32464 GNDA.n2194 GNDA.n2190 0.0217373
R32465 GNDA.n685 GNDA.n683 0.0217373
R32466 GNDA.n683 GNDA.n681 0.0217373
R32467 GNDA.n5489 GNDA.n5488 0.0217373
R32468 GNDA.n5493 GNDA.n659 0.0217373
R32469 GNDA.n5494 GNDA.n5493 0.0217373
R32470 GNDA.n5498 GNDA.n654 0.0217373
R32471 GNDA.n5499 GNDA.n5498 0.0217373
R32472 GNDA.n5502 GNDA.n5501 0.0217373
R32473 GNDA.n5504 GNDA.n648 0.0217373
R32474 GNDA.n3613 GNDA.n3611 0.0217373
R32475 GNDA.n3614 GNDA.n3613 0.0217373
R32476 GNDA.n5487 GNDA.n664 0.0217373
R32477 GNDA.n5490 GNDA.n5489 0.0217373
R32478 GNDA.n5491 GNDA.n659 0.0217373
R32479 GNDA.n5495 GNDA.n5494 0.0217373
R32480 GNDA.n5492 GNDA.n656 0.0217373
R32481 GNDA.n5496 GNDA.n654 0.0217373
R32482 GNDA.n5500 GNDA.n5499 0.0217373
R32483 GNDA.n5497 GNDA.n651 0.0217373
R32484 GNDA.n3611 GNDA.n649 0.0217373
R32485 GNDA.n3612 GNDA.n3610 0.0217373
R32486 GNDA.n5502 GNDA.n646 0.0217373
R32487 GNDA.n648 GNDA.n646 0.0217373
R32488 GNDA.n601 GNDA.n580 0.0217373
R32489 GNDA.n5533 GNDA.n5532 0.0217373
R32490 GNDA.n5539 GNDA.n5538 0.0217373
R32491 GNDA.n5531 GNDA.n29 0.0217373
R32492 GNDA.n5534 GNDA.n5533 0.0217373
R32493 GNDA.n5537 GNDA.n26 0.0217373
R32494 GNDA.n5540 GNDA.n5539 0.0217373
R32495 GNDA.n356 GNDA.n271 0.0217373
R32496 GNDA.n354 GNDA.n271 0.0217373
R32497 GNDA.n269 GNDA.n184 0.0217373
R32498 GNDA.n270 GNDA.n184 0.0217373
R32499 GNDA.n182 GNDA.n98 0.0217373
R32500 GNDA.n183 GNDA.n98 0.0217373
R32501 GNDA.n448 GNDA.n370 0.0217373
R32502 GNDA.n449 GNDA.n448 0.0217373
R32503 GNDA.n444 GNDA.n375 0.0217373
R32504 GNDA.n369 GNDA.n97 0.0217373
R32505 GNDA.n366 GNDA.n365 0.0217373
R32506 GNDA.n362 GNDA.n361 0.0217373
R32507 GNDA.n358 GNDA.n357 0.0217373
R32508 GNDA.n374 GNDA.n373 0.0217373
R32509 GNDA.n375 GNDA.n374 0.0217373
R32510 GNDA.n446 GNDA.n370 0.0217373
R32511 GNDA.n450 GNDA.n449 0.0217373
R32512 GNDA.n447 GNDA.n97 0.0217373
R32513 GNDA.n182 GNDA.n99 0.0217373
R32514 GNDA.n183 GNDA.n181 0.0217373
R32515 GNDA.n367 GNDA.n366 0.0217373
R32516 GNDA.n269 GNDA.n185 0.0217373
R32517 GNDA.n270 GNDA.n268 0.0217373
R32518 GNDA.n363 GNDA.n362 0.0217373
R32519 GNDA.n356 GNDA.n272 0.0217373
R32520 GNDA.n355 GNDA.n354 0.0217373
R32521 GNDA.n359 GNDA.n358 0.0217373
R32522 GNDA.n605 GNDA.n602 0.0217373
R32523 GNDA.n606 GNDA.n605 0.0217373
R32524 GNDA.n608 GNDA.n43 0.0217373
R32525 GNDA.n611 GNDA.n44 0.0217373
R32526 GNDA.n603 GNDA.n602 0.0217373
R32527 GNDA.n607 GNDA.n606 0.0217373
R32528 GNDA.n604 GNDA.n580 0.0217373
R32529 GNDA.n579 GNDA.n43 0.0217373
R32530 GNDA.n579 GNDA.n44 0.0217373
R32531 GNDA.n4912 GNDA.n947 0.0217373
R32532 GNDA.n4905 GNDA.n4904 0.0217373
R32533 GNDA.n4908 GNDA.n948 0.0217373
R32534 GNDA.n4903 GNDA.n949 0.0217373
R32535 GNDA.n4906 GNDA.n4905 0.0217373
R32536 GNDA.n4907 GNDA.n947 0.0217373
R32537 GNDA.n2215 GNDA.n2213 0.0217373
R32538 GNDA.n2216 GNDA.n2214 0.0217373
R32539 GNDA.n3631 GNDA.n3629 0.0217373
R32540 GNDA.n3632 GNDA.n3630 0.0217373
R32541 GNDA.n3638 GNDA.n3637 0.0217373
R32542 GNDA.n3637 GNDA.n3627 0.0217373
R32543 GNDA.n5053 GNDA.n5051 0.0217373
R32544 GNDA.n5149 GNDA.n5052 0.0217373
R32545 GNDA.n5150 GNDA.n5149 0.0217373
R32546 GNDA.n5064 GNDA.n5051 0.0217373
R32547 GNDA.n5152 GNDA.n5048 0.0217373
R32548 GNDA.n766 GNDA.n764 0.0217373
R32549 GNDA.n5049 GNDA.n5048 0.0217373
R32550 GNDA.n5322 GNDA.n765 0.0217373
R32551 GNDA.n5323 GNDA.n5322 0.0217373
R32552 GNDA.n5319 GNDA.n764 0.0217373
R32553 GNDA.n4886 GNDA.n1108 0.0217373
R32554 GNDA.n4889 GNDA.n1108 0.0217373
R32555 GNDA.n3396 GNDA.n3394 0.0217373
R32556 GNDA.n4185 GNDA.n1973 0.0217373
R32557 GNDA.n4180 GNDA.n3512 0.0217373
R32558 GNDA.n4176 GNDA.n3597 0.0217373
R32559 GNDA.n4172 GNDA.n3602 0.0217373
R32560 GNDA.n4164 GNDA.n3644 0.0217373
R32561 GNDA.n4160 GNDA.n3649 0.0217373
R32562 GNDA.n4156 GNDA.n3654 0.0217373
R32563 GNDA.n4152 GNDA.n3659 0.0217373
R32564 GNDA.n3595 GNDA.n3512 0.0217373
R32565 GNDA.n3600 GNDA.n3597 0.0217373
R32566 GNDA.n3605 GNDA.n3602 0.0217373
R32567 GNDA.n4185 GNDA.n3510 0.0217373
R32568 GNDA.n3647 GNDA.n3644 0.0217373
R32569 GNDA.n3652 GNDA.n3649 0.0217373
R32570 GNDA.n3657 GNDA.n3654 0.0217373
R32571 GNDA.n4148 GNDA.n3659 0.0217373
R32572 GNDA.n3397 GNDA.n3395 0.0217373
R32573 GNDA.n2684 GNDA.n2683 0.0217373
R32574 GNDA.n2230 GNDA.n2226 0.0217373
R32575 GNDA.n2683 GNDA.n2681 0.0217373
R32576 GNDA.n2227 GNDA.n2226 0.0217373
R32577 GNDA.n2197 GNDA.n2190 0.0217373
R32578 GNDA.n695 GNDA.n693 0.0217373
R32579 GNDA.n5429 GNDA.n5428 0.0217373
R32580 GNDA.n5430 GNDA.n5427 0.0217373
R32581 GNDA.n5428 GNDA.n5422 0.0217373
R32582 GNDA.n692 GNDA.n690 0.0217373
R32583 GNDA.n5439 GNDA.n5435 0.0217373
R32584 GNDA.n5436 GNDA.n5435 0.0217373
R32585 GNDA.n5445 GNDA.n689 0.0217373
R32586 GNDA.n5447 GNDA.n680 0.0217373
R32587 GNDA.n5441 GNDA.n691 0.0217373
R32588 GNDA.n5412 GNDA.n694 0.0217373
R32589 GNDA.n2195 GNDA.n2193 0.0217373
R32590 GNDA.n5447 GNDA.n5446 0.0217373
R32591 GNDA.n5442 GNDA.n5441 0.0217373
R32592 GNDA.n5413 GNDA.n5412 0.0217373
R32593 GNDA.n2196 GNDA.n2195 0.0217373
R32594 GNDA.n2198 GNDA.n2197 0.0217373
R32595 GNDA.n687 GNDA.n686 0.0217373
R32596 GNDA.n5487 GNDA.n5486 0.0217373
R32597 GNDA.n686 GNDA.n684 0.0217373
R32598 GNDA.n5488 GNDA.n5485 0.0217373
R32599 GNDA.n5486 GNDA.n5484 0.0217373
R32600 GNDA.n5505 GNDA.n647 0.0217373
R32601 GNDA.n650 GNDA.n647 0.0217373
R32602 GNDA.n5537 GNDA.n5536 0.0217373
R32603 GNDA.n5531 GNDA.n5530 0.0217373
R32604 GNDA.n5532 GNDA.n5529 0.0217373
R32605 GNDA.n5538 GNDA.n28 0.0217373
R32606 GNDA.n5530 GNDA.n5528 0.0217373
R32607 GNDA.n5535 GNDA.n28 0.0217373
R32608 GNDA.n5536 GNDA.n27 0.0217373
R32609 GNDA.n372 GNDA.n45 0.0217373
R32610 GNDA.n372 GNDA.n371 0.0217373
R32611 GNDA.n610 GNDA.n609 0.0217373
R32612 GNDA.n609 GNDA.n42 0.0217373
R32613 GNDA.n4909 GNDA.n4907 0.0217373
R32614 GNDA.n4903 GNDA.n950 0.0217373
R32615 GNDA.n4904 GNDA.n4902 0.0217373
R32616 GNDA.n4911 GNDA.n948 0.0217373
R32617 GNDA.n4902 GNDA.n4901 0.0217373
R32618 GNDA.n4911 GNDA.n4910 0.0217373
R32619 GNDA.n4188 GNDA.n3509 0.0181756
R32620 GNDA.n4186 GNDA.n4184 0.0181756
R32621 GNDA.n4184 GNDA.n3509 0.0181756
R32622 GNDA.n3290 GNDA.n2117 0.0181756
R32623 GNDA.n3291 GNDA.n2117 0.0181756
R32624 GNDA.n3290 GNDA.n2118 0.0181756
R32625 GNDA.n3291 GNDA.n3289 0.0181756
R32626 GNDA.n2817 GNDA.n2741 0.0107812
R32627 GNDA.n2817 GNDA.n2161 0.0107812
R32628 GNDA.n2975 GNDA.n2161 0.0107812
R32629 GNDA.n3051 GNDA.n2975 0.0107812
R32630 GNDA.n3051 GNDA.n2122 0.0107812
R32631 GNDA.n3209 GNDA.n2122 0.0107812
R32632 GNDA.n3285 GNDA.n3209 0.0107812
R32633 GNDA.n3285 GNDA.n2003 0.0107812
R32634 GNDA.n3368 GNDA.n2003 0.0107812
R32635 GNDA.n4237 GNDA.n3457 0.0107812
R32636 GNDA.n4237 GNDA.n4236 0.0107812
R32637 GNDA.n4236 GNDA.n3486 0.0107812
R32638 GNDA.n3770 GNDA.n3486 0.0107812
R32639 GNDA.n3851 GNDA.n3770 0.0107812
R32640 GNDA.n3932 GNDA.n3851 0.0107812
R32641 GNDA.n4013 GNDA.n3932 0.0107812
R32642 GNDA.n4094 GNDA.n4013 0.0107812
R32643 GNDA.n4111 GNDA.n4094 0.0107812
R32644 GNDA.n574 GNDA.n509 0.0107812
R32645 GNDA.n509 GNDA.n508 0.0107812
R32646 GNDA.n508 GNDA.n84 0.0107812
R32647 GNDA.n264 GNDA.n84 0.0107812
R32648 GNDA.n264 GNDA.n0 0.0107812
R32649 GNDA.n5599 GNDA.n0 0.0107812
R32650 GNDA.n2651 GNDA.n2342 0.00182188
R32651 GNDA.n2649 GNDA.n2648 0.00182188
R32652 GNDA.n2543 GNDA.n2474 0.00182188
R32653 GNDA.n2610 GNDA.n2376 0.00182188
R32654 GNDA.n2649 GNDA.n2325 0.00166081
R32655 GNDA.n2648 GNDA.n2617 0.00166081
R32656 GNDA.n2323 GNDA.n2280 0.00166081
R32657 GNDA.n2618 GNDA.n2280 0.00166081
R32658 GNDA.n2321 GNDA.n2281 0.00166081
R32659 GNDA.n2619 GNDA.n2281 0.00166081
R32660 GNDA.n2319 GNDA.n2282 0.00166081
R32661 GNDA.n2620 GNDA.n2282 0.00166081
R32662 GNDA.n2317 GNDA.n2283 0.00166081
R32663 GNDA.n2621 GNDA.n2283 0.00166081
R32664 GNDA.n2315 GNDA.n2284 0.00166081
R32665 GNDA.n2622 GNDA.n2284 0.00166081
R32666 GNDA.n2313 GNDA.n2285 0.00166081
R32667 GNDA.n2623 GNDA.n2285 0.00166081
R32668 GNDA.n2311 GNDA.n2286 0.00166081
R32669 GNDA.n2624 GNDA.n2286 0.00166081
R32670 GNDA.n2309 GNDA.n2287 0.00166081
R32671 GNDA.n2625 GNDA.n2287 0.00166081
R32672 GNDA.n2307 GNDA.n2288 0.00166081
R32673 GNDA.n2626 GNDA.n2288 0.00166081
R32674 GNDA.n2305 GNDA.n2289 0.00166081
R32675 GNDA.n2627 GNDA.n2289 0.00166081
R32676 GNDA.n2303 GNDA.n2290 0.00166081
R32677 GNDA.n2628 GNDA.n2290 0.00166081
R32678 GNDA.n2301 GNDA.n2291 0.00166081
R32679 GNDA.n2629 GNDA.n2291 0.00166081
R32680 GNDA.n2299 GNDA.n2292 0.00166081
R32681 GNDA.n2630 GNDA.n2292 0.00166081
R32682 GNDA.n2297 GNDA.n2293 0.00166081
R32683 GNDA.n2631 GNDA.n2293 0.00166081
R32684 GNDA.n2295 GNDA.n2294 0.00166081
R32685 GNDA.n2294 GNDA.n2262 0.00166081
R32686 GNDA.n2475 GNDA.n2474 0.00166081
R32687 GNDA.n2458 GNDA.n2410 0.00166081
R32688 GNDA.n2476 GNDA.n2410 0.00166081
R32689 GNDA.n2459 GNDA.n2411 0.00166081
R32690 GNDA.n2477 GNDA.n2411 0.00166081
R32691 GNDA.n2460 GNDA.n2412 0.00166081
R32692 GNDA.n2478 GNDA.n2412 0.00166081
R32693 GNDA.n2461 GNDA.n2413 0.00166081
R32694 GNDA.n2479 GNDA.n2413 0.00166081
R32695 GNDA.n2462 GNDA.n2414 0.00166081
R32696 GNDA.n2480 GNDA.n2414 0.00166081
R32697 GNDA.n2463 GNDA.n2415 0.00166081
R32698 GNDA.n2481 GNDA.n2415 0.00166081
R32699 GNDA.n2464 GNDA.n2416 0.00166081
R32700 GNDA.n2482 GNDA.n2416 0.00166081
R32701 GNDA.n2465 GNDA.n2417 0.00166081
R32702 GNDA.n2483 GNDA.n2417 0.00166081
R32703 GNDA.n2466 GNDA.n2418 0.00166081
R32704 GNDA.n2484 GNDA.n2418 0.00166081
R32705 GNDA.n2467 GNDA.n2419 0.00166081
R32706 GNDA.n2485 GNDA.n2419 0.00166081
R32707 GNDA.n2468 GNDA.n2420 0.00166081
R32708 GNDA.n2486 GNDA.n2420 0.00166081
R32709 GNDA.n2469 GNDA.n2421 0.00166081
R32710 GNDA.n2487 GNDA.n2421 0.00166081
R32711 GNDA.n2470 GNDA.n2422 0.00166081
R32712 GNDA.n2488 GNDA.n2422 0.00166081
R32713 GNDA.n2471 GNDA.n2423 0.00166081
R32714 GNDA.n2489 GNDA.n2423 0.00166081
R32715 GNDA.n2472 GNDA.n2424 0.00166081
R32716 GNDA.n2490 GNDA.n2424 0.00166081
R32717 GNDA.n2540 GNDA.n2539 0.00166081
R32718 GNDA.n2425 GNDA.n954 0.00166081
R32719 GNDA.n2491 GNDA.n2473 0.00166081
R32720 GNDA.n2495 GNDA.n2493 0.00166081
R32721 GNDA.n2494 GNDA.n2457 0.00166081
R32722 GNDA.n2498 GNDA.n2496 0.00166081
R32723 GNDA.n2497 GNDA.n2456 0.00166081
R32724 GNDA.n2501 GNDA.n2499 0.00166081
R32725 GNDA.n2500 GNDA.n2455 0.00166081
R32726 GNDA.n2504 GNDA.n2502 0.00166081
R32727 GNDA.n2503 GNDA.n2454 0.00166081
R32728 GNDA.n2507 GNDA.n2505 0.00166081
R32729 GNDA.n2506 GNDA.n2453 0.00166081
R32730 GNDA.n2510 GNDA.n2508 0.00166081
R32731 GNDA.n2509 GNDA.n2452 0.00166081
R32732 GNDA.n2513 GNDA.n2511 0.00166081
R32733 GNDA.n2512 GNDA.n2451 0.00166081
R32734 GNDA.n2516 GNDA.n2514 0.00166081
R32735 GNDA.n2515 GNDA.n2450 0.00166081
R32736 GNDA.n2519 GNDA.n2517 0.00166081
R32737 GNDA.n2518 GNDA.n2449 0.00166081
R32738 GNDA.n2522 GNDA.n2520 0.00166081
R32739 GNDA.n2521 GNDA.n2448 0.00166081
R32740 GNDA.n2525 GNDA.n2523 0.00166081
R32741 GNDA.n2524 GNDA.n2447 0.00166081
R32742 GNDA.n2528 GNDA.n2526 0.00166081
R32743 GNDA.n2527 GNDA.n2446 0.00166081
R32744 GNDA.n2531 GNDA.n2529 0.00166081
R32745 GNDA.n2530 GNDA.n2445 0.00166081
R32746 GNDA.n2534 GNDA.n2532 0.00166081
R32747 GNDA.n2533 GNDA.n2444 0.00166081
R32748 GNDA.n2537 GNDA.n2535 0.00166081
R32749 GNDA.n2536 GNDA.n2443 0.00166081
R32750 GNDA.n2542 GNDA.n2538 0.00166081
R32751 GNDA.n2541 GNDA.n2442 0.00166081
R32752 GNDA.n2544 GNDA.n2409 0.00166081
R32753 GNDA.n2562 GNDA.n2561 0.00166081
R32754 GNDA.n2595 GNDA.n2566 0.00166081
R32755 GNDA.n2564 GNDA.n2392 0.00166081
R32756 GNDA.n2596 GNDA.n2568 0.00166081
R32757 GNDA.n2567 GNDA.n2391 0.00166081
R32758 GNDA.n2597 GNDA.n2570 0.00166081
R32759 GNDA.n2569 GNDA.n2390 0.00166081
R32760 GNDA.n2598 GNDA.n2572 0.00166081
R32761 GNDA.n2571 GNDA.n2389 0.00166081
R32762 GNDA.n2599 GNDA.n2574 0.00166081
R32763 GNDA.n2573 GNDA.n2388 0.00166081
R32764 GNDA.n2600 GNDA.n2576 0.00166081
R32765 GNDA.n2575 GNDA.n2387 0.00166081
R32766 GNDA.n2601 GNDA.n2578 0.00166081
R32767 GNDA.n2577 GNDA.n2386 0.00166081
R32768 GNDA.n2602 GNDA.n2580 0.00166081
R32769 GNDA.n2579 GNDA.n2385 0.00166081
R32770 GNDA.n2603 GNDA.n2582 0.00166081
R32771 GNDA.n2581 GNDA.n2384 0.00166081
R32772 GNDA.n2604 GNDA.n2584 0.00166081
R32773 GNDA.n2583 GNDA.n2383 0.00166081
R32774 GNDA.n2605 GNDA.n2586 0.00166081
R32775 GNDA.n2585 GNDA.n2382 0.00166081
R32776 GNDA.n2606 GNDA.n2588 0.00166081
R32777 GNDA.n2587 GNDA.n2381 0.00166081
R32778 GNDA.n2607 GNDA.n2590 0.00166081
R32779 GNDA.n2589 GNDA.n2380 0.00166081
R32780 GNDA.n2608 GNDA.n2592 0.00166081
R32781 GNDA.n2591 GNDA.n2379 0.00166081
R32782 GNDA.n2609 GNDA.n2594 0.00166081
R32783 GNDA.n2593 GNDA.n2378 0.00166081
R32784 GNDA.n2613 GNDA.n2611 0.00166081
R32785 GNDA.n2612 GNDA.n2377 0.00166081
R32786 GNDA.n2615 GNDA.n2343 0.00166081
R32787 GNDA.n2616 GNDA.n2261 0.00166081
R32788 GNDA.n2632 GNDA.n2263 0.00166081
R32789 GNDA.n2341 GNDA.n2260 0.00166081
R32790 GNDA.n2633 GNDA.n2264 0.00166081
R32791 GNDA.n2340 GNDA.n2259 0.00166081
R32792 GNDA.n2634 GNDA.n2265 0.00166081
R32793 GNDA.n2339 GNDA.n2258 0.00166081
R32794 GNDA.n2635 GNDA.n2266 0.00166081
R32795 GNDA.n2338 GNDA.n2257 0.00166081
R32796 GNDA.n2636 GNDA.n2267 0.00166081
R32797 GNDA.n2337 GNDA.n2256 0.00166081
R32798 GNDA.n2637 GNDA.n2268 0.00166081
R32799 GNDA.n2336 GNDA.n2255 0.00166081
R32800 GNDA.n2638 GNDA.n2269 0.00166081
R32801 GNDA.n2335 GNDA.n2254 0.00166081
R32802 GNDA.n2639 GNDA.n2270 0.00166081
R32803 GNDA.n2334 GNDA.n2253 0.00166081
R32804 GNDA.n2640 GNDA.n2271 0.00166081
R32805 GNDA.n2333 GNDA.n2252 0.00166081
R32806 GNDA.n2641 GNDA.n2272 0.00166081
R32807 GNDA.n2332 GNDA.n2251 0.00166081
R32808 GNDA.n2642 GNDA.n2273 0.00166081
R32809 GNDA.n2331 GNDA.n2250 0.00166081
R32810 GNDA.n2643 GNDA.n2274 0.00166081
R32811 GNDA.n2330 GNDA.n2249 0.00166081
R32812 GNDA.n2644 GNDA.n2275 0.00166081
R32813 GNDA.n2329 GNDA.n2248 0.00166081
R32814 GNDA.n2645 GNDA.n2276 0.00166081
R32815 GNDA.n2328 GNDA.n2247 0.00166081
R32816 GNDA.n2646 GNDA.n2277 0.00166081
R32817 GNDA.n2327 GNDA.n2246 0.00166081
R32818 GNDA.n2647 GNDA.n2278 0.00166081
R32819 GNDA.n2326 GNDA.n2245 0.00166081
R32820 GNDA.n2652 GNDA.n2279 0.00166081
R32821 GNDA.n2492 GNDA.n2491 0.00166081
R32822 GNDA.n2490 GNDA.n2426 0.00166081
R32823 GNDA.n2489 GNDA.n2427 0.00166081
R32824 GNDA.n2488 GNDA.n2428 0.00166081
R32825 GNDA.n2487 GNDA.n2429 0.00166081
R32826 GNDA.n2486 GNDA.n2430 0.00166081
R32827 GNDA.n2485 GNDA.n2431 0.00166081
R32828 GNDA.n2484 GNDA.n2432 0.00166081
R32829 GNDA.n2483 GNDA.n2433 0.00166081
R32830 GNDA.n2482 GNDA.n2434 0.00166081
R32831 GNDA.n2481 GNDA.n2435 0.00166081
R32832 GNDA.n2480 GNDA.n2436 0.00166081
R32833 GNDA.n2479 GNDA.n2437 0.00166081
R32834 GNDA.n2478 GNDA.n2438 0.00166081
R32835 GNDA.n2477 GNDA.n2439 0.00166081
R32836 GNDA.n2476 GNDA.n2440 0.00166081
R32837 GNDA.n2475 GNDA.n2441 0.00166081
R32838 GNDA.n2539 GNDA.n2426 0.00166081
R32839 GNDA.n2472 GNDA.n2427 0.00166081
R32840 GNDA.n2471 GNDA.n2428 0.00166081
R32841 GNDA.n2470 GNDA.n2429 0.00166081
R32842 GNDA.n2469 GNDA.n2430 0.00166081
R32843 GNDA.n2468 GNDA.n2431 0.00166081
R32844 GNDA.n2467 GNDA.n2432 0.00166081
R32845 GNDA.n2466 GNDA.n2433 0.00166081
R32846 GNDA.n2465 GNDA.n2434 0.00166081
R32847 GNDA.n2464 GNDA.n2435 0.00166081
R32848 GNDA.n2463 GNDA.n2436 0.00166081
R32849 GNDA.n2462 GNDA.n2437 0.00166081
R32850 GNDA.n2461 GNDA.n2438 0.00166081
R32851 GNDA.n2460 GNDA.n2439 0.00166081
R32852 GNDA.n2459 GNDA.n2440 0.00166081
R32853 GNDA.n2458 GNDA.n2441 0.00166081
R32854 GNDA.n2493 GNDA.n2473 0.00166081
R32855 GNDA.n2495 GNDA.n2494 0.00166081
R32856 GNDA.n2496 GNDA.n2457 0.00166081
R32857 GNDA.n2498 GNDA.n2497 0.00166081
R32858 GNDA.n2499 GNDA.n2456 0.00166081
R32859 GNDA.n2501 GNDA.n2500 0.00166081
R32860 GNDA.n2502 GNDA.n2455 0.00166081
R32861 GNDA.n2504 GNDA.n2503 0.00166081
R32862 GNDA.n2505 GNDA.n2454 0.00166081
R32863 GNDA.n2507 GNDA.n2506 0.00166081
R32864 GNDA.n2508 GNDA.n2453 0.00166081
R32865 GNDA.n2510 GNDA.n2509 0.00166081
R32866 GNDA.n2511 GNDA.n2452 0.00166081
R32867 GNDA.n2513 GNDA.n2512 0.00166081
R32868 GNDA.n2514 GNDA.n2451 0.00166081
R32869 GNDA.n2516 GNDA.n2515 0.00166081
R32870 GNDA.n2517 GNDA.n2450 0.00166081
R32871 GNDA.n2519 GNDA.n2518 0.00166081
R32872 GNDA.n2520 GNDA.n2449 0.00166081
R32873 GNDA.n2522 GNDA.n2521 0.00166081
R32874 GNDA.n2523 GNDA.n2448 0.00166081
R32875 GNDA.n2525 GNDA.n2524 0.00166081
R32876 GNDA.n2526 GNDA.n2447 0.00166081
R32877 GNDA.n2528 GNDA.n2527 0.00166081
R32878 GNDA.n2529 GNDA.n2446 0.00166081
R32879 GNDA.n2531 GNDA.n2530 0.00166081
R32880 GNDA.n2532 GNDA.n2445 0.00166081
R32881 GNDA.n2534 GNDA.n2533 0.00166081
R32882 GNDA.n2535 GNDA.n2444 0.00166081
R32883 GNDA.n2537 GNDA.n2536 0.00166081
R32884 GNDA.n2538 GNDA.n2443 0.00166081
R32885 GNDA.n2542 GNDA.n2541 0.00166081
R32886 GNDA.n2442 GNDA.n2409 0.00166081
R32887 GNDA.n2540 GNDA.n2425 0.00166081
R32888 GNDA.n2653 GNDA.n2262 0.00166081
R32889 GNDA.n2631 GNDA.n2296 0.00166081
R32890 GNDA.n2630 GNDA.n2298 0.00166081
R32891 GNDA.n2629 GNDA.n2300 0.00166081
R32892 GNDA.n2628 GNDA.n2302 0.00166081
R32893 GNDA.n2627 GNDA.n2304 0.00166081
R32894 GNDA.n2626 GNDA.n2306 0.00166081
R32895 GNDA.n2625 GNDA.n2308 0.00166081
R32896 GNDA.n2624 GNDA.n2310 0.00166081
R32897 GNDA.n2623 GNDA.n2312 0.00166081
R32898 GNDA.n2622 GNDA.n2314 0.00166081
R32899 GNDA.n2621 GNDA.n2316 0.00166081
R32900 GNDA.n2620 GNDA.n2318 0.00166081
R32901 GNDA.n2619 GNDA.n2320 0.00166081
R32902 GNDA.n2618 GNDA.n2322 0.00166081
R32903 GNDA.n2617 GNDA.n2324 0.00166081
R32904 GNDA.n2650 GNDA.n2616 0.00166081
R32905 GNDA.n2296 GNDA.n2295 0.00166081
R32906 GNDA.n2298 GNDA.n2297 0.00166081
R32907 GNDA.n2300 GNDA.n2299 0.00166081
R32908 GNDA.n2302 GNDA.n2301 0.00166081
R32909 GNDA.n2304 GNDA.n2303 0.00166081
R32910 GNDA.n2306 GNDA.n2305 0.00166081
R32911 GNDA.n2308 GNDA.n2307 0.00166081
R32912 GNDA.n2310 GNDA.n2309 0.00166081
R32913 GNDA.n2312 GNDA.n2311 0.00166081
R32914 GNDA.n2314 GNDA.n2313 0.00166081
R32915 GNDA.n2316 GNDA.n2315 0.00166081
R32916 GNDA.n2318 GNDA.n2317 0.00166081
R32917 GNDA.n2320 GNDA.n2319 0.00166081
R32918 GNDA.n2322 GNDA.n2321 0.00166081
R32919 GNDA.n2324 GNDA.n2323 0.00166081
R32920 GNDA.n2632 GNDA.n2261 0.00166081
R32921 GNDA.n2341 GNDA.n2263 0.00166081
R32922 GNDA.n2633 GNDA.n2260 0.00166081
R32923 GNDA.n2340 GNDA.n2264 0.00166081
R32924 GNDA.n2634 GNDA.n2259 0.00166081
R32925 GNDA.n2339 GNDA.n2265 0.00166081
R32926 GNDA.n2635 GNDA.n2258 0.00166081
R32927 GNDA.n2338 GNDA.n2266 0.00166081
R32928 GNDA.n2636 GNDA.n2257 0.00166081
R32929 GNDA.n2337 GNDA.n2267 0.00166081
R32930 GNDA.n2637 GNDA.n2256 0.00166081
R32931 GNDA.n2336 GNDA.n2268 0.00166081
R32932 GNDA.n2638 GNDA.n2255 0.00166081
R32933 GNDA.n2335 GNDA.n2269 0.00166081
R32934 GNDA.n2639 GNDA.n2254 0.00166081
R32935 GNDA.n2334 GNDA.n2270 0.00166081
R32936 GNDA.n2640 GNDA.n2253 0.00166081
R32937 GNDA.n2333 GNDA.n2271 0.00166081
R32938 GNDA.n2641 GNDA.n2252 0.00166081
R32939 GNDA.n2332 GNDA.n2272 0.00166081
R32940 GNDA.n2642 GNDA.n2251 0.00166081
R32941 GNDA.n2331 GNDA.n2273 0.00166081
R32942 GNDA.n2643 GNDA.n2250 0.00166081
R32943 GNDA.n2330 GNDA.n2274 0.00166081
R32944 GNDA.n2644 GNDA.n2249 0.00166081
R32945 GNDA.n2329 GNDA.n2275 0.00166081
R32946 GNDA.n2645 GNDA.n2248 0.00166081
R32947 GNDA.n2328 GNDA.n2276 0.00166081
R32948 GNDA.n2646 GNDA.n2247 0.00166081
R32949 GNDA.n2327 GNDA.n2277 0.00166081
R32950 GNDA.n2647 GNDA.n2246 0.00166081
R32951 GNDA.n2326 GNDA.n2278 0.00166081
R32952 GNDA.n2279 GNDA.n2245 0.00166081
R32953 GNDA.n2342 GNDA.n2325 0.00166081
R32954 GNDA.n2614 GNDA.n2563 0.00166081
R32955 GNDA.n2545 GNDA.n2376 0.00166081
R32956 GNDA.n2393 GNDA.n2344 0.00166081
R32957 GNDA.n2546 GNDA.n2375 0.00166081
R32958 GNDA.n2394 GNDA.n2345 0.00166081
R32959 GNDA.n2547 GNDA.n2374 0.00166081
R32960 GNDA.n2395 GNDA.n2346 0.00166081
R32961 GNDA.n2548 GNDA.n2373 0.00166081
R32962 GNDA.n2396 GNDA.n2347 0.00166081
R32963 GNDA.n2549 GNDA.n2372 0.00166081
R32964 GNDA.n2397 GNDA.n2348 0.00166081
R32965 GNDA.n2550 GNDA.n2371 0.00166081
R32966 GNDA.n2398 GNDA.n2349 0.00166081
R32967 GNDA.n2551 GNDA.n2370 0.00166081
R32968 GNDA.n2399 GNDA.n2350 0.00166081
R32969 GNDA.n2552 GNDA.n2369 0.00166081
R32970 GNDA.n2400 GNDA.n2351 0.00166081
R32971 GNDA.n2553 GNDA.n2368 0.00166081
R32972 GNDA.n2401 GNDA.n2352 0.00166081
R32973 GNDA.n2554 GNDA.n2367 0.00166081
R32974 GNDA.n2402 GNDA.n2353 0.00166081
R32975 GNDA.n2555 GNDA.n2366 0.00166081
R32976 GNDA.n2403 GNDA.n2354 0.00166081
R32977 GNDA.n2556 GNDA.n2365 0.00166081
R32978 GNDA.n2404 GNDA.n2355 0.00166081
R32979 GNDA.n2557 GNDA.n2364 0.00166081
R32980 GNDA.n2405 GNDA.n2356 0.00166081
R32981 GNDA.n2558 GNDA.n2363 0.00166081
R32982 GNDA.n2406 GNDA.n2357 0.00166081
R32983 GNDA.n2559 GNDA.n2362 0.00166081
R32984 GNDA.n2407 GNDA.n2358 0.00166081
R32985 GNDA.n2560 GNDA.n2361 0.00166081
R32986 GNDA.n2565 GNDA.n2359 0.00166081
R32987 GNDA.n2560 GNDA.n2359 0.00166081
R32988 GNDA.n2559 GNDA.n2358 0.00166081
R32989 GNDA.n2558 GNDA.n2357 0.00166081
R32990 GNDA.n2557 GNDA.n2356 0.00166081
R32991 GNDA.n2556 GNDA.n2355 0.00166081
R32992 GNDA.n2555 GNDA.n2354 0.00166081
R32993 GNDA.n2554 GNDA.n2353 0.00166081
R32994 GNDA.n2553 GNDA.n2352 0.00166081
R32995 GNDA.n2552 GNDA.n2351 0.00166081
R32996 GNDA.n2551 GNDA.n2350 0.00166081
R32997 GNDA.n2550 GNDA.n2349 0.00166081
R32998 GNDA.n2549 GNDA.n2348 0.00166081
R32999 GNDA.n2548 GNDA.n2347 0.00166081
R33000 GNDA.n2547 GNDA.n2346 0.00166081
R33001 GNDA.n2546 GNDA.n2345 0.00166081
R33002 GNDA.n2545 GNDA.n2344 0.00166081
R33003 GNDA.n2610 GNDA.n2563 0.00166081
R33004 GNDA.n2561 GNDA.n2408 0.00166081
R33005 GNDA.n2407 GNDA.n2361 0.00166081
R33006 GNDA.n2406 GNDA.n2362 0.00166081
R33007 GNDA.n2405 GNDA.n2363 0.00166081
R33008 GNDA.n2404 GNDA.n2364 0.00166081
R33009 GNDA.n2403 GNDA.n2365 0.00166081
R33010 GNDA.n2402 GNDA.n2366 0.00166081
R33011 GNDA.n2401 GNDA.n2367 0.00166081
R33012 GNDA.n2400 GNDA.n2368 0.00166081
R33013 GNDA.n2399 GNDA.n2369 0.00166081
R33014 GNDA.n2398 GNDA.n2370 0.00166081
R33015 GNDA.n2397 GNDA.n2371 0.00166081
R33016 GNDA.n2396 GNDA.n2372 0.00166081
R33017 GNDA.n2395 GNDA.n2373 0.00166081
R33018 GNDA.n2394 GNDA.n2374 0.00166081
R33019 GNDA.n2393 GNDA.n2375 0.00166081
R33020 GNDA.n2595 GNDA.n2408 0.00166081
R33021 GNDA.n2565 GNDA.n2360 0.00166081
R33022 GNDA.n2566 GNDA.n2564 0.00166081
R33023 GNDA.n2596 GNDA.n2392 0.00166081
R33024 GNDA.n2568 GNDA.n2567 0.00166081
R33025 GNDA.n2597 GNDA.n2391 0.00166081
R33026 GNDA.n2570 GNDA.n2569 0.00166081
R33027 GNDA.n2598 GNDA.n2390 0.00166081
R33028 GNDA.n2572 GNDA.n2571 0.00166081
R33029 GNDA.n2599 GNDA.n2389 0.00166081
R33030 GNDA.n2574 GNDA.n2573 0.00166081
R33031 GNDA.n2600 GNDA.n2388 0.00166081
R33032 GNDA.n2576 GNDA.n2575 0.00166081
R33033 GNDA.n2601 GNDA.n2387 0.00166081
R33034 GNDA.n2578 GNDA.n2577 0.00166081
R33035 GNDA.n2602 GNDA.n2386 0.00166081
R33036 GNDA.n2580 GNDA.n2579 0.00166081
R33037 GNDA.n2603 GNDA.n2385 0.00166081
R33038 GNDA.n2582 GNDA.n2581 0.00166081
R33039 GNDA.n2604 GNDA.n2384 0.00166081
R33040 GNDA.n2584 GNDA.n2583 0.00166081
R33041 GNDA.n2605 GNDA.n2383 0.00166081
R33042 GNDA.n2586 GNDA.n2585 0.00166081
R33043 GNDA.n2606 GNDA.n2382 0.00166081
R33044 GNDA.n2588 GNDA.n2587 0.00166081
R33045 GNDA.n2607 GNDA.n2381 0.00166081
R33046 GNDA.n2590 GNDA.n2589 0.00166081
R33047 GNDA.n2608 GNDA.n2380 0.00166081
R33048 GNDA.n2592 GNDA.n2591 0.00166081
R33049 GNDA.n2609 GNDA.n2379 0.00166081
R33050 GNDA.n2594 GNDA.n2593 0.00166081
R33051 GNDA.n2611 GNDA.n2378 0.00166081
R33052 GNDA.n2613 GNDA.n2612 0.00166081
R33053 GNDA.n2377 GNDA.n2343 0.00166081
C0 two_stage_opamp_dummy_magic_29_0.Vb1 VDDA 0.743962f
C1 two_stage_opamp_dummy_magic_29_0.Vb1 two_stage_opamp_dummy_magic_29_0.V_tail_gate 3.74348f
C2 two_stage_opamp_dummy_magic_29_0.Y VDDA 7.31689f
C3 bgr_11_0.Vin+ VDDA 1.72765f
C4 bgr_11_0.V_CUR_REF_REG two_stage_opamp_dummy_magic_29_0.Vb1 0.051644f
C5 bgr_11_0.Vin+ two_stage_opamp_dummy_magic_29_0.V_tail_gate 0.014649f
C6 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3 VOUT- 0.014192f
C7 bgr_11_0.Vin+ bgr_11_0.V_CUR_REF_REG 1.57077f
C8 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref two_stage_opamp_dummy_magic_29_0.cap_res_Y 0.143283f
C9 two_stage_opamp_dummy_magic_29_0.Vb1 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage 0.167852f
C10 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref two_stage_opamp_dummy_magic_29_0.V_err_gate 0.804531f
C11 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref two_stage_opamp_dummy_magic_29_0.X 0.010624f
C12 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2 bgr_11_0.1st_Vout_1 1.93991f
C13 two_stage_opamp_dummy_magic_29_0.Vb1 VDDA_2 10.021099f
C14 two_stage_opamp_dummy_magic_29_0.V_source VOUT+ 0.052538f
C15 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref bgr_11_0.START_UP 1.39993f
C16 bgr_11_0.V_TOP VDDA 16.3418f
C17 two_stage_opamp_dummy_magic_29_0.cap_res_X two_stage_opamp_dummy_magic_29_0.V_source 0.073057f
C18 bgr_11_0.V_TOP two_stage_opamp_dummy_magic_29_0.V_tail_gate 0.028061f
C19 bgr_11_0.V_CUR_REF_REG bgr_11_0.V_TOP 0.308375f
C20 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter VDDA 0.023423f
C21 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_11_0.V_CUR_REF_REG 0.779503f
C22 two_stage_opamp_dummy_magic_29_0.V_err_gate two_stage_opamp_dummy_magic_29_0.V_CMFB_S1 0.066208f
C23 two_stage_opamp_dummy_magic_29_0.V_tot VOUT+ 0.210263f
C24 bgr_11_0.Vin+ two_stage_opamp_dummy_magic_29_0.V_CMFB_S2 0.055084f
C25 two_stage_opamp_dummy_magic_29_0.Vb1 VOUT+ 0.068172f
C26 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1 two_stage_opamp_dummy_magic_29_0.X 0.90004f
C27 two_stage_opamp_dummy_magic_29_0.V_source VOUT- 0.054787f
C28 two_stage_opamp_dummy_magic_29_0.Y VOUT+ 3.91972f
C29 two_stage_opamp_dummy_magic_29_0.cap_res_Y VDDA 1.28042f
C30 two_stage_opamp_dummy_magic_29_0.V_err_gate VDDA 2.05908f
C31 two_stage_opamp_dummy_magic_29_0.V_tail_gate two_stage_opamp_dummy_magic_29_0.cap_res_Y 2.02177f
C32 two_stage_opamp_dummy_magic_29_0.V_err_gate two_stage_opamp_dummy_magic_29_0.V_tail_gate 0.271999f
C33 two_stage_opamp_dummy_magic_29_0.Vb1 two_stage_opamp_dummy_magic_29_0.cap_res_X 0.228543f
C34 two_stage_opamp_dummy_magic_29_0.V_tail_gate two_stage_opamp_dummy_magic_29_0.VD1 0.021061f
C35 bgr_11_0.V_CUR_REF_REG two_stage_opamp_dummy_magic_29_0.V_err_gate 0.375039f
C36 two_stage_opamp_dummy_magic_29_0.err_amp_out two_stage_opamp_dummy_magic_29_0.V_source 0.184635f
C37 two_stage_opamp_dummy_magic_29_0.X VDDA 7.32388f
C38 two_stage_opamp_dummy_magic_29_0.V_tail_gate two_stage_opamp_dummy_magic_29_0.VD2 0.02134f
C39 two_stage_opamp_dummy_magic_29_0.VD4 two_stage_opamp_dummy_magic_29_0.Y 7.95637f
C40 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3 two_stage_opamp_dummy_magic_29_0.Vb1 0.010591f
C41 two_stage_opamp_dummy_magic_29_0.V_tot VOUT- 0.210256f
C42 bgr_11_0.START_UP VDDA 2.29037f
C43 bgr_11_0.PFET_GATE_10uA two_stage_opamp_dummy_magic_29_0.Vb1 0.091713f
C44 two_stage_opamp_dummy_magic_29_0.Vb1 VOUT- 0.062068f
C45 two_stage_opamp_dummy_magic_29_0.V_tot two_stage_opamp_dummy_magic_29_0.err_amp_out 3.37378f
C46 two_stage_opamp_dummy_magic_29_0.V_source VIN+ 0.523933f
C47 two_stage_opamp_dummy_magic_29_0.cap_res_Y VDDA_2 0.025574f
C48 bgr_11_0.V_TOP two_stage_opamp_dummy_magic_29_0.V_CMFB_S2 0.230311f
C49 two_stage_opamp_dummy_magic_29_0.Vb1 two_stage_opamp_dummy_magic_29_0.err_amp_out 2.98002f
C50 VIN+ VIN- 0.096614f
C51 two_stage_opamp_dummy_magic_29_0.V_tot VIN+ 0.020171f
C52 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2 two_stage_opamp_dummy_magic_29_0.V_err_gate 0.774203f
C53 two_stage_opamp_dummy_magic_29_0.V_source VIN- 0.524384f
C54 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref VDDA 5.14397f
C55 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref two_stage_opamp_dummy_magic_29_0.V_tail_gate 0.169754f
C56 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2 two_stage_opamp_dummy_magic_29_0.X 1.27179f
C57 two_stage_opamp_dummy_magic_29_0.cap_res_Y VOUT+ 52.8086f
C58 bgr_11_0.PFET_GATE_10uA bgr_11_0.V_TOP 0.198375f
C59 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref bgr_11_0.V_CUR_REF_REG 2.48263f
C60 two_stage_opamp_dummy_magic_29_0.cap_res_Y two_stage_opamp_dummy_magic_29_0.cap_res_X 0.477735f
C61 m2_4090_4530# VDDA 0.012155f
C62 two_stage_opamp_dummy_magic_29_0.V_err_gate two_stage_opamp_dummy_magic_29_0.cap_res_X 0.162955f
C63 two_stage_opamp_dummy_magic_29_0.V_tot two_stage_opamp_dummy_magic_29_0.V_source 0.040248f
C64 two_stage_opamp_dummy_magic_29_0.X two_stage_opamp_dummy_magic_29_0.cap_res_X 0.058941f
C65 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2 bgr_11_0.START_UP 0.011661f
C66 two_stage_opamp_dummy_magic_29_0.VD3 two_stage_opamp_dummy_magic_29_0.X 7.95637f
C67 two_stage_opamp_dummy_magic_29_0.VD4 two_stage_opamp_dummy_magic_29_0.cap_res_Y 0.168036f
C68 two_stage_opamp_dummy_magic_29_0.Vb1 two_stage_opamp_dummy_magic_29_0.V_source 1.30282f
C69 two_stage_opamp_dummy_magic_29_0.V_tot VIN- 0.020171f
C70 bgr_11_0.Vin+ bgr_11_0.1st_Vout_1 0.275724f
C71 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3 two_stage_opamp_dummy_magic_29_0.V_err_gate 0.274513f
C72 two_stage_opamp_dummy_magic_29_0.V_tot two_stage_opamp_dummy_magic_29_0.V_err_mir_p 0.047221f
C73 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref VDDA_2 1.07798f
C74 two_stage_opamp_dummy_magic_29_0.cap_res_Y VOUT- 0.02055f
C75 two_stage_opamp_dummy_magic_29_0.V_err_gate VOUT- 0.022554f
C76 bgr_11_0.START_UP_NFET1 bgr_11_0.START_UP 0.145663f
C77 two_stage_opamp_dummy_magic_29_0.V_err_gate two_stage_opamp_dummy_magic_29_0.err_amp_out 0.068782f
C78 two_stage_opamp_dummy_magic_29_0.X VOUT- 3.91972f
C79 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1 VDDA 4.27737f
C80 two_stage_opamp_dummy_magic_29_0.V_tail_gate two_stage_opamp_dummy_magic_29_0.V_CMFB_S1 0.728199f
C81 two_stage_opamp_dummy_magic_29_0.Vb1 two_stage_opamp_dummy_magic_29_0.V_tot 1.87985f
C82 two_stage_opamp_dummy_magic_29_0.Y two_stage_opamp_dummy_magic_29_0.V_tot 0.803388f
C83 bgr_11_0.V_CUR_REF_REG two_stage_opamp_dummy_magic_29_0.V_CMFB_S1 0.295226f
C84 two_stage_opamp_dummy_magic_29_0.err_amp_out two_stage_opamp_dummy_magic_29_0.X 1.31029f
C85 two_stage_opamp_dummy_magic_29_0.Vb1 two_stage_opamp_dummy_magic_29_0.Y 2.31404f
C86 two_stage_opamp_dummy_magic_29_0.V_tail_gate VDDA 5.07347f
C87 bgr_11_0.V_CUR_REF_REG VDDA 3.22107f
C88 bgr_11_0.V_CUR_REF_REG two_stage_opamp_dummy_magic_29_0.V_tail_gate 0.403953f
C89 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref VOUT+ 0.02251f
C90 bgr_11_0.V_TOP bgr_11_0.1st_Vout_1 2.62306f
C91 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage VDDA 0.015355f
C92 two_stage_opamp_dummy_magic_29_0.V_tail_gate two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage 5.93798f
C93 two_stage_opamp_dummy_magic_29_0.VD2 VIN+ 0.532103f
C94 VDDA VDDA_2 23.9878f
C95 two_stage_opamp_dummy_magic_29_0.V_tail_gate VDDA_2 0.297195f
C96 two_stage_opamp_dummy_magic_29_0.cap_res_Y two_stage_opamp_dummy_magic_29_0.V_source 0.066068f
C97 bgr_11_0.V_CUR_REF_REG VDDA_2 0.611124f
C98 two_stage_opamp_dummy_magic_29_0.VD1 two_stage_opamp_dummy_magic_29_0.V_source 5.0157f
C99 two_stage_opamp_dummy_magic_29_0.V_err_gate bgr_11_0.1st_Vout_1 0.131319f
C100 bgr_11_0.PFET_GATE_10uA two_stage_opamp_dummy_magic_29_0.V_err_amp_ref 0.792332f
C101 bgr_11_0.Vin+ bgr_11_0.V_TOP 1.8967f
C102 two_stage_opamp_dummy_magic_29_0.VD1 VIN- 0.532103f
C103 two_stage_opamp_dummy_magic_29_0.VD2 two_stage_opamp_dummy_magic_29_0.V_source 5.01421f
C104 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1 3.51695f
C105 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref two_stage_opamp_dummy_magic_29_0.err_amp_out 0.158625f
C106 two_stage_opamp_dummy_magic_29_0.V_err_gate two_stage_opamp_dummy_magic_29_0.V_err_mir_p 0.429395f
C107 bgr_11_0.Vin+ bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 1.06291f
C108 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2 VDDA 9.2851f
C109 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2 two_stage_opamp_dummy_magic_29_0.V_tail_gate 0.461222f
C110 two_stage_opamp_dummy_magic_29_0.V_source two_stage_opamp_dummy_magic_29_0.Vb1_2 0.443345f
C111 two_stage_opamp_dummy_magic_29_0.V_err_gate two_stage_opamp_dummy_magic_29_0.V_tot 0.611029f
C112 bgr_11_0.V_CUR_REF_REG two_stage_opamp_dummy_magic_29_0.V_CMFB_S2 0.160792f
C113 two_stage_opamp_dummy_magic_29_0.V_tot two_stage_opamp_dummy_magic_29_0.VD1 0.222452f
C114 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1 two_stage_opamp_dummy_magic_29_0.cap_res_X 1.1249f
C115 bgr_11_0.START_UP bgr_11_0.1st_Vout_1 0.13011f
C116 VDDA VOUT+ 13.9096f
C117 two_stage_opamp_dummy_magic_29_0.Vb1 two_stage_opamp_dummy_magic_29_0.cap_res_Y 0.235025f
C118 two_stage_opamp_dummy_magic_29_0.V_err_gate two_stage_opamp_dummy_magic_29_0.Vb1 1.62727f
C119 two_stage_opamp_dummy_magic_29_0.V_tail_gate VOUT+ 1.55356f
C120 two_stage_opamp_dummy_magic_29_0.V_tot two_stage_opamp_dummy_magic_29_0.X 0.518118f
C121 two_stage_opamp_dummy_magic_29_0.Y two_stage_opamp_dummy_magic_29_0.cap_res_Y 0.058941f
C122 two_stage_opamp_dummy_magic_29_0.Vb1 two_stage_opamp_dummy_magic_29_0.VD1 0.556757f
C123 bgr_11_0.Vin+ two_stage_opamp_dummy_magic_29_0.V_err_gate 0.066808f
C124 two_stage_opamp_dummy_magic_29_0.V_tot two_stage_opamp_dummy_magic_29_0.VD2 0.222452f
C125 two_stage_opamp_dummy_magic_29_0.cap_res_X VDDA 1.32028f
C126 two_stage_opamp_dummy_magic_29_0.V_tail_gate two_stage_opamp_dummy_magic_29_0.cap_res_X 2.02142f
C127 two_stage_opamp_dummy_magic_29_0.Vb1 two_stage_opamp_dummy_magic_29_0.X 2.28638f
C128 two_stage_opamp_dummy_magic_29_0.VD3 VDDA 8.70244f
C129 two_stage_opamp_dummy_magic_29_0.Vb1 two_stage_opamp_dummy_magic_29_0.VD2 0.556757f
C130 two_stage_opamp_dummy_magic_29_0.Y two_stage_opamp_dummy_magic_29_0.X 0.056155f
C131 bgr_11_0.START_UP_NFET1 VDDA 0.18791f
C132 two_stage_opamp_dummy_magic_29_0.Y two_stage_opamp_dummy_magic_29_0.VD2 4.15353f
C133 two_stage_opamp_dummy_magic_29_0.VD4 VDDA 8.70244f
C134 bgr_11_0.PFET_GATE_10uA two_stage_opamp_dummy_magic_29_0.V_CMFB_S1 0.329697f
C135 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage VOUT+ 4.69775f
C136 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1 VOUT- 1.16944f
C137 two_stage_opamp_dummy_magic_29_0.Vb1 two_stage_opamp_dummy_magic_29_0.Vb1_2 2.00615f
C138 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3 VDDA 1.83425f
C139 bgr_11_0.PFET_GATE_10uA VDDA 9.597219f
C140 bgr_11_0.Vin+ bgr_11_0.START_UP 0.170134f
C141 bgr_11_0.PFET_GATE_10uA two_stage_opamp_dummy_magic_29_0.V_tail_gate 0.573668f
C142 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_11_0.V_TOP 0.04106f
C143 VDDA VOUT- 13.919099f
C144 bgr_11_0.PFET_GATE_10uA bgr_11_0.V_CUR_REF_REG 0.344267f
C145 two_stage_opamp_dummy_magic_29_0.V_tail_gate VOUT- 1.55483f
C146 two_stage_opamp_dummy_magic_29_0.err_amp_out VDDA 0.228909f
C147 two_stage_opamp_dummy_magic_29_0.V_tail_gate two_stage_opamp_dummy_magic_29_0.err_amp_out 0.168894f
C148 bgr_11_0.V_TOP two_stage_opamp_dummy_magic_29_0.V_err_gate 0.103375f
C149 m2_4090_4530# m2_4000_4420# 0.065657f
C150 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage VOUT- 4.67194f
C151 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref two_stage_opamp_dummy_magic_29_0.V_err_mir_p 0.047283f
C152 two_stage_opamp_dummy_magic_29_0.err_amp_out two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage 0.328005f
C153 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref two_stage_opamp_dummy_magic_29_0.V_tot 1.21201f
C154 bgr_11_0.PFET_GATE_10uA VDDA_2 0.806656f
C155 two_stage_opamp_dummy_magic_29_0.V_tail_gate VIN+ 0.060774f
C156 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref two_stage_opamp_dummy_magic_29_0.Vb1 2.55536f
C157 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2 two_stage_opamp_dummy_magic_29_0.cap_res_X 1.00943f
C158 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref two_stage_opamp_dummy_magic_29_0.Y 0.043425f
C159 two_stage_opamp_dummy_magic_29_0.VD3 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2 0.421441f
C160 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref bgr_11_0.Vin+ 0.25235f
C161 bgr_11_0.V_TOP bgr_11_0.START_UP 1.37378f
C162 two_stage_opamp_dummy_magic_29_0.cap_res_X VOUT+ 0.02055f
C163 two_stage_opamp_dummy_magic_29_0.X two_stage_opamp_dummy_magic_29_0.VD1 4.15353f
C164 two_stage_opamp_dummy_magic_29_0.VD3 two_stage_opamp_dummy_magic_29_0.cap_res_X 0.167711f
C165 two_stage_opamp_dummy_magic_29_0.VD2 two_stage_opamp_dummy_magic_29_0.VD1 0.068381f
C166 two_stage_opamp_dummy_magic_29_0.VD4 VOUT+ 0.034338f
C167 two_stage_opamp_dummy_magic_29_0.V_tail_gate two_stage_opamp_dummy_magic_29_0.V_source 3.43886f
C168 bgr_11_0.1st_Vout_1 VDDA 2.66764f
C169 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2 VOUT- 0.666476f
C170 two_stage_opamp_dummy_magic_29_0.V_err_gate bgr_11_0.START_UP 0.743841f
C171 two_stage_opamp_dummy_magic_29_0.V_tail_gate VIN- 0.058275f
C172 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3 two_stage_opamp_dummy_magic_29_0.cap_res_X 0.063357f
C173 VOUT+ VOUT- 0.213277f
C174 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1 two_stage_opamp_dummy_magic_29_0.V_tot 0.438905f
C175 two_stage_opamp_dummy_magic_29_0.V_err_mir_p VDDA 0.661231f
C176 two_stage_opamp_dummy_magic_29_0.cap_res_X VOUT- 52.7123f
C177 two_stage_opamp_dummy_magic_29_0.V_source two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage 1.17205f
C178 bgr_11_0.PFET_GATE_10uA bgr_11_0.START_UP_NFET1 0.010791f
C179 two_stage_opamp_dummy_magic_29_0.VD3 VOUT- 0.027349f
C180 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref bgr_11_0.V_TOP 0.939477f
C181 two_stage_opamp_dummy_magic_29_0.V_tot VDDA 0.140302f
C182 two_stage_opamp_dummy_magic_29_0.V_tail_gate two_stage_opamp_dummy_magic_29_0.V_tot 4.4704f
C183 VIN- GNDA_2 2.03908f
C184 VIN+ GNDA_2 2.04027f
C185 VOUT- GNDA_2 27.286724f
C186 VOUT+ GNDA_2 27.276207f
C187 VDDA_2 GNDA_2 85.74283f
C188 VDDA GNDA_2 0.218829p
C189 m2_4000_4420# GNDA_2 0.039661f $ **FLOATING
C190 m2_4090_4530# GNDA_2 0.122312f $ **FLOATING
C191 two_stage_opamp_dummy_magic_29_0.Vb1_2 GNDA_2 2.88117f
C192 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage GNDA_2 10.256769f
C193 two_stage_opamp_dummy_magic_29_0.V_source GNDA_2 25.211973f
C194 two_stage_opamp_dummy_magic_29_0.VD1 GNDA_2 4.927533f
C195 two_stage_opamp_dummy_magic_29_0.VD2 GNDA_2 4.928203f
C196 two_stage_opamp_dummy_magic_29_0.cap_res_X GNDA_2 44.17326f
C197 two_stage_opamp_dummy_magic_29_0.cap_res_Y GNDA_2 44.14844f
C198 two_stage_opamp_dummy_magic_29_0.X GNDA_2 12.037578f
C199 two_stage_opamp_dummy_magic_29_0.err_amp_out GNDA_2 7.38754f
C200 two_stage_opamp_dummy_magic_29_0.V_err_mir_p GNDA_2 0.117954f
C201 two_stage_opamp_dummy_magic_29_0.V_tot GNDA_2 12.801761f
C202 two_stage_opamp_dummy_magic_29_0.Y GNDA_2 12.153778f
C203 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1 GNDA_2 15.270994f
C204 two_stage_opamp_dummy_magic_29_0.V_tail_gate GNDA_2 31.905264f
C205 two_stage_opamp_dummy_magic_29_0.Vb1 GNDA_2 37.60854f
C206 bgr_11_0.1st_Vout_1 GNDA_2 12.002972f
C207 bgr_11_0.START_UP GNDA_2 6.619071f
C208 bgr_11_0.START_UP_NFET1 GNDA_2 5.23862f
C209 two_stage_opamp_dummy_magic_29_0.V_err_gate GNDA_2 10.51149f
C210 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2 GNDA_2 20.303059f
C211 bgr_11_0.V_TOP GNDA_2 11.556623f
C212 bgr_11_0.V_CUR_REF_REG GNDA_2 4.79155f
C213 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter GNDA_2 16.8453f
C214 bgr_11_0.Vin+ GNDA_2 4.646547f
C215 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref GNDA_2 10.617849f
C216 bgr_11_0.PFET_GATE_10uA GNDA_2 8.560524f
C217 two_stage_opamp_dummy_magic_29_0.VD3 GNDA_2 5.799711f
C218 two_stage_opamp_dummy_magic_29_0.VD4 GNDA_2 5.821531f
C219 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3 GNDA_2 2.394186f
C220 bgr_11_0.V_CUR_REF_REG.t3 GNDA_2 0.06039f
C221 bgr_11_0.V_CUR_REF_REG.t0 GNDA_2 0.409222f
C222 bgr_11_0.V_CUR_REF_REG.t1 GNDA_2 0.011813f
C223 bgr_11_0.V_CUR_REF_REG.t2 GNDA_2 0.011813f
C224 bgr_11_0.V_CUR_REF_REG.n0 GNDA_2 0.090497f
C225 bgr_11_0.V_CUR_REF_REG.n1 GNDA_2 4.64964f
C226 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.t1 GNDA_2 0.038831f
C227 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.n0 GNDA_2 0.08326f
C228 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.t3 GNDA_2 0.078001f
C229 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.n1 GNDA_2 0.249488f
C230 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.t2 GNDA_2 0.186912f
C231 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.t9 GNDA_2 0.146604f
C232 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.t5 GNDA_2 0.186912f
C233 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.t7 GNDA_2 0.078001f
C234 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.n2 GNDA_2 0.249488f
C235 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.t4 GNDA_2 0.038831f
C236 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.n3 GNDA_2 0.08202f
C237 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.n4 GNDA_2 0.040176f
C238 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.n5 GNDA_2 0.062249f
C239 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.t10 GNDA_2 0.021928f
C240 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.t6 GNDA_2 0.021928f
C241 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.n6 GNDA_2 0.044856f
C242 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.n7 GNDA_2 0.16213f
C243 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.t0 GNDA_2 0.021928f
C244 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.t8 GNDA_2 0.021928f
C245 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.n8 GNDA_2 0.044856f
C246 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.n9 GNDA_2 0.210199f
C247 VDDA_2.n1 GNDA_2 0.033877f
C248 VDDA_2.n2 GNDA_2 0.033877f
C249 VDDA_2.n3 GNDA_2 0.033877f
C250 VDDA_2.n4 GNDA_2 0.033877f
C251 VDDA_2.n5 GNDA_2 0.033877f
C252 VDDA_2.n6 GNDA_2 0.033877f
C253 VDDA_2.n7 GNDA_2 0.033877f
C254 VDDA_2.n8 GNDA_2 0.033877f
C255 VDDA_2.n9 GNDA_2 0.033877f
C256 VDDA_2.n10 GNDA_2 0.033877f
C257 VDDA_2.n11 GNDA_2 0.033877f
C258 VDDA_2.n12 GNDA_2 0.033877f
C259 VDDA_2.n13 GNDA_2 0.033877f
C260 VDDA_2.n14 GNDA_2 0.033877f
C261 VDDA_2.n15 GNDA_2 0.033877f
C262 VDDA_2.n17 GNDA_2 0.033877f
C263 VDDA_2.n18 GNDA_2 0.033877f
C264 VDDA_2.n19 GNDA_2 0.033877f
C265 VDDA_2.n20 GNDA_2 0.033877f
C266 VDDA_2.n21 GNDA_2 0.033877f
C267 VDDA_2.n22 GNDA_2 0.033877f
C268 VDDA_2.n23 GNDA_2 0.033877f
C269 VDDA_2.n24 GNDA_2 0.033877f
C270 VDDA_2.n25 GNDA_2 0.033877f
C271 VDDA_2.n26 GNDA_2 0.033877f
C272 VDDA_2.n27 GNDA_2 0.033877f
C273 VDDA_2.n28 GNDA_2 0.033877f
C274 VDDA_2.n29 GNDA_2 0.033877f
C275 VDDA_2.n30 GNDA_2 0.033877f
C276 VDDA_2.n31 GNDA_2 0.033877f
C277 VDDA_2.n32 GNDA_2 0.033877f
C278 VDDA_2.n33 GNDA_2 0.06399f
C279 VDDA_2.n74 GNDA_2 0.029614f
C280 VDDA_2.n75 GNDA_2 0.011836f
C281 VDDA_2.n86 GNDA_2 0.060226f
C282 VDDA_2.n161 GNDA_2 0.024947f
C283 VDDA_2.n162 GNDA_2 0.02421f
C284 VDDA_2.n172 GNDA_2 0.013923f
C285 VDDA_2.t1 GNDA_2 0.020475f
C286 VDDA_2.t4 GNDA_2 0.021105f
C287 VDDA_2.n174 GNDA_2 0.014699f
C288 VDDA_2.n184 GNDA_2 0.023695f
C289 VDDA_2.n185 GNDA_2 0.047989f
C290 VDDA_2.n233 GNDA_2 0.010646f
C291 VDDA_2.n236 GNDA_2 15.230701f
C292 VDDA_2.n237 GNDA_2 0.035083f
C293 VDDA_2.n238 GNDA_2 0.035083f
C294 VDDA_2.n239 GNDA_2 0.035083f
C295 VDDA_2.n240 GNDA_2 0.035083f
C296 VDDA_2.n241 GNDA_2 0.035083f
C297 VDDA_2.n242 GNDA_2 0.035083f
C298 VDDA_2.n243 GNDA_2 0.035083f
C299 VDDA_2.n244 GNDA_2 0.035083f
C300 VDDA_2.n245 GNDA_2 0.035083f
C301 VDDA_2.n246 GNDA_2 0.035083f
C302 VDDA_2.n247 GNDA_2 0.035083f
C303 VDDA_2.n248 GNDA_2 0.035083f
C304 VDDA_2.n249 GNDA_2 0.035083f
C305 VDDA_2.n250 GNDA_2 0.035083f
C306 VDDA_2.n251 GNDA_2 0.035083f
C307 VDDA_2.n252 GNDA_2 0.035083f
C308 VDDA_2.n268 GNDA_2 0.038981f
C309 VDDA_2.n269 GNDA_2 0.033877f
C310 VDDA_2.n286 GNDA_2 0.035083f
C311 VDDA_2.n288 GNDA_2 0.035083f
C312 VDDA_2.n290 GNDA_2 0.035083f
C313 VDDA_2.n292 GNDA_2 0.035083f
C314 VDDA_2.n294 GNDA_2 0.035083f
C315 VDDA_2.n296 GNDA_2 0.035083f
C316 VDDA_2.n298 GNDA_2 0.035083f
C317 VDDA_2.n300 GNDA_2 0.035083f
C318 VDDA_2.n302 GNDA_2 0.035083f
C319 VDDA_2.n304 GNDA_2 0.035083f
C320 VDDA_2.n306 GNDA_2 0.035083f
C321 VDDA_2.n308 GNDA_2 0.035083f
C322 VDDA_2.n310 GNDA_2 0.035083f
C323 VDDA_2.n312 GNDA_2 0.035083f
C324 VDDA_2.n314 GNDA_2 0.035083f
C325 VDDA_2.n317 GNDA_2 0.033877f
C326 VDDA_2.n333 GNDA_2 0.041405f
C327 VDDA_2.n335 GNDA_2 0.035083f
C328 VDDA_2.n336 GNDA_2 15.225f
C329 VDDA_2.n337 GNDA_2 0.223168f
C330 bgr_11_0.Vin-.n0 GNDA_2 0.07858f
C331 bgr_11_0.Vin-.n1 GNDA_2 0.088293f
C332 bgr_11_0.Vin-.n2 GNDA_2 0.12735f
C333 bgr_11_0.Vin-.t4 GNDA_2 0.294736f
C334 bgr_11_0.Vin-.t3 GNDA_2 0.030534f
C335 bgr_11_0.Vin-.t0 GNDA_2 0.030534f
C336 bgr_11_0.Vin-.n3 GNDA_2 0.085799f
C337 bgr_11_0.Vin-.t1 GNDA_2 0.030534f
C338 bgr_11_0.Vin-.t2 GNDA_2 0.030534f
C339 bgr_11_0.Vin-.n4 GNDA_2 0.074088f
C340 bgr_11_0.Vin-.n5 GNDA_2 0.633984f
C341 bgr_11_0.Vin-.t7 GNDA_2 0.010178f
C342 bgr_11_0.Vin-.t6 GNDA_2 0.010178f
C343 bgr_11_0.Vin-.n6 GNDA_2 0.031534f
C344 bgr_11_0.Vin-.n7 GNDA_2 0.428495f
C345 bgr_11_0.Vin-.t8 GNDA_2 0.049457f
C346 bgr_11_0.Vin-.n8 GNDA_2 0.623119f
C347 bgr_11_0.Vin-.t5 GNDA_2 0.128901f
C348 bgr_11_0.Vin-.n9 GNDA_2 0.734405f
C349 bgr_11_0.Vin-.n10 GNDA_2 1.36082f
C350 bgr_11_0.Vin-.n11 GNDA_2 0.531118f
C351 bgr_11_0.Vin-.n12 GNDA_2 0.079463f
C352 bgr_11_0.Vin-.n13 GNDA_2 0.13464f
C353 bgr_11_0.Vin-.n14 GNDA_2 0.078726f
C354 bgr_11_0.Vin-.n15 GNDA_2 0.155721f
C355 bgr_11_0.Vin-.n16 GNDA_2 0.155721f
C356 bgr_11_0.Vin-.n17 GNDA_2 -0.303656f
C357 bgr_11_0.Vin-.n18 GNDA_2 0.501878f
C358 bgr_11_0.Vin-.n19 GNDA_2 0.240599f
C359 bgr_11_0.Vin-.n20 GNDA_2 0.454563f
C360 bgr_11_0.Vin-.n21 GNDA_2 0.043263f
C361 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_23.Emitter GNDA_2 0.045912f
C362 bgr_11_0.START_UP.t4 GNDA_2 1.72724f
C363 bgr_11_0.START_UP.t5 GNDA_2 0.045404f
C364 bgr_11_0.START_UP.n0 GNDA_2 1.15615f
C365 bgr_11_0.START_UP.t0 GNDA_2 0.04333f
C366 bgr_11_0.START_UP.t2 GNDA_2 0.04333f
C367 bgr_11_0.START_UP.n1 GNDA_2 0.135247f
C368 bgr_11_0.START_UP.t1 GNDA_2 0.04333f
C369 bgr_11_0.START_UP.t3 GNDA_2 0.04333f
C370 bgr_11_0.START_UP.n2 GNDA_2 0.106737f
C371 bgr_11_0.START_UP.n3 GNDA_2 1.0283f
C372 bgr_11_0.START_UP.t6 GNDA_2 0.016282f
C373 bgr_11_0.START_UP.t7 GNDA_2 0.016282f
C374 bgr_11_0.START_UP.n4 GNDA_2 0.046713f
C375 bgr_11_0.START_UP.n5 GNDA_2 0.477587f
C376 two_stage_opamp_dummy_magic_29_0.VD1.t11 GNDA_2 0.033932f
C377 two_stage_opamp_dummy_magic_29_0.VD1.t18 GNDA_2 0.033932f
C378 two_stage_opamp_dummy_magic_29_0.VD1.n0 GNDA_2 0.075122f
C379 two_stage_opamp_dummy_magic_29_0.VD1.n1 GNDA_2 0.564997f
C380 two_stage_opamp_dummy_magic_29_0.VD1.n2 GNDA_2 0.050916f
C381 two_stage_opamp_dummy_magic_29_0.VD1.n3 GNDA_2 0.222536f
C382 two_stage_opamp_dummy_magic_29_0.VD1.t7 GNDA_2 0.033932f
C383 two_stage_opamp_dummy_magic_29_0.VD1.t4 GNDA_2 0.033932f
C384 two_stage_opamp_dummy_magic_29_0.VD1.n4 GNDA_2 0.073831f
C385 two_stage_opamp_dummy_magic_29_0.VD1.n5 GNDA_2 0.284467f
C386 two_stage_opamp_dummy_magic_29_0.VD1.n6 GNDA_2 0.072163f
C387 two_stage_opamp_dummy_magic_29_0.VD1.t3 GNDA_2 0.033932f
C388 two_stage_opamp_dummy_magic_29_0.VD1.t5 GNDA_2 0.033932f
C389 two_stage_opamp_dummy_magic_29_0.VD1.n7 GNDA_2 0.073831f
C390 two_stage_opamp_dummy_magic_29_0.VD1.n8 GNDA_2 0.292399f
C391 two_stage_opamp_dummy_magic_29_0.VD1.t10 GNDA_2 0.033932f
C392 two_stage_opamp_dummy_magic_29_0.VD1.t15 GNDA_2 0.033932f
C393 two_stage_opamp_dummy_magic_29_0.VD1.n9 GNDA_2 0.075122f
C394 two_stage_opamp_dummy_magic_29_0.VD1.t14 GNDA_2 0.033932f
C395 two_stage_opamp_dummy_magic_29_0.VD1.t19 GNDA_2 0.033932f
C396 two_stage_opamp_dummy_magic_29_0.VD1.n10 GNDA_2 0.075122f
C397 two_stage_opamp_dummy_magic_29_0.VD1.n11 GNDA_2 0.767242f
C398 two_stage_opamp_dummy_magic_29_0.VD1.t13 GNDA_2 0.033932f
C399 two_stage_opamp_dummy_magic_29_0.VD1.t17 GNDA_2 0.033932f
C400 two_stage_opamp_dummy_magic_29_0.VD1.n12 GNDA_2 0.075122f
C401 two_stage_opamp_dummy_magic_29_0.VD1.n13 GNDA_2 0.268181f
C402 two_stage_opamp_dummy_magic_29_0.VD1.t6 GNDA_2 0.033932f
C403 two_stage_opamp_dummy_magic_29_0.VD1.t8 GNDA_2 0.033932f
C404 two_stage_opamp_dummy_magic_29_0.VD1.n14 GNDA_2 0.073831f
C405 two_stage_opamp_dummy_magic_29_0.VD1.n15 GNDA_2 0.292399f
C406 two_stage_opamp_dummy_magic_29_0.VD1.n16 GNDA_2 0.122664f
C407 two_stage_opamp_dummy_magic_29_0.VD1.t20 GNDA_2 0.033932f
C408 two_stage_opamp_dummy_magic_29_0.VD1.t0 GNDA_2 0.033932f
C409 two_stage_opamp_dummy_magic_29_0.VD1.n17 GNDA_2 0.073831f
C410 two_stage_opamp_dummy_magic_29_0.VD1.n18 GNDA_2 0.284467f
C411 two_stage_opamp_dummy_magic_29_0.VD1.n19 GNDA_2 0.050916f
C412 two_stage_opamp_dummy_magic_29_0.VD1.n20 GNDA_2 0.222536f
C413 two_stage_opamp_dummy_magic_29_0.VD1.n21 GNDA_2 0.761461f
C414 two_stage_opamp_dummy_magic_29_0.VD1.n22 GNDA_2 0.114111f
C415 two_stage_opamp_dummy_magic_29_0.VD1.n23 GNDA_2 0.067863f
C416 two_stage_opamp_dummy_magic_29_0.VD1.t12 GNDA_2 0.033932f
C417 two_stage_opamp_dummy_magic_29_0.VD1.t16 GNDA_2 0.033932f
C418 two_stage_opamp_dummy_magic_29_0.VD1.n24 GNDA_2 0.075122f
C419 two_stage_opamp_dummy_magic_29_0.VD1.n25 GNDA_2 0.761461f
C420 two_stage_opamp_dummy_magic_29_0.VD1.n26 GNDA_2 0.114111f
C421 two_stage_opamp_dummy_magic_29_0.VD1.n27 GNDA_2 0.767242f
C422 two_stage_opamp_dummy_magic_29_0.VD1.n28 GNDA_2 0.268181f
C423 two_stage_opamp_dummy_magic_29_0.VD1.n29 GNDA_2 0.050916f
C424 two_stage_opamp_dummy_magic_29_0.VD1.t2 GNDA_2 0.033932f
C425 two_stage_opamp_dummy_magic_29_0.VD1.t21 GNDA_2 0.033932f
C426 two_stage_opamp_dummy_magic_29_0.VD1.n30 GNDA_2 0.073831f
C427 two_stage_opamp_dummy_magic_29_0.VD1.n31 GNDA_2 0.284467f
C428 two_stage_opamp_dummy_magic_29_0.VD1.n32 GNDA_2 0.122664f
C429 two_stage_opamp_dummy_magic_29_0.VD1.n33 GNDA_2 0.072163f
C430 two_stage_opamp_dummy_magic_29_0.VD1.t9 GNDA_2 0.033932f
C431 two_stage_opamp_dummy_magic_29_0.VD1.t1 GNDA_2 0.033932f
C432 two_stage_opamp_dummy_magic_29_0.VD1.n34 GNDA_2 0.073831f
C433 two_stage_opamp_dummy_magic_29_0.VD1.n35 GNDA_2 0.284467f
C434 two_stage_opamp_dummy_magic_29_0.VD1.n36 GNDA_2 0.050916f
C435 two_stage_opamp_dummy_magic_29_0.VD1.n37 GNDA_2 0.039407f
C436 two_stage_opamp_dummy_magic_29_0.err_amp_out.t5 GNDA_2 0.072503f
C437 two_stage_opamp_dummy_magic_29_0.err_amp_out.t4 GNDA_2 0.084623f
C438 two_stage_opamp_dummy_magic_29_0.err_amp_out.n0 GNDA_2 0.280015f
C439 two_stage_opamp_dummy_magic_29_0.err_amp_out.t1 GNDA_2 0.068078f
C440 two_stage_opamp_dummy_magic_29_0.err_amp_out.t3 GNDA_2 0.068078f
C441 two_stage_opamp_dummy_magic_29_0.err_amp_out.n1 GNDA_2 0.220809f
C442 two_stage_opamp_dummy_magic_29_0.err_amp_out.t2 GNDA_2 0.068078f
C443 two_stage_opamp_dummy_magic_29_0.err_amp_out.t0 GNDA_2 0.068078f
C444 two_stage_opamp_dummy_magic_29_0.err_amp_out.n2 GNDA_2 0.22061f
C445 two_stage_opamp_dummy_magic_29_0.err_amp_out.n3 GNDA_2 1.20062f
C446 bgr_11_0.cap_res2.t4 GNDA_2 0.334798f
C447 bgr_11_0.cap_res2.t10 GNDA_2 0.336011f
C448 bgr_11_0.cap_res2.t20 GNDA_2 0.318043f
C449 bgr_11_0.cap_res2.t9 GNDA_2 0.334798f
C450 bgr_11_0.cap_res2.t14 GNDA_2 0.336011f
C451 bgr_11_0.cap_res2.t5 GNDA_2 0.318043f
C452 bgr_11_0.cap_res2.t3 GNDA_2 0.334798f
C453 bgr_11_0.cap_res2.t8 GNDA_2 0.336011f
C454 bgr_11_0.cap_res2.t18 GNDA_2 0.318043f
C455 bgr_11_0.cap_res2.t16 GNDA_2 0.334798f
C456 bgr_11_0.cap_res2.t2 GNDA_2 0.336011f
C457 bgr_11_0.cap_res2.t12 GNDA_2 0.318043f
C458 bgr_11_0.cap_res2.t1 GNDA_2 0.334798f
C459 bgr_11_0.cap_res2.t6 GNDA_2 0.336011f
C460 bgr_11_0.cap_res2.t17 GNDA_2 0.318043f
C461 bgr_11_0.cap_res2.n0 GNDA_2 0.224415f
C462 bgr_11_0.cap_res2.t11 GNDA_2 0.178714f
C463 bgr_11_0.cap_res2.n1 GNDA_2 0.243496f
C464 bgr_11_0.cap_res2.t7 GNDA_2 0.178714f
C465 bgr_11_0.cap_res2.n2 GNDA_2 0.243496f
C466 bgr_11_0.cap_res2.t13 GNDA_2 0.178714f
C467 bgr_11_0.cap_res2.n3 GNDA_2 0.243496f
C468 bgr_11_0.cap_res2.t19 GNDA_2 0.178714f
C469 bgr_11_0.cap_res2.n4 GNDA_2 0.243496f
C470 bgr_11_0.cap_res2.t15 GNDA_2 0.360089f
C471 bgr_11_0.cap_res2.t0 GNDA_2 0.082395f
C472 two_stage_opamp_dummy_magic_29_0.V_tot.t1 GNDA_2 0.164539f
C473 two_stage_opamp_dummy_magic_29_0.V_tot.t3 GNDA_2 0.154461f
C474 two_stage_opamp_dummy_magic_29_0.V_tot.n0 GNDA_2 1.65862f
C475 two_stage_opamp_dummy_magic_29_0.V_tot.t2 GNDA_2 0.164539f
C476 two_stage_opamp_dummy_magic_29_0.V_tot.t0 GNDA_2 0.154461f
C477 two_stage_opamp_dummy_magic_29_0.V_tot.n1 GNDA_2 1.74658f
C478 two_stage_opamp_dummy_magic_29_0.V_tot.t4 GNDA_2 0.046802f
C479 two_stage_opamp_dummy_magic_29_0.V_tot.n2 GNDA_2 1.83779f
C480 two_stage_opamp_dummy_magic_29_0.V_tot.t5 GNDA_2 0.046802f
C481 two_stage_opamp_dummy_magic_29_0.V_tot.n3 GNDA_2 0.322038f
C482 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n0 GNDA_2 6.90355f
C483 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n1 GNDA_2 10.6261f
C484 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n2 GNDA_2 0.160409f
C485 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n3 GNDA_2 6.52288f
C486 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t2 GNDA_2 0.010902f
C487 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t0 GNDA_2 0.010902f
C488 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n4 GNDA_2 0.024129f
C489 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n5 GNDA_2 0.113606f
C490 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t28 GNDA_2 0.019352f
C491 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t17 GNDA_2 0.019352f
C492 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t26 GNDA_2 0.019352f
C493 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t16 GNDA_2 0.019352f
C494 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t25 GNDA_2 0.019352f
C495 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t14 GNDA_2 0.019352f
C496 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t23 GNDA_2 0.019352f
C497 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t27 GNDA_2 0.022587f
C498 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n6 GNDA_2 0.021296f
C499 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n7 GNDA_2 0.013356f
C500 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n8 GNDA_2 0.013356f
C501 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n9 GNDA_2 0.013356f
C502 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n10 GNDA_2 0.013356f
C503 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n11 GNDA_2 0.013356f
C504 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n12 GNDA_2 0.012498f
C505 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n13 GNDA_2 0.011317f
C506 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n14 GNDA_2 0.014537f
C507 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n15 GNDA_2 0.014537f
C508 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n16 GNDA_2 0.026396f
C509 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n17 GNDA_2 0.083229f
C510 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n18 GNDA_2 0.014537f
C511 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n19 GNDA_2 0.159989f
C512 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n20 GNDA_2 0.083229f
C513 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n21 GNDA_2 0.014537f
C514 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n22 GNDA_2 0.160419f
C515 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t3 GNDA_2 0.010902f
C516 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t1 GNDA_2 0.010902f
C517 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n23 GNDA_2 0.024129f
C518 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n24 GNDA_2 0.122073f
C519 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t22 GNDA_2 0.019352f
C520 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t19 GNDA_2 0.019352f
C521 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n25 GNDA_2 0.012498f
C522 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n26 GNDA_2 0.012498f
C523 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t13 GNDA_2 0.019352f
C524 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t30 GNDA_2 0.019352f
C525 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t20 GNDA_2 0.019352f
C526 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t31 GNDA_2 0.019352f
C527 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t21 GNDA_2 0.019352f
C528 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t12 GNDA_2 0.019352f
C529 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t24 GNDA_2 0.019352f
C530 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t15 GNDA_2 0.019352f
C531 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t18 GNDA_2 0.019352f
C532 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t29 GNDA_2 0.022587f
C533 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n27 GNDA_2 0.021296f
C534 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n28 GNDA_2 0.013356f
C535 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n29 GNDA_2 0.013356f
C536 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n30 GNDA_2 0.013356f
C537 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n31 GNDA_2 0.013356f
C538 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n32 GNDA_2 0.013356f
C539 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n33 GNDA_2 0.013356f
C540 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n34 GNDA_2 0.013356f
C541 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n35 GNDA_2 0.012498f
C542 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n36 GNDA_2 0.011317f
C543 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n37 GNDA_2 0.119304f
C544 two_stage_opamp_dummy_magic_29_0.V_source.n0 GNDA_2 0.339486f
C545 two_stage_opamp_dummy_magic_29_0.V_source.n1 GNDA_2 0.304203f
C546 two_stage_opamp_dummy_magic_29_0.V_source.n2 GNDA_2 0.540854f
C547 two_stage_opamp_dummy_magic_29_0.V_source.n3 GNDA_2 0.586883f
C548 two_stage_opamp_dummy_magic_29_0.V_source.t40 GNDA_2 0.021514f
C549 two_stage_opamp_dummy_magic_29_0.V_source.t22 GNDA_2 0.021514f
C550 two_stage_opamp_dummy_magic_29_0.V_source.n4 GNDA_2 0.045993f
C551 two_stage_opamp_dummy_magic_29_0.V_source.n5 GNDA_2 0.199232f
C552 two_stage_opamp_dummy_magic_29_0.V_source.n6 GNDA_2 0.04198f
C553 two_stage_opamp_dummy_magic_29_0.V_source.t21 GNDA_2 0.021514f
C554 two_stage_opamp_dummy_magic_29_0.V_source.t27 GNDA_2 0.021514f
C555 two_stage_opamp_dummy_magic_29_0.V_source.n7 GNDA_2 0.045993f
C556 two_stage_opamp_dummy_magic_29_0.V_source.n8 GNDA_2 0.164071f
C557 two_stage_opamp_dummy_magic_29_0.V_source.n9 GNDA_2 0.153086f
C558 two_stage_opamp_dummy_magic_29_0.V_source.n10 GNDA_2 0.153086f
C559 two_stage_opamp_dummy_magic_29_0.V_source.n11 GNDA_2 0.147729f
C560 two_stage_opamp_dummy_magic_29_0.V_source.n12 GNDA_2 0.069673f
C561 two_stage_opamp_dummy_magic_29_0.V_source.n13 GNDA_2 0.046931f
C562 two_stage_opamp_dummy_magic_29_0.V_source.t15 GNDA_2 0.012908f
C563 two_stage_opamp_dummy_magic_29_0.V_source.t24 GNDA_2 0.012908f
C564 two_stage_opamp_dummy_magic_29_0.V_source.n14 GNDA_2 0.028087f
C565 two_stage_opamp_dummy_magic_29_0.V_source.n15 GNDA_2 0.117879f
C566 two_stage_opamp_dummy_magic_29_0.V_source.t3 GNDA_2 0.012908f
C567 two_stage_opamp_dummy_magic_29_0.V_source.t14 GNDA_2 0.012908f
C568 two_stage_opamp_dummy_magic_29_0.V_source.n16 GNDA_2 0.028087f
C569 two_stage_opamp_dummy_magic_29_0.V_source.n17 GNDA_2 0.113801f
C570 two_stage_opamp_dummy_magic_29_0.V_source.n18 GNDA_2 0.069673f
C571 two_stage_opamp_dummy_magic_29_0.V_source.n19 GNDA_2 0.054121f
C572 two_stage_opamp_dummy_magic_29_0.V_source.t10 GNDA_2 0.012908f
C573 two_stage_opamp_dummy_magic_29_0.V_source.t19 GNDA_2 0.012908f
C574 two_stage_opamp_dummy_magic_29_0.V_source.n20 GNDA_2 0.028087f
C575 two_stage_opamp_dummy_magic_29_0.V_source.n21 GNDA_2 0.113801f
C576 two_stage_opamp_dummy_magic_29_0.V_source.n22 GNDA_2 0.027589f
C577 two_stage_opamp_dummy_magic_29_0.V_source.n23 GNDA_2 0.027589f
C578 two_stage_opamp_dummy_magic_29_0.V_source.t4 GNDA_2 0.012908f
C579 two_stage_opamp_dummy_magic_29_0.V_source.t6 GNDA_2 0.012908f
C580 two_stage_opamp_dummy_magic_29_0.V_source.n24 GNDA_2 0.028087f
C581 two_stage_opamp_dummy_magic_29_0.V_source.n25 GNDA_2 0.085239f
C582 two_stage_opamp_dummy_magic_29_0.V_source.t39 GNDA_2 0.012908f
C583 two_stage_opamp_dummy_magic_29_0.V_source.t9 GNDA_2 0.012908f
C584 two_stage_opamp_dummy_magic_29_0.V_source.n26 GNDA_2 0.028087f
C585 two_stage_opamp_dummy_magic_29_0.V_source.n27 GNDA_2 0.085239f
C586 two_stage_opamp_dummy_magic_29_0.V_source.n28 GNDA_2 0.069756f
C587 two_stage_opamp_dummy_magic_29_0.V_source.t30 GNDA_2 0.012908f
C588 two_stage_opamp_dummy_magic_29_0.V_source.t35 GNDA_2 0.012908f
C589 two_stage_opamp_dummy_magic_29_0.V_source.n29 GNDA_2 0.028087f
C590 two_stage_opamp_dummy_magic_29_0.V_source.n30 GNDA_2 0.085239f
C591 two_stage_opamp_dummy_magic_29_0.V_source.n31 GNDA_2 0.069756f
C592 two_stage_opamp_dummy_magic_29_0.V_source.t28 GNDA_2 0.012908f
C593 two_stage_opamp_dummy_magic_29_0.V_source.t31 GNDA_2 0.012908f
C594 two_stage_opamp_dummy_magic_29_0.V_source.n32 GNDA_2 0.028087f
C595 two_stage_opamp_dummy_magic_29_0.V_source.n33 GNDA_2 0.085239f
C596 two_stage_opamp_dummy_magic_29_0.V_source.n34 GNDA_2 0.027589f
C597 two_stage_opamp_dummy_magic_29_0.V_source.t36 GNDA_2 0.012908f
C598 two_stage_opamp_dummy_magic_29_0.V_source.t32 GNDA_2 0.012908f
C599 two_stage_opamp_dummy_magic_29_0.V_source.n35 GNDA_2 0.028087f
C600 two_stage_opamp_dummy_magic_29_0.V_source.n36 GNDA_2 0.117879f
C601 two_stage_opamp_dummy_magic_29_0.V_source.t37 GNDA_2 0.012908f
C602 two_stage_opamp_dummy_magic_29_0.V_source.t33 GNDA_2 0.012908f
C603 two_stage_opamp_dummy_magic_29_0.V_source.n37 GNDA_2 0.028087f
C604 two_stage_opamp_dummy_magic_29_0.V_source.n38 GNDA_2 0.113801f
C605 two_stage_opamp_dummy_magic_29_0.V_source.n39 GNDA_2 0.046931f
C606 two_stage_opamp_dummy_magic_29_0.V_source.n40 GNDA_2 0.027589f
C607 two_stage_opamp_dummy_magic_29_0.V_source.t29 GNDA_2 0.012908f
C608 two_stage_opamp_dummy_magic_29_0.V_source.t34 GNDA_2 0.012908f
C609 two_stage_opamp_dummy_magic_29_0.V_source.n41 GNDA_2 0.028087f
C610 two_stage_opamp_dummy_magic_29_0.V_source.n42 GNDA_2 0.113801f
C611 two_stage_opamp_dummy_magic_29_0.V_source.n43 GNDA_2 0.054121f
C612 two_stage_opamp_dummy_magic_29_0.V_source.n44 GNDA_2 0.147729f
C613 two_stage_opamp_dummy_magic_29_0.V_source.t16 GNDA_2 0.021514f
C614 two_stage_opamp_dummy_magic_29_0.V_source.t25 GNDA_2 0.021514f
C615 two_stage_opamp_dummy_magic_29_0.V_source.n45 GNDA_2 0.045993f
C616 two_stage_opamp_dummy_magic_29_0.V_source.n46 GNDA_2 0.164071f
C617 two_stage_opamp_dummy_magic_29_0.V_source.t8 GNDA_2 0.021514f
C618 two_stage_opamp_dummy_magic_29_0.V_source.t38 GNDA_2 0.021514f
C619 two_stage_opamp_dummy_magic_29_0.V_source.n47 GNDA_2 0.045993f
C620 two_stage_opamp_dummy_magic_29_0.V_source.n48 GNDA_2 0.164071f
C621 two_stage_opamp_dummy_magic_29_0.V_source.t11 GNDA_2 0.021514f
C622 two_stage_opamp_dummy_magic_29_0.V_source.t20 GNDA_2 0.021514f
C623 two_stage_opamp_dummy_magic_29_0.V_source.n49 GNDA_2 0.045993f
C624 two_stage_opamp_dummy_magic_29_0.V_source.n50 GNDA_2 0.164071f
C625 two_stage_opamp_dummy_magic_29_0.V_source.n51 GNDA_2 0.153086f
C626 two_stage_opamp_dummy_magic_29_0.V_source.t18 GNDA_2 0.021514f
C627 two_stage_opamp_dummy_magic_29_0.V_source.t2 GNDA_2 0.021514f
C628 two_stage_opamp_dummy_magic_29_0.V_source.n52 GNDA_2 0.045993f
C629 two_stage_opamp_dummy_magic_29_0.V_source.n53 GNDA_2 0.164071f
C630 two_stage_opamp_dummy_magic_29_0.V_source.n54 GNDA_2 0.153086f
C631 two_stage_opamp_dummy_magic_29_0.V_source.n55 GNDA_2 0.956519f
C632 two_stage_opamp_dummy_magic_29_0.V_source.t23 GNDA_2 0.047788f
C633 two_stage_opamp_dummy_magic_29_0.V_source.n56 GNDA_2 2.31891f
C634 two_stage_opamp_dummy_magic_29_0.V_source.n57 GNDA_2 1.17166f
C635 two_stage_opamp_dummy_magic_29_0.V_source.n58 GNDA_2 0.153086f
C636 two_stage_opamp_dummy_magic_29_0.V_source.t17 GNDA_2 0.021514f
C637 two_stage_opamp_dummy_magic_29_0.V_source.t12 GNDA_2 0.021514f
C638 two_stage_opamp_dummy_magic_29_0.V_source.n59 GNDA_2 0.045993f
C639 two_stage_opamp_dummy_magic_29_0.V_source.n60 GNDA_2 0.164071f
C640 two_stage_opamp_dummy_magic_29_0.V_source.n61 GNDA_2 0.118148f
C641 two_stage_opamp_dummy_magic_29_0.V_source.t13 GNDA_2 0.021514f
C642 two_stage_opamp_dummy_magic_29_0.V_source.t1 GNDA_2 0.021514f
C643 two_stage_opamp_dummy_magic_29_0.V_source.n62 GNDA_2 0.045993f
C644 two_stage_opamp_dummy_magic_29_0.V_source.n63 GNDA_2 0.193086f
C645 two_stage_opamp_dummy_magic_29_0.V_source.n64 GNDA_2 0.153086f
C646 two_stage_opamp_dummy_magic_29_0.V_source.t7 GNDA_2 0.021514f
C647 two_stage_opamp_dummy_magic_29_0.V_source.t26 GNDA_2 0.021514f
C648 two_stage_opamp_dummy_magic_29_0.V_source.n65 GNDA_2 0.045993f
C649 two_stage_opamp_dummy_magic_29_0.V_source.n66 GNDA_2 0.193086f
C650 two_stage_opamp_dummy_magic_29_0.V_source.n67 GNDA_2 0.153086f
C651 two_stage_opamp_dummy_magic_29_0.V_source.n68 GNDA_2 0.153086f
C652 two_stage_opamp_dummy_magic_29_0.V_source.t5 GNDA_2 0.021514f
C653 two_stage_opamp_dummy_magic_29_0.V_source.t0 GNDA_2 0.021514f
C654 two_stage_opamp_dummy_magic_29_0.V_source.n69 GNDA_2 0.045993f
C655 two_stage_opamp_dummy_magic_29_0.V_source.n70 GNDA_2 0.193086f
C656 two_stage_opamp_dummy_magic_29_0.V_source.n71 GNDA_2 0.066185f
C657 two_stage_opamp_dummy_magic_29_0.V_source.n72 GNDA_2 0.113174f
C658 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n0 GNDA_2 0.029703f
C659 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n1 GNDA_2 0.02026f
C660 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n2 GNDA_2 0.664294f
C661 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.t1 GNDA_2 0.113706f
C662 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n3 GNDA_2 0.046075f
C663 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n4 GNDA_2 0.056526f
C664 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.t13 GNDA_2 0.028335f
C665 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.t6 GNDA_2 0.028335f
C666 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n5 GNDA_2 0.060602f
C667 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n6 GNDA_2 0.189038f
C668 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.t10 GNDA_2 0.028335f
C669 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.t5 GNDA_2 0.028335f
C670 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n7 GNDA_2 0.060602f
C671 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n8 GNDA_2 0.184429f
C672 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n9 GNDA_2 0.076885f
C673 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n10 GNDA_2 0.046075f
C674 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.t9 GNDA_2 0.028335f
C675 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.t14 GNDA_2 0.028335f
C676 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n11 GNDA_2 0.060602f
C677 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n12 GNDA_2 0.184429f
C678 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n13 GNDA_2 0.032852f
C679 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.t12 GNDA_2 0.028335f
C680 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.t8 GNDA_2 0.028335f
C681 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n14 GNDA_2 0.060602f
C682 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n15 GNDA_2 0.184429f
C683 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n16 GNDA_2 0.056526f
C684 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.t11 GNDA_2 0.028335f
C685 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.t7 GNDA_2 0.028335f
C686 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n17 GNDA_2 0.060602f
C687 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n18 GNDA_2 0.186996f
C688 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n19 GNDA_2 0.130351f
C689 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n20 GNDA_2 6.67459f
C690 bgr_11_0.V_CMFB_S4 GNDA_2 2.9987f
C691 two_stage_opamp_dummy_magic_29_0.V_err_gate.t1 GNDA_2 0.019449f
C692 two_stage_opamp_dummy_magic_29_0.V_err_gate.t2 GNDA_2 0.019449f
C693 two_stage_opamp_dummy_magic_29_0.V_err_gate.n0 GNDA_2 0.238208f
C694 two_stage_opamp_dummy_magic_29_0.V_err_gate.t0 GNDA_2 0.048624f
C695 two_stage_opamp_dummy_magic_29_0.V_err_gate.t4 GNDA_2 0.048624f
C696 two_stage_opamp_dummy_magic_29_0.V_err_gate.n1 GNDA_2 0.154108f
C697 two_stage_opamp_dummy_magic_29_0.V_err_gate.t9 GNDA_2 0.054296f
C698 two_stage_opamp_dummy_magic_29_0.V_err_gate.t7 GNDA_2 0.054296f
C699 two_stage_opamp_dummy_magic_29_0.V_err_gate.n2 GNDA_2 0.081557f
C700 two_stage_opamp_dummy_magic_29_0.V_err_gate.n3 GNDA_2 0.295866f
C701 two_stage_opamp_dummy_magic_29_0.V_err_gate.t3 GNDA_2 0.048624f
C702 two_stage_opamp_dummy_magic_29_0.V_err_gate.t5 GNDA_2 0.048624f
C703 two_stage_opamp_dummy_magic_29_0.V_err_gate.n4 GNDA_2 0.153478f
C704 two_stage_opamp_dummy_magic_29_0.V_err_gate.n5 GNDA_2 0.225156f
C705 two_stage_opamp_dummy_magic_29_0.V_err_gate.t8 GNDA_2 0.054296f
C706 two_stage_opamp_dummy_magic_29_0.V_err_gate.t6 GNDA_2 0.054296f
C707 two_stage_opamp_dummy_magic_29_0.V_err_gate.n6 GNDA_2 0.081557f
C708 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n0 GNDA_2 0.011962f
C709 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n1 GNDA_2 0.081192f
C710 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n2 GNDA_2 0.012656f
C711 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n3 GNDA_2 0.086961f
C712 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n4 GNDA_2 0.011962f
C713 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n5 GNDA_2 0.395797f
C714 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n7 GNDA_2 0.028116f
C715 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n8 GNDA_2 0.028116f
C716 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n11 GNDA_2 0.028116f
C717 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n12 GNDA_2 0.028116f
C718 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.t0 GNDA_2 0.071178f
C719 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n13 GNDA_2 0.026704f
C720 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n14 GNDA_2 0.03273f
C721 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.t14 GNDA_2 0.011715f
C722 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.t7 GNDA_2 0.011715f
C723 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n15 GNDA_2 0.023952f
C724 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n16 GNDA_2 0.080191f
C725 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.t11 GNDA_2 0.011715f
C726 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.t16 GNDA_2 0.011715f
C727 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n17 GNDA_2 0.023952f
C728 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n18 GNDA_2 0.077479f
C729 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n19 GNDA_2 0.044027f
C730 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n20 GNDA_2 0.026704f
C731 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.t10 GNDA_2 0.011715f
C732 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.t15 GNDA_2 0.011715f
C733 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n21 GNDA_2 0.023952f
C734 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n22 GNDA_2 0.077479f
C735 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n23 GNDA_2 0.01918f
C736 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.t13 GNDA_2 0.011715f
C737 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.t9 GNDA_2 0.011715f
C738 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n24 GNDA_2 0.023952f
C739 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n25 GNDA_2 0.077479f
C740 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n26 GNDA_2 0.03273f
C741 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.t12 GNDA_2 0.011715f
C742 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.t8 GNDA_2 0.011715f
C743 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n27 GNDA_2 0.023952f
C744 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n28 GNDA_2 0.07901f
C745 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n29 GNDA_2 0.106722f
C746 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n30 GNDA_2 0.710297f
C747 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n31 GNDA_2 0.170453f
C748 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n33 GNDA_2 0.028116f
C749 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n34 GNDA_2 0.027852f
C750 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n35 GNDA_2 0.040417f
C751 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n36 GNDA_2 0.040417f
C752 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n37 GNDA_2 0.028116f
C753 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n38 GNDA_2 0.028116f
C754 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n40 GNDA_2 3.14455f
C755 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n41 GNDA_2 1.49923f
C756 bgr_11_0.V_CMFB_S3 GNDA_2 0.345498f
C757 bgr_11_0.Vin+.t4 GNDA_2 0.221779f
C758 bgr_11_0.Vin+.t5 GNDA_2 0.096124f
C759 bgr_11_0.Vin+.n0 GNDA_2 1.46352f
C760 bgr_11_0.Vin+.t0 GNDA_2 0.033039f
C761 bgr_11_0.Vin+.t3 GNDA_2 0.033039f
C762 bgr_11_0.Vin+.n1 GNDA_2 0.084276f
C763 bgr_11_0.Vin+.t2 GNDA_2 0.033039f
C764 bgr_11_0.Vin+.t1 GNDA_2 0.033039f
C765 bgr_11_0.Vin+.n2 GNDA_2 0.078979f
C766 bgr_11_0.Vin+.n3 GNDA_2 0.79622f
C767 bgr_11_0.Vin+.n4 GNDA_2 0.652102f
C768 bgr_11_0.Vin+.t6 GNDA_2 0.052809f
C769 two_stage_opamp_dummy_magic_29_0.Vb3.n0 GNDA_2 0.201673f
C770 two_stage_opamp_dummy_magic_29_0.Vb3.n1 GNDA_2 0.210233f
C771 two_stage_opamp_dummy_magic_29_0.Vb3.n2 GNDA_2 0.068292f
C772 two_stage_opamp_dummy_magic_29_0.Vb3.n3 GNDA_2 0.159849f
C773 two_stage_opamp_dummy_magic_29_0.Vb3.n4 GNDA_2 0.210233f
C774 two_stage_opamp_dummy_magic_29_0.Vb3.n5 GNDA_2 0.486246f
C775 two_stage_opamp_dummy_magic_29_0.Vb3.n6 GNDA_2 0.139263f
C776 two_stage_opamp_dummy_magic_29_0.Vb3.n7 GNDA_2 0.210233f
C777 two_stage_opamp_dummy_magic_29_0.Vb3.n8 GNDA_2 0.139263f
C778 two_stage_opamp_dummy_magic_29_0.Vb3.n9 GNDA_2 0.30679f
C779 two_stage_opamp_dummy_magic_29_0.Vb3.t0 GNDA_2 0.014227f
C780 two_stage_opamp_dummy_magic_29_0.Vb3.t3 GNDA_2 0.014227f
C781 two_stage_opamp_dummy_magic_29_0.Vb3.n10 GNDA_2 0.045828f
C782 two_stage_opamp_dummy_magic_29_0.Vb3.t1 GNDA_2 0.014227f
C783 two_stage_opamp_dummy_magic_29_0.Vb3.t2 GNDA_2 0.014227f
C784 two_stage_opamp_dummy_magic_29_0.Vb3.n11 GNDA_2 0.045828f
C785 two_stage_opamp_dummy_magic_29_0.Vb3.n12 GNDA_2 0.252648f
C786 two_stage_opamp_dummy_magic_29_0.Vb3.t5 GNDA_2 0.014227f
C787 two_stage_opamp_dummy_magic_29_0.Vb3.t4 GNDA_2 0.014227f
C788 two_stage_opamp_dummy_magic_29_0.Vb3.n13 GNDA_2 0.042973f
C789 two_stage_opamp_dummy_magic_29_0.Vb3.n14 GNDA_2 0.806482f
C790 two_stage_opamp_dummy_magic_29_0.Vb3.t28 GNDA_2 0.091246f
C791 two_stage_opamp_dummy_magic_29_0.Vb3.t23 GNDA_2 0.091222f
C792 two_stage_opamp_dummy_magic_29_0.Vb3.t15 GNDA_2 0.091222f
C793 two_stage_opamp_dummy_magic_29_0.Vb3.t12 GNDA_2 0.091222f
C794 two_stage_opamp_dummy_magic_29_0.Vb3.t10 GNDA_2 0.090805f
C795 two_stage_opamp_dummy_magic_29_0.Vb3.t9 GNDA_2 0.090805f
C796 two_stage_opamp_dummy_magic_29_0.Vb3.t27 GNDA_2 0.091222f
C797 two_stage_opamp_dummy_magic_29_0.Vb3.t21 GNDA_2 0.091222f
C798 two_stage_opamp_dummy_magic_29_0.Vb3.t24 GNDA_2 0.091222f
C799 two_stage_opamp_dummy_magic_29_0.Vb3.t17 GNDA_2 0.091222f
C800 two_stage_opamp_dummy_magic_29_0.Vb3.t6 GNDA_2 0.049796f
C801 two_stage_opamp_dummy_magic_29_0.Vb3.t7 GNDA_2 0.049796f
C802 two_stage_opamp_dummy_magic_29_0.Vb3.n15 GNDA_2 0.134068f
C803 two_stage_opamp_dummy_magic_29_0.Vb3.t19 GNDA_2 0.093507f
C804 two_stage_opamp_dummy_magic_29_0.Vb3.n16 GNDA_2 0.936585f
C805 two_stage_opamp_dummy_magic_29_0.Vb3.n17 GNDA_2 1.06421f
C806 two_stage_opamp_dummy_magic_29_0.Vb3.t22 GNDA_2 0.091246f
C807 two_stage_opamp_dummy_magic_29_0.Vb3.t18 GNDA_2 0.091222f
C808 two_stage_opamp_dummy_magic_29_0.Vb3.t25 GNDA_2 0.091222f
C809 two_stage_opamp_dummy_magic_29_0.Vb3.t11 GNDA_2 0.091222f
C810 two_stage_opamp_dummy_magic_29_0.Vb3.t16 GNDA_2 0.090795f
C811 two_stage_opamp_dummy_magic_29_0.Vb3.t13 GNDA_2 0.090795f
C812 two_stage_opamp_dummy_magic_29_0.Vb3.n18 GNDA_2 0.079934f
C813 two_stage_opamp_dummy_magic_29_0.Vb3.n19 GNDA_2 0.079934f
C814 two_stage_opamp_dummy_magic_29_0.Vb3.t14 GNDA_2 0.091222f
C815 two_stage_opamp_dummy_magic_29_0.Vb3.t20 GNDA_2 0.091222f
C816 two_stage_opamp_dummy_magic_29_0.Vb3.t26 GNDA_2 0.091222f
C817 two_stage_opamp_dummy_magic_29_0.Vb3.t8 GNDA_2 0.091222f
C818 two_stage_opamp_dummy_magic_29_0.Vb3.n20 GNDA_2 0.146376f
C819 two_stage_opamp_dummy_magic_29_0.Vb3.n21 GNDA_2 1.25819f
C820 bgr_11_0.VB3_CUR_BIAS GNDA_2 1.7736f
C821 two_stage_opamp_dummy_magic_29_0.VD3.n0 GNDA_2 1.11096f
C822 two_stage_opamp_dummy_magic_29_0.VD3.n1 GNDA_2 0.20151f
C823 two_stage_opamp_dummy_magic_29_0.VD3.n2 GNDA_2 0.378259f
C824 two_stage_opamp_dummy_magic_29_0.VD3.t3 GNDA_2 0.078836f
C825 two_stage_opamp_dummy_magic_29_0.VD3.n3 GNDA_2 0.149757f
C826 two_stage_opamp_dummy_magic_29_0.VD3.t12 GNDA_2 0.045031f
C827 two_stage_opamp_dummy_magic_29_0.VD3.t15 GNDA_2 0.045031f
C828 two_stage_opamp_dummy_magic_29_0.VD3.n4 GNDA_2 0.092115f
C829 two_stage_opamp_dummy_magic_29_0.VD3.n5 GNDA_2 0.260153f
C830 two_stage_opamp_dummy_magic_29_0.VD3.t22 GNDA_2 0.045031f
C831 two_stage_opamp_dummy_magic_29_0.VD3.t18 GNDA_2 0.045031f
C832 two_stage_opamp_dummy_magic_29_0.VD3.n6 GNDA_2 0.095624f
C833 two_stage_opamp_dummy_magic_29_0.VD3.t14 GNDA_2 0.045031f
C834 two_stage_opamp_dummy_magic_29_0.VD3.t2 GNDA_2 0.045031f
C835 two_stage_opamp_dummy_magic_29_0.VD3.n7 GNDA_2 0.092115f
C836 two_stage_opamp_dummy_magic_29_0.VD3.n8 GNDA_2 0.25692f
C837 two_stage_opamp_dummy_magic_29_0.VD3.t1 GNDA_2 0.045031f
C838 two_stage_opamp_dummy_magic_29_0.VD3.t10 GNDA_2 0.045031f
C839 two_stage_opamp_dummy_magic_29_0.VD3.n9 GNDA_2 0.092115f
C840 two_stage_opamp_dummy_magic_29_0.VD3.n10 GNDA_2 0.25692f
C841 two_stage_opamp_dummy_magic_29_0.VD3.t26 GNDA_2 0.045031f
C842 two_stage_opamp_dummy_magic_29_0.VD3.t28 GNDA_2 0.045031f
C843 two_stage_opamp_dummy_magic_29_0.VD3.n11 GNDA_2 0.095624f
C844 two_stage_opamp_dummy_magic_29_0.VD3.n12 GNDA_2 0.76157f
C845 two_stage_opamp_dummy_magic_29_0.VD3.t5 GNDA_2 0.160181f
C846 two_stage_opamp_dummy_magic_29_0.VD3.n13 GNDA_2 0.51334f
C847 two_stage_opamp_dummy_magic_29_0.VD3.t4 GNDA_2 0.383839f
C848 two_stage_opamp_dummy_magic_29_0.VD3.t17 GNDA_2 0.301063f
C849 two_stage_opamp_dummy_magic_29_0.VD3.t21 GNDA_2 0.301063f
C850 two_stage_opamp_dummy_magic_29_0.VD3.t35 GNDA_2 0.301063f
C851 two_stage_opamp_dummy_magic_29_0.VD3.t31 GNDA_2 0.301063f
C852 two_stage_opamp_dummy_magic_29_0.VD3.t27 GNDA_2 0.301063f
C853 two_stage_opamp_dummy_magic_29_0.VD3.t25 GNDA_2 0.301063f
C854 two_stage_opamp_dummy_magic_29_0.VD3.t23 GNDA_2 0.301063f
C855 two_stage_opamp_dummy_magic_29_0.VD3.t19 GNDA_2 0.301063f
C856 two_stage_opamp_dummy_magic_29_0.VD3.t33 GNDA_2 0.301063f
C857 two_stage_opamp_dummy_magic_29_0.VD3.t29 GNDA_2 0.301063f
C858 two_stage_opamp_dummy_magic_29_0.VD3.t7 GNDA_2 0.383839f
C859 two_stage_opamp_dummy_magic_29_0.VD3.t8 GNDA_2 0.160181f
C860 two_stage_opamp_dummy_magic_29_0.VD3.n14 GNDA_2 0.51334f
C861 two_stage_opamp_dummy_magic_29_0.VD3.t6 GNDA_2 0.078836f
C862 two_stage_opamp_dummy_magic_29_0.VD3.n15 GNDA_2 0.215181f
C863 two_stage_opamp_dummy_magic_29_0.VD3.t20 GNDA_2 0.045031f
C864 two_stage_opamp_dummy_magic_29_0.VD3.t24 GNDA_2 0.045031f
C865 two_stage_opamp_dummy_magic_29_0.VD3.n16 GNDA_2 0.095624f
C866 two_stage_opamp_dummy_magic_29_0.VD3.t37 GNDA_2 0.045031f
C867 two_stage_opamp_dummy_magic_29_0.VD3.t11 GNDA_2 0.045031f
C868 two_stage_opamp_dummy_magic_29_0.VD3.n17 GNDA_2 0.092115f
C869 two_stage_opamp_dummy_magic_29_0.VD3.n18 GNDA_2 0.25692f
C870 two_stage_opamp_dummy_magic_29_0.VD3.t30 GNDA_2 0.045031f
C871 two_stage_opamp_dummy_magic_29_0.VD3.t34 GNDA_2 0.045031f
C872 two_stage_opamp_dummy_magic_29_0.VD3.n19 GNDA_2 0.095624f
C873 two_stage_opamp_dummy_magic_29_0.VD3.n20 GNDA_2 0.115041f
C874 two_stage_opamp_dummy_magic_29_0.VD3.n21 GNDA_2 0.069429f
C875 two_stage_opamp_dummy_magic_29_0.VD3.t13 GNDA_2 0.045031f
C876 two_stage_opamp_dummy_magic_29_0.VD3.t9 GNDA_2 0.045031f
C877 two_stage_opamp_dummy_magic_29_0.VD3.n22 GNDA_2 0.092115f
C878 two_stage_opamp_dummy_magic_29_0.VD3.n23 GNDA_2 0.25692f
C879 two_stage_opamp_dummy_magic_29_0.VD3.n24 GNDA_2 0.069429f
C880 two_stage_opamp_dummy_magic_29_0.VD3.n25 GNDA_2 0.115041f
C881 two_stage_opamp_dummy_magic_29_0.VD3.t16 GNDA_2 0.045031f
C882 two_stage_opamp_dummy_magic_29_0.VD3.t0 GNDA_2 0.045031f
C883 two_stage_opamp_dummy_magic_29_0.VD3.n26 GNDA_2 0.092115f
C884 two_stage_opamp_dummy_magic_29_0.VD3.n27 GNDA_2 0.260153f
C885 two_stage_opamp_dummy_magic_29_0.VD3.n28 GNDA_2 0.76157f
C886 two_stage_opamp_dummy_magic_29_0.VD3.n29 GNDA_2 1.26178f
C887 two_stage_opamp_dummy_magic_29_0.VD3.n30 GNDA_2 0.432296f
C888 two_stage_opamp_dummy_magic_29_0.VD3.t32 GNDA_2 0.045031f
C889 two_stage_opamp_dummy_magic_29_0.VD3.t36 GNDA_2 0.045031f
C890 two_stage_opamp_dummy_magic_29_0.VD3.n31 GNDA_2 0.095624f
C891 two_stage_opamp_dummy_magic_29_0.VD3.n32 GNDA_2 0.76157f
C892 two_stage_opamp_dummy_magic_29_0.VD3.n33 GNDA_2 0.76157f
C893 two_stage_opamp_dummy_magic_29_0.VD3.n34 GNDA_2 0.342878f
C894 two_stage_opamp_dummy_magic_29_0.VD2.t10 GNDA_2 0.033932f
C895 two_stage_opamp_dummy_magic_29_0.VD2.t15 GNDA_2 0.033932f
C896 two_stage_opamp_dummy_magic_29_0.VD2.n0 GNDA_2 0.075122f
C897 two_stage_opamp_dummy_magic_29_0.VD2.n1 GNDA_2 0.564997f
C898 two_stage_opamp_dummy_magic_29_0.VD2.n2 GNDA_2 0.050916f
C899 two_stage_opamp_dummy_magic_29_0.VD2.n3 GNDA_2 0.222536f
C900 two_stage_opamp_dummy_magic_29_0.VD2.t19 GNDA_2 0.033932f
C901 two_stage_opamp_dummy_magic_29_0.VD2.t4 GNDA_2 0.033932f
C902 two_stage_opamp_dummy_magic_29_0.VD2.n4 GNDA_2 0.073831f
C903 two_stage_opamp_dummy_magic_29_0.VD2.n5 GNDA_2 0.284467f
C904 two_stage_opamp_dummy_magic_29_0.VD2.n6 GNDA_2 0.072163f
C905 two_stage_opamp_dummy_magic_29_0.VD2.t1 GNDA_2 0.033932f
C906 two_stage_opamp_dummy_magic_29_0.VD2.t3 GNDA_2 0.033932f
C907 two_stage_opamp_dummy_magic_29_0.VD2.n7 GNDA_2 0.073831f
C908 two_stage_opamp_dummy_magic_29_0.VD2.n8 GNDA_2 0.292399f
C909 two_stage_opamp_dummy_magic_29_0.VD2.t7 GNDA_2 0.033932f
C910 two_stage_opamp_dummy_magic_29_0.VD2.t13 GNDA_2 0.033932f
C911 two_stage_opamp_dummy_magic_29_0.VD2.n9 GNDA_2 0.075122f
C912 two_stage_opamp_dummy_magic_29_0.VD2.t11 GNDA_2 0.033932f
C913 two_stage_opamp_dummy_magic_29_0.VD2.t6 GNDA_2 0.033932f
C914 two_stage_opamp_dummy_magic_29_0.VD2.n10 GNDA_2 0.075122f
C915 two_stage_opamp_dummy_magic_29_0.VD2.n11 GNDA_2 0.767242f
C916 two_stage_opamp_dummy_magic_29_0.VD2.t9 GNDA_2 0.033932f
C917 two_stage_opamp_dummy_magic_29_0.VD2.t12 GNDA_2 0.033932f
C918 two_stage_opamp_dummy_magic_29_0.VD2.n12 GNDA_2 0.075122f
C919 two_stage_opamp_dummy_magic_29_0.VD2.n13 GNDA_2 0.268181f
C920 two_stage_opamp_dummy_magic_29_0.VD2.t2 GNDA_2 0.033932f
C921 two_stage_opamp_dummy_magic_29_0.VD2.t17 GNDA_2 0.033932f
C922 two_stage_opamp_dummy_magic_29_0.VD2.n14 GNDA_2 0.073831f
C923 two_stage_opamp_dummy_magic_29_0.VD2.n15 GNDA_2 0.292399f
C924 two_stage_opamp_dummy_magic_29_0.VD2.n16 GNDA_2 0.122664f
C925 two_stage_opamp_dummy_magic_29_0.VD2.t18 GNDA_2 0.033932f
C926 two_stage_opamp_dummy_magic_29_0.VD2.t16 GNDA_2 0.033932f
C927 two_stage_opamp_dummy_magic_29_0.VD2.n17 GNDA_2 0.073831f
C928 two_stage_opamp_dummy_magic_29_0.VD2.n18 GNDA_2 0.284467f
C929 two_stage_opamp_dummy_magic_29_0.VD2.n19 GNDA_2 0.050916f
C930 two_stage_opamp_dummy_magic_29_0.VD2.n20 GNDA_2 0.222536f
C931 two_stage_opamp_dummy_magic_29_0.VD2.n21 GNDA_2 0.761461f
C932 two_stage_opamp_dummy_magic_29_0.VD2.n22 GNDA_2 0.114111f
C933 two_stage_opamp_dummy_magic_29_0.VD2.n23 GNDA_2 0.067863f
C934 two_stage_opamp_dummy_magic_29_0.VD2.t8 GNDA_2 0.033932f
C935 two_stage_opamp_dummy_magic_29_0.VD2.t14 GNDA_2 0.033932f
C936 two_stage_opamp_dummy_magic_29_0.VD2.n24 GNDA_2 0.075122f
C937 two_stage_opamp_dummy_magic_29_0.VD2.n25 GNDA_2 0.761461f
C938 two_stage_opamp_dummy_magic_29_0.VD2.n26 GNDA_2 0.114111f
C939 two_stage_opamp_dummy_magic_29_0.VD2.n27 GNDA_2 0.767242f
C940 two_stage_opamp_dummy_magic_29_0.VD2.n28 GNDA_2 0.268181f
C941 two_stage_opamp_dummy_magic_29_0.VD2.n29 GNDA_2 0.050916f
C942 two_stage_opamp_dummy_magic_29_0.VD2.t20 GNDA_2 0.033932f
C943 two_stage_opamp_dummy_magic_29_0.VD2.t5 GNDA_2 0.033932f
C944 two_stage_opamp_dummy_magic_29_0.VD2.n30 GNDA_2 0.073831f
C945 two_stage_opamp_dummy_magic_29_0.VD2.n31 GNDA_2 0.284467f
C946 two_stage_opamp_dummy_magic_29_0.VD2.n32 GNDA_2 0.122664f
C947 two_stage_opamp_dummy_magic_29_0.VD2.n33 GNDA_2 0.072163f
C948 two_stage_opamp_dummy_magic_29_0.VD2.t21 GNDA_2 0.033932f
C949 two_stage_opamp_dummy_magic_29_0.VD2.t0 GNDA_2 0.033932f
C950 two_stage_opamp_dummy_magic_29_0.VD2.n34 GNDA_2 0.073831f
C951 two_stage_opamp_dummy_magic_29_0.VD2.n35 GNDA_2 0.284467f
C952 two_stage_opamp_dummy_magic_29_0.VD2.n36 GNDA_2 0.050916f
C953 two_stage_opamp_dummy_magic_29_0.VD2.n37 GNDA_2 0.039407f
C954 two_stage_opamp_dummy_magic_29_0.Vb1_2.t2 GNDA_2 0.029732f
C955 two_stage_opamp_dummy_magic_29_0.Vb1_2.t0 GNDA_2 0.029732f
C956 two_stage_opamp_dummy_magic_29_0.Vb1_2.n0 GNDA_2 0.087151f
C957 two_stage_opamp_dummy_magic_29_0.Vb1_2.t4 GNDA_2 0.189479f
C958 two_stage_opamp_dummy_magic_29_0.Vb1_2.t1 GNDA_2 0.029732f
C959 two_stage_opamp_dummy_magic_29_0.Vb1_2.t3 GNDA_2 0.029732f
C960 two_stage_opamp_dummy_magic_29_0.Vb1_2.n1 GNDA_2 0.086354f
C961 two_stage_opamp_dummy_magic_29_0.Vb1.n0 GNDA_2 1.88534f
C962 two_stage_opamp_dummy_magic_29_0.Vb1.n1 GNDA_2 0.234861f
C963 two_stage_opamp_dummy_magic_29_0.Vb1.n2 GNDA_2 1.99634f
C964 two_stage_opamp_dummy_magic_29_0.Vb1.n3 GNDA_2 0.486012f
C965 two_stage_opamp_dummy_magic_29_0.Vb1.n4 GNDA_2 0.573498f
C966 two_stage_opamp_dummy_magic_29_0.Vb1.n5 GNDA_2 0.486012f
C967 two_stage_opamp_dummy_magic_29_0.Vb1.n6 GNDA_2 1.75333f
C968 two_stage_opamp_dummy_magic_29_0.Vb1.n7 GNDA_2 0.330492f
C969 two_stage_opamp_dummy_magic_29_0.Vb1.t20 GNDA_2 0.047637f
C970 two_stage_opamp_dummy_magic_29_0.Vb1.t5 GNDA_2 0.030922f
C971 two_stage_opamp_dummy_magic_29_0.Vb1.t3 GNDA_2 0.040107f
C972 two_stage_opamp_dummy_magic_29_0.Vb1.n8 GNDA_2 0.041235f
C973 two_stage_opamp_dummy_magic_29_0.Vb1.t7 GNDA_2 0.030922f
C974 two_stage_opamp_dummy_magic_29_0.Vb1.t9 GNDA_2 0.040107f
C975 two_stage_opamp_dummy_magic_29_0.Vb1.n9 GNDA_2 0.041235f
C976 two_stage_opamp_dummy_magic_29_0.Vb1.n10 GNDA_2 0.030737f
C977 two_stage_opamp_dummy_magic_29_0.Vb1.t6 GNDA_2 0.030168f
C978 two_stage_opamp_dummy_magic_29_0.Vb1.t8 GNDA_2 0.030168f
C979 two_stage_opamp_dummy_magic_29_0.Vb1.n11 GNDA_2 0.065642f
C980 two_stage_opamp_dummy_magic_29_0.Vb1.t31 GNDA_2 0.93909f
C981 two_stage_opamp_dummy_magic_29_0.Vb1.n12 GNDA_2 0.110397f
C982 two_stage_opamp_dummy_magic_29_0.Vb1.t30 GNDA_2 0.047637f
C983 two_stage_opamp_dummy_magic_29_0.Vb1.t19 GNDA_2 0.047637f
C984 two_stage_opamp_dummy_magic_29_0.Vb1.t28 GNDA_2 0.047637f
C985 two_stage_opamp_dummy_magic_29_0.Vb1.t16 GNDA_2 0.047637f
C986 two_stage_opamp_dummy_magic_29_0.Vb1.t29 GNDA_2 0.047637f
C987 two_stage_opamp_dummy_magic_29_0.Vb1.t17 GNDA_2 0.047637f
C988 two_stage_opamp_dummy_magic_29_0.Vb1.t27 GNDA_2 0.047637f
C989 two_stage_opamp_dummy_magic_29_0.Vb1.t14 GNDA_2 0.047637f
C990 two_stage_opamp_dummy_magic_29_0.Vb1.t21 GNDA_2 0.047637f
C991 two_stage_opamp_dummy_magic_29_0.Vb1.n13 GNDA_2 1.79685f
C992 two_stage_opamp_dummy_magic_29_0.Vb1.t0 GNDA_2 0.030168f
C993 two_stage_opamp_dummy_magic_29_0.Vb1.t4 GNDA_2 0.030168f
C994 two_stage_opamp_dummy_magic_29_0.Vb1.n14 GNDA_2 0.065642f
C995 two_stage_opamp_dummy_magic_29_0.Vb1.n15 GNDA_2 0.246742f
C996 two_stage_opamp_dummy_magic_29_0.Vb1.n16 GNDA_2 0.242154f
C997 two_stage_opamp_dummy_magic_29_0.Vb1.t10 GNDA_2 0.030168f
C998 two_stage_opamp_dummy_magic_29_0.Vb1.t1 GNDA_2 0.030168f
C999 two_stage_opamp_dummy_magic_29_0.Vb1.n17 GNDA_2 0.065642f
C1000 two_stage_opamp_dummy_magic_29_0.Vb1.n18 GNDA_2 0.246742f
C1001 two_stage_opamp_dummy_magic_29_0.Vb1.t15 GNDA_2 0.047637f
C1002 two_stage_opamp_dummy_magic_29_0.Vb1.t26 GNDA_2 0.047637f
C1003 two_stage_opamp_dummy_magic_29_0.Vb1.t13 GNDA_2 0.047637f
C1004 two_stage_opamp_dummy_magic_29_0.Vb1.t25 GNDA_2 0.047637f
C1005 two_stage_opamp_dummy_magic_29_0.Vb1.t12 GNDA_2 0.047637f
C1006 two_stage_opamp_dummy_magic_29_0.Vb1.t23 GNDA_2 0.047637f
C1007 two_stage_opamp_dummy_magic_29_0.Vb1.t18 GNDA_2 0.047637f
C1008 two_stage_opamp_dummy_magic_29_0.Vb1.t24 GNDA_2 0.047637f
C1009 two_stage_opamp_dummy_magic_29_0.Vb1.t32 GNDA_2 0.047637f
C1010 two_stage_opamp_dummy_magic_29_0.Vb1.t22 GNDA_2 0.047637f
C1011 two_stage_opamp_dummy_magic_29_0.Vb1.t2 GNDA_2 0.040224f
C1012 two_stage_opamp_dummy_magic_29_0.Vb1.t11 GNDA_2 0.040224f
C1013 two_stage_opamp_dummy_magic_29_0.Vb1.n19 GNDA_2 0.091512f
C1014 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.t3 GNDA_2 0.011168f
C1015 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.t0 GNDA_2 0.011168f
C1016 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n0 GNDA_2 0.035122f
C1017 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.t1 GNDA_2 0.011168f
C1018 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.t2 GNDA_2 0.011168f
C1019 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n1 GNDA_2 0.023956f
C1020 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n2 GNDA_2 1.0883f
C1021 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.t14 GNDA_2 0.134451f
C1022 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n3 GNDA_2 0.054481f
C1023 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n4 GNDA_2 0.066839f
C1024 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.t7 GNDA_2 0.033504f
C1025 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.t12 GNDA_2 0.033504f
C1026 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n5 GNDA_2 0.071659f
C1027 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n6 GNDA_2 0.223527f
C1028 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.t8 GNDA_2 0.033504f
C1029 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.t13 GNDA_2 0.033504f
C1030 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n7 GNDA_2 0.071659f
C1031 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n8 GNDA_2 0.218077f
C1032 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n9 GNDA_2 0.090913f
C1033 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n10 GNDA_2 0.054481f
C1034 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.t10 GNDA_2 0.033504f
C1035 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.t4 GNDA_2 0.033504f
C1036 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n11 GNDA_2 0.071659f
C1037 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n12 GNDA_2 0.218077f
C1038 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n13 GNDA_2 0.038846f
C1039 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.t9 GNDA_2 0.033504f
C1040 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.t6 GNDA_2 0.033504f
C1041 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n14 GNDA_2 0.071659f
C1042 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n15 GNDA_2 0.218077f
C1043 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n16 GNDA_2 0.066839f
C1044 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.t11 GNDA_2 0.033504f
C1045 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.t5 GNDA_2 0.033504f
C1046 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n17 GNDA_2 0.071659f
C1047 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n18 GNDA_2 0.221113f
C1048 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n19 GNDA_2 0.154135f
C1049 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n20 GNDA_2 0.739467f
C1050 two_stage_opamp_dummy_magic_29_0.VD4.n0 GNDA_2 1.1096f
C1051 two_stage_opamp_dummy_magic_29_0.VD4.n1 GNDA_2 0.201538f
C1052 two_stage_opamp_dummy_magic_29_0.VD4.n2 GNDA_2 0.342878f
C1053 two_stage_opamp_dummy_magic_29_0.VD4.n3 GNDA_2 0.432296f
C1054 two_stage_opamp_dummy_magic_29_0.VD4.t6 GNDA_2 0.045031f
C1055 two_stage_opamp_dummy_magic_29_0.VD4.t9 GNDA_2 0.045031f
C1056 two_stage_opamp_dummy_magic_29_0.VD4.n4 GNDA_2 0.092115f
C1057 two_stage_opamp_dummy_magic_29_0.VD4.n5 GNDA_2 0.25692f
C1058 two_stage_opamp_dummy_magic_29_0.VD4.t25 GNDA_2 0.045031f
C1059 two_stage_opamp_dummy_magic_29_0.VD4.t21 GNDA_2 0.045031f
C1060 two_stage_opamp_dummy_magic_29_0.VD4.n6 GNDA_2 0.095624f
C1061 two_stage_opamp_dummy_magic_29_0.VD4.t2 GNDA_2 0.045031f
C1062 two_stage_opamp_dummy_magic_29_0.VD4.t0 GNDA_2 0.045031f
C1063 two_stage_opamp_dummy_magic_29_0.VD4.n7 GNDA_2 0.092115f
C1064 two_stage_opamp_dummy_magic_29_0.VD4.n8 GNDA_2 0.25692f
C1065 two_stage_opamp_dummy_magic_29_0.VD4.t27 GNDA_2 0.045031f
C1066 two_stage_opamp_dummy_magic_29_0.VD4.t29 GNDA_2 0.045031f
C1067 two_stage_opamp_dummy_magic_29_0.VD4.n9 GNDA_2 0.095624f
C1068 two_stage_opamp_dummy_magic_29_0.VD4.t7 GNDA_2 0.045031f
C1069 two_stage_opamp_dummy_magic_29_0.VD4.t1 GNDA_2 0.045031f
C1070 two_stage_opamp_dummy_magic_29_0.VD4.n10 GNDA_2 0.092115f
C1071 two_stage_opamp_dummy_magic_29_0.VD4.n11 GNDA_2 0.25692f
C1072 two_stage_opamp_dummy_magic_29_0.VD4.t13 GNDA_2 0.045031f
C1073 two_stage_opamp_dummy_magic_29_0.VD4.t19 GNDA_2 0.045031f
C1074 two_stage_opamp_dummy_magic_29_0.VD4.n12 GNDA_2 0.095624f
C1075 two_stage_opamp_dummy_magic_29_0.VD4.n13 GNDA_2 0.76157f
C1076 two_stage_opamp_dummy_magic_29_0.VD4.t34 GNDA_2 0.160181f
C1077 two_stage_opamp_dummy_magic_29_0.VD4.t35 GNDA_2 0.078836f
C1078 two_stage_opamp_dummy_magic_29_0.VD4.n14 GNDA_2 0.149757f
C1079 two_stage_opamp_dummy_magic_29_0.VD4.t37 GNDA_2 0.160181f
C1080 two_stage_opamp_dummy_magic_29_0.VD4.n15 GNDA_2 0.51334f
C1081 two_stage_opamp_dummy_magic_29_0.VD4.t36 GNDA_2 0.383839f
C1082 two_stage_opamp_dummy_magic_29_0.VD4.t30 GNDA_2 0.301063f
C1083 two_stage_opamp_dummy_magic_29_0.VD4.t16 GNDA_2 0.301063f
C1084 two_stage_opamp_dummy_magic_29_0.VD4.t24 GNDA_2 0.301063f
C1085 two_stage_opamp_dummy_magic_29_0.VD4.t20 GNDA_2 0.301063f
C1086 two_stage_opamp_dummy_magic_29_0.VD4.t26 GNDA_2 0.301063f
C1087 two_stage_opamp_dummy_magic_29_0.VD4.t28 GNDA_2 0.301063f
C1088 two_stage_opamp_dummy_magic_29_0.VD4.t12 GNDA_2 0.301063f
C1089 two_stage_opamp_dummy_magic_29_0.VD4.t18 GNDA_2 0.301063f
C1090 two_stage_opamp_dummy_magic_29_0.VD4.t14 GNDA_2 0.301063f
C1091 two_stage_opamp_dummy_magic_29_0.VD4.t22 GNDA_2 0.301063f
C1092 two_stage_opamp_dummy_magic_29_0.VD4.t33 GNDA_2 0.383839f
C1093 two_stage_opamp_dummy_magic_29_0.VD4.n16 GNDA_2 0.51334f
C1094 two_stage_opamp_dummy_magic_29_0.VD4.t32 GNDA_2 0.078836f
C1095 two_stage_opamp_dummy_magic_29_0.VD4.n17 GNDA_2 0.216535f
C1096 two_stage_opamp_dummy_magic_29_0.VD4.t15 GNDA_2 0.045031f
C1097 two_stage_opamp_dummy_magic_29_0.VD4.t23 GNDA_2 0.045031f
C1098 two_stage_opamp_dummy_magic_29_0.VD4.n18 GNDA_2 0.095624f
C1099 two_stage_opamp_dummy_magic_29_0.VD4.t11 GNDA_2 0.045031f
C1100 two_stage_opamp_dummy_magic_29_0.VD4.t5 GNDA_2 0.045031f
C1101 two_stage_opamp_dummy_magic_29_0.VD4.n19 GNDA_2 0.092115f
C1102 two_stage_opamp_dummy_magic_29_0.VD4.n20 GNDA_2 0.260153f
C1103 two_stage_opamp_dummy_magic_29_0.VD4.n21 GNDA_2 0.115041f
C1104 two_stage_opamp_dummy_magic_29_0.VD4.n22 GNDA_2 0.069429f
C1105 two_stage_opamp_dummy_magic_29_0.VD4.n23 GNDA_2 0.069429f
C1106 two_stage_opamp_dummy_magic_29_0.VD4.t8 GNDA_2 0.045031f
C1107 two_stage_opamp_dummy_magic_29_0.VD4.t3 GNDA_2 0.045031f
C1108 two_stage_opamp_dummy_magic_29_0.VD4.n24 GNDA_2 0.092115f
C1109 two_stage_opamp_dummy_magic_29_0.VD4.n25 GNDA_2 0.25692f
C1110 two_stage_opamp_dummy_magic_29_0.VD4.n26 GNDA_2 0.115041f
C1111 two_stage_opamp_dummy_magic_29_0.VD4.t4 GNDA_2 0.045031f
C1112 two_stage_opamp_dummy_magic_29_0.VD4.t10 GNDA_2 0.045031f
C1113 two_stage_opamp_dummy_magic_29_0.VD4.n27 GNDA_2 0.092115f
C1114 two_stage_opamp_dummy_magic_29_0.VD4.n28 GNDA_2 0.260153f
C1115 two_stage_opamp_dummy_magic_29_0.VD4.n29 GNDA_2 1.26176f
C1116 two_stage_opamp_dummy_magic_29_0.VD4.n30 GNDA_2 0.76157f
C1117 two_stage_opamp_dummy_magic_29_0.VD4.n31 GNDA_2 0.76157f
C1118 two_stage_opamp_dummy_magic_29_0.VD4.t31 GNDA_2 0.045031f
C1119 two_stage_opamp_dummy_magic_29_0.VD4.t17 GNDA_2 0.045031f
C1120 two_stage_opamp_dummy_magic_29_0.VD4.n32 GNDA_2 0.095624f
C1121 two_stage_opamp_dummy_magic_29_0.VD4.n33 GNDA_2 0.76157f
C1122 two_stage_opamp_dummy_magic_29_0.VD4.n34 GNDA_2 0.378259f
C1123 bgr_11_0.cap_res1.t5 GNDA_2 0.339883f
C1124 bgr_11_0.cap_res1.t17 GNDA_2 0.357788f
C1125 bgr_11_0.cap_res1.t9 GNDA_2 0.359085f
C1126 bgr_11_0.cap_res1.t12 GNDA_2 0.339883f
C1127 bgr_11_0.cap_res1.t19 GNDA_2 0.357788f
C1128 bgr_11_0.cap_res1.t16 GNDA_2 0.359085f
C1129 bgr_11_0.cap_res1.t4 GNDA_2 0.339883f
C1130 bgr_11_0.cap_res1.t15 GNDA_2 0.357788f
C1131 bgr_11_0.cap_res1.t8 GNDA_2 0.359085f
C1132 bgr_11_0.cap_res1.t0 GNDA_2 0.339883f
C1133 bgr_11_0.cap_res1.t7 GNDA_2 0.357788f
C1134 bgr_11_0.cap_res1.t1 GNDA_2 0.359085f
C1135 bgr_11_0.cap_res1.t2 GNDA_2 0.339883f
C1136 bgr_11_0.cap_res1.t14 GNDA_2 0.357788f
C1137 bgr_11_0.cap_res1.t6 GNDA_2 0.359085f
C1138 bgr_11_0.cap_res1.n0 GNDA_2 0.239826f
C1139 bgr_11_0.cap_res1.t10 GNDA_2 0.190986f
C1140 bgr_11_0.cap_res1.n1 GNDA_2 0.260216f
C1141 bgr_11_0.cap_res1.t3 GNDA_2 0.190986f
C1142 bgr_11_0.cap_res1.n2 GNDA_2 0.260216f
C1143 bgr_11_0.cap_res1.t11 GNDA_2 0.190986f
C1144 bgr_11_0.cap_res1.n3 GNDA_2 0.260216f
C1145 bgr_11_0.cap_res1.t18 GNDA_2 0.190986f
C1146 bgr_11_0.cap_res1.n4 GNDA_2 0.260216f
C1147 bgr_11_0.cap_res1.t13 GNDA_2 0.383393f
C1148 bgr_11_0.cap_res1.t20 GNDA_2 0.088196f
C1149 bgr_11_0.1st_Vout_1.n0 GNDA_2 0.191219f
C1150 bgr_11_0.1st_Vout_1.t27 GNDA_2 0.240974f
C1151 bgr_11_0.1st_Vout_1.t18 GNDA_2 0.236938f
C1152 bgr_11_0.1st_Vout_1.t14 GNDA_2 0.240974f
C1153 bgr_11_0.1st_Vout_1.t23 GNDA_2 0.236938f
C1154 bgr_11_0.1st_Vout_1.n1 GNDA_2 0.158859f
C1155 bgr_11_0.1st_Vout_1.n2 GNDA_2 0.203285f
C1156 bgr_11_0.1st_Vout_1.t32 GNDA_2 0.240974f
C1157 bgr_11_0.1st_Vout_1.t26 GNDA_2 0.236938f
C1158 bgr_11_0.1st_Vout_1.t22 GNDA_2 0.240974f
C1159 bgr_11_0.1st_Vout_1.t31 GNDA_2 0.236938f
C1160 bgr_11_0.1st_Vout_1.n3 GNDA_2 0.158859f
C1161 bgr_11_0.1st_Vout_1.n4 GNDA_2 0.247711f
C1162 bgr_11_0.1st_Vout_1.t25 GNDA_2 0.240974f
C1163 bgr_11_0.1st_Vout_1.t17 GNDA_2 0.236938f
C1164 bgr_11_0.1st_Vout_1.t12 GNDA_2 0.240974f
C1165 bgr_11_0.1st_Vout_1.t21 GNDA_2 0.236938f
C1166 bgr_11_0.1st_Vout_1.n5 GNDA_2 0.158859f
C1167 bgr_11_0.1st_Vout_1.n6 GNDA_2 0.247711f
C1168 bgr_11_0.1st_Vout_1.t16 GNDA_2 0.240974f
C1169 bgr_11_0.1st_Vout_1.t8 GNDA_2 0.236938f
C1170 bgr_11_0.1st_Vout_1.t7 GNDA_2 0.240974f
C1171 bgr_11_0.1st_Vout_1.t11 GNDA_2 0.236938f
C1172 bgr_11_0.1st_Vout_1.n7 GNDA_2 0.158859f
C1173 bgr_11_0.1st_Vout_1.n8 GNDA_2 0.247711f
C1174 bgr_11_0.1st_Vout_1.t24 GNDA_2 0.240974f
C1175 bgr_11_0.1st_Vout_1.t15 GNDA_2 0.236938f
C1176 bgr_11_0.1st_Vout_1.n9 GNDA_2 0.203285f
C1177 bgr_11_0.1st_Vout_1.t20 GNDA_2 0.236938f
C1178 bgr_11_0.1st_Vout_1.n10 GNDA_2 0.10366f
C1179 bgr_11_0.1st_Vout_1.t9 GNDA_2 0.236938f
C1180 bgr_11_0.1st_Vout_1.n11 GNDA_2 2.00975f
C1181 bgr_11_0.1st_Vout_1.t29 GNDA_2 0.01424f
C1182 bgr_11_0.1st_Vout_1.n12 GNDA_2 3.07165f
C1183 bgr_11_0.1st_Vout_1.n13 GNDA_2 0.012548f
C1184 bgr_11_0.1st_Vout_1.n14 GNDA_2 0.191219f
C1185 bgr_11_0.1st_Vout_1.n15 GNDA_2 0.017467f
C1186 bgr_11_0.1st_Vout_1.n16 GNDA_2 0.173289f
C1187 bgr_11_0.1st_Vout_1.n17 GNDA_2 0.012189f
C1188 bgr_11_0.1st_Vout_1.t3 GNDA_2 0.054022f
C1189 bgr_11_0.1st_Vout_1.n18 GNDA_2 0.173688f
C1190 bgr_11_0.1st_Vout_1.n19 GNDA_2 0.127946f
C1191 bgr_11_0.1st_Vout_1.n20 GNDA_2 0.017467f
C1192 bgr_11_0.1st_Vout_1.n21 GNDA_2 0.173289f
C1193 bgr_11_0.1st_Vout_1.n22 GNDA_2 0.012548f
C1194 bgr_11_0.1st_Vout_1.t13 GNDA_2 0.013988f
C1195 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n0 GNDA_2 0.028048f
C1196 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n1 GNDA_2 0.028314f
C1197 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n4 GNDA_2 0.028314f
C1198 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n5 GNDA_2 0.012047f
C1199 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n6 GNDA_2 0.371229f
C1200 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n7 GNDA_2 0.012745f
C1201 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n8 GNDA_2 0.087573f
C1202 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n9 GNDA_2 0.012047f
C1203 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n10 GNDA_2 0.360362f
C1204 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n11 GNDA_2 1.56671f
C1205 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n12 GNDA_2 3.15981f
C1206 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n14 GNDA_2 0.028314f
C1207 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n15 GNDA_2 0.028314f
C1208 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n16 GNDA_2 0.040701f
C1209 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n17 GNDA_2 0.040701f
C1210 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n18 GNDA_2 0.028314f
C1211 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n20 GNDA_2 0.028314f
C1212 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n21 GNDA_2 0.028314f
C1213 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n23 GNDA_2 0.164574f
C1214 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.t0 GNDA_2 0.071678f
C1215 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n24 GNDA_2 0.026892f
C1216 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n25 GNDA_2 0.03296f
C1217 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.t3 GNDA_2 0.011797f
C1218 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.t8 GNDA_2 0.011797f
C1219 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n26 GNDA_2 0.024121f
C1220 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n27 GNDA_2 0.081021f
C1221 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.t4 GNDA_2 0.011797f
C1222 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.t9 GNDA_2 0.011797f
C1223 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n28 GNDA_2 0.024121f
C1224 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n29 GNDA_2 0.078024f
C1225 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n30 GNDA_2 0.035812f
C1226 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n31 GNDA_2 0.026892f
C1227 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.t6 GNDA_2 0.011797f
C1228 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.t10 GNDA_2 0.011797f
C1229 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n32 GNDA_2 0.024121f
C1230 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n33 GNDA_2 0.078024f
C1231 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n34 GNDA_2 0.019315f
C1232 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.t5 GNDA_2 0.011797f
C1233 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.t2 GNDA_2 0.011797f
C1234 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n35 GNDA_2 0.024121f
C1235 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n36 GNDA_2 0.078024f
C1236 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n37 GNDA_2 0.03296f
C1237 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.t7 GNDA_2 0.011797f
C1238 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.t1 GNDA_2 0.011797f
C1239 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n38 GNDA_2 0.024121f
C1240 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n39 GNDA_2 0.079565f
C1241 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n40 GNDA_2 0.107479f
C1242 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n41 GNDA_2 0.56487f
C1243 two_stage_opamp_dummy_magic_29_0.X.n0 GNDA_2 0.162105f
C1244 two_stage_opamp_dummy_magic_29_0.X.n1 GNDA_2 0.237753f
C1245 two_stage_opamp_dummy_magic_29_0.X.n2 GNDA_2 0.417266f
C1246 two_stage_opamp_dummy_magic_29_0.X.n3 GNDA_2 0.388675f
C1247 two_stage_opamp_dummy_magic_29_0.X.n4 GNDA_2 0.237753f
C1248 two_stage_opamp_dummy_magic_29_0.X.n5 GNDA_2 0.237753f
C1249 two_stage_opamp_dummy_magic_29_0.X.n9 GNDA_2 0.074105f
C1250 two_stage_opamp_dummy_magic_29_0.X.n10 GNDA_2 0.083312f
C1251 two_stage_opamp_dummy_magic_29_0.X.n11 GNDA_2 0.083312f
C1252 two_stage_opamp_dummy_magic_29_0.X.t2 GNDA_2 0.054035f
C1253 two_stage_opamp_dummy_magic_29_0.X.t20 GNDA_2 0.054035f
C1254 two_stage_opamp_dummy_magic_29_0.X.n12 GNDA_2 0.110534f
C1255 two_stage_opamp_dummy_magic_29_0.X.n13 GNDA_2 0.35586f
C1256 two_stage_opamp_dummy_magic_29_0.X.n14 GNDA_2 0.138043f
C1257 two_stage_opamp_dummy_magic_29_0.X.t15 GNDA_2 0.054035f
C1258 two_stage_opamp_dummy_magic_29_0.X.t21 GNDA_2 0.054035f
C1259 two_stage_opamp_dummy_magic_29_0.X.n15 GNDA_2 0.110534f
C1260 two_stage_opamp_dummy_magic_29_0.X.n16 GNDA_2 0.348103f
C1261 two_stage_opamp_dummy_magic_29_0.X.n17 GNDA_2 0.138043f
C1262 two_stage_opamp_dummy_magic_29_0.X.t19 GNDA_2 0.054035f
C1263 two_stage_opamp_dummy_magic_29_0.X.t18 GNDA_2 0.054035f
C1264 two_stage_opamp_dummy_magic_29_0.X.n18 GNDA_2 0.110534f
C1265 two_stage_opamp_dummy_magic_29_0.X.n19 GNDA_2 0.348103f
C1266 two_stage_opamp_dummy_magic_29_0.X.n20 GNDA_2 0.083312f
C1267 two_stage_opamp_dummy_magic_29_0.X.n21 GNDA_2 0.083312f
C1268 two_stage_opamp_dummy_magic_29_0.X.t13 GNDA_2 0.054035f
C1269 two_stage_opamp_dummy_magic_29_0.X.t16 GNDA_2 0.054035f
C1270 two_stage_opamp_dummy_magic_29_0.X.n22 GNDA_2 0.110534f
C1271 two_stage_opamp_dummy_magic_29_0.X.n23 GNDA_2 0.348103f
C1272 two_stage_opamp_dummy_magic_29_0.X.n24 GNDA_2 0.083312f
C1273 two_stage_opamp_dummy_magic_29_0.X.t17 GNDA_2 0.054035f
C1274 two_stage_opamp_dummy_magic_29_0.X.t14 GNDA_2 0.054035f
C1275 two_stage_opamp_dummy_magic_29_0.X.n25 GNDA_2 0.110534f
C1276 two_stage_opamp_dummy_magic_29_0.X.n26 GNDA_2 0.348103f
C1277 two_stage_opamp_dummy_magic_29_0.X.n27 GNDA_2 0.138043f
C1278 two_stage_opamp_dummy_magic_29_0.X.t12 GNDA_2 0.054035f
C1279 two_stage_opamp_dummy_magic_29_0.X.t23 GNDA_2 0.054035f
C1280 two_stage_opamp_dummy_magic_29_0.X.n28 GNDA_2 0.110534f
C1281 two_stage_opamp_dummy_magic_29_0.X.n29 GNDA_2 0.351981f
C1282 two_stage_opamp_dummy_magic_29_0.X.n30 GNDA_2 0.220124f
C1283 two_stage_opamp_dummy_magic_29_0.X.n31 GNDA_2 0.172911f
C1284 two_stage_opamp_dummy_magic_29_0.X.n33 GNDA_2 0.074105f
C1285 two_stage_opamp_dummy_magic_29_0.X.n34 GNDA_2 0.074105f
C1286 two_stage_opamp_dummy_magic_29_0.X.t44 GNDA_2 0.049789f
C1287 two_stage_opamp_dummy_magic_29_0.X.t29 GNDA_2 0.056602f
C1288 two_stage_opamp_dummy_magic_29_0.X.n36 GNDA_2 0.046161f
C1289 two_stage_opamp_dummy_magic_29_0.X.t26 GNDA_2 0.049789f
C1290 two_stage_opamp_dummy_magic_29_0.X.t40 GNDA_2 0.049789f
C1291 two_stage_opamp_dummy_magic_29_0.X.t52 GNDA_2 0.049789f
C1292 two_stage_opamp_dummy_magic_29_0.X.t35 GNDA_2 0.049789f
C1293 two_stage_opamp_dummy_magic_29_0.X.t48 GNDA_2 0.049789f
C1294 two_stage_opamp_dummy_magic_29_0.X.t36 GNDA_2 0.049789f
C1295 two_stage_opamp_dummy_magic_29_0.X.t49 GNDA_2 0.049789f
C1296 two_stage_opamp_dummy_magic_29_0.X.t33 GNDA_2 0.056602f
C1297 two_stage_opamp_dummy_magic_29_0.X.n37 GNDA_2 0.051082f
C1298 two_stage_opamp_dummy_magic_29_0.X.n38 GNDA_2 0.031263f
C1299 two_stage_opamp_dummy_magic_29_0.X.n39 GNDA_2 0.031263f
C1300 two_stage_opamp_dummy_magic_29_0.X.n40 GNDA_2 0.031263f
C1301 two_stage_opamp_dummy_magic_29_0.X.n41 GNDA_2 0.031263f
C1302 two_stage_opamp_dummy_magic_29_0.X.n42 GNDA_2 0.031263f
C1303 two_stage_opamp_dummy_magic_29_0.X.n43 GNDA_2 0.026342f
C1304 two_stage_opamp_dummy_magic_29_0.X.n44 GNDA_2 0.012791f
C1305 two_stage_opamp_dummy_magic_29_0.X.t46 GNDA_2 0.032421f
C1306 two_stage_opamp_dummy_magic_29_0.X.t31 GNDA_2 0.039368f
C1307 two_stage_opamp_dummy_magic_29_0.X.n45 GNDA_2 0.034447f
C1308 two_stage_opamp_dummy_magic_29_0.X.t28 GNDA_2 0.032421f
C1309 two_stage_opamp_dummy_magic_29_0.X.t43 GNDA_2 0.032421f
C1310 two_stage_opamp_dummy_magic_29_0.X.t25 GNDA_2 0.032421f
C1311 two_stage_opamp_dummy_magic_29_0.X.t38 GNDA_2 0.032421f
C1312 two_stage_opamp_dummy_magic_29_0.X.t50 GNDA_2 0.032421f
C1313 two_stage_opamp_dummy_magic_29_0.X.t39 GNDA_2 0.032421f
C1314 two_stage_opamp_dummy_magic_29_0.X.t51 GNDA_2 0.032421f
C1315 two_stage_opamp_dummy_magic_29_0.X.t34 GNDA_2 0.039368f
C1316 two_stage_opamp_dummy_magic_29_0.X.n46 GNDA_2 0.039368f
C1317 two_stage_opamp_dummy_magic_29_0.X.n47 GNDA_2 0.025474f
C1318 two_stage_opamp_dummy_magic_29_0.X.n48 GNDA_2 0.025474f
C1319 two_stage_opamp_dummy_magic_29_0.X.n49 GNDA_2 0.025474f
C1320 two_stage_opamp_dummy_magic_29_0.X.n50 GNDA_2 0.025474f
C1321 two_stage_opamp_dummy_magic_29_0.X.n51 GNDA_2 0.025474f
C1322 two_stage_opamp_dummy_magic_29_0.X.n52 GNDA_2 0.020552f
C1323 two_stage_opamp_dummy_magic_29_0.X.n53 GNDA_2 0.012791f
C1324 two_stage_opamp_dummy_magic_29_0.X.n54 GNDA_2 0.079789f
C1325 two_stage_opamp_dummy_magic_29_0.X.n56 GNDA_2 0.074105f
C1326 two_stage_opamp_dummy_magic_29_0.X.t8 GNDA_2 0.640789f
C1327 two_stage_opamp_dummy_magic_29_0.X.n57 GNDA_2 0.074105f
C1328 two_stage_opamp_dummy_magic_29_0.X.n58 GNDA_2 0.074105f
C1329 two_stage_opamp_dummy_magic_29_0.X.n59 GNDA_2 0.073409f
C1330 two_stage_opamp_dummy_magic_29_0.X.n60 GNDA_2 0.687542f
C1331 two_stage_opamp_dummy_magic_29_0.X.n62 GNDA_2 0.643787f
C1332 two_stage_opamp_dummy_magic_29_0.X.n63 GNDA_2 0.024538f
C1333 two_stage_opamp_dummy_magic_29_0.X.n64 GNDA_2 0.024702f
C1334 two_stage_opamp_dummy_magic_29_0.X.n65 GNDA_2 0.024702f
C1335 two_stage_opamp_dummy_magic_29_0.X.t27 GNDA_2 0.101894f
C1336 two_stage_opamp_dummy_magic_29_0.X.t45 GNDA_2 0.101894f
C1337 two_stage_opamp_dummy_magic_29_0.X.t30 GNDA_2 0.101894f
C1338 two_stage_opamp_dummy_magic_29_0.X.t47 GNDA_2 0.101894f
C1339 two_stage_opamp_dummy_magic_29_0.X.t32 GNDA_2 0.108524f
C1340 two_stage_opamp_dummy_magic_29_0.X.n66 GNDA_2 0.086001f
C1341 two_stage_opamp_dummy_magic_29_0.X.n67 GNDA_2 0.048631f
C1342 two_stage_opamp_dummy_magic_29_0.X.n68 GNDA_2 0.048631f
C1343 two_stage_opamp_dummy_magic_29_0.X.n69 GNDA_2 0.04371f
C1344 two_stage_opamp_dummy_magic_29_0.X.t41 GNDA_2 0.101894f
C1345 two_stage_opamp_dummy_magic_29_0.X.t53 GNDA_2 0.101894f
C1346 two_stage_opamp_dummy_magic_29_0.X.t42 GNDA_2 0.101894f
C1347 two_stage_opamp_dummy_magic_29_0.X.t54 GNDA_2 0.101894f
C1348 two_stage_opamp_dummy_magic_29_0.X.t37 GNDA_2 0.108524f
C1349 two_stage_opamp_dummy_magic_29_0.X.n70 GNDA_2 0.086001f
C1350 two_stage_opamp_dummy_magic_29_0.X.n71 GNDA_2 0.048631f
C1351 two_stage_opamp_dummy_magic_29_0.X.n72 GNDA_2 0.048631f
C1352 two_stage_opamp_dummy_magic_29_0.X.n73 GNDA_2 0.04371f
C1353 two_stage_opamp_dummy_magic_29_0.X.n74 GNDA_2 0.010496f
C1354 two_stage_opamp_dummy_magic_29_0.X.n75 GNDA_2 0.024866f
C1355 two_stage_opamp_dummy_magic_29_0.X.n76 GNDA_2 0.058532f
C1356 two_stage_opamp_dummy_magic_29_0.X.n77 GNDA_2 0.033384f
C1357 two_stage_opamp_dummy_magic_29_0.X.n78 GNDA_2 0.037886f
C1358 two_stage_opamp_dummy_magic_29_0.X.n79 GNDA_2 1.02357f
C1359 two_stage_opamp_dummy_magic_29_0.X.n80 GNDA_2 0.453893f
C1360 two_stage_opamp_dummy_magic_29_0.X.n81 GNDA_2 2.18995f
C1361 two_stage_opamp_dummy_magic_29_0.X.n82 GNDA_2 0.074105f
C1362 two_stage_opamp_dummy_magic_29_0.X.n84 GNDA_2 0.463156f
C1363 two_stage_opamp_dummy_magic_29_0.X.n85 GNDA_2 0.463156f
C1364 two_stage_opamp_dummy_magic_29_0.X.n86 GNDA_2 0.074105f
C1365 two_stage_opamp_dummy_magic_29_0.X.n88 GNDA_2 0.074105f
C1366 two_stage_opamp_dummy_magic_29_0.X.n90 GNDA_2 0.074105f
C1367 two_stage_opamp_dummy_magic_29_0.X.n92 GNDA_2 0.074105f
C1368 two_stage_opamp_dummy_magic_29_0.X.n93 GNDA_2 0.172911f
C1369 two_stage_opamp_dummy_magic_29_0.X.n95 GNDA_2 0.619675f
C1370 two_stage_opamp_dummy_magic_29_0.X.n97 GNDA_2 1.3941f
C1371 two_stage_opamp_dummy_magic_29_0.X.n98 GNDA_2 1.42652f
C1372 two_stage_opamp_dummy_magic_29_0.X.n99 GNDA_2 0.237753f
C1373 two_stage_opamp_dummy_magic_29_0.X.n100 GNDA_2 0.237753f
C1374 two_stage_opamp_dummy_magic_29_0.X.n101 GNDA_2 0.237753f
C1375 two_stage_opamp_dummy_magic_29_0.X.n102 GNDA_2 0.417266f
C1376 two_stage_opamp_dummy_magic_29_0.X.n103 GNDA_2 0.146616f
C1377 two_stage_opamp_dummy_magic_29_0.X.n104 GNDA_2 0.08603f
C1378 two_stage_opamp_dummy_magic_29_0.X.n105 GNDA_2 0.08603f
C1379 two_stage_opamp_dummy_magic_29_0.X.n106 GNDA_2 0.496725f
C1380 two_stage_opamp_dummy_magic_29_0.X.n107 GNDA_2 0.08603f
C1381 two_stage_opamp_dummy_magic_29_0.X.t7 GNDA_2 0.023158f
C1382 two_stage_opamp_dummy_magic_29_0.X.t10 GNDA_2 0.023158f
C1383 two_stage_opamp_dummy_magic_29_0.X.n108 GNDA_2 0.068053f
C1384 two_stage_opamp_dummy_magic_29_0.X.t11 GNDA_2 0.023158f
C1385 two_stage_opamp_dummy_magic_29_0.X.t9 GNDA_2 0.023158f
C1386 two_stage_opamp_dummy_magic_29_0.X.n109 GNDA_2 0.066733f
C1387 two_stage_opamp_dummy_magic_29_0.X.n110 GNDA_2 0.44107f
C1388 two_stage_opamp_dummy_magic_29_0.X.t24 GNDA_2 0.023158f
C1389 two_stage_opamp_dummy_magic_29_0.X.t3 GNDA_2 0.023158f
C1390 two_stage_opamp_dummy_magic_29_0.X.n111 GNDA_2 0.066733f
C1391 two_stage_opamp_dummy_magic_29_0.X.n112 GNDA_2 0.232002f
C1392 two_stage_opamp_dummy_magic_29_0.X.t4 GNDA_2 0.023158f
C1393 two_stage_opamp_dummy_magic_29_0.X.t5 GNDA_2 0.023158f
C1394 two_stage_opamp_dummy_magic_29_0.X.n113 GNDA_2 0.066733f
C1395 two_stage_opamp_dummy_magic_29_0.X.n114 GNDA_2 0.232002f
C1396 two_stage_opamp_dummy_magic_29_0.X.t1 GNDA_2 0.023158f
C1397 two_stage_opamp_dummy_magic_29_0.X.t22 GNDA_2 0.023158f
C1398 two_stage_opamp_dummy_magic_29_0.X.n115 GNDA_2 0.066733f
C1399 two_stage_opamp_dummy_magic_29_0.X.n116 GNDA_2 0.232002f
C1400 two_stage_opamp_dummy_magic_29_0.X.t0 GNDA_2 0.023158f
C1401 two_stage_opamp_dummy_magic_29_0.X.t6 GNDA_2 0.023158f
C1402 two_stage_opamp_dummy_magic_29_0.X.n117 GNDA_2 0.066733f
C1403 two_stage_opamp_dummy_magic_29_0.X.n118 GNDA_2 0.431159f
C1404 two_stage_opamp_dummy_magic_29_0.X.n119 GNDA_2 0.287483f
C1405 two_stage_opamp_dummy_magic_29_0.X.n120 GNDA_2 0.644415f
C1406 two_stage_opamp_dummy_magic_29_0.X.n121 GNDA_2 0.815021f
C1407 two_stage_opamp_dummy_magic_29_0.X.n122 GNDA_2 0.237753f
C1408 two_stage_opamp_dummy_magic_29_0.X.n123 GNDA_2 0.417266f
C1409 two_stage_opamp_dummy_magic_29_0.X.n124 GNDA_2 0.237753f
C1410 two_stage_opamp_dummy_magic_29_0.X.n125 GNDA_2 0.194525f
C1411 two_stage_opamp_dummy_magic_29_0.cap_res_X.t97 GNDA_2 0.358056f
C1412 two_stage_opamp_dummy_magic_29_0.cap_res_X.t75 GNDA_2 0.359353f
C1413 two_stage_opamp_dummy_magic_29_0.cap_res_X.t63 GNDA_2 0.358056f
C1414 two_stage_opamp_dummy_magic_29_0.cap_res_X.t37 GNDA_2 0.359353f
C1415 two_stage_opamp_dummy_magic_29_0.cap_res_X.t92 GNDA_2 0.358056f
C1416 two_stage_opamp_dummy_magic_29_0.cap_res_X.t117 GNDA_2 0.359353f
C1417 two_stage_opamp_dummy_magic_29_0.cap_res_X.t20 GNDA_2 0.358056f
C1418 two_stage_opamp_dummy_magic_29_0.cap_res_X.t72 GNDA_2 0.359353f
C1419 two_stage_opamp_dummy_magic_29_0.cap_res_X.t52 GNDA_2 0.358056f
C1420 two_stage_opamp_dummy_magic_29_0.cap_res_X.t141 GNDA_2 0.359353f
C1421 two_stage_opamp_dummy_magic_29_0.cap_res_X.t60 GNDA_2 0.358056f
C1422 two_stage_opamp_dummy_magic_29_0.cap_res_X.t110 GNDA_2 0.359353f
C1423 two_stage_opamp_dummy_magic_29_0.cap_res_X.t89 GNDA_2 0.358056f
C1424 two_stage_opamp_dummy_magic_29_0.cap_res_X.t38 GNDA_2 0.359353f
C1425 two_stage_opamp_dummy_magic_29_0.cap_res_X.t23 GNDA_2 0.358056f
C1426 two_stage_opamp_dummy_magic_29_0.cap_res_X.t77 GNDA_2 0.359353f
C1427 two_stage_opamp_dummy_magic_29_0.cap_res_X.t58 GNDA_2 0.358056f
C1428 two_stage_opamp_dummy_magic_29_0.cap_res_X.t2 GNDA_2 0.359353f
C1429 two_stage_opamp_dummy_magic_29_0.cap_res_X.t65 GNDA_2 0.358056f
C1430 two_stage_opamp_dummy_magic_29_0.cap_res_X.t116 GNDA_2 0.359353f
C1431 two_stage_opamp_dummy_magic_29_0.cap_res_X.t96 GNDA_2 0.358056f
C1432 two_stage_opamp_dummy_magic_29_0.cap_res_X.t43 GNDA_2 0.359353f
C1433 two_stage_opamp_dummy_magic_29_0.cap_res_X.t105 GNDA_2 0.358056f
C1434 two_stage_opamp_dummy_magic_29_0.cap_res_X.t16 GNDA_2 0.359353f
C1435 two_stage_opamp_dummy_magic_29_0.cap_res_X.t135 GNDA_2 0.358056f
C1436 two_stage_opamp_dummy_magic_29_0.cap_res_X.t84 GNDA_2 0.359353f
C1437 two_stage_opamp_dummy_magic_29_0.cap_res_X.t71 GNDA_2 0.358056f
C1438 two_stage_opamp_dummy_magic_29_0.cap_res_X.t121 GNDA_2 0.359353f
C1439 two_stage_opamp_dummy_magic_29_0.cap_res_X.t103 GNDA_2 0.358056f
C1440 two_stage_opamp_dummy_magic_29_0.cap_res_X.t51 GNDA_2 0.359353f
C1441 two_stage_opamp_dummy_magic_29_0.cap_res_X.t108 GNDA_2 0.358056f
C1442 two_stage_opamp_dummy_magic_29_0.cap_res_X.t21 GNDA_2 0.359353f
C1443 two_stage_opamp_dummy_magic_29_0.cap_res_X.t142 GNDA_2 0.358056f
C1444 two_stage_opamp_dummy_magic_29_0.cap_res_X.t88 GNDA_2 0.359353f
C1445 two_stage_opamp_dummy_magic_29_0.cap_res_X.t7 GNDA_2 0.358056f
C1446 two_stage_opamp_dummy_magic_29_0.cap_res_X.t61 GNDA_2 0.359353f
C1447 two_stage_opamp_dummy_magic_29_0.cap_res_X.t40 GNDA_2 0.358056f
C1448 two_stage_opamp_dummy_magic_29_0.cap_res_X.t127 GNDA_2 0.359353f
C1449 two_stage_opamp_dummy_magic_29_0.cap_res_X.t48 GNDA_2 0.358056f
C1450 two_stage_opamp_dummy_magic_29_0.cap_res_X.t100 GNDA_2 0.359353f
C1451 two_stage_opamp_dummy_magic_29_0.cap_res_X.t81 GNDA_2 0.358056f
C1452 two_stage_opamp_dummy_magic_29_0.cap_res_X.t27 GNDA_2 0.359353f
C1453 two_stage_opamp_dummy_magic_29_0.cap_res_X.t13 GNDA_2 0.358056f
C1454 two_stage_opamp_dummy_magic_29_0.cap_res_X.t68 GNDA_2 0.359353f
C1455 two_stage_opamp_dummy_magic_29_0.cap_res_X.t45 GNDA_2 0.358056f
C1456 two_stage_opamp_dummy_magic_29_0.cap_res_X.t134 GNDA_2 0.359353f
C1457 two_stage_opamp_dummy_magic_29_0.cap_res_X.t54 GNDA_2 0.358056f
C1458 two_stage_opamp_dummy_magic_29_0.cap_res_X.t106 GNDA_2 0.359353f
C1459 two_stage_opamp_dummy_magic_29_0.cap_res_X.t85 GNDA_2 0.358056f
C1460 two_stage_opamp_dummy_magic_29_0.cap_res_X.t34 GNDA_2 0.359353f
C1461 two_stage_opamp_dummy_magic_29_0.cap_res_X.t93 GNDA_2 0.358056f
C1462 two_stage_opamp_dummy_magic_29_0.cap_res_X.t0 GNDA_2 0.359353f
C1463 two_stage_opamp_dummy_magic_29_0.cap_res_X.t125 GNDA_2 0.358056f
C1464 two_stage_opamp_dummy_magic_29_0.cap_res_X.t76 GNDA_2 0.359353f
C1465 two_stage_opamp_dummy_magic_29_0.cap_res_X.t59 GNDA_2 0.358056f
C1466 two_stage_opamp_dummy_magic_29_0.cap_res_X.t111 GNDA_2 0.359353f
C1467 two_stage_opamp_dummy_magic_29_0.cap_res_X.t90 GNDA_2 0.358056f
C1468 two_stage_opamp_dummy_magic_29_0.cap_res_X.t39 GNDA_2 0.359353f
C1469 two_stage_opamp_dummy_magic_29_0.cap_res_X.t74 GNDA_2 0.358056f
C1470 two_stage_opamp_dummy_magic_29_0.cap_res_X.t115 GNDA_2 0.359353f
C1471 two_stage_opamp_dummy_magic_29_0.cap_res_X.t57 GNDA_2 0.358056f
C1472 two_stage_opamp_dummy_magic_29_0.cap_res_X.t12 GNDA_2 0.359353f
C1473 two_stage_opamp_dummy_magic_29_0.cap_res_X.t87 GNDA_2 0.358056f
C1474 two_stage_opamp_dummy_magic_29_0.cap_res_X.t138 GNDA_2 0.359353f
C1475 two_stage_opamp_dummy_magic_29_0.cap_res_X.t120 GNDA_2 0.358056f
C1476 two_stage_opamp_dummy_magic_29_0.cap_res_X.t70 GNDA_2 0.359353f
C1477 two_stage_opamp_dummy_magic_29_0.cap_res_X.t124 GNDA_2 0.358056f
C1478 two_stage_opamp_dummy_magic_29_0.cap_res_X.t32 GNDA_2 0.359353f
C1479 two_stage_opamp_dummy_magic_29_0.cap_res_X.t14 GNDA_2 0.358056f
C1480 two_stage_opamp_dummy_magic_29_0.cap_res_X.t104 GNDA_2 0.359353f
C1481 two_stage_opamp_dummy_magic_29_0.cap_res_X.t118 GNDA_2 0.358056f
C1482 two_stage_opamp_dummy_magic_29_0.cap_res_X.t95 GNDA_2 0.359353f
C1483 two_stage_opamp_dummy_magic_29_0.cap_res_X.t6 GNDA_2 0.358056f
C1484 two_stage_opamp_dummy_magic_29_0.cap_res_X.t47 GNDA_2 0.375611f
C1485 two_stage_opamp_dummy_magic_29_0.cap_res_X.t28 GNDA_2 0.358056f
C1486 two_stage_opamp_dummy_magic_29_0.cap_res_X.t73 GNDA_2 0.192319f
C1487 two_stage_opamp_dummy_magic_29_0.cap_res_X.n0 GNDA_2 0.205829f
C1488 two_stage_opamp_dummy_magic_29_0.cap_res_X.t11 GNDA_2 0.358056f
C1489 two_stage_opamp_dummy_magic_29_0.cap_res_X.t53 GNDA_2 0.192319f
C1490 two_stage_opamp_dummy_magic_29_0.cap_res_X.n1 GNDA_2 0.204169f
C1491 two_stage_opamp_dummy_magic_29_0.cap_res_X.t114 GNDA_2 0.358056f
C1492 two_stage_opamp_dummy_magic_29_0.cap_res_X.t15 GNDA_2 0.192319f
C1493 two_stage_opamp_dummy_magic_29_0.cap_res_X.n2 GNDA_2 0.204169f
C1494 two_stage_opamp_dummy_magic_29_0.cap_res_X.t136 GNDA_2 0.358056f
C1495 two_stage_opamp_dummy_magic_29_0.cap_res_X.t35 GNDA_2 0.192319f
C1496 two_stage_opamp_dummy_magic_29_0.cap_res_X.n3 GNDA_2 0.204169f
C1497 two_stage_opamp_dummy_magic_29_0.cap_res_X.t98 GNDA_2 0.358056f
C1498 two_stage_opamp_dummy_magic_29_0.cap_res_X.t139 GNDA_2 0.192319f
C1499 two_stage_opamp_dummy_magic_29_0.cap_res_X.n4 GNDA_2 0.204169f
C1500 two_stage_opamp_dummy_magic_29_0.cap_res_X.t62 GNDA_2 0.358056f
C1501 two_stage_opamp_dummy_magic_29_0.cap_res_X.t102 GNDA_2 0.192319f
C1502 two_stage_opamp_dummy_magic_29_0.cap_res_X.n5 GNDA_2 0.204169f
C1503 two_stage_opamp_dummy_magic_29_0.cap_res_X.t22 GNDA_2 0.358056f
C1504 two_stage_opamp_dummy_magic_29_0.cap_res_X.t64 GNDA_2 0.192319f
C1505 two_stage_opamp_dummy_magic_29_0.cap_res_X.n6 GNDA_2 0.204169f
C1506 two_stage_opamp_dummy_magic_29_0.cap_res_X.t42 GNDA_2 0.358056f
C1507 two_stage_opamp_dummy_magic_29_0.cap_res_X.t83 GNDA_2 0.192319f
C1508 two_stage_opamp_dummy_magic_29_0.cap_res_X.n7 GNDA_2 0.204169f
C1509 two_stage_opamp_dummy_magic_29_0.cap_res_X.t4 GNDA_2 0.358056f
C1510 two_stage_opamp_dummy_magic_29_0.cap_res_X.t46 GNDA_2 0.192319f
C1511 two_stage_opamp_dummy_magic_29_0.cap_res_X.n8 GNDA_2 0.204169f
C1512 two_stage_opamp_dummy_magic_29_0.cap_res_X.t109 GNDA_2 0.358056f
C1513 two_stage_opamp_dummy_magic_29_0.cap_res_X.t8 GNDA_2 0.192319f
C1514 two_stage_opamp_dummy_magic_29_0.cap_res_X.n9 GNDA_2 0.204169f
C1515 two_stage_opamp_dummy_magic_29_0.cap_res_X.t128 GNDA_2 0.358056f
C1516 two_stage_opamp_dummy_magic_29_0.cap_res_X.t29 GNDA_2 0.192319f
C1517 two_stage_opamp_dummy_magic_29_0.cap_res_X.n10 GNDA_2 0.204169f
C1518 two_stage_opamp_dummy_magic_29_0.cap_res_X.t78 GNDA_2 0.358056f
C1519 two_stage_opamp_dummy_magic_29_0.cap_res_X.t56 GNDA_2 0.359353f
C1520 two_stage_opamp_dummy_magic_29_0.cap_res_X.t91 GNDA_2 0.173103f
C1521 two_stage_opamp_dummy_magic_29_0.cap_res_X.n11 GNDA_2 0.223277f
C1522 two_stage_opamp_dummy_magic_29_0.cap_res_X.t130 GNDA_2 0.191129f
C1523 two_stage_opamp_dummy_magic_29_0.cap_res_X.n12 GNDA_2 0.242493f
C1524 two_stage_opamp_dummy_magic_29_0.cap_res_X.t69 GNDA_2 0.191129f
C1525 two_stage_opamp_dummy_magic_29_0.cap_res_X.n13 GNDA_2 0.260411f
C1526 two_stage_opamp_dummy_magic_29_0.cap_res_X.t33 GNDA_2 0.191129f
C1527 two_stage_opamp_dummy_magic_29_0.cap_res_X.n14 GNDA_2 0.260411f
C1528 two_stage_opamp_dummy_magic_29_0.cap_res_X.t66 GNDA_2 0.191129f
C1529 two_stage_opamp_dummy_magic_29_0.cap_res_X.n15 GNDA_2 0.260411f
C1530 two_stage_opamp_dummy_magic_29_0.cap_res_X.t3 GNDA_2 0.191129f
C1531 two_stage_opamp_dummy_magic_29_0.cap_res_X.n16 GNDA_2 0.260411f
C1532 two_stage_opamp_dummy_magic_29_0.cap_res_X.t36 GNDA_2 0.191129f
C1533 two_stage_opamp_dummy_magic_29_0.cap_res_X.n17 GNDA_2 0.260411f
C1534 two_stage_opamp_dummy_magic_29_0.cap_res_X.t140 GNDA_2 0.191129f
C1535 two_stage_opamp_dummy_magic_29_0.cap_res_X.n18 GNDA_2 0.260411f
C1536 two_stage_opamp_dummy_magic_29_0.cap_res_X.t101 GNDA_2 0.191129f
C1537 two_stage_opamp_dummy_magic_29_0.cap_res_X.n19 GNDA_2 0.260411f
C1538 two_stage_opamp_dummy_magic_29_0.cap_res_X.t133 GNDA_2 0.191129f
C1539 two_stage_opamp_dummy_magic_29_0.cap_res_X.n20 GNDA_2 0.260411f
C1540 two_stage_opamp_dummy_magic_29_0.cap_res_X.t94 GNDA_2 0.191129f
C1541 two_stage_opamp_dummy_magic_29_0.cap_res_X.n21 GNDA_2 0.260411f
C1542 two_stage_opamp_dummy_magic_29_0.cap_res_X.t55 GNDA_2 0.191129f
C1543 two_stage_opamp_dummy_magic_29_0.cap_res_X.n22 GNDA_2 0.260411f
C1544 two_stage_opamp_dummy_magic_29_0.cap_res_X.t17 GNDA_2 0.191129f
C1545 two_stage_opamp_dummy_magic_29_0.cap_res_X.n23 GNDA_2 0.260411f
C1546 two_stage_opamp_dummy_magic_29_0.cap_res_X.t49 GNDA_2 0.191129f
C1547 two_stage_opamp_dummy_magic_29_0.cap_res_X.n24 GNDA_2 0.260411f
C1548 two_stage_opamp_dummy_magic_29_0.cap_res_X.t9 GNDA_2 0.191129f
C1549 two_stage_opamp_dummy_magic_29_0.cap_res_X.n25 GNDA_2 0.260411f
C1550 two_stage_opamp_dummy_magic_29_0.cap_res_X.t112 GNDA_2 0.191129f
C1551 two_stage_opamp_dummy_magic_29_0.cap_res_X.n26 GNDA_2 0.260411f
C1552 two_stage_opamp_dummy_magic_29_0.cap_res_X.t1 GNDA_2 0.191129f
C1553 two_stage_opamp_dummy_magic_29_0.cap_res_X.n27 GNDA_2 0.260411f
C1554 two_stage_opamp_dummy_magic_29_0.cap_res_X.t107 GNDA_2 0.191129f
C1555 two_stage_opamp_dummy_magic_29_0.cap_res_X.n28 GNDA_2 0.260411f
C1556 two_stage_opamp_dummy_magic_29_0.cap_res_X.t79 GNDA_2 0.191129f
C1557 two_stage_opamp_dummy_magic_29_0.cap_res_X.n29 GNDA_2 0.260411f
C1558 two_stage_opamp_dummy_magic_29_0.cap_res_X.t113 GNDA_2 0.191129f
C1559 two_stage_opamp_dummy_magic_29_0.cap_res_X.n30 GNDA_2 0.240005f
C1560 two_stage_opamp_dummy_magic_29_0.cap_res_X.t10 GNDA_2 0.359353f
C1561 two_stage_opamp_dummy_magic_29_0.cap_res_X.t126 GNDA_2 0.359353f
C1562 two_stage_opamp_dummy_magic_29_0.cap_res_X.t86 GNDA_2 0.358056f
C1563 two_stage_opamp_dummy_magic_29_0.cap_res_X.t129 GNDA_2 0.377272f
C1564 two_stage_opamp_dummy_magic_29_0.cap_res_X.t24 GNDA_2 0.192319f
C1565 two_stage_opamp_dummy_magic_29_0.cap_res_X.n31 GNDA_2 0.222087f
C1566 two_stage_opamp_dummy_magic_29_0.cap_res_X.t122 GNDA_2 0.358056f
C1567 two_stage_opamp_dummy_magic_29_0.cap_res_X.t26 GNDA_2 0.377272f
C1568 two_stage_opamp_dummy_magic_29_0.cap_res_X.t67 GNDA_2 0.192319f
C1569 two_stage_opamp_dummy_magic_29_0.cap_res_X.n32 GNDA_2 0.204169f
C1570 two_stage_opamp_dummy_magic_29_0.cap_res_X.t131 GNDA_2 0.358056f
C1571 two_stage_opamp_dummy_magic_29_0.cap_res_X.t25 GNDA_2 0.375611f
C1572 two_stage_opamp_dummy_magic_29_0.cap_res_X.t18 GNDA_2 0.358056f
C1573 two_stage_opamp_dummy_magic_29_0.cap_res_X.t50 GNDA_2 0.192319f
C1574 two_stage_opamp_dummy_magic_29_0.cap_res_X.n33 GNDA_2 0.205829f
C1575 two_stage_opamp_dummy_magic_29_0.cap_res_X.t137 GNDA_2 0.358056f
C1576 two_stage_opamp_dummy_magic_29_0.cap_res_X.t31 GNDA_2 0.192319f
C1577 two_stage_opamp_dummy_magic_29_0.cap_res_X.n34 GNDA_2 0.204169f
C1578 two_stage_opamp_dummy_magic_29_0.cap_res_X.t99 GNDA_2 0.358056f
C1579 two_stage_opamp_dummy_magic_29_0.cap_res_X.t132 GNDA_2 0.192319f
C1580 two_stage_opamp_dummy_magic_29_0.cap_res_X.n35 GNDA_2 0.204169f
C1581 two_stage_opamp_dummy_magic_29_0.cap_res_X.t123 GNDA_2 0.358056f
C1582 two_stage_opamp_dummy_magic_29_0.cap_res_X.t19 GNDA_2 0.192319f
C1583 two_stage_opamp_dummy_magic_29_0.cap_res_X.n36 GNDA_2 0.204169f
C1584 two_stage_opamp_dummy_magic_29_0.cap_res_X.t82 GNDA_2 0.358056f
C1585 two_stage_opamp_dummy_magic_29_0.cap_res_X.t119 GNDA_2 0.192319f
C1586 two_stage_opamp_dummy_magic_29_0.cap_res_X.n37 GNDA_2 0.204169f
C1587 two_stage_opamp_dummy_magic_29_0.cap_res_X.t44 GNDA_2 0.358056f
C1588 two_stage_opamp_dummy_magic_29_0.cap_res_X.t80 GNDA_2 0.192319f
C1589 two_stage_opamp_dummy_magic_29_0.cap_res_X.n38 GNDA_2 0.204169f
C1590 two_stage_opamp_dummy_magic_29_0.cap_res_X.n39 GNDA_2 0.204169f
C1591 two_stage_opamp_dummy_magic_29_0.cap_res_X.t41 GNDA_2 0.192319f
C1592 two_stage_opamp_dummy_magic_29_0.cap_res_X.t5 GNDA_2 0.377272f
C1593 two_stage_opamp_dummy_magic_29_0.cap_res_X.t30 GNDA_2 0.453363f
C1594 two_stage_opamp_dummy_magic_29_0.cap_res_X.t143 GNDA_2 0.317057f
C1595 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref.t4 GNDA_2 0.322909f
C1596 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref.t9 GNDA_2 0.102139f
C1597 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref.n0 GNDA_2 3.32123f
C1598 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref.t5 GNDA_2 0.061102f
C1599 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref.t1 GNDA_2 0.061102f
C1600 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref.n1 GNDA_2 0.170444f
C1601 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref.t3 GNDA_2 0.061102f
C1602 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref.t0 GNDA_2 0.061102f
C1603 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref.n2 GNDA_2 0.153411f
C1604 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref.n3 GNDA_2 1.88397f
C1605 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref.t2 GNDA_2 0.061102f
C1606 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref.t6 GNDA_2 0.061102f
C1607 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref.n4 GNDA_2 0.153411f
C1608 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref.n5 GNDA_2 1.40074f
C1609 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref.n6 GNDA_2 0.894007f
C1610 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref.t7 GNDA_2 0.070166f
C1611 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref.t8 GNDA_2 0.068986f
C1612 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref.n7 GNDA_2 0.499932f
C1613 bgr_11_0.V_TOP.n0 GNDA_2 0.016831f
C1614 bgr_11_0.V_TOP.t29 GNDA_2 0.128711f
C1615 bgr_11_0.V_TOP.t37 GNDA_2 0.128973f
C1616 bgr_11_0.V_TOP.t38 GNDA_2 0.129529f
C1617 bgr_11_0.V_TOP.n1 GNDA_2 0.162971f
C1618 bgr_11_0.V_TOP.t23 GNDA_2 0.129529f
C1619 bgr_11_0.V_TOP.n2 GNDA_2 0.089272f
C1620 bgr_11_0.V_TOP.t48 GNDA_2 0.129529f
C1621 bgr_11_0.V_TOP.n3 GNDA_2 0.089272f
C1622 bgr_11_0.V_TOP.t39 GNDA_2 0.129529f
C1623 bgr_11_0.V_TOP.n4 GNDA_2 0.089272f
C1624 bgr_11_0.V_TOP.t27 GNDA_2 0.129529f
C1625 bgr_11_0.V_TOP.n5 GNDA_2 0.089272f
C1626 bgr_11_0.V_TOP.n6 GNDA_2 0.025246f
C1627 bgr_11_0.V_TOP.n7 GNDA_2 0.057364f
C1628 bgr_11_0.V_TOP.t8 GNDA_2 0.129887f
C1629 bgr_11_0.V_TOP.t20 GNDA_2 0.374019f
C1630 bgr_11_0.V_TOP.t24 GNDA_2 0.38039f
C1631 bgr_11_0.V_TOP.t32 GNDA_2 0.374019f
C1632 bgr_11_0.V_TOP.n8 GNDA_2 0.250768f
C1633 bgr_11_0.V_TOP.t19 GNDA_2 0.374019f
C1634 bgr_11_0.V_TOP.t46 GNDA_2 0.38039f
C1635 bgr_11_0.V_TOP.n9 GNDA_2 0.320897f
C1636 bgr_11_0.V_TOP.t34 GNDA_2 0.38039f
C1637 bgr_11_0.V_TOP.t40 GNDA_2 0.374019f
C1638 bgr_11_0.V_TOP.n10 GNDA_2 0.250768f
C1639 bgr_11_0.V_TOP.t31 GNDA_2 0.374019f
C1640 bgr_11_0.V_TOP.t18 GNDA_2 0.38039f
C1641 bgr_11_0.V_TOP.n11 GNDA_2 0.391025f
C1642 bgr_11_0.V_TOP.t22 GNDA_2 0.38039f
C1643 bgr_11_0.V_TOP.t30 GNDA_2 0.374019f
C1644 bgr_11_0.V_TOP.n12 GNDA_2 0.250768f
C1645 bgr_11_0.V_TOP.t17 GNDA_2 0.374019f
C1646 bgr_11_0.V_TOP.t44 GNDA_2 0.38039f
C1647 bgr_11_0.V_TOP.n13 GNDA_2 0.391025f
C1648 bgr_11_0.V_TOP.t47 GNDA_2 0.38039f
C1649 bgr_11_0.V_TOP.t16 GNDA_2 0.374019f
C1650 bgr_11_0.V_TOP.n14 GNDA_2 0.250768f
C1651 bgr_11_0.V_TOP.t43 GNDA_2 0.374019f
C1652 bgr_11_0.V_TOP.t35 GNDA_2 0.38039f
C1653 bgr_11_0.V_TOP.n15 GNDA_2 0.391025f
C1654 bgr_11_0.V_TOP.t41 GNDA_2 0.38039f
C1655 bgr_11_0.V_TOP.t15 GNDA_2 0.374019f
C1656 bgr_11_0.V_TOP.n16 GNDA_2 0.320897f
C1657 bgr_11_0.V_TOP.t28 GNDA_2 0.374019f
C1658 bgr_11_0.V_TOP.n17 GNDA_2 0.163634f
C1659 bgr_11_0.V_TOP.n18 GNDA_2 0.875119f
C1660 bgr_11_0.V_TOP.t13 GNDA_2 0.105245f
C1661 bgr_11_0.V_TOP.n19 GNDA_2 1.42428f
C1662 bgr_11_0.V_TOP.n20 GNDA_2 0.019145f
C1663 bgr_11_0.V_TOP.n21 GNDA_2 0.024925f
C1664 bgr_11_0.V_TOP.n22 GNDA_2 0.022551f
C1665 bgr_11_0.V_TOP.n23 GNDA_2 0.25922f
C1666 bgr_11_0.V_TOP.n24 GNDA_2 0.158514f
C1667 bgr_11_0.V_TOP.n25 GNDA_2 0.655866f
C1668 bgr_11_0.V_TOP.n26 GNDA_2 0.020198f
C1669 bgr_11_0.V_TOP.n27 GNDA_2 0.198604f
C1670 bgr_11_0.V_TOP.n28 GNDA_2 0.020198f
C1671 bgr_11_0.V_TOP.n29 GNDA_2 0.204214f
C1672 bgr_11_0.V_TOP.n30 GNDA_2 0.020198f
C1673 bgr_11_0.V_TOP.n31 GNDA_2 0.190361f
C1674 bgr_11_0.V_TOP.n32 GNDA_2 0.391697f
C1675 bgr_11_0.V_TOP.n33 GNDA_2 0.089765f
C1676 bgr_11_0.V_TOP.t14 GNDA_2 0.127788f
C1677 bgr_11_0.V_TOP.n34 GNDA_2 0.052677f
C1678 bgr_11_0.V_TOP.n35 GNDA_2 0.025246f
C1679 bgr_11_0.V_TOP.t45 GNDA_2 0.128533f
C1680 bgr_11_0.V_TOP.n36 GNDA_2 0.084658f
C1681 bgr_11_0.V_TOP.t36 GNDA_2 0.129529f
C1682 bgr_11_0.V_TOP.n37 GNDA_2 0.089272f
C1683 bgr_11_0.V_TOP.t25 GNDA_2 0.129529f
C1684 bgr_11_0.V_TOP.n38 GNDA_2 0.089272f
C1685 bgr_11_0.V_TOP.t26 GNDA_2 0.129529f
C1686 bgr_11_0.V_TOP.n39 GNDA_2 0.089272f
C1687 bgr_11_0.V_TOP.t49 GNDA_2 0.129529f
C1688 bgr_11_0.V_TOP.n40 GNDA_2 0.089272f
C1689 bgr_11_0.V_TOP.t42 GNDA_2 0.129529f
C1690 bgr_11_0.V_TOP.n41 GNDA_2 0.089272f
C1691 bgr_11_0.V_TOP.t33 GNDA_2 0.129529f
C1692 bgr_11_0.V_TOP.n42 GNDA_2 0.080857f
C1693 bgr_11_0.V_TOP.t21 GNDA_2 0.128562f
C1694 VOUT-.n1 GNDA_2 0.074623f
C1695 VOUT-.n4 GNDA_2 0.055967f
C1696 VOUT-.n5 GNDA_2 0.093278f
C1697 VOUT-.n6 GNDA_2 0.055967f
C1698 VOUT-.n7 GNDA_2 0.055967f
C1699 VOUT-.n9 GNDA_2 0.038057f
C1700 VOUT-.n11 GNDA_2 0.038057f
C1701 VOUT-.n13 GNDA_2 0.074623f
C1702 VOUT-.n14 GNDA_2 0.038057f
C1703 VOUT-.n16 GNDA_2 0.038057f
C1704 VOUT-.n18 GNDA_2 0.049251f
C1705 VOUT-.n19 GNDA_2 0.071057f
C1706 VOUT-.n20 GNDA_2 0.06915f
C1707 VOUT-.n21 GNDA_2 0.049251f
C1708 VOUT-.n22 GNDA_2 0.049251f
C1709 VOUT-.n23 GNDA_2 0.06915f
C1710 VOUT-.n24 GNDA_2 0.06915f
C1711 VOUT-.n25 GNDA_2 0.049251f
C1712 VOUT-.n26 GNDA_2 0.078847f
C1713 VOUT-.t17 GNDA_2 0.044774f
C1714 VOUT-.t14 GNDA_2 0.044774f
C1715 VOUT-.n27 GNDA_2 0.091741f
C1716 VOUT-.n28 GNDA_2 0.236811f
C1717 VOUT-.t0 GNDA_2 0.044774f
C1718 VOUT-.t3 GNDA_2 0.044774f
C1719 VOUT-.n29 GNDA_2 0.091741f
C1720 VOUT-.n30 GNDA_2 0.234424f
C1721 VOUT-.n31 GNDA_2 0.056934f
C1722 VOUT-.t12 GNDA_2 0.044774f
C1723 VOUT-.t15 GNDA_2 0.044774f
C1724 VOUT-.n32 GNDA_2 0.091741f
C1725 VOUT-.n33 GNDA_2 0.234424f
C1726 VOUT-.n34 GNDA_2 0.032272f
C1727 VOUT-.t1 GNDA_2 0.044774f
C1728 VOUT-.t13 GNDA_2 0.044774f
C1729 VOUT-.n35 GNDA_2 0.091741f
C1730 VOUT-.n36 GNDA_2 0.234424f
C1731 VOUT-.n37 GNDA_2 0.032272f
C1732 VOUT-.t11 GNDA_2 0.044774f
C1733 VOUT-.t18 GNDA_2 0.044774f
C1734 VOUT-.n38 GNDA_2 0.091741f
C1735 VOUT-.n39 GNDA_2 0.236811f
C1736 VOUT-.n40 GNDA_2 0.056934f
C1737 VOUT-.t2 GNDA_2 0.044774f
C1738 VOUT-.t16 GNDA_2 0.044774f
C1739 VOUT-.n41 GNDA_2 0.091741f
C1740 VOUT-.n42 GNDA_2 0.234424f
C1741 VOUT-.n43 GNDA_2 0.037643f
C1742 VOUT-.n44 GNDA_2 0.022387f
C1743 VOUT-.n45 GNDA_2 0.022387f
C1744 VOUT-.n46 GNDA_2 0.037643f
C1745 VOUT-.n47 GNDA_2 0.06915f
C1746 VOUT-.n48 GNDA_2 0.096796f
C1747 VOUT-.n49 GNDA_2 0.120613f
C1748 VOUT-.n50 GNDA_2 0.168809f
C1749 VOUT-.n51 GNDA_2 0.049251f
C1750 VOUT-.n52 GNDA_2 0.080592f
C1751 VOUT-.n53 GNDA_2 0.049251f
C1752 VOUT-.n54 GNDA_2 0.080592f
C1753 VOUT-.n55 GNDA_2 0.049251f
C1754 VOUT-.n56 GNDA_2 0.049251f
C1755 VOUT-.n57 GNDA_2 0.049251f
C1756 VOUT-.n58 GNDA_2 0.080592f
C1757 VOUT-.n59 GNDA_2 0.049251f
C1758 VOUT-.n60 GNDA_2 0.073876f
C1759 VOUT-.n61 GNDA_2 0.394007f
C1760 VOUT-.n62 GNDA_2 0.387291f
C1761 VOUT-.n64 GNDA_2 0.074623f
C1762 VOUT-.n65 GNDA_2 0.035819f
C1763 VOUT-.n66 GNDA_2 0.494375f
C1764 VOUT-.n69 GNDA_2 0.055967f
C1765 VOUT-.n70 GNDA_2 0.055967f
C1766 VOUT-.t83 GNDA_2 0.303574f
C1767 VOUT-.t105 GNDA_2 0.29849f
C1768 VOUT-.n71 GNDA_2 0.200128f
C1769 VOUT-.t70 GNDA_2 0.29849f
C1770 VOUT-.n72 GNDA_2 0.13059f
C1771 VOUT-.t43 GNDA_2 0.303574f
C1772 VOUT-.t66 GNDA_2 0.29849f
C1773 VOUT-.n73 GNDA_2 0.200128f
C1774 VOUT-.t31 GNDA_2 0.29849f
C1775 VOUT-.t33 GNDA_2 0.302938f
C1776 VOUT-.t52 GNDA_2 0.302938f
C1777 VOUT-.t157 GNDA_2 0.302938f
C1778 VOUT-.t119 GNDA_2 0.302938f
C1779 VOUT-.t139 GNDA_2 0.302938f
C1780 VOUT-.t99 GNDA_2 0.302938f
C1781 VOUT-.t63 GNDA_2 0.302938f
C1782 VOUT-.t25 GNDA_2 0.302938f
C1783 VOUT-.t47 GNDA_2 0.302938f
C1784 VOUT-.t150 GNDA_2 0.302938f
C1785 VOUT-.t133 GNDA_2 0.302938f
C1786 VOUT-.t155 GNDA_2 0.302938f
C1787 VOUT-.t114 GNDA_2 0.29849f
C1788 VOUT-.n74 GNDA_2 0.200765f
C1789 VOUT-.t88 GNDA_2 0.29849f
C1790 VOUT-.n75 GNDA_2 0.256732f
C1791 VOUT-.t108 GNDA_2 0.29849f
C1792 VOUT-.n76 GNDA_2 0.256732f
C1793 VOUT-.t146 GNDA_2 0.29849f
C1794 VOUT-.n77 GNDA_2 0.256732f
C1795 VOUT-.t126 GNDA_2 0.29849f
C1796 VOUT-.n78 GNDA_2 0.256732f
C1797 VOUT-.t22 GNDA_2 0.29849f
C1798 VOUT-.n79 GNDA_2 0.256732f
C1799 VOUT-.t59 GNDA_2 0.29849f
C1800 VOUT-.n80 GNDA_2 0.256732f
C1801 VOUT-.t97 GNDA_2 0.29849f
C1802 VOUT-.n81 GNDA_2 0.256732f
C1803 VOUT-.t78 GNDA_2 0.29849f
C1804 VOUT-.n82 GNDA_2 0.256732f
C1805 VOUT-.t115 GNDA_2 0.29849f
C1806 VOUT-.n83 GNDA_2 0.256732f
C1807 VOUT-.t153 GNDA_2 0.29849f
C1808 VOUT-.n84 GNDA_2 0.256732f
C1809 VOUT-.t132 GNDA_2 0.29849f
C1810 VOUT-.n85 GNDA_2 0.256732f
C1811 VOUT-.n86 GNDA_2 0.242523f
C1812 VOUT-.t37 GNDA_2 0.303574f
C1813 VOUT-.t129 GNDA_2 0.29849f
C1814 VOUT-.n87 GNDA_2 0.200128f
C1815 VOUT-.t92 GNDA_2 0.29849f
C1816 VOUT-.t147 GNDA_2 0.303574f
C1817 VOUT-.t57 GNDA_2 0.29849f
C1818 VOUT-.n88 GNDA_2 0.200128f
C1819 VOUT-.n89 GNDA_2 0.242523f
C1820 VOUT-.t74 GNDA_2 0.303574f
C1821 VOUT-.t23 GNDA_2 0.29849f
C1822 VOUT-.n90 GNDA_2 0.200128f
C1823 VOUT-.t128 GNDA_2 0.29849f
C1824 VOUT-.t41 GNDA_2 0.303574f
C1825 VOUT-.t91 GNDA_2 0.29849f
C1826 VOUT-.n91 GNDA_2 0.200128f
C1827 VOUT-.n92 GNDA_2 0.242523f
C1828 VOUT-.t87 GNDA_2 0.303574f
C1829 VOUT-.t46 GNDA_2 0.29849f
C1830 VOUT-.n93 GNDA_2 0.200128f
C1831 VOUT-.t95 GNDA_2 0.29849f
C1832 VOUT-.t104 GNDA_2 0.303574f
C1833 VOUT-.t149 GNDA_2 0.29849f
C1834 VOUT-.n94 GNDA_2 0.200128f
C1835 VOUT-.n95 GNDA_2 0.242523f
C1836 VOUT-.t102 GNDA_2 0.303574f
C1837 VOUT-.t50 GNDA_2 0.29849f
C1838 VOUT-.n96 GNDA_2 0.200128f
C1839 VOUT-.t158 GNDA_2 0.29849f
C1840 VOUT-.t71 GNDA_2 0.303574f
C1841 VOUT-.t122 GNDA_2 0.29849f
C1842 VOUT-.n97 GNDA_2 0.200128f
C1843 VOUT-.n98 GNDA_2 0.242523f
C1844 VOUT-.t68 GNDA_2 0.303574f
C1845 VOUT-.t161 GNDA_2 0.29849f
C1846 VOUT-.n99 GNDA_2 0.200128f
C1847 VOUT-.t125 GNDA_2 0.29849f
C1848 VOUT-.t36 GNDA_2 0.303574f
C1849 VOUT-.t85 GNDA_2 0.29849f
C1850 VOUT-.n100 GNDA_2 0.200128f
C1851 VOUT-.n101 GNDA_2 0.242523f
C1852 VOUT-.t107 GNDA_2 0.303574f
C1853 VOUT-.t55 GNDA_2 0.29849f
C1854 VOUT-.n102 GNDA_2 0.200128f
C1855 VOUT-.t21 GNDA_2 0.29849f
C1856 VOUT-.t76 GNDA_2 0.303574f
C1857 VOUT-.t127 GNDA_2 0.29849f
C1858 VOUT-.n103 GNDA_2 0.200128f
C1859 VOUT-.n104 GNDA_2 0.242523f
C1860 VOUT-.t148 GNDA_2 0.303574f
C1861 VOUT-.t93 GNDA_2 0.29849f
C1862 VOUT-.n105 GNDA_2 0.200128f
C1863 VOUT-.t60 GNDA_2 0.29849f
C1864 VOUT-.t116 GNDA_2 0.303574f
C1865 VOUT-.t27 GNDA_2 0.29849f
C1866 VOUT-.n106 GNDA_2 0.200128f
C1867 VOUT-.n107 GNDA_2 0.242523f
C1868 VOUT-.t64 GNDA_2 0.303574f
C1869 VOUT-.t86 GNDA_2 0.29849f
C1870 VOUT-.n108 GNDA_2 0.200128f
C1871 VOUT-.t48 GNDA_2 0.29849f
C1872 VOUT-.t75 GNDA_2 0.303574f
C1873 VOUT-.t32 GNDA_2 0.29849f
C1874 VOUT-.n109 GNDA_2 0.195464f
C1875 VOUT-.t39 GNDA_2 0.303574f
C1876 VOUT-.t135 GNDA_2 0.29849f
C1877 VOUT-.n110 GNDA_2 0.195464f
C1878 VOUT-.t131 GNDA_2 0.303574f
C1879 VOUT-.t156 GNDA_2 0.29849f
C1880 VOUT-.n111 GNDA_2 0.195464f
C1881 VOUT-.t117 GNDA_2 0.302938f
C1882 VOUT-.t79 GNDA_2 0.302938f
C1883 VOUT-.t38 GNDA_2 0.302943f
C1884 VOUT-.t62 GNDA_2 0.303188f
C1885 VOUT-.t24 GNDA_2 0.302938f
C1886 VOUT-.t143 GNDA_2 0.302943f
C1887 VOUT-.t30 GNDA_2 0.303188f
C1888 VOUT-.t136 GNDA_2 0.29849f
C1889 VOUT-.n112 GNDA_2 0.204246f
C1890 VOUT-.t111 GNDA_2 0.29849f
C1891 VOUT-.n113 GNDA_2 0.256727f
C1892 VOUT-.t130 GNDA_2 0.29849f
C1893 VOUT-.n114 GNDA_2 0.256732f
C1894 VOUT-.t29 GNDA_2 0.29849f
C1895 VOUT-.n115 GNDA_2 0.260213f
C1896 VOUT-.t142 GNDA_2 0.29849f
C1897 VOUT-.n116 GNDA_2 0.256727f
C1898 VOUT-.t42 GNDA_2 0.29849f
C1899 VOUT-.n117 GNDA_2 0.256732f
C1900 VOUT-.t81 GNDA_2 0.29849f
C1901 VOUT-.n118 GNDA_2 0.256732f
C1902 VOUT-.t120 GNDA_2 0.29849f
C1903 VOUT-.n119 GNDA_2 0.19122f
C1904 VOUT-.t94 GNDA_2 0.29849f
C1905 VOUT-.n120 GNDA_2 0.19122f
C1906 VOUT-.t137 GNDA_2 0.29849f
C1907 VOUT-.n121 GNDA_2 0.19122f
C1908 VOUT-.t35 GNDA_2 0.29849f
C1909 VOUT-.n122 GNDA_2 0.13059f
C1910 VOUT-.t151 GNDA_2 0.29849f
C1911 VOUT-.n123 GNDA_2 0.13059f
C1912 VOUT-.n124 GNDA_2 0.186556f
C1913 VOUT-.t98 GNDA_2 0.303574f
C1914 VOUT-.t124 GNDA_2 0.29849f
C1915 VOUT-.n125 GNDA_2 0.200128f
C1916 VOUT-.t82 GNDA_2 0.29849f
C1917 VOUT-.t69 GNDA_2 0.303574f
C1918 VOUT-.t44 GNDA_2 0.29849f
C1919 VOUT-.n126 GNDA_2 0.200128f
C1920 VOUT-.n127 GNDA_2 0.242523f
C1921 VOUT-.t141 GNDA_2 0.303574f
C1922 VOUT-.t89 GNDA_2 0.29849f
C1923 VOUT-.n128 GNDA_2 0.200128f
C1924 VOUT-.t54 GNDA_2 0.29849f
C1925 VOUT-.t109 GNDA_2 0.303574f
C1926 VOUT-.t20 GNDA_2 0.29849f
C1927 VOUT-.n129 GNDA_2 0.200128f
C1928 VOUT-.n130 GNDA_2 0.242523f
C1929 VOUT-.t101 GNDA_2 0.303574f
C1930 VOUT-.t51 GNDA_2 0.29849f
C1931 VOUT-.n131 GNDA_2 0.200128f
C1932 VOUT-.t160 GNDA_2 0.29849f
C1933 VOUT-.t72 GNDA_2 0.303574f
C1934 VOUT-.t123 GNDA_2 0.29849f
C1935 VOUT-.n132 GNDA_2 0.200128f
C1936 VOUT-.n133 GNDA_2 0.242523f
C1937 VOUT-.t138 GNDA_2 0.303574f
C1938 VOUT-.t84 GNDA_2 0.29849f
C1939 VOUT-.n134 GNDA_2 0.200128f
C1940 VOUT-.t49 GNDA_2 0.29849f
C1941 VOUT-.t103 GNDA_2 0.303574f
C1942 VOUT-.t159 GNDA_2 0.29849f
C1943 VOUT-.n135 GNDA_2 0.200128f
C1944 VOUT-.n136 GNDA_2 0.242523f
C1945 VOUT-.t96 GNDA_2 0.303574f
C1946 VOUT-.t45 GNDA_2 0.29849f
C1947 VOUT-.n137 GNDA_2 0.200128f
C1948 VOUT-.t152 GNDA_2 0.29849f
C1949 VOUT-.t65 GNDA_2 0.303574f
C1950 VOUT-.t118 GNDA_2 0.29849f
C1951 VOUT-.n138 GNDA_2 0.200128f
C1952 VOUT-.n139 GNDA_2 0.242523f
C1953 VOUT-.t56 GNDA_2 0.303574f
C1954 VOUT-.t145 GNDA_2 0.29849f
C1955 VOUT-.n140 GNDA_2 0.200128f
C1956 VOUT-.t112 GNDA_2 0.29849f
C1957 VOUT-.t26 GNDA_2 0.303574f
C1958 VOUT-.t77 GNDA_2 0.29849f
C1959 VOUT-.n141 GNDA_2 0.200128f
C1960 VOUT-.n142 GNDA_2 0.242523f
C1961 VOUT-.t90 GNDA_2 0.303574f
C1962 VOUT-.t40 GNDA_2 0.29849f
C1963 VOUT-.n143 GNDA_2 0.200128f
C1964 VOUT-.t144 GNDA_2 0.29849f
C1965 VOUT-.t58 GNDA_2 0.303574f
C1966 VOUT-.t110 GNDA_2 0.29849f
C1967 VOUT-.n144 GNDA_2 0.200128f
C1968 VOUT-.n145 GNDA_2 0.242523f
C1969 VOUT-.t53 GNDA_2 0.303574f
C1970 VOUT-.t140 GNDA_2 0.29849f
C1971 VOUT-.n146 GNDA_2 0.200128f
C1972 VOUT-.t106 GNDA_2 0.29849f
C1973 VOUT-.t19 GNDA_2 0.303574f
C1974 VOUT-.t73 GNDA_2 0.29849f
C1975 VOUT-.n147 GNDA_2 0.200128f
C1976 VOUT-.n148 GNDA_2 0.242523f
C1977 VOUT-.t154 GNDA_2 0.303574f
C1978 VOUT-.t100 GNDA_2 0.29849f
C1979 VOUT-.n149 GNDA_2 0.200128f
C1980 VOUT-.t67 GNDA_2 0.29849f
C1981 VOUT-.t121 GNDA_2 0.303574f
C1982 VOUT-.t34 GNDA_2 0.29849f
C1983 VOUT-.n150 GNDA_2 0.200128f
C1984 VOUT-.n151 GNDA_2 0.242523f
C1985 VOUT-.t113 GNDA_2 0.303574f
C1986 VOUT-.t61 GNDA_2 0.29849f
C1987 VOUT-.n152 GNDA_2 0.200128f
C1988 VOUT-.t28 GNDA_2 0.29849f
C1989 VOUT-.n153 GNDA_2 0.242523f
C1990 VOUT-.t134 GNDA_2 0.29849f
C1991 VOUT-.n154 GNDA_2 0.127311f
C1992 VOUT-.t80 GNDA_2 0.29849f
C1993 VOUT-.n155 GNDA_2 0.337215f
C1994 VOUT-.n156 GNDA_2 0.274238f
C1995 VOUT-.n157 GNDA_2 0.055967f
C1996 VOUT-.n158 GNDA_2 0.055967f
C1997 VOUT-.n159 GNDA_2 0.055967f
C1998 VOUT-.n160 GNDA_2 0.16416f
C1999 VOUT-.n161 GNDA_2 0.059295f
C2000 VOUT-.n162 GNDA_2 0.05638f
C2001 VOUT-.n164 GNDA_2 0.503703f
C2002 VOUT-.n165 GNDA_2 0.055967f
C2003 VOUT-.n166 GNDA_2 1.06337f
C2004 VOUT-.n170 GNDA_2 0.038057f
C2005 VOUT-.n171 GNDA_2 0.038057f
C2006 VOUT-.n172 GNDA_2 0.035819f
C2007 VOUT-.n173 GNDA_2 0.074623f
C2008 VOUT-.n174 GNDA_2 0.038057f
C2009 VOUT-.n175 GNDA_2 0.038057f
C2010 VOUT-.n177 GNDA_2 1.05404f
C2011 VOUT-.n178 GNDA_2 0.257448f
C2012 VOUT-.t10 GNDA_2 0.085506f
C2013 VOUT-.n179 GNDA_2 0.419876f
C2014 VOUT-.n180 GNDA_2 0.035819f
C2015 VOUT-.t5 GNDA_2 0.052236f
C2016 VOUT-.t8 GNDA_2 0.052236f
C2017 VOUT-.n181 GNDA_2 0.112235f
C2018 VOUT-.n182 GNDA_2 0.275519f
C2019 VOUT-.n183 GNDA_2 0.035819f
C2020 VOUT-.n184 GNDA_2 0.237647f
C2021 VOUT-.t7 GNDA_2 0.052236f
C2022 VOUT-.t4 GNDA_2 0.052236f
C2023 VOUT-.n185 GNDA_2 0.112235f
C2024 VOUT-.n186 GNDA_2 0.284206f
C2025 VOUT-.n187 GNDA_2 0.159675f
C2026 VOUT-.t9 GNDA_2 0.052236f
C2027 VOUT-.t6 GNDA_2 0.052236f
C2028 VOUT-.n188 GNDA_2 0.112235f
C2029 VOUT-.n189 GNDA_2 0.270977f
C2030 VOUT-.n190 GNDA_2 0.127387f
C2031 VOUT-.n191 GNDA_2 0.035819f
C2032 VOUT-.n192 GNDA_2 0.184829f
C2033 VOUT-.n193 GNDA_2 0.035819f
C2034 VOUT-.n194 GNDA_2 0.035819f
C2035 VOUT-.n195 GNDA_2 0.035819f
C2036 VOUT-.n196 GNDA_2 0.035819f
C2037 VOUT-.n197 GNDA_2 0.082271f
C2038 VOUT-.n198 GNDA_2 0.096263f
C2039 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.t1 GNDA_2 0.245842f
C2040 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.t5 GNDA_2 0.773204f
C2041 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.t7 GNDA_2 0.772991f
C2042 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.n0 GNDA_2 0.636556f
C2043 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.t2 GNDA_2 0.772991f
C2044 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.n1 GNDA_2 0.331481f
C2045 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.t3 GNDA_2 0.772991f
C2046 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.n2 GNDA_2 0.667625f
C2047 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.n3 GNDA_2 0.790892f
C2048 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.t0 GNDA_2 0.245842f
C2049 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.n4 GNDA_2 0.431779f
C2050 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.t9 GNDA_2 0.667922f
C2051 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.t4 GNDA_2 0.667922f
C2052 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.t6 GNDA_2 0.667922f
C2053 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.t8 GNDA_2 0.722234f
C2054 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.n5 GNDA_2 0.241787f
C2055 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.n6 GNDA_2 0.300709f
C2056 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.n7 GNDA_2 0.300709f
C2057 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.n8 GNDA_2 0.294161f
C2058 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.n9 GNDA_2 0.489447f
C2059 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.n10 GNDA_2 1.39879f
C2060 two_stage_opamp_dummy_magic_29_0.Y.n0 GNDA_2 0.194525f
C2061 two_stage_opamp_dummy_magic_29_0.Y.n1 GNDA_2 0.08603f
C2062 two_stage_opamp_dummy_magic_29_0.Y.n2 GNDA_2 0.237753f
C2063 two_stage_opamp_dummy_magic_29_0.Y.n3 GNDA_2 0.815021f
C2064 two_stage_opamp_dummy_magic_29_0.Y.n4 GNDA_2 0.08603f
C2065 two_stage_opamp_dummy_magic_29_0.Y.n5 GNDA_2 0.08603f
C2066 two_stage_opamp_dummy_magic_29_0.Y.t5 GNDA_2 0.023158f
C2067 two_stage_opamp_dummy_magic_29_0.Y.t4 GNDA_2 0.023158f
C2068 two_stage_opamp_dummy_magic_29_0.Y.n6 GNDA_2 0.068053f
C2069 two_stage_opamp_dummy_magic_29_0.Y.t1 GNDA_2 0.023158f
C2070 two_stage_opamp_dummy_magic_29_0.Y.t6 GNDA_2 0.023158f
C2071 two_stage_opamp_dummy_magic_29_0.Y.n7 GNDA_2 0.066733f
C2072 two_stage_opamp_dummy_magic_29_0.Y.n8 GNDA_2 0.441071f
C2073 two_stage_opamp_dummy_magic_29_0.Y.t7 GNDA_2 0.023158f
C2074 two_stage_opamp_dummy_magic_29_0.Y.t12 GNDA_2 0.023158f
C2075 two_stage_opamp_dummy_magic_29_0.Y.n9 GNDA_2 0.066733f
C2076 two_stage_opamp_dummy_magic_29_0.Y.n10 GNDA_2 0.232002f
C2077 two_stage_opamp_dummy_magic_29_0.Y.t10 GNDA_2 0.023158f
C2078 two_stage_opamp_dummy_magic_29_0.Y.t8 GNDA_2 0.023158f
C2079 two_stage_opamp_dummy_magic_29_0.Y.n11 GNDA_2 0.066733f
C2080 two_stage_opamp_dummy_magic_29_0.Y.n12 GNDA_2 0.232002f
C2081 two_stage_opamp_dummy_magic_29_0.Y.t23 GNDA_2 0.023158f
C2082 two_stage_opamp_dummy_magic_29_0.Y.t11 GNDA_2 0.023158f
C2083 two_stage_opamp_dummy_magic_29_0.Y.n13 GNDA_2 0.066733f
C2084 two_stage_opamp_dummy_magic_29_0.Y.n14 GNDA_2 0.232002f
C2085 two_stage_opamp_dummy_magic_29_0.Y.t3 GNDA_2 0.023158f
C2086 two_stage_opamp_dummy_magic_29_0.Y.t9 GNDA_2 0.023158f
C2087 two_stage_opamp_dummy_magic_29_0.Y.n15 GNDA_2 0.066733f
C2088 two_stage_opamp_dummy_magic_29_0.Y.n16 GNDA_2 0.431159f
C2089 two_stage_opamp_dummy_magic_29_0.Y.n17 GNDA_2 0.287483f
C2090 two_stage_opamp_dummy_magic_29_0.Y.n18 GNDA_2 0.644415f
C2091 two_stage_opamp_dummy_magic_29_0.Y.n19 GNDA_2 0.496725f
C2092 two_stage_opamp_dummy_magic_29_0.Y.n20 GNDA_2 0.237753f
C2093 two_stage_opamp_dummy_magic_29_0.Y.n21 GNDA_2 0.417266f
C2094 two_stage_opamp_dummy_magic_29_0.Y.n22 GNDA_2 0.237753f
C2095 two_stage_opamp_dummy_magic_29_0.Y.n23 GNDA_2 0.237753f
C2096 two_stage_opamp_dummy_magic_29_0.Y.n24 GNDA_2 0.237753f
C2097 two_stage_opamp_dummy_magic_29_0.Y.n25 GNDA_2 0.146616f
C2098 two_stage_opamp_dummy_magic_29_0.Y.n27 GNDA_2 0.074105f
C2099 two_stage_opamp_dummy_magic_29_0.Y.n28 GNDA_2 0.074105f
C2100 two_stage_opamp_dummy_magic_29_0.Y.n30 GNDA_2 0.074105f
C2101 two_stage_opamp_dummy_magic_29_0.Y.n32 GNDA_2 0.074105f
C2102 two_stage_opamp_dummy_magic_29_0.Y.n34 GNDA_2 0.172912f
C2103 two_stage_opamp_dummy_magic_29_0.Y.n36 GNDA_2 0.074105f
C2104 two_stage_opamp_dummy_magic_29_0.Y.n37 GNDA_2 0.074105f
C2105 two_stage_opamp_dummy_magic_29_0.Y.n38 GNDA_2 0.073409f
C2106 two_stage_opamp_dummy_magic_29_0.Y.n39 GNDA_2 0.074105f
C2107 two_stage_opamp_dummy_magic_29_0.Y.t2 GNDA_2 0.640789f
C2108 two_stage_opamp_dummy_magic_29_0.Y.n40 GNDA_2 0.074105f
C2109 two_stage_opamp_dummy_magic_29_0.Y.n41 GNDA_2 0.074105f
C2110 two_stage_opamp_dummy_magic_29_0.Y.n43 GNDA_2 0.687542f
C2111 two_stage_opamp_dummy_magic_29_0.Y.n45 GNDA_2 0.643787f
C2112 two_stage_opamp_dummy_magic_29_0.Y.n46 GNDA_2 0.024538f
C2113 two_stage_opamp_dummy_magic_29_0.Y.n47 GNDA_2 0.024702f
C2114 two_stage_opamp_dummy_magic_29_0.Y.n48 GNDA_2 0.024702f
C2115 two_stage_opamp_dummy_magic_29_0.Y.t32 GNDA_2 0.101894f
C2116 two_stage_opamp_dummy_magic_29_0.Y.t38 GNDA_2 0.101894f
C2117 two_stage_opamp_dummy_magic_29_0.Y.t51 GNDA_2 0.101894f
C2118 two_stage_opamp_dummy_magic_29_0.Y.t41 GNDA_2 0.101894f
C2119 two_stage_opamp_dummy_magic_29_0.Y.t25 GNDA_2 0.108524f
C2120 two_stage_opamp_dummy_magic_29_0.Y.n49 GNDA_2 0.086001f
C2121 two_stage_opamp_dummy_magic_29_0.Y.n50 GNDA_2 0.048631f
C2122 two_stage_opamp_dummy_magic_29_0.Y.n51 GNDA_2 0.048631f
C2123 two_stage_opamp_dummy_magic_29_0.Y.n52 GNDA_2 0.04371f
C2124 two_stage_opamp_dummy_magic_29_0.Y.t46 GNDA_2 0.101894f
C2125 two_stage_opamp_dummy_magic_29_0.Y.t29 GNDA_2 0.101894f
C2126 two_stage_opamp_dummy_magic_29_0.Y.t44 GNDA_2 0.101894f
C2127 two_stage_opamp_dummy_magic_29_0.Y.t26 GNDA_2 0.101894f
C2128 two_stage_opamp_dummy_magic_29_0.Y.t34 GNDA_2 0.108524f
C2129 two_stage_opamp_dummy_magic_29_0.Y.n53 GNDA_2 0.086001f
C2130 two_stage_opamp_dummy_magic_29_0.Y.n54 GNDA_2 0.048631f
C2131 two_stage_opamp_dummy_magic_29_0.Y.n55 GNDA_2 0.048631f
C2132 two_stage_opamp_dummy_magic_29_0.Y.n56 GNDA_2 0.04371f
C2133 two_stage_opamp_dummy_magic_29_0.Y.n57 GNDA_2 0.010496f
C2134 two_stage_opamp_dummy_magic_29_0.Y.n58 GNDA_2 0.024866f
C2135 two_stage_opamp_dummy_magic_29_0.Y.n59 GNDA_2 0.058532f
C2136 two_stage_opamp_dummy_magic_29_0.Y.n60 GNDA_2 0.033384f
C2137 two_stage_opamp_dummy_magic_29_0.Y.n61 GNDA_2 0.037886f
C2138 two_stage_opamp_dummy_magic_29_0.Y.n62 GNDA_2 1.02357f
C2139 two_stage_opamp_dummy_magic_29_0.Y.t40 GNDA_2 0.049789f
C2140 two_stage_opamp_dummy_magic_29_0.Y.t54 GNDA_2 0.049789f
C2141 two_stage_opamp_dummy_magic_29_0.Y.t43 GNDA_2 0.049789f
C2142 two_stage_opamp_dummy_magic_29_0.Y.t28 GNDA_2 0.049789f
C2143 two_stage_opamp_dummy_magic_29_0.Y.t35 GNDA_2 0.049789f
C2144 two_stage_opamp_dummy_magic_29_0.Y.t47 GNDA_2 0.049789f
C2145 two_stage_opamp_dummy_magic_29_0.Y.t37 GNDA_2 0.049789f
C2146 two_stage_opamp_dummy_magic_29_0.Y.t49 GNDA_2 0.056602f
C2147 two_stage_opamp_dummy_magic_29_0.Y.n64 GNDA_2 0.051082f
C2148 two_stage_opamp_dummy_magic_29_0.Y.n65 GNDA_2 0.031263f
C2149 two_stage_opamp_dummy_magic_29_0.Y.n66 GNDA_2 0.031263f
C2150 two_stage_opamp_dummy_magic_29_0.Y.n67 GNDA_2 0.031263f
C2151 two_stage_opamp_dummy_magic_29_0.Y.n68 GNDA_2 0.031263f
C2152 two_stage_opamp_dummy_magic_29_0.Y.n69 GNDA_2 0.031263f
C2153 two_stage_opamp_dummy_magic_29_0.Y.n70 GNDA_2 0.026342f
C2154 two_stage_opamp_dummy_magic_29_0.Y.t50 GNDA_2 0.049789f
C2155 two_stage_opamp_dummy_magic_29_0.Y.t30 GNDA_2 0.056602f
C2156 two_stage_opamp_dummy_magic_29_0.Y.n71 GNDA_2 0.046161f
C2157 two_stage_opamp_dummy_magic_29_0.Y.n72 GNDA_2 0.012791f
C2158 two_stage_opamp_dummy_magic_29_0.Y.t42 GNDA_2 0.032421f
C2159 two_stage_opamp_dummy_magic_29_0.Y.t27 GNDA_2 0.032421f
C2160 two_stage_opamp_dummy_magic_29_0.Y.t45 GNDA_2 0.032421f
C2161 two_stage_opamp_dummy_magic_29_0.Y.t31 GNDA_2 0.032421f
C2162 two_stage_opamp_dummy_magic_29_0.Y.t36 GNDA_2 0.032421f
C2163 two_stage_opamp_dummy_magic_29_0.Y.t48 GNDA_2 0.032421f
C2164 two_stage_opamp_dummy_magic_29_0.Y.t39 GNDA_2 0.032421f
C2165 two_stage_opamp_dummy_magic_29_0.Y.t52 GNDA_2 0.039368f
C2166 two_stage_opamp_dummy_magic_29_0.Y.n73 GNDA_2 0.039368f
C2167 two_stage_opamp_dummy_magic_29_0.Y.n74 GNDA_2 0.025474f
C2168 two_stage_opamp_dummy_magic_29_0.Y.n75 GNDA_2 0.025474f
C2169 two_stage_opamp_dummy_magic_29_0.Y.n76 GNDA_2 0.025474f
C2170 two_stage_opamp_dummy_magic_29_0.Y.n77 GNDA_2 0.025474f
C2171 two_stage_opamp_dummy_magic_29_0.Y.n78 GNDA_2 0.025474f
C2172 two_stage_opamp_dummy_magic_29_0.Y.n79 GNDA_2 0.020552f
C2173 two_stage_opamp_dummy_magic_29_0.Y.t53 GNDA_2 0.032421f
C2174 two_stage_opamp_dummy_magic_29_0.Y.t33 GNDA_2 0.039368f
C2175 two_stage_opamp_dummy_magic_29_0.Y.n80 GNDA_2 0.034447f
C2176 two_stage_opamp_dummy_magic_29_0.Y.n81 GNDA_2 0.012791f
C2177 two_stage_opamp_dummy_magic_29_0.Y.n82 GNDA_2 0.079795f
C2178 two_stage_opamp_dummy_magic_29_0.Y.n83 GNDA_2 0.074105f
C2179 two_stage_opamp_dummy_magic_29_0.Y.n84 GNDA_2 2.18995f
C2180 two_stage_opamp_dummy_magic_29_0.Y.n85 GNDA_2 0.453893f
C2181 two_stage_opamp_dummy_magic_29_0.Y.n87 GNDA_2 0.463156f
C2182 two_stage_opamp_dummy_magic_29_0.Y.n88 GNDA_2 0.463156f
C2183 two_stage_opamp_dummy_magic_29_0.Y.n91 GNDA_2 0.083312f
C2184 two_stage_opamp_dummy_magic_29_0.Y.n92 GNDA_2 0.083312f
C2185 two_stage_opamp_dummy_magic_29_0.Y.t13 GNDA_2 0.054035f
C2186 two_stage_opamp_dummy_magic_29_0.Y.t0 GNDA_2 0.054035f
C2187 two_stage_opamp_dummy_magic_29_0.Y.n93 GNDA_2 0.110534f
C2188 two_stage_opamp_dummy_magic_29_0.Y.n94 GNDA_2 0.35586f
C2189 two_stage_opamp_dummy_magic_29_0.Y.n95 GNDA_2 0.138043f
C2190 two_stage_opamp_dummy_magic_29_0.Y.t19 GNDA_2 0.054035f
C2191 two_stage_opamp_dummy_magic_29_0.Y.t21 GNDA_2 0.054035f
C2192 two_stage_opamp_dummy_magic_29_0.Y.n96 GNDA_2 0.110534f
C2193 two_stage_opamp_dummy_magic_29_0.Y.n97 GNDA_2 0.348103f
C2194 two_stage_opamp_dummy_magic_29_0.Y.n98 GNDA_2 0.138043f
C2195 two_stage_opamp_dummy_magic_29_0.Y.t16 GNDA_2 0.054035f
C2196 two_stage_opamp_dummy_magic_29_0.Y.t14 GNDA_2 0.054035f
C2197 two_stage_opamp_dummy_magic_29_0.Y.n99 GNDA_2 0.110534f
C2198 two_stage_opamp_dummy_magic_29_0.Y.n100 GNDA_2 0.348103f
C2199 two_stage_opamp_dummy_magic_29_0.Y.n101 GNDA_2 0.083312f
C2200 two_stage_opamp_dummy_magic_29_0.Y.n102 GNDA_2 0.083312f
C2201 two_stage_opamp_dummy_magic_29_0.Y.t20 GNDA_2 0.054035f
C2202 two_stage_opamp_dummy_magic_29_0.Y.t18 GNDA_2 0.054035f
C2203 two_stage_opamp_dummy_magic_29_0.Y.n103 GNDA_2 0.110534f
C2204 two_stage_opamp_dummy_magic_29_0.Y.n104 GNDA_2 0.348103f
C2205 two_stage_opamp_dummy_magic_29_0.Y.n105 GNDA_2 0.083312f
C2206 two_stage_opamp_dummy_magic_29_0.Y.t22 GNDA_2 0.054035f
C2207 two_stage_opamp_dummy_magic_29_0.Y.t15 GNDA_2 0.054035f
C2208 two_stage_opamp_dummy_magic_29_0.Y.n106 GNDA_2 0.110534f
C2209 two_stage_opamp_dummy_magic_29_0.Y.n107 GNDA_2 0.348103f
C2210 two_stage_opamp_dummy_magic_29_0.Y.n108 GNDA_2 0.138043f
C2211 two_stage_opamp_dummy_magic_29_0.Y.t24 GNDA_2 0.054035f
C2212 two_stage_opamp_dummy_magic_29_0.Y.t17 GNDA_2 0.054035f
C2213 two_stage_opamp_dummy_magic_29_0.Y.n109 GNDA_2 0.110534f
C2214 two_stage_opamp_dummy_magic_29_0.Y.n110 GNDA_2 0.351981f
C2215 two_stage_opamp_dummy_magic_29_0.Y.n111 GNDA_2 0.220104f
C2216 two_stage_opamp_dummy_magic_29_0.Y.n112 GNDA_2 0.619696f
C2217 two_stage_opamp_dummy_magic_29_0.Y.n114 GNDA_2 0.172912f
C2218 two_stage_opamp_dummy_magic_29_0.Y.n116 GNDA_2 0.074105f
C2219 two_stage_opamp_dummy_magic_29_0.Y.n117 GNDA_2 1.3941f
C2220 two_stage_opamp_dummy_magic_29_0.Y.n118 GNDA_2 1.42652f
C2221 two_stage_opamp_dummy_magic_29_0.Y.n119 GNDA_2 0.388675f
C2222 two_stage_opamp_dummy_magic_29_0.Y.n120 GNDA_2 0.237753f
C2223 two_stage_opamp_dummy_magic_29_0.Y.n121 GNDA_2 0.417266f
C2224 two_stage_opamp_dummy_magic_29_0.Y.n122 GNDA_2 0.237753f
C2225 two_stage_opamp_dummy_magic_29_0.Y.n123 GNDA_2 0.237753f
C2226 two_stage_opamp_dummy_magic_29_0.Y.n124 GNDA_2 0.237753f
C2227 two_stage_opamp_dummy_magic_29_0.Y.n125 GNDA_2 0.341617f
C2228 two_stage_opamp_dummy_magic_29_0.Vb2.n0 GNDA_2 0.528073f
C2229 two_stage_opamp_dummy_magic_29_0.Vb2.n1 GNDA_2 0.539048f
C2230 two_stage_opamp_dummy_magic_29_0.Vb2.n2 GNDA_2 0.393311f
C2231 two_stage_opamp_dummy_magic_29_0.Vb2.n3 GNDA_2 0.539048f
C2232 two_stage_opamp_dummy_magic_29_0.Vb2.n4 GNDA_2 0.953442f
C2233 two_stage_opamp_dummy_magic_29_0.Vb2.n5 GNDA_2 0.784984f
C2234 two_stage_opamp_dummy_magic_29_0.Vb2.t1 GNDA_2 0.01824f
C2235 two_stage_opamp_dummy_magic_29_0.Vb2.t2 GNDA_2 0.01824f
C2236 two_stage_opamp_dummy_magic_29_0.Vb2.n6 GNDA_2 0.061156f
C2237 two_stage_opamp_dummy_magic_29_0.Vb2.t0 GNDA_2 0.01824f
C2238 two_stage_opamp_dummy_magic_29_0.Vb2.t5 GNDA_2 0.01824f
C2239 two_stage_opamp_dummy_magic_29_0.Vb2.n7 GNDA_2 0.059478f
C2240 two_stage_opamp_dummy_magic_29_0.Vb2.n8 GNDA_2 0.55333f
C2241 two_stage_opamp_dummy_magic_29_0.Vb2.t4 GNDA_2 0.01824f
C2242 two_stage_opamp_dummy_magic_29_0.Vb2.t6 GNDA_2 0.01824f
C2243 two_stage_opamp_dummy_magic_29_0.Vb2.n9 GNDA_2 0.059478f
C2244 two_stage_opamp_dummy_magic_29_0.Vb2.n10 GNDA_2 0.366423f
C2245 two_stage_opamp_dummy_magic_29_0.Vb2.t3 GNDA_2 0.01824f
C2246 two_stage_opamp_dummy_magic_29_0.Vb2.t7 GNDA_2 0.01824f
C2247 two_stage_opamp_dummy_magic_29_0.Vb2.n11 GNDA_2 0.059478f
C2248 two_stage_opamp_dummy_magic_29_0.Vb2.n12 GNDA_2 1.13805f
C2249 two_stage_opamp_dummy_magic_29_0.Vb2.t15 GNDA_2 0.11698f
C2250 two_stage_opamp_dummy_magic_29_0.Vb2.t13 GNDA_2 0.116949f
C2251 two_stage_opamp_dummy_magic_29_0.Vb2.t29 GNDA_2 0.116949f
C2252 two_stage_opamp_dummy_magic_29_0.Vb2.t23 GNDA_2 0.116949f
C2253 two_stage_opamp_dummy_magic_29_0.Vb2.t19 GNDA_2 0.116949f
C2254 two_stage_opamp_dummy_magic_29_0.Vb2.t16 GNDA_2 0.116949f
C2255 two_stage_opamp_dummy_magic_29_0.Vb2.t14 GNDA_2 0.116949f
C2256 two_stage_opamp_dummy_magic_29_0.Vb2.t12 GNDA_2 0.116949f
C2257 two_stage_opamp_dummy_magic_29_0.Vb2.t27 GNDA_2 0.116949f
C2258 two_stage_opamp_dummy_magic_29_0.Vb2.t31 GNDA_2 0.116949f
C2259 two_stage_opamp_dummy_magic_29_0.Vb2.t22 GNDA_2 0.11698f
C2260 two_stage_opamp_dummy_magic_29_0.Vb2.t28 GNDA_2 0.116949f
C2261 two_stage_opamp_dummy_magic_29_0.Vb2.t25 GNDA_2 0.116949f
C2262 two_stage_opamp_dummy_magic_29_0.Vb2.t32 GNDA_2 0.116949f
C2263 two_stage_opamp_dummy_magic_29_0.Vb2.t18 GNDA_2 0.116949f
C2264 two_stage_opamp_dummy_magic_29_0.Vb2.t20 GNDA_2 0.116949f
C2265 two_stage_opamp_dummy_magic_29_0.Vb2.t24 GNDA_2 0.116949f
C2266 two_stage_opamp_dummy_magic_29_0.Vb2.t21 GNDA_2 0.116949f
C2267 two_stage_opamp_dummy_magic_29_0.Vb2.t26 GNDA_2 0.116949f
C2268 two_stage_opamp_dummy_magic_29_0.Vb2.t11 GNDA_2 0.116949f
C2269 two_stage_opamp_dummy_magic_29_0.Vb2.t9 GNDA_2 0.06384f
C2270 two_stage_opamp_dummy_magic_29_0.Vb2.t10 GNDA_2 0.06384f
C2271 two_stage_opamp_dummy_magic_29_0.Vb2.n13 GNDA_2 0.135818f
C2272 two_stage_opamp_dummy_magic_29_0.Vb2.t8 GNDA_2 0.120795f
C2273 two_stage_opamp_dummy_magic_29_0.Vb2.n14 GNDA_2 0.516758f
C2274 two_stage_opamp_dummy_magic_29_0.Vb2.n15 GNDA_2 0.711221f
C2275 two_stage_opamp_dummy_magic_29_0.Vb2.t30 GNDA_2 0.073327f
C2276 two_stage_opamp_dummy_magic_29_0.Vb2.n16 GNDA_2 0.668033f
C2277 two_stage_opamp_dummy_magic_29_0.Vb2.t17 GNDA_2 0.117333f
C2278 two_stage_opamp_dummy_magic_29_0.Vb2.n17 GNDA_2 0.642085f
C2279 two_stage_opamp_dummy_magic_29_0.Vb2.n18 GNDA_2 1.87158f
C2280 bgr_11_0.VB2_CUR_BIAS GNDA_2 4.99512f
C2281 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t18 GNDA_2 0.35871f
C2282 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t51 GNDA_2 0.376298f
C2283 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t54 GNDA_2 0.35871f
C2284 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t94 GNDA_2 0.19267f
C2285 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n0 GNDA_2 0.206205f
C2286 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t37 GNDA_2 0.35871f
C2287 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t65 GNDA_2 0.19267f
C2288 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n1 GNDA_2 0.204542f
C2289 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t70 GNDA_2 0.35871f
C2290 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t108 GNDA_2 0.19267f
C2291 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n2 GNDA_2 0.204542f
C2292 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t109 GNDA_2 0.35871f
C2293 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t8 GNDA_2 0.19267f
C2294 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n3 GNDA_2 0.204542f
C2295 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t10 GNDA_2 0.35871f
C2296 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t43 GNDA_2 0.19267f
C2297 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n4 GNDA_2 0.204542f
C2298 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t137 GNDA_2 0.35871f
C2299 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t21 GNDA_2 0.19267f
C2300 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n5 GNDA_2 0.204542f
C2301 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t129 GNDA_2 0.35871f
C2302 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t17 GNDA_2 0.36001f
C2303 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t79 GNDA_2 0.35871f
C2304 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t85 GNDA_2 0.36001f
C2305 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t91 GNDA_2 0.35871f
C2306 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t130 GNDA_2 0.36001f
C2307 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t55 GNDA_2 0.35871f
C2308 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t84 GNDA_2 0.36001f
C2309 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t83 GNDA_2 0.35871f
C2310 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t139 GNDA_2 0.36001f
C2311 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t99 GNDA_2 0.35871f
C2312 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t127 GNDA_2 0.36001f
C2313 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t124 GNDA_2 0.35871f
C2314 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t30 GNDA_2 0.36001f
C2315 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t58 GNDA_2 0.35871f
C2316 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t89 GNDA_2 0.36001f
C2317 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t88 GNDA_2 0.35871f
C2318 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t2 GNDA_2 0.36001f
C2319 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t103 GNDA_2 0.35871f
C2320 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t136 GNDA_2 0.36001f
C2321 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t135 GNDA_2 0.35871f
C2322 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t35 GNDA_2 0.36001f
C2323 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t6 GNDA_2 0.35871f
C2324 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t29 GNDA_2 0.36001f
C2325 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t28 GNDA_2 0.35871f
C2326 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t71 GNDA_2 0.36001f
C2327 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t107 GNDA_2 0.35871f
C2328 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t142 GNDA_2 0.36001f
C2329 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t141 GNDA_2 0.35871f
C2330 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t39 GNDA_2 0.36001f
C2331 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t9 GNDA_2 0.35871f
C2332 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t34 GNDA_2 0.36001f
C2333 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t33 GNDA_2 0.35871f
C2334 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t80 GNDA_2 0.36001f
C2335 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t47 GNDA_2 0.35871f
C2336 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t68 GNDA_2 0.36001f
C2337 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t67 GNDA_2 0.35871f
C2338 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t122 GNDA_2 0.36001f
C2339 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t90 GNDA_2 0.35871f
C2340 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t113 GNDA_2 0.36001f
C2341 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t111 GNDA_2 0.35871f
C2342 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t19 GNDA_2 0.36001f
C2343 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t50 GNDA_2 0.35871f
C2344 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t77 GNDA_2 0.36001f
C2345 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t76 GNDA_2 0.35871f
C2346 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t131 GNDA_2 0.36001f
C2347 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t95 GNDA_2 0.35871f
C2348 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t119 GNDA_2 0.36001f
C2349 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t118 GNDA_2 0.35871f
C2350 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t23 GNDA_2 0.36001f
C2351 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t143 GNDA_2 0.35871f
C2352 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t16 GNDA_2 0.36001f
C2353 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t15 GNDA_2 0.35871f
C2354 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t61 GNDA_2 0.36001f
C2355 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t100 GNDA_2 0.35871f
C2356 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t128 GNDA_2 0.36001f
C2357 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t126 GNDA_2 0.35871f
C2358 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t31 GNDA_2 0.36001f
C2359 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t64 GNDA_2 0.35871f
C2360 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t105 GNDA_2 0.36001f
C2361 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t60 GNDA_2 0.35871f
C2362 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t115 GNDA_2 0.36001f
C2363 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t132 GNDA_2 0.35871f
C2364 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t12 GNDA_2 0.36001f
C2365 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t13 GNDA_2 0.35871f
C2366 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t56 GNDA_2 0.36001f
C2367 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t20 GNDA_2 0.35871f
C2368 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t46 GNDA_2 0.36001f
C2369 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t45 GNDA_2 0.35871f
C2370 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t96 GNDA_2 0.36001f
C2371 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t36 GNDA_2 0.35871f
C2372 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t72 GNDA_2 0.376298f
C2373 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t69 GNDA_2 0.35871f
C2374 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t114 GNDA_2 0.19267f
C2375 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n6 GNDA_2 0.206205f
C2376 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t48 GNDA_2 0.35871f
C2377 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t93 GNDA_2 0.19267f
C2378 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n7 GNDA_2 0.204542f
C2379 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t92 GNDA_2 0.35871f
C2380 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t138 GNDA_2 0.19267f
C2381 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n8 GNDA_2 0.204542f
C2382 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t133 GNDA_2 0.35871f
C2383 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t26 GNDA_2 0.19267f
C2384 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n9 GNDA_2 0.204542f
C2385 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t24 GNDA_2 0.35871f
C2386 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t62 GNDA_2 0.19267f
C2387 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n10 GNDA_2 0.204542f
C2388 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t5 GNDA_2 0.35871f
C2389 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t42 GNDA_2 0.19267f
C2390 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n11 GNDA_2 0.204542f
C2391 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t40 GNDA_2 0.35871f
C2392 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t81 GNDA_2 0.19267f
C2393 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n12 GNDA_2 0.204542f
C2394 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t78 GNDA_2 0.35871f
C2395 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t120 GNDA_2 0.19267f
C2396 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n13 GNDA_2 0.204542f
C2397 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t53 GNDA_2 0.35871f
C2398 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t98 GNDA_2 0.19267f
C2399 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n14 GNDA_2 0.204542f
C2400 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t97 GNDA_2 0.35871f
C2401 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t1 GNDA_2 0.19267f
C2402 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n15 GNDA_2 0.204542f
C2403 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t102 GNDA_2 0.35871f
C2404 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t4 GNDA_2 0.19267f
C2405 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n16 GNDA_2 0.204542f
C2406 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t7 GNDA_2 0.35871f
C2407 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t38 GNDA_2 0.36001f
C2408 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t104 GNDA_2 0.35871f
C2409 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t3 GNDA_2 0.36001f
C2410 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t63 GNDA_2 0.173419f
C2411 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n17 GNDA_2 0.223685f
C2412 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t106 GNDA_2 0.191478f
C2413 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n18 GNDA_2 0.242936f
C2414 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t44 GNDA_2 0.191478f
C2415 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n19 GNDA_2 0.260887f
C2416 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t11 GNDA_2 0.191478f
C2417 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n20 GNDA_2 0.260887f
C2418 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t52 GNDA_2 0.191478f
C2419 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n21 GNDA_2 0.260887f
C2420 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t123 GNDA_2 0.191478f
C2421 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n22 GNDA_2 0.260887f
C2422 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t14 GNDA_2 0.191478f
C2423 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n23 GNDA_2 0.260887f
C2424 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t117 GNDA_2 0.191478f
C2425 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n24 GNDA_2 0.260887f
C2426 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t75 GNDA_2 0.191478f
C2427 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n25 GNDA_2 0.260887f
C2428 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t110 GNDA_2 0.191478f
C2429 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n26 GNDA_2 0.260887f
C2430 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t66 GNDA_2 0.191478f
C2431 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n27 GNDA_2 0.260887f
C2432 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t32 GNDA_2 0.191478f
C2433 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n28 GNDA_2 0.260887f
C2434 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t140 GNDA_2 0.191478f
C2435 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n29 GNDA_2 0.260887f
C2436 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t27 GNDA_2 0.191478f
C2437 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n30 GNDA_2 0.260887f
C2438 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t134 GNDA_2 0.191478f
C2439 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n31 GNDA_2 0.260887f
C2440 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t87 GNDA_2 0.191478f
C2441 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n32 GNDA_2 0.260887f
C2442 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t125 GNDA_2 0.191478f
C2443 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n33 GNDA_2 0.260887f
C2444 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t82 GNDA_2 0.191478f
C2445 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n34 GNDA_2 0.260887f
C2446 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t49 GNDA_2 0.191478f
C2447 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n35 GNDA_2 0.260887f
C2448 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t86 GNDA_2 0.191478f
C2449 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n36 GNDA_2 0.240444f
C2450 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t121 GNDA_2 0.36001f
C2451 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t116 GNDA_2 0.36001f
C2452 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t22 GNDA_2 0.35871f
C2453 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t41 GNDA_2 0.377961f
C2454 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t73 GNDA_2 0.19267f
C2455 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n37 GNDA_2 0.222493f
C2456 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t112 GNDA_2 0.35871f
C2457 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t59 GNDA_2 0.377961f
C2458 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t101 GNDA_2 0.19267f
C2459 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n38 GNDA_2 0.204542f
C2460 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n39 GNDA_2 0.204542f
C2461 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t57 GNDA_2 0.19267f
C2462 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t25 GNDA_2 0.377961f
C2463 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t74 GNDA_2 0.454191f
C2464 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t0 GNDA_2 0.317638f
C2465 VOUT+.n0 GNDA_2 0.035859f
C2466 VOUT+.t7 GNDA_2 0.052295f
C2467 VOUT+.t18 GNDA_2 0.052295f
C2468 VOUT+.n1 GNDA_2 0.112362f
C2469 VOUT+.n2 GNDA_2 0.275831f
C2470 VOUT+.n3 GNDA_2 0.035859f
C2471 VOUT+.n4 GNDA_2 0.237916f
C2472 VOUT+.t14 GNDA_2 0.052295f
C2473 VOUT+.t1 GNDA_2 0.052295f
C2474 VOUT+.n5 GNDA_2 0.112362f
C2475 VOUT+.n6 GNDA_2 0.284527f
C2476 VOUT+.n7 GNDA_2 0.159855f
C2477 VOUT+.t13 GNDA_2 0.052295f
C2478 VOUT+.t4 GNDA_2 0.052295f
C2479 VOUT+.n8 GNDA_2 0.112362f
C2480 VOUT+.n9 GNDA_2 0.271284f
C2481 VOUT+.n10 GNDA_2 0.127531f
C2482 VOUT+.n11 GNDA_2 0.035859f
C2483 VOUT+.n12 GNDA_2 0.185038f
C2484 VOUT+.n13 GNDA_2 0.035859f
C2485 VOUT+.n14 GNDA_2 0.035859f
C2486 VOUT+.n15 GNDA_2 0.035859f
C2487 VOUT+.n16 GNDA_2 0.035859f
C2488 VOUT+.n17 GNDA_2 0.082365f
C2489 VOUT+.n18 GNDA_2 0.096372f
C2490 VOUT+.n19 GNDA_2 0.074707f
C2491 VOUT+.n22 GNDA_2 0.038101f
C2492 VOUT+.n24 GNDA_2 0.038101f
C2493 VOUT+.n27 GNDA_2 0.05603f
C2494 VOUT+.n28 GNDA_2 0.093384f
C2495 VOUT+.n29 GNDA_2 0.059362f
C2496 VOUT+.n30 GNDA_2 0.05603f
C2497 VOUT+.n32 GNDA_2 0.038101f
C2498 VOUT+.n33 GNDA_2 0.035523f
C2499 VOUT+.n34 GNDA_2 0.038101f
C2500 VOUT+.n35 GNDA_2 0.049307f
C2501 VOUT+.n36 GNDA_2 0.071138f
C2502 VOUT+.n37 GNDA_2 0.069229f
C2503 VOUT+.n38 GNDA_2 0.049307f
C2504 VOUT+.n39 GNDA_2 0.049307f
C2505 VOUT+.n40 GNDA_2 0.069229f
C2506 VOUT+.n41 GNDA_2 0.069229f
C2507 VOUT+.n42 GNDA_2 0.049307f
C2508 VOUT+.n43 GNDA_2 0.078936f
C2509 VOUT+.t10 GNDA_2 0.044824f
C2510 VOUT+.t16 GNDA_2 0.044824f
C2511 VOUT+.n44 GNDA_2 0.091845f
C2512 VOUT+.n45 GNDA_2 0.237078f
C2513 VOUT+.t0 GNDA_2 0.044824f
C2514 VOUT+.t11 GNDA_2 0.044824f
C2515 VOUT+.n46 GNDA_2 0.091845f
C2516 VOUT+.n47 GNDA_2 0.237078f
C2517 VOUT+.t9 GNDA_2 0.044824f
C2518 VOUT+.t2 GNDA_2 0.044824f
C2519 VOUT+.n48 GNDA_2 0.091845f
C2520 VOUT+.n49 GNDA_2 0.234689f
C2521 VOUT+.n50 GNDA_2 0.056999f
C2522 VOUT+.t6 GNDA_2 0.044824f
C2523 VOUT+.t8 GNDA_2 0.044824f
C2524 VOUT+.n51 GNDA_2 0.091845f
C2525 VOUT+.n52 GNDA_2 0.234689f
C2526 VOUT+.n53 GNDA_2 0.032309f
C2527 VOUT+.t15 GNDA_2 0.044824f
C2528 VOUT+.t17 GNDA_2 0.044824f
C2529 VOUT+.n54 GNDA_2 0.091845f
C2530 VOUT+.n55 GNDA_2 0.234689f
C2531 VOUT+.n56 GNDA_2 0.032309f
C2532 VOUT+.n57 GNDA_2 0.056999f
C2533 VOUT+.t5 GNDA_2 0.044824f
C2534 VOUT+.t12 GNDA_2 0.044824f
C2535 VOUT+.n58 GNDA_2 0.091845f
C2536 VOUT+.n59 GNDA_2 0.234689f
C2537 VOUT+.n60 GNDA_2 0.037686f
C2538 VOUT+.n61 GNDA_2 0.022412f
C2539 VOUT+.n62 GNDA_2 0.022412f
C2540 VOUT+.n63 GNDA_2 0.037686f
C2541 VOUT+.n64 GNDA_2 0.069229f
C2542 VOUT+.n65 GNDA_2 0.096906f
C2543 VOUT+.n66 GNDA_2 0.120749f
C2544 VOUT+.n67 GNDA_2 0.169f
C2545 VOUT+.n68 GNDA_2 0.049307f
C2546 VOUT+.n69 GNDA_2 0.080684f
C2547 VOUT+.n70 GNDA_2 0.049307f
C2548 VOUT+.n71 GNDA_2 0.080684f
C2549 VOUT+.n72 GNDA_2 0.049307f
C2550 VOUT+.n73 GNDA_2 0.049307f
C2551 VOUT+.n74 GNDA_2 0.049307f
C2552 VOUT+.n75 GNDA_2 0.080684f
C2553 VOUT+.n76 GNDA_2 0.049307f
C2554 VOUT+.n77 GNDA_2 0.07396f
C2555 VOUT+.n78 GNDA_2 0.394453f
C2556 VOUT+.n80 GNDA_2 0.074707f
C2557 VOUT+.n81 GNDA_2 0.038101f
C2558 VOUT+.n83 GNDA_2 0.038101f
C2559 VOUT+.n86 GNDA_2 0.074707f
C2560 VOUT+.n87 GNDA_2 0.387729f
C2561 VOUT+.n88 GNDA_2 0.494934f
C2562 VOUT+.n91 GNDA_2 0.05603f
C2563 VOUT+.n92 GNDA_2 0.05603f
C2564 VOUT+.n93 GNDA_2 0.05603f
C2565 VOUT+.n94 GNDA_2 0.05603f
C2566 VOUT+.n95 GNDA_2 0.164346f
C2567 VOUT+.n96 GNDA_2 0.05603f
C2568 VOUT+.t99 GNDA_2 0.298828f
C2569 VOUT+.t58 GNDA_2 0.303918f
C2570 VOUT+.t159 GNDA_2 0.298828f
C2571 VOUT+.n97 GNDA_2 0.200354f
C2572 VOUT+.n98 GNDA_2 0.130737f
C2573 VOUT+.t60 GNDA_2 0.303281f
C2574 VOUT+.t65 GNDA_2 0.303281f
C2575 VOUT+.t109 GNDA_2 0.303281f
C2576 VOUT+.t84 GNDA_2 0.303281f
C2577 VOUT+.t122 GNDA_2 0.303281f
C2578 VOUT+.t157 GNDA_2 0.303281f
C2579 VOUT+.t138 GNDA_2 0.303281f
C2580 VOUT+.t29 GNDA_2 0.303281f
C2581 VOUT+.t70 GNDA_2 0.303281f
C2582 VOUT+.t114 GNDA_2 0.303281f
C2583 VOUT+.t93 GNDA_2 0.303281f
C2584 VOUT+.t126 GNDA_2 0.303281f
C2585 VOUT+.t90 GNDA_2 0.298828f
C2586 VOUT+.n99 GNDA_2 0.200992f
C2587 VOUT+.t48 GNDA_2 0.298828f
C2588 VOUT+.n100 GNDA_2 0.257022f
C2589 VOUT+.t69 GNDA_2 0.298828f
C2590 VOUT+.n101 GNDA_2 0.257022f
C2591 VOUT+.t24 GNDA_2 0.298828f
C2592 VOUT+.n102 GNDA_2 0.257022f
C2593 VOUT+.t136 GNDA_2 0.298828f
C2594 VOUT+.n103 GNDA_2 0.257022f
C2595 VOUT+.t100 GNDA_2 0.298828f
C2596 VOUT+.n104 GNDA_2 0.257022f
C2597 VOUT+.t120 GNDA_2 0.298828f
C2598 VOUT+.n105 GNDA_2 0.257022f
C2599 VOUT+.t81 GNDA_2 0.298828f
C2600 VOUT+.n106 GNDA_2 0.257022f
C2601 VOUT+.t42 GNDA_2 0.298828f
C2602 VOUT+.n107 GNDA_2 0.257022f
C2603 VOUT+.t64 GNDA_2 0.298828f
C2604 VOUT+.n108 GNDA_2 0.257022f
C2605 VOUT+.t161 GNDA_2 0.298828f
C2606 VOUT+.n109 GNDA_2 0.257022f
C2607 VOUT+.t158 GNDA_2 0.298828f
C2608 VOUT+.n110 GNDA_2 0.257022f
C2609 VOUT+.t56 GNDA_2 0.298828f
C2610 VOUT+.t155 GNDA_2 0.303918f
C2611 VOUT+.t124 GNDA_2 0.298828f
C2612 VOUT+.n111 GNDA_2 0.200354f
C2613 VOUT+.n112 GNDA_2 0.242798f
C2614 VOUT+.t142 GNDA_2 0.303918f
C2615 VOUT+.t116 GNDA_2 0.298828f
C2616 VOUT+.n113 GNDA_2 0.200354f
C2617 VOUT+.t118 GNDA_2 0.298828f
C2618 VOUT+.t117 GNDA_2 0.303918f
C2619 VOUT+.t66 GNDA_2 0.298828f
C2620 VOUT+.n114 GNDA_2 0.200354f
C2621 VOUT+.n115 GNDA_2 0.242798f
C2622 VOUT+.t30 GNDA_2 0.303918f
C2623 VOUT+.t150 GNDA_2 0.298828f
C2624 VOUT+.n116 GNDA_2 0.200354f
C2625 VOUT+.t151 GNDA_2 0.298828f
C2626 VOUT+.t149 GNDA_2 0.303918f
C2627 VOUT+.t106 GNDA_2 0.298828f
C2628 VOUT+.n117 GNDA_2 0.200354f
C2629 VOUT+.n118 GNDA_2 0.242798f
C2630 VOUT+.t98 GNDA_2 0.303918f
C2631 VOUT+.t57 GNDA_2 0.298828f
C2632 VOUT+.n119 GNDA_2 0.200354f
C2633 VOUT+.t110 GNDA_2 0.298828f
C2634 VOUT+.t102 GNDA_2 0.303918f
C2635 VOUT+.t47 GNDA_2 0.298828f
C2636 VOUT+.n120 GNDA_2 0.200354f
C2637 VOUT+.n121 GNDA_2 0.242798f
C2638 VOUT+.t62 GNDA_2 0.303918f
C2639 VOUT+.t34 GNDA_2 0.298828f
C2640 VOUT+.n122 GNDA_2 0.200354f
C2641 VOUT+.t39 GNDA_2 0.298828f
C2642 VOUT+.t36 GNDA_2 0.303918f
C2643 VOUT+.t131 GNDA_2 0.298828f
C2644 VOUT+.n123 GNDA_2 0.200354f
C2645 VOUT+.n124 GNDA_2 0.242798f
C2646 VOUT+.t19 GNDA_2 0.303918f
C2647 VOUT+.t146 GNDA_2 0.298828f
C2648 VOUT+.n125 GNDA_2 0.200354f
C2649 VOUT+.t148 GNDA_2 0.298828f
C2650 VOUT+.t147 GNDA_2 0.303918f
C2651 VOUT+.t101 GNDA_2 0.298828f
C2652 VOUT+.n126 GNDA_2 0.200354f
C2653 VOUT+.n127 GNDA_2 0.242798f
C2654 VOUT+.t67 GNDA_2 0.303918f
C2655 VOUT+.t43 GNDA_2 0.298828f
C2656 VOUT+.n128 GNDA_2 0.200354f
C2657 VOUT+.t45 GNDA_2 0.298828f
C2658 VOUT+.t44 GNDA_2 0.303918f
C2659 VOUT+.t139 GNDA_2 0.298828f
C2660 VOUT+.n129 GNDA_2 0.200354f
C2661 VOUT+.n130 GNDA_2 0.242798f
C2662 VOUT+.t112 GNDA_2 0.303918f
C2663 VOUT+.t85 GNDA_2 0.298828f
C2664 VOUT+.n131 GNDA_2 0.200354f
C2665 VOUT+.t87 GNDA_2 0.298828f
C2666 VOUT+.t86 GNDA_2 0.303918f
C2667 VOUT+.t31 GNDA_2 0.298828f
C2668 VOUT+.n132 GNDA_2 0.200354f
C2669 VOUT+.n133 GNDA_2 0.242798f
C2670 VOUT+.t140 GNDA_2 0.303918f
C2671 VOUT+.t121 GNDA_2 0.298828f
C2672 VOUT+.n134 GNDA_2 0.195685f
C2673 VOUT+.t50 GNDA_2 0.303918f
C2674 VOUT+.t103 GNDA_2 0.298828f
C2675 VOUT+.n135 GNDA_2 0.195685f
C2676 VOUT+.t88 GNDA_2 0.303918f
C2677 VOUT+.t137 GNDA_2 0.298828f
C2678 VOUT+.n136 GNDA_2 0.195685f
C2679 VOUT+.t25 GNDA_2 0.303518f
C2680 VOUT+.t152 GNDA_2 0.303518f
C2681 VOUT+.t53 GNDA_2 0.303531f
C2682 VOUT+.t92 GNDA_2 0.303531f
C2683 VOUT+.t125 GNDA_2 0.303518f
C2684 VOUT+.t108 GNDA_2 0.303531f
C2685 VOUT+.t144 GNDA_2 0.303531f
C2686 VOUT+.t111 GNDA_2 0.298828f
C2687 VOUT+.n137 GNDA_2 0.204477f
C2688 VOUT+.t68 GNDA_2 0.298828f
C2689 VOUT+.n138 GNDA_2 0.260507f
C2690 VOUT+.t97 GNDA_2 0.298828f
C2691 VOUT+.n139 GNDA_2 0.26052f
C2692 VOUT+.t54 GNDA_2 0.298828f
C2693 VOUT+.n140 GNDA_2 0.260507f
C2694 VOUT+.t154 GNDA_2 0.298828f
C2695 VOUT+.n141 GNDA_2 0.260507f
C2696 VOUT+.t119 GNDA_2 0.298828f
C2697 VOUT+.n142 GNDA_2 0.26052f
C2698 VOUT+.t141 GNDA_2 0.298828f
C2699 VOUT+.n143 GNDA_2 0.26052f
C2700 VOUT+.t105 GNDA_2 0.298828f
C2701 VOUT+.n144 GNDA_2 0.191437f
C2702 VOUT+.t61 GNDA_2 0.298828f
C2703 VOUT+.n145 GNDA_2 0.191437f
C2704 VOUT+.t89 GNDA_2 0.298828f
C2705 VOUT+.n146 GNDA_2 0.191437f
C2706 VOUT+.t46 GNDA_2 0.298828f
C2707 VOUT+.n147 GNDA_2 0.130737f
C2708 VOUT+.t41 GNDA_2 0.298828f
C2709 VOUT+.n148 GNDA_2 0.130737f
C2710 VOUT+.t76 GNDA_2 0.298828f
C2711 VOUT+.t33 GNDA_2 0.303918f
C2712 VOUT+.t145 GNDA_2 0.298828f
C2713 VOUT+.n149 GNDA_2 0.200354f
C2714 VOUT+.n150 GNDA_2 0.186768f
C2715 VOUT+.t83 GNDA_2 0.303918f
C2716 VOUT+.t77 GNDA_2 0.298828f
C2717 VOUT+.n151 GNDA_2 0.200354f
C2718 VOUT+.t113 GNDA_2 0.298828f
C2719 VOUT+.t71 GNDA_2 0.303918f
C2720 VOUT+.t32 GNDA_2 0.298828f
C2721 VOUT+.n152 GNDA_2 0.200354f
C2722 VOUT+.n153 GNDA_2 0.242798f
C2723 VOUT+.t107 GNDA_2 0.303918f
C2724 VOUT+.t78 GNDA_2 0.298828f
C2725 VOUT+.n154 GNDA_2 0.200354f
C2726 VOUT+.t80 GNDA_2 0.298828f
C2727 VOUT+.t79 GNDA_2 0.303918f
C2728 VOUT+.t23 GNDA_2 0.298828f
C2729 VOUT+.n155 GNDA_2 0.200354f
C2730 VOUT+.n156 GNDA_2 0.242798f
C2731 VOUT+.t63 GNDA_2 0.303918f
C2732 VOUT+.t35 GNDA_2 0.298828f
C2733 VOUT+.n157 GNDA_2 0.200354f
C2734 VOUT+.t37 GNDA_2 0.298828f
C2735 VOUT+.t38 GNDA_2 0.303918f
C2736 VOUT+.t132 GNDA_2 0.298828f
C2737 VOUT+.n158 GNDA_2 0.200354f
C2738 VOUT+.n159 GNDA_2 0.242798f
C2739 VOUT+.t104 GNDA_2 0.303918f
C2740 VOUT+.t73 GNDA_2 0.298828f
C2741 VOUT+.n160 GNDA_2 0.200354f
C2742 VOUT+.t75 GNDA_2 0.298828f
C2743 VOUT+.t74 GNDA_2 0.303918f
C2744 VOUT+.t160 GNDA_2 0.298828f
C2745 VOUT+.n161 GNDA_2 0.200354f
C2746 VOUT+.n162 GNDA_2 0.242798f
C2747 VOUT+.t59 GNDA_2 0.303918f
C2748 VOUT+.t26 GNDA_2 0.298828f
C2749 VOUT+.n163 GNDA_2 0.200354f
C2750 VOUT+.t28 GNDA_2 0.298828f
C2751 VOUT+.t27 GNDA_2 0.303918f
C2752 VOUT+.t127 GNDA_2 0.298828f
C2753 VOUT+.n164 GNDA_2 0.200354f
C2754 VOUT+.n165 GNDA_2 0.242798f
C2755 VOUT+.t156 GNDA_2 0.303918f
C2756 VOUT+.t133 GNDA_2 0.298828f
C2757 VOUT+.n166 GNDA_2 0.200354f
C2758 VOUT+.t135 GNDA_2 0.298828f
C2759 VOUT+.t134 GNDA_2 0.303918f
C2760 VOUT+.t91 GNDA_2 0.298828f
C2761 VOUT+.n167 GNDA_2 0.200354f
C2762 VOUT+.n168 GNDA_2 0.242798f
C2763 VOUT+.t55 GNDA_2 0.303918f
C2764 VOUT+.t20 GNDA_2 0.298828f
C2765 VOUT+.n169 GNDA_2 0.200354f
C2766 VOUT+.t22 GNDA_2 0.298828f
C2767 VOUT+.t21 GNDA_2 0.303918f
C2768 VOUT+.t123 GNDA_2 0.298828f
C2769 VOUT+.n170 GNDA_2 0.200354f
C2770 VOUT+.n171 GNDA_2 0.242798f
C2771 VOUT+.t153 GNDA_2 0.303918f
C2772 VOUT+.t128 GNDA_2 0.298828f
C2773 VOUT+.n172 GNDA_2 0.200354f
C2774 VOUT+.t130 GNDA_2 0.298828f
C2775 VOUT+.t129 GNDA_2 0.303918f
C2776 VOUT+.t82 GNDA_2 0.298828f
C2777 VOUT+.n173 GNDA_2 0.200354f
C2778 VOUT+.n174 GNDA_2 0.242798f
C2779 VOUT+.t115 GNDA_2 0.303918f
C2780 VOUT+.t94 GNDA_2 0.298828f
C2781 VOUT+.n175 GNDA_2 0.200354f
C2782 VOUT+.t96 GNDA_2 0.298828f
C2783 VOUT+.t95 GNDA_2 0.303918f
C2784 VOUT+.t40 GNDA_2 0.298828f
C2785 VOUT+.n176 GNDA_2 0.200354f
C2786 VOUT+.n177 GNDA_2 0.242798f
C2787 VOUT+.t51 GNDA_2 0.303918f
C2788 VOUT+.t143 GNDA_2 0.298828f
C2789 VOUT+.n178 GNDA_2 0.200354f
C2790 VOUT+.t52 GNDA_2 0.298828f
C2791 VOUT+.n179 GNDA_2 0.242798f
C2792 VOUT+.t49 GNDA_2 0.298828f
C2793 VOUT+.n180 GNDA_2 0.127936f
C2794 VOUT+.t72 GNDA_2 0.298828f
C2795 VOUT+.n181 GNDA_2 0.33338f
C2796 VOUT+.n182 GNDA_2 0.274548f
C2797 VOUT+.n183 GNDA_2 0.05603f
C2798 VOUT+.n184 GNDA_2 0.05603f
C2799 VOUT+.n186 GNDA_2 0.504272f
C2800 VOUT+.n187 GNDA_2 0.056444f
C2801 VOUT+.n188 GNDA_2 1.06457f
C2802 VOUT+.n189 GNDA_2 0.038101f
C2803 VOUT+.n191 GNDA_2 0.035859f
C2804 VOUT+.n192 GNDA_2 1.05524f
C2805 VOUT+.n194 GNDA_2 0.038101f
C2806 VOUT+.n195 GNDA_2 0.074707f
C2807 VOUT+.n196 GNDA_2 0.257739f
C2808 VOUT+.t3 GNDA_2 0.085603f
C2809 VOUT+.n197 GNDA_2 0.42035f
C2810 VDDA.n16 GNDA_2 0.126984f
C2811 VDDA.n17 GNDA_2 0.155202f
C2812 VDDA.n18 GNDA_2 0.126984f
C2813 VDDA.n32 GNDA_2 0.014794f
C2814 VDDA.n34 GNDA_2 0.015342f
C2815 VDDA.n36 GNDA_2 0.013698f
C2816 VDDA.n38 GNDA_2 0.014794f
C2817 VDDA.n40 GNDA_2 0.015342f
C2818 VDDA.t395 GNDA_2 0.102098f
C2819 VDDA.t382 GNDA_2 0.102468f
C2820 VDDA.t18 GNDA_2 0.096989f
C2821 VDDA.t108 GNDA_2 0.102098f
C2822 VDDA.t87 GNDA_2 0.102468f
C2823 VDDA.t410 GNDA_2 0.096989f
C2824 VDDA.t379 GNDA_2 0.102098f
C2825 VDDA.t143 GNDA_2 0.102468f
C2826 VDDA.t171 GNDA_2 0.096989f
C2827 VDDA.t409 GNDA_2 0.102098f
C2828 VDDA.t17 GNDA_2 0.102468f
C2829 VDDA.t81 GNDA_2 0.096989f
C2830 VDDA.t101 GNDA_2 0.102098f
C2831 VDDA.t104 GNDA_2 0.102468f
C2832 VDDA.t107 GNDA_2 0.096989f
C2833 VDDA.n42 GNDA_2 0.068437f
C2834 VDDA.t82 GNDA_2 0.0545f
C2835 VDDA.n43 GNDA_2 0.074255f
C2836 VDDA.t144 GNDA_2 0.0545f
C2837 VDDA.n44 GNDA_2 0.074255f
C2838 VDDA.t88 GNDA_2 0.0545f
C2839 VDDA.n45 GNDA_2 0.074255f
C2840 VDDA.t151 GNDA_2 0.0545f
C2841 VDDA.n46 GNDA_2 0.074255f
C2842 VDDA.t369 GNDA_2 0.292019f
C2843 VDDA.n48 GNDA_2 1.23658f
C2844 VDDA.n49 GNDA_2 0.014794f
C2845 VDDA.n50 GNDA_2 0.015342f
C2846 VDDA.n58 GNDA_2 0.014794f
C2847 VDDA.n59 GNDA_2 0.013698f
C2848 VDDA.n60 GNDA_2 0.013698f
C2849 VDDA.n68 GNDA_2 0.015342f
C2850 VDDA.n69 GNDA_2 0.015342f
C2851 VDDA.n70 GNDA_2 0.014794f
C2852 VDDA.n78 GNDA_2 0.013698f
C2853 VDDA.n79 GNDA_2 0.014794f
C2854 VDDA.n80 GNDA_2 0.015342f
C2855 VDDA.n88 GNDA_2 0.014794f
C2856 VDDA.n89 GNDA_2 0.013698f
C2857 VDDA.n90 GNDA_2 0.013698f
C2858 VDDA.n98 GNDA_2 0.045863f
C2859 VDDA.n101 GNDA_2 7.59079f
C2860 VDDA.n115 GNDA_2 0.014794f
C2861 VDDA.n119 GNDA_2 0.015342f
C2862 VDDA.n123 GNDA_2 0.013698f
C2863 VDDA.n127 GNDA_2 0.014794f
C2864 VDDA.n131 GNDA_2 0.015342f
C2865 VDDA.n136 GNDA_2 0.042737f
C2866 VDDA.n142 GNDA_2 0.014794f
C2867 VDDA.n143 GNDA_2 0.013698f
C2868 VDDA.n144 GNDA_2 0.013698f
C2869 VDDA.n150 GNDA_2 0.015342f
C2870 VDDA.n151 GNDA_2 0.015342f
C2871 VDDA.n152 GNDA_2 0.014794f
C2872 VDDA.n158 GNDA_2 0.013698f
C2873 VDDA.n159 GNDA_2 0.014794f
C2874 VDDA.n160 GNDA_2 0.015342f
C2875 VDDA.n166 GNDA_2 0.014794f
C2876 VDDA.n167 GNDA_2 0.013698f
C2877 VDDA.n168 GNDA_2 0.013698f
C2878 VDDA.n174 GNDA_2 0.015342f
C2879 VDDA.n175 GNDA_2 0.015342f
C2880 VDDA.t54 GNDA_2 0.010959f
C2881 VDDA.t20 GNDA_2 0.010959f
C2882 VDDA.n180 GNDA_2 0.028292f
C2883 VDDA.n181 GNDA_2 0.096637f
C2884 VDDA.t305 GNDA_2 0.038566f
C2885 VDDA.n186 GNDA_2 0.016587f
C2886 VDDA.n187 GNDA_2 0.053731f
C2887 VDDA.t283 GNDA_2 0.016358f
C2888 VDDA.t337 GNDA_2 0.032442f
C2889 VDDA.n192 GNDA_2 0.016059f
C2890 VDDA.n193 GNDA_2 0.046771f
C2891 VDDA.t363 GNDA_2 0.022739f
C2892 VDDA.t361 GNDA_2 0.01132f
C2893 VDDA.n194 GNDA_2 0.016059f
C2894 VDDA.n195 GNDA_2 0.046771f
C2895 VDDA.n196 GNDA_2 0.016059f
C2896 VDDA.n197 GNDA_2 0.046771f
C2897 VDDA.n198 GNDA_2 0.016059f
C2898 VDDA.n199 GNDA_2 0.046771f
C2899 VDDA.n200 GNDA_2 0.016059f
C2900 VDDA.n201 GNDA_2 0.052166f
C2901 VDDA.n202 GNDA_2 0.024187f
C2902 VDDA.n203 GNDA_2 0.072732f
C2903 VDDA.t362 GNDA_2 0.05449f
C2904 VDDA.t11 GNDA_2 0.042739f
C2905 VDDA.t393 GNDA_2 0.042739f
C2906 VDDA.t95 GNDA_2 0.042739f
C2907 VDDA.t180 GNDA_2 0.042739f
C2908 VDDA.t83 GNDA_2 0.042739f
C2909 VDDA.t35 GNDA_2 0.042739f
C2910 VDDA.t89 GNDA_2 0.042739f
C2911 VDDA.t204 GNDA_2 0.042739f
C2912 VDDA.t50 GNDA_2 0.042739f
C2913 VDDA.t156 GNDA_2 0.042739f
C2914 VDDA.t328 GNDA_2 0.05449f
C2915 VDDA.t329 GNDA_2 0.022739f
C2916 VDDA.n204 GNDA_2 0.072732f
C2917 VDDA.t327 GNDA_2 0.01132f
C2918 VDDA.n205 GNDA_2 0.023738f
C2919 VDDA.n206 GNDA_2 0.025487f
C2920 VDDA.n218 GNDA_2 0.015458f
C2921 VDDA.n219 GNDA_2 0.015219f
C2922 VDDA.n220 GNDA_2 0.119457f
C2923 VDDA.n221 GNDA_2 0.015219f
C2924 VDDA.n222 GNDA_2 0.063683f
C2925 VDDA.n223 GNDA_2 0.015219f
C2926 VDDA.n224 GNDA_2 0.063683f
C2927 VDDA.n225 GNDA_2 0.015219f
C2928 VDDA.n226 GNDA_2 0.063683f
C2929 VDDA.n227 GNDA_2 0.015219f
C2930 VDDA.n228 GNDA_2 0.085601f
C2931 VDDA.n229 GNDA_2 0.038355f
C2932 VDDA.n233 GNDA_2 0.11671f
C2933 VDDA.n234 GNDA_2 0.047461f
C2934 VDDA.t277 GNDA_2 0.013032f
C2935 VDDA.n235 GNDA_2 0.040036f
C2936 VDDA.t276 GNDA_2 0.032467f
C2937 VDDA.t76 GNDA_2 0.024109f
C2938 VDDA.t118 GNDA_2 0.024109f
C2939 VDDA.t74 GNDA_2 0.024109f
C2940 VDDA.t97 GNDA_2 0.024109f
C2941 VDDA.t128 GNDA_2 0.024109f
C2942 VDDA.t75 GNDA_2 0.024109f
C2943 VDDA.t185 GNDA_2 0.024109f
C2944 VDDA.t113 GNDA_2 0.024109f
C2945 VDDA.t43 GNDA_2 0.024109f
C2946 VDDA.t32 GNDA_2 0.024109f
C2947 VDDA.t301 GNDA_2 0.032467f
C2948 VDDA.t302 GNDA_2 0.013032f
C2949 VDDA.n236 GNDA_2 0.040036f
C2950 VDDA.n237 GNDA_2 0.028696f
C2951 VDDA.n238 GNDA_2 0.166566f
C2952 VDDA.n239 GNDA_2 0.032328f
C2953 VDDA.n241 GNDA_2 0.11671f
C2954 VDDA.n244 GNDA_2 0.124929f
C2955 VDDA.t203 GNDA_2 0.010959f
C2956 VDDA.t130 GNDA_2 0.010959f
C2957 VDDA.n245 GNDA_2 0.028292f
C2958 VDDA.n246 GNDA_2 0.096637f
C2959 VDDA.t265 GNDA_2 0.038566f
C2960 VDDA.n249 GNDA_2 0.015342f
C2961 VDDA.n262 GNDA_2 0.012978f
C2962 VDDA.n265 GNDA_2 0.014794f
C2963 VDDA.n267 GNDA_2 0.015342f
C2964 VDDA.n269 GNDA_2 0.013698f
C2965 VDDA.n271 GNDA_2 0.014794f
C2966 VDDA.n273 GNDA_2 0.015342f
C2967 VDDA.n274 GNDA_2 0.014038f
C2968 VDDA.t412 GNDA_2 0.215762f
C2969 VDDA.t414 GNDA_2 0.215762f
C2970 VDDA.t415 GNDA_2 0.204985f
C2971 VDDA.n283 GNDA_2 0.39674f
C2972 VDDA.n284 GNDA_2 0.209478f
C2973 VDDA.t413 GNDA_2 0.202486f
C2974 VDDA.n285 GNDA_2 0.271825f
C2975 VDDA.n286 GNDA_2 0.143743f
C2976 VDDA.n291 GNDA_2 0.103559f
C2977 VDDA.n292 GNDA_2 0.103559f
C2978 VDDA.n294 GNDA_2 0.048826f
C2979 VDDA.n298 GNDA_2 0.048826f
C2980 VDDA.n300 GNDA_2 0.048826f
C2981 VDDA.n302 GNDA_2 0.048826f
C2982 VDDA.n304 GNDA_2 0.048826f
C2983 VDDA.n306 GNDA_2 0.048826f
C2984 VDDA.n308 GNDA_2 0.048826f
C2985 VDDA.n310 GNDA_2 0.048826f
C2986 VDDA.n312 GNDA_2 0.048826f
C2987 VDDA.n314 GNDA_2 0.048826f
C2988 VDDA.n318 GNDA_2 0.048826f
C2989 VDDA.n320 GNDA_2 0.048826f
C2990 VDDA.n322 GNDA_2 0.048826f
C2991 VDDA.n324 GNDA_2 0.048826f
C2992 VDDA.n326 GNDA_2 0.048826f
C2993 VDDA.n328 GNDA_2 0.048826f
C2994 VDDA.n330 GNDA_2 0.048826f
C2995 VDDA.n332 GNDA_2 0.066533f
C2996 VDDA.n333 GNDA_2 0.021353f
C2997 VDDA.n336 GNDA_2 0.022514f
C2998 VDDA.t258 GNDA_2 0.018955f
C2999 VDDA.t210 GNDA_2 0.015342f
C3000 VDDA.t188 GNDA_2 0.015342f
C3001 VDDA.t77 GNDA_2 0.015342f
C3002 VDDA.t13 GNDA_2 0.015342f
C3003 VDDA.t62 GNDA_2 0.015342f
C3004 VDDA.t206 GNDA_2 0.015342f
C3005 VDDA.t214 GNDA_2 0.015342f
C3006 VDDA.t37 GNDA_2 0.015342f
C3007 VDDA.t114 GNDA_2 0.015342f
C3008 VDDA.t194 GNDA_2 0.015342f
C3009 VDDA.t126 GNDA_2 0.015342f
C3010 VDDA.t208 GNDA_2 0.015342f
C3011 VDDA.t216 GNDA_2 0.015342f
C3012 VDDA.t162 GNDA_2 0.015342f
C3013 VDDA.t376 GNDA_2 0.015342f
C3014 VDDA.t186 GNDA_2 0.015342f
C3015 VDDA.t29 GNDA_2 0.015342f
C3016 VDDA.t212 GNDA_2 0.015342f
C3017 VDDA.t295 GNDA_2 0.023313f
C3018 VDDA.n337 GNDA_2 0.019434f
C3019 VDDA.n340 GNDA_2 0.01508f
C3020 VDDA.n341 GNDA_2 0.049636f
C3021 VDDA.n342 GNDA_2 0.049636f
C3022 VDDA.n343 GNDA_2 0.020108f
C3023 VDDA.n346 GNDA_2 0.023637f
C3024 VDDA.t261 GNDA_2 0.01911f
C3025 VDDA.t154 GNDA_2 0.015342f
C3026 VDDA.t158 GNDA_2 0.015342f
C3027 VDDA.t64 GNDA_2 0.015342f
C3028 VDDA.t192 GNDA_2 0.015342f
C3029 VDDA.t365 GNDA_2 0.015342f
C3030 VDDA.t66 GNDA_2 0.015342f
C3031 VDDA.t68 GNDA_2 0.015342f
C3032 VDDA.t7 GNDA_2 0.015342f
C3033 VDDA.t15 GNDA_2 0.015342f
C3034 VDDA.t46 GNDA_2 0.015342f
C3035 VDDA.t39 GNDA_2 0.015342f
C3036 VDDA.t5 GNDA_2 0.015342f
C3037 VDDA.t70 GNDA_2 0.015342f
C3038 VDDA.t160 GNDA_2 0.015342f
C3039 VDDA.t190 GNDA_2 0.015342f
C3040 VDDA.t1 GNDA_2 0.015342f
C3041 VDDA.t196 GNDA_2 0.015342f
C3042 VDDA.t33 GNDA_2 0.015342f
C3043 VDDA.t343 GNDA_2 0.022957f
C3044 VDDA.n347 GNDA_2 0.018511f
C3045 VDDA.n350 GNDA_2 0.01508f
C3046 VDDA.n351 GNDA_2 0.105525f
C3047 VDDA.n352 GNDA_2 0.09534f
C3048 VDDA.n357 GNDA_2 0.075067f
C3049 VDDA.n358 GNDA_2 0.075067f
C3050 VDDA.t278 GNDA_2 0.026128f
C3051 VDDA.n359 GNDA_2 0.010016f
C3052 VDDA.n360 GNDA_2 0.02132f
C3053 VDDA.n361 GNDA_2 0.02132f
C3054 VDDA.n362 GNDA_2 0.02132f
C3055 VDDA.n363 GNDA_2 0.02132f
C3056 VDDA.n364 GNDA_2 0.02132f
C3057 VDDA.n365 GNDA_2 0.02132f
C3058 VDDA.n366 GNDA_2 0.02132f
C3059 VDDA.n367 GNDA_2 0.02132f
C3060 VDDA.n393 GNDA_2 0.051232f
C3061 VDDA.t279 GNDA_2 0.054337f
C3062 VDDA.t387 GNDA_2 0.055889f
C3063 VDDA.t145 GNDA_2 0.055889f
C3064 VDDA.t380 GNDA_2 0.055889f
C3065 VDDA.t119 GNDA_2 0.055889f
C3066 VDDA.t147 GNDA_2 0.055889f
C3067 VDDA.t407 GNDA_2 0.055889f
C3068 VDDA.t383 GNDA_2 0.055889f
C3069 VDDA.t367 GNDA_2 0.055889f
C3070 VDDA.t172 GNDA_2 0.055889f
C3071 VDDA.t385 GNDA_2 0.055889f
C3072 VDDA.t102 GNDA_2 0.055889f
C3073 VDDA.t405 GNDA_2 0.055889f
C3074 VDDA.t121 GNDA_2 0.055889f
C3075 VDDA.t149 GNDA_2 0.055889f
C3076 VDDA.t105 GNDA_2 0.055889f
C3077 VDDA.t396 GNDA_2 0.055889f
C3078 VDDA.t356 GNDA_2 0.054337f
C3079 VDDA.n410 GNDA_2 0.051232f
C3080 VDDA.t355 GNDA_2 0.026128f
C3081 VDDA.n413 GNDA_2 0.010553f
C3082 VDDA.n414 GNDA_2 0.104418f
C3083 VDDA.n415 GNDA_2 0.07329f
C3084 VDDA.n416 GNDA_2 0.07329f
C3085 VDDA.n417 GNDA_2 0.07329f
C3086 VDDA.n418 GNDA_2 0.07329f
C3087 VDDA.n419 GNDA_2 0.07329f
C3088 VDDA.n420 GNDA_2 0.07329f
C3089 VDDA.n421 GNDA_2 0.07329f
C3090 VDDA.n422 GNDA_2 0.061802f
C3091 VDDA.n423 GNDA_2 0.07047f
C3092 VDDA.n425 GNDA_2 0.033519f
C3093 VDDA.t350 GNDA_2 0.02265f
C3094 VDDA.t164 GNDA_2 0.014064f
C3095 VDDA.t152 GNDA_2 0.014064f
C3096 VDDA.t319 GNDA_2 0.022163f
C3097 VDDA.n426 GNDA_2 0.032005f
C3098 VDDA.n428 GNDA_2 0.128551f
C3099 VDDA.n429 GNDA_2 0.096984f
C3100 VDDA.n434 GNDA_2 0.035068f
C3101 VDDA.n435 GNDA_2 0.035068f
C3102 VDDA.n438 GNDA_2 0.031828f
C3103 VDDA.t340 GNDA_2 0.022161f
C3104 VDDA.t232 GNDA_2 0.014064f
C3105 VDDA.t218 GNDA_2 0.014064f
C3106 VDDA.t255 GNDA_2 0.022161f
C3107 VDDA.n439 GNDA_2 0.031828f
C3108 VDDA.n441 GNDA_2 0.019375f
C3109 VDDA.n442 GNDA_2 0.019537f
C3110 VDDA.t285 GNDA_2 0.02015f
C3111 VDDA.t224 GNDA_2 0.014064f
C3112 VDDA.t246 GNDA_2 0.014064f
C3113 VDDA.t238 GNDA_2 0.014064f
C3114 VDDA.t222 GNDA_2 0.014064f
C3115 VDDA.t359 GNDA_2 0.02015f
C3116 VDDA.n443 GNDA_2 0.019537f
C3117 VDDA.n444 GNDA_2 0.019375f
C3118 VDDA.n451 GNDA_2 0.031828f
C3119 VDDA.t331 GNDA_2 0.022161f
C3120 VDDA.t228 GNDA_2 0.014064f
C3121 VDDA.t248 GNDA_2 0.014064f
C3122 VDDA.t240 GNDA_2 0.014064f
C3123 VDDA.t226 GNDA_2 0.014064f
C3124 VDDA.t244 GNDA_2 0.014064f
C3125 VDDA.t234 GNDA_2 0.014064f
C3126 VDDA.t236 GNDA_2 0.014064f
C3127 VDDA.t220 GNDA_2 0.014064f
C3128 VDDA.t346 GNDA_2 0.022161f
C3129 VDDA.n452 GNDA_2 0.031828f
C3130 VDDA.n454 GNDA_2 0.019375f
C3131 VDDA.n455 GNDA_2 0.019537f
C3132 VDDA.t298 GNDA_2 0.02015f
C3133 VDDA.t252 GNDA_2 0.014064f
C3134 VDDA.t242 GNDA_2 0.014064f
C3135 VDDA.t230 GNDA_2 0.014064f
C3136 VDDA.t250 GNDA_2 0.014064f
C3137 VDDA.t334 GNDA_2 0.02015f
C3138 VDDA.n456 GNDA_2 0.019537f
C3139 VDDA.n457 GNDA_2 0.02052f
C3140 VDDA.n459 GNDA_2 0.059321f
C3141 VDDA.n461 GNDA_2 0.043646f
C3142 VDDA.n462 GNDA_2 0.043121f
C3143 VDDA.n463 GNDA_2 0.045364f
C3144 VDDA.n464 GNDA_2 0.035701f
C3145 VDDA.n465 GNDA_2 0.040632f
C3146 VDDA.n466 GNDA_2 0.040632f
C3147 VDDA.n467 GNDA_2 0.040632f
C3148 VDDA.n468 GNDA_2 0.035701f
C3149 VDDA.n469 GNDA_2 0.045364f
C3150 VDDA.n470 GNDA_2 0.043121f
C3151 VDDA.n472 GNDA_2 0.043646f
C3152 VDDA.n474 GNDA_2 0.043646f
C3153 VDDA.n475 GNDA_2 0.043121f
C3154 VDDA.n476 GNDA_2 0.051391f
C3155 VDDA.n477 GNDA_2 0.042824f
C3156 VDDA.n478 GNDA_2 0.105636f
C3157 VDDA.n479 GNDA_2 0.089313f
C3158 VDDA.n484 GNDA_2 0.051506f
C3159 VDDA.n485 GNDA_2 0.054793f
C3160 VDDA.n486 GNDA_2 0.015342f
C3161 VDDA.n493 GNDA_2 0.014794f
C3162 VDDA.n494 GNDA_2 0.013698f
C3163 VDDA.n495 GNDA_2 0.013698f
C3164 VDDA.n503 GNDA_2 0.015342f
C3165 VDDA.n504 GNDA_2 0.015342f
C3166 VDDA.n505 GNDA_2 0.014794f
C3167 VDDA.n513 GNDA_2 0.013698f
C3168 VDDA.n514 GNDA_2 0.014794f
C3169 VDDA.n515 GNDA_2 0.015342f
C3170 VDDA.n523 GNDA_2 0.014794f
C3171 VDDA.n524 GNDA_2 0.013698f
C3172 VDDA.n525 GNDA_2 0.013698f
C3173 VDDA.n533 GNDA_2 0.045863f
C3174 VDDA.n536 GNDA_2 7.58379f
C3175 VDDA.n549 GNDA_2 0.042737f
C3176 VDDA.n550 GNDA_2 0.015342f
C3177 VDDA.n551 GNDA_2 0.014794f
C3178 VDDA.n552 GNDA_2 0.013698f
C3179 VDDA.n553 GNDA_2 0.013698f
C3180 VDDA.n554 GNDA_2 0.014794f
C3181 VDDA.n555 GNDA_2 0.015342f
C3182 VDDA.n556 GNDA_2 0.015342f
C3183 VDDA.n557 GNDA_2 0.014794f
C3184 VDDA.n558 GNDA_2 0.013698f
C3185 VDDA.n559 GNDA_2 0.013698f
C3186 VDDA.n560 GNDA_2 0.014794f
C3187 VDDA.n561 GNDA_2 0.015342f
C3188 VDDA.n562 GNDA_2 0.015342f
C3189 VDDA.n563 GNDA_2 0.014794f
C3190 VDDA.n564 GNDA_2 0.013698f
C3191 VDDA.n565 GNDA_2 0.013698f
C3192 VDDA.n566 GNDA_2 0.014794f
C3193 VDDA.n567 GNDA_2 0.015342f
C3194 VDDA.n608 GNDA_2 1.46737f
C3195 VDDA.n611 GNDA_2 0.489852f
C3196 VDDA.n615 GNDA_2 0.486565f
C3197 VDDA.n617 GNDA_2 0.097532f
C3198 VDDA.t168 GNDA_2 0.010959f
C3199 VDDA.t49 GNDA_2 0.010959f
C3200 VDDA.n618 GNDA_2 0.028292f
C3201 VDDA.n619 GNDA_2 0.096637f
C3202 VDDA.t199 GNDA_2 0.010959f
C3203 VDDA.t45 GNDA_2 0.010959f
C3204 VDDA.n620 GNDA_2 0.028292f
C3205 VDDA.n621 GNDA_2 0.096637f
C3206 VDDA.t57 GNDA_2 0.010959f
C3207 VDDA.t133 GNDA_2 0.010959f
C3208 VDDA.n622 GNDA_2 0.028292f
C3209 VDDA.n623 GNDA_2 0.096637f
C3210 VDDA.t176 GNDA_2 0.010959f
C3211 VDDA.t42 GNDA_2 0.010959f
C3212 VDDA.n624 GNDA_2 0.028292f
C3213 VDDA.n625 GNDA_2 0.096637f
C3214 VDDA.n626 GNDA_2 0.10717f
C3215 VDDA.t263 GNDA_2 0.013296f
C3216 VDDA.n627 GNDA_2 0.034789f
C3217 VDDA.n628 GNDA_2 0.129008f
C3218 VDDA.t264 GNDA_2 0.083555f
C3219 VDDA.t175 GNDA_2 0.064291f
C3220 VDDA.t41 GNDA_2 0.063884f
C3221 VDDA.t56 GNDA_2 0.063419f
C3222 VDDA.t132 GNDA_2 0.064291f
C3223 VDDA.t198 GNDA_2 0.064291f
C3224 VDDA.t44 GNDA_2 0.064291f
C3225 VDDA.t167 GNDA_2 0.064291f
C3226 VDDA.t48 GNDA_2 0.064291f
C3227 VDDA.t202 GNDA_2 0.064291f
C3228 VDDA.t129 GNDA_2 0.064291f
C3229 VDDA.t292 GNDA_2 0.083555f
C3230 VDDA.t293 GNDA_2 0.038566f
C3231 VDDA.n629 GNDA_2 0.129008f
C3232 VDDA.t291 GNDA_2 0.013296f
C3233 VDDA.n630 GNDA_2 0.034789f
C3234 VDDA.n631 GNDA_2 0.041966f
C3235 VDDA.n632 GNDA_2 0.032328f
C3236 VDDA.n633 GNDA_2 0.124929f
C3237 VDDA.n636 GNDA_2 0.056437f
C3238 VDDA.n637 GNDA_2 0.056437f
C3239 VDDA.n640 GNDA_2 0.072776f
C3240 VDDA.n642 GNDA_2 0.102464f
C3241 VDDA.t375 GNDA_2 0.029132f
C3242 VDDA.t58 GNDA_2 0.029132f
C3243 VDDA.t27 GNDA_2 0.029132f
C3244 VDDA.t378 GNDA_2 0.029132f
C3245 VDDA.t307 GNDA_2 0.038969f
C3246 VDDA.t308 GNDA_2 0.016358f
C3247 VDDA.n643 GNDA_2 0.046145f
C3248 VDDA.n644 GNDA_2 0.012817f
C3249 VDDA.n645 GNDA_2 0.123718f
C3250 VDDA.n646 GNDA_2 0.016587f
C3251 VDDA.n647 GNDA_2 0.053731f
C3252 VDDA.n648 GNDA_2 0.026849f
C3253 VDDA.n653 GNDA_2 0.075982f
C3254 VDDA.t321 GNDA_2 0.01132f
C3255 VDDA.n654 GNDA_2 0.014556f
C3256 VDDA.t274 GNDA_2 0.029132f
C3257 VDDA.t272 GNDA_2 0.01132f
C3258 VDDA.n655 GNDA_2 0.029636f
C3259 VDDA.n656 GNDA_2 0.072732f
C3260 VDDA.t273 GNDA_2 0.05449f
C3261 VDDA.t85 GNDA_2 0.042739f
C3262 VDDA.t322 GNDA_2 0.05449f
C3263 VDDA.t323 GNDA_2 0.022739f
C3264 VDDA.n657 GNDA_2 0.072732f
C3265 VDDA.n658 GNDA_2 0.029202f
C3266 VDDA.n659 GNDA_2 0.035996f
C3267 VDDA.n663 GNDA_2 0.026849f
C3268 VDDA.n665 GNDA_2 0.014246f
C3269 VDDA.n667 GNDA_2 0.058629f
C3270 VDDA.n668 GNDA_2 0.023915f
C3271 VDDA.t290 GNDA_2 0.011866f
C3272 VDDA.n669 GNDA_2 0.035728f
C3273 VDDA.t288 GNDA_2 0.031808f
C3274 VDDA.t134 GNDA_2 0.024109f
C3275 VDDA.t270 GNDA_2 0.031808f
C3276 VDDA.t271 GNDA_2 0.011866f
C3277 VDDA.n670 GNDA_2 0.035728f
C3278 VDDA.n671 GNDA_2 0.023481f
C3279 VDDA.n672 GNDA_2 0.035996f
C3280 VDDA.n673 GNDA_2 0.026849f
C3281 VDDA.n675 GNDA_2 0.014246f
C3282 VDDA.n679 GNDA_2 0.048218f
C3283 VDDA.n680 GNDA_2 0.048218f
C3284 VDDA.n682 GNDA_2 0.026849f
C3285 VDDA.n685 GNDA_2 0.01564f
C3286 VDDA.t268 GNDA_2 0.016358f
C3287 VDDA.t338 GNDA_2 0.016358f
C3288 VDDA.n686 GNDA_2 0.030844f
C3289 VDDA.n687 GNDA_2 0.02662f
C3290 VDDA.t267 GNDA_2 0.032442f
C3291 VDDA.t372 GNDA_2 0.029132f
C3292 VDDA.t373 GNDA_2 0.029132f
C3293 VDDA.t25 GNDA_2 0.029132f
C3294 VDDA.t72 GNDA_2 0.029132f
C3295 VDDA.t282 GNDA_2 0.038969f
C3296 VDDA.n688 GNDA_2 0.046145f
C3297 VDDA.n689 GNDA_2 0.012817f
C3298 VDDA.n690 GNDA_2 0.123719f
C3299 VDDA.n693 GNDA_2 0.016059f
C3300 VDDA.n694 GNDA_2 0.046771f
C3301 VDDA.t312 GNDA_2 0.01132f
C3302 VDDA.n695 GNDA_2 0.016059f
C3303 VDDA.n696 GNDA_2 0.046771f
C3304 VDDA.n697 GNDA_2 0.016059f
C3305 VDDA.n698 GNDA_2 0.046771f
C3306 VDDA.n699 GNDA_2 0.016059f
C3307 VDDA.n700 GNDA_2 0.046771f
C3308 VDDA.n701 GNDA_2 0.016059f
C3309 VDDA.n702 GNDA_2 0.052166f
C3310 VDDA.n703 GNDA_2 0.024187f
C3311 VDDA.t314 GNDA_2 0.022739f
C3312 VDDA.n704 GNDA_2 0.072732f
C3313 VDDA.t313 GNDA_2 0.05449f
C3314 VDDA.t99 GNDA_2 0.042739f
C3315 VDDA.t79 GNDA_2 0.042739f
C3316 VDDA.t182 GNDA_2 0.042739f
C3317 VDDA.t9 GNDA_2 0.042739f
C3318 VDDA.t178 GNDA_2 0.042739f
C3319 VDDA.t3 GNDA_2 0.042739f
C3320 VDDA.t60 GNDA_2 0.042739f
C3321 VDDA.t200 GNDA_2 0.042739f
C3322 VDDA.t169 GNDA_2 0.042739f
C3323 VDDA.t116 GNDA_2 0.042739f
C3324 VDDA.t353 GNDA_2 0.05449f
C3325 VDDA.t354 GNDA_2 0.022739f
C3326 VDDA.n705 GNDA_2 0.072732f
C3327 VDDA.t352 GNDA_2 0.01132f
C3328 VDDA.n706 GNDA_2 0.023738f
C3329 VDDA.n707 GNDA_2 0.025484f
C3330 VDDA.n709 GNDA_2 0.072778f
C3331 VDDA.n711 GNDA_2 0.102464f
C3332 VDDA.n712 GNDA_2 0.056437f
C3333 VDDA.n722 GNDA_2 0.015458f
C3334 VDDA.n723 GNDA_2 0.015219f
C3335 VDDA.n724 GNDA_2 0.119457f
C3336 VDDA.n725 GNDA_2 0.015219f
C3337 VDDA.n726 GNDA_2 0.063683f
C3338 VDDA.n727 GNDA_2 0.015219f
C3339 VDDA.n728 GNDA_2 0.063683f
C3340 VDDA.n729 GNDA_2 0.015219f
C3341 VDDA.n730 GNDA_2 0.063683f
C3342 VDDA.n731 GNDA_2 0.015219f
C3343 VDDA.n732 GNDA_2 0.085601f
C3344 VDDA.n733 GNDA_2 0.038355f
C3345 VDDA.n735 GNDA_2 0.11671f
C3346 VDDA.n737 GNDA_2 0.11671f
C3347 VDDA.n739 GNDA_2 0.047461f
C3348 VDDA.t326 GNDA_2 0.013032f
C3349 VDDA.n740 GNDA_2 0.040036f
C3350 VDDA.t325 GNDA_2 0.032467f
C3351 VDDA.t142 GNDA_2 0.024109f
C3352 VDDA.t174 GNDA_2 0.024109f
C3353 VDDA.t21 GNDA_2 0.024109f
C3354 VDDA.t0 GNDA_2 0.024109f
C3355 VDDA.t52 GNDA_2 0.024109f
C3356 VDDA.t398 GNDA_2 0.024109f
C3357 VDDA.t165 GNDA_2 0.024109f
C3358 VDDA.t125 GNDA_2 0.024109f
C3359 VDDA.t98 GNDA_2 0.024109f
C3360 VDDA.t112 GNDA_2 0.024109f
C3361 VDDA.t310 GNDA_2 0.032467f
C3362 VDDA.t311 GNDA_2 0.013032f
C3363 VDDA.n741 GNDA_2 0.040036f
C3364 VDDA.n742 GNDA_2 0.028696f
C3365 VDDA.n743 GNDA_2 0.166566f
C3366 VDDA.n744 GNDA_2 0.032328f
C3367 VDDA.n746 GNDA_2 0.124929f
C3368 VDDA.n747 GNDA_2 0.124929f
C3369 VDDA.n750 GNDA_2 0.056437f
C3370 VDDA.n752 GNDA_2 0.032328f
C3371 VDDA.t138 GNDA_2 0.010959f
C3372 VDDA.t141 GNDA_2 0.010959f
C3373 VDDA.n753 GNDA_2 0.028292f
C3374 VDDA.n754 GNDA_2 0.096637f
C3375 VDDA.t400 GNDA_2 0.010959f
C3376 VDDA.t124 GNDA_2 0.010959f
C3377 VDDA.n755 GNDA_2 0.028292f
C3378 VDDA.n756 GNDA_2 0.096637f
C3379 VDDA.t371 GNDA_2 0.010959f
C3380 VDDA.t390 GNDA_2 0.010959f
C3381 VDDA.n757 GNDA_2 0.028292f
C3382 VDDA.n758 GNDA_2 0.096637f
C3383 VDDA.t392 GNDA_2 0.010959f
C3384 VDDA.t111 GNDA_2 0.010959f
C3385 VDDA.n759 GNDA_2 0.028292f
C3386 VDDA.n760 GNDA_2 0.096637f
C3387 VDDA.n761 GNDA_2 0.041966f
C3388 VDDA.t303 GNDA_2 0.013296f
C3389 VDDA.n762 GNDA_2 0.034789f
C3390 VDDA.n763 GNDA_2 0.129008f
C3391 VDDA.t304 GNDA_2 0.083555f
C3392 VDDA.t391 GNDA_2 0.064291f
C3393 VDDA.t110 GNDA_2 0.064291f
C3394 VDDA.t370 GNDA_2 0.064291f
C3395 VDDA.t389 GNDA_2 0.064291f
C3396 VDDA.t399 GNDA_2 0.064291f
C3397 VDDA.t123 GNDA_2 0.064291f
C3398 VDDA.t137 GNDA_2 0.064291f
C3399 VDDA.t140 GNDA_2 0.064291f
C3400 VDDA.t53 GNDA_2 0.064291f
C3401 VDDA.t19 GNDA_2 0.064291f
C3402 VDDA.t316 GNDA_2 0.083555f
C3403 VDDA.t317 GNDA_2 0.038566f
C3404 VDDA.n764 GNDA_2 0.129008f
C3405 VDDA.t315 GNDA_2 0.013296f
C3406 VDDA.n765 GNDA_2 0.034789f
C3407 VDDA.n766 GNDA_2 0.10717f
C3408 VDDA.n767 GNDA_2 0.097532f
C3409 VDDA.n771 GNDA_2 0.486565f
C3410 VDDA.n772 GNDA_2 0.489852f
C3411 VDDA.n775 GNDA_2 55.692898f
C3412 VDDA.n776 GNDA_2 0.131504f
C3413 VDDA.n777 GNDA_2 0.131504f
C3414 VDDA.n778 GNDA_2 0.131504f
C3415 VDDA.n779 GNDA_2 0.131504f
C3416 VDDA.n780 GNDA_2 0.131504f
C3417 VDDA.n781 GNDA_2 0.131504f
C3418 VDDA.n782 GNDA_2 0.131504f
C3419 VDDA.n783 GNDA_2 0.131504f
C3420 VDDA.n784 GNDA_2 0.131504f
C3421 VDDA.n785 GNDA_2 0.131504f
C3422 VDDA.n786 GNDA_2 0.131504f
C3423 VDDA.n787 GNDA_2 0.131504f
C3424 VDDA.n788 GNDA_2 0.131504f
C3425 VDDA.n789 GNDA_2 0.131504f
C3426 VDDA.n790 GNDA_2 0.131504f
C3427 VDDA.n791 GNDA_2 0.131504f
C3428 VDDA.n792 GNDA_2 0.126984f
C3429 VDDA.n794 GNDA_2 0.131504f
C3430 VDDA.n797 GNDA_2 0.131504f
C3431 VDDA.n800 GNDA_2 0.131504f
C3432 VDDA.n803 GNDA_2 0.131504f
C3433 VDDA.n806 GNDA_2 0.131504f
C3434 VDDA.n809 GNDA_2 0.131504f
C3435 VDDA.n812 GNDA_2 0.131504f
C3436 VDDA.n815 GNDA_2 0.131504f
C3437 VDDA.n818 GNDA_2 0.131504f
C3438 VDDA.n821 GNDA_2 0.131504f
C3439 VDDA.n824 GNDA_2 0.131504f
C3440 VDDA.n827 GNDA_2 0.131504f
C3441 VDDA.n830 GNDA_2 0.131504f
C3442 VDDA.n833 GNDA_2 0.131504f
C3443 VDDA.n836 GNDA_2 0.131504f
C3444 VDDA.n839 GNDA_2 0.131504f
C3445 VDDA.n842 GNDA_2 0.126984f
C3446 VDDA.n843 GNDA_2 0.126984f
C3447 VDDA.n844 GNDA_2 0.126984f
C3448 VDDA.n845 GNDA_2 0.126984f
C3449 VDDA.n846 GNDA_2 0.126984f
C3450 VDDA.n847 GNDA_2 0.126984f
C3451 VDDA.n848 GNDA_2 0.126984f
C3452 VDDA.n849 GNDA_2 0.126984f
C3453 VDDA.n850 GNDA_2 0.126984f
C3454 VDDA.n851 GNDA_2 0.126984f
C3455 VDDA.n852 GNDA_2 0.126984f
C3456 VDDA.n853 GNDA_2 0.126984f
C3457 VDDA.n854 GNDA_2 0.126984f
C3458 VDDA.n855 GNDA_2 0.126984f
C3459 VDDA.n856 GNDA_2 0.126984f
C3460 VDDA.n859 GNDA_2 0.126984f
C3461 VDDA.n861 GNDA_2 0.126984f
C3462 VDDA.n863 GNDA_2 0.126984f
C3463 VDDA.n865 GNDA_2 0.126984f
C3464 VDDA.n867 GNDA_2 0.126984f
C3465 VDDA.n869 GNDA_2 0.126984f
C3466 VDDA.n871 GNDA_2 0.126984f
C3467 VDDA.n873 GNDA_2 0.126984f
C3468 VDDA.n875 GNDA_2 0.126984f
C3469 VDDA.n877 GNDA_2 0.126984f
C3470 VDDA.n879 GNDA_2 0.126984f
C3471 VDDA.n881 GNDA_2 0.126984f
C3472 VDDA.n883 GNDA_2 0.126984f
C3473 VDDA.n885 GNDA_2 0.126984f
C3474 VDDA.n887 GNDA_2 0.126984f
C3475 VDDA.n888 GNDA_2 0.131504f
C3476 VDDA.n889 GNDA_2 54.4512f
C3477 VDDA.n890 GNDA_2 0.858429f
C3478 bgr_11_0.PFET_GATE_10uA.t28 GNDA_2 0.022652f
C3479 bgr_11_0.PFET_GATE_10uA.t20 GNDA_2 0.022652f
C3480 bgr_11_0.PFET_GATE_10uA.n0 GNDA_2 0.079313f
C3481 bgr_11_0.PFET_GATE_10uA.t13 GNDA_2 0.019516f
C3482 bgr_11_0.PFET_GATE_10uA.t24 GNDA_2 0.02885f
C3483 bgr_11_0.PFET_GATE_10uA.n1 GNDA_2 0.031789f
C3484 bgr_11_0.PFET_GATE_10uA.t17 GNDA_2 0.019516f
C3485 bgr_11_0.PFET_GATE_10uA.t25 GNDA_2 0.02885f
C3486 bgr_11_0.PFET_GATE_10uA.n2 GNDA_2 0.031789f
C3487 bgr_11_0.PFET_GATE_10uA.n3 GNDA_2 0.031141f
C3488 bgr_11_0.PFET_GATE_10uA.n4 GNDA_2 0.992009f
C3489 bgr_11_0.PFET_GATE_10uA.t0 GNDA_2 0.348615f
C3490 bgr_11_0.PFET_GATE_10uA.t1 GNDA_2 0.310845f
C3491 bgr_11_0.PFET_GATE_10uA.t9 GNDA_2 0.020017f
C3492 bgr_11_0.PFET_GATE_10uA.t2 GNDA_2 0.020017f
C3493 bgr_11_0.PFET_GATE_10uA.n5 GNDA_2 0.043237f
C3494 bgr_11_0.PFET_GATE_10uA.n6 GNDA_2 1.07309f
C3495 bgr_11_0.PFET_GATE_10uA.t5 GNDA_2 0.020017f
C3496 bgr_11_0.PFET_GATE_10uA.t7 GNDA_2 0.020017f
C3497 bgr_11_0.PFET_GATE_10uA.n7 GNDA_2 0.043237f
C3498 bgr_11_0.PFET_GATE_10uA.n8 GNDA_2 0.437158f
C3499 bgr_11_0.PFET_GATE_10uA.t3 GNDA_2 0.020017f
C3500 bgr_11_0.PFET_GATE_10uA.t6 GNDA_2 0.020017f
C3501 bgr_11_0.PFET_GATE_10uA.n9 GNDA_2 0.043237f
C3502 bgr_11_0.PFET_GATE_10uA.n10 GNDA_2 0.428151f
C3503 bgr_11_0.PFET_GATE_10uA.t4 GNDA_2 0.020017f
C3504 bgr_11_0.PFET_GATE_10uA.t8 GNDA_2 0.020017f
C3505 bgr_11_0.PFET_GATE_10uA.n11 GNDA_2 0.043237f
C3506 bgr_11_0.PFET_GATE_10uA.n12 GNDA_2 0.672012f
C3507 bgr_11_0.PFET_GATE_10uA.n13 GNDA_2 2.87808f
C3508 bgr_11_0.PFET_GATE_10uA.t26 GNDA_2 0.066817f
C3509 bgr_11_0.PFET_GATE_10uA.n14 GNDA_2 1.52702f
C3510 bgr_11_0.PFET_GATE_10uA.t15 GNDA_2 0.019516f
C3511 bgr_11_0.PFET_GATE_10uA.t10 GNDA_2 0.02885f
C3512 bgr_11_0.PFET_GATE_10uA.n15 GNDA_2 0.031789f
C3513 bgr_11_0.PFET_GATE_10uA.t21 GNDA_2 0.019516f
C3514 bgr_11_0.PFET_GATE_10uA.t11 GNDA_2 0.02885f
C3515 bgr_11_0.PFET_GATE_10uA.n16 GNDA_2 0.031789f
C3516 bgr_11_0.PFET_GATE_10uA.n17 GNDA_2 0.031141f
C3517 bgr_11_0.PFET_GATE_10uA.n18 GNDA_2 1.24671f
C3518 bgr_11_0.PFET_GATE_10uA.t14 GNDA_2 0.019516f
C3519 bgr_11_0.PFET_GATE_10uA.t19 GNDA_2 0.019516f
C3520 bgr_11_0.PFET_GATE_10uA.t18 GNDA_2 0.019516f
C3521 bgr_11_0.PFET_GATE_10uA.t27 GNDA_2 0.02885f
C3522 bgr_11_0.PFET_GATE_10uA.n19 GNDA_2 0.035703f
C3523 bgr_11_0.PFET_GATE_10uA.n20 GNDA_2 0.025521f
C3524 bgr_11_0.PFET_GATE_10uA.n21 GNDA_2 0.019891f
C3525 bgr_11_0.PFET_GATE_10uA.t23 GNDA_2 0.019516f
C3526 bgr_11_0.PFET_GATE_10uA.t16 GNDA_2 0.019516f
C3527 bgr_11_0.PFET_GATE_10uA.t12 GNDA_2 0.019516f
C3528 bgr_11_0.PFET_GATE_10uA.t22 GNDA_2 0.02885f
C3529 bgr_11_0.PFET_GATE_10uA.n22 GNDA_2 0.035703f
C3530 bgr_11_0.PFET_GATE_10uA.n23 GNDA_2 0.025521f
C3531 bgr_11_0.PFET_GATE_10uA.n24 GNDA_2 0.019891f
C3532 bgr_11_0.PFET_GATE_10uA.n25 GNDA_2 0.056627f
C3533 bgr_11_0.1st_Vout_2.n0 GNDA_2 1.07305f
C3534 bgr_11_0.1st_Vout_2.n1 GNDA_2 0.297625f
C3535 bgr_11_0.1st_Vout_2.n2 GNDA_2 0.668271f
C3536 bgr_11_0.1st_Vout_2.n3 GNDA_2 0.091542f
C3537 bgr_11_0.1st_Vout_2.n4 GNDA_2 0.158156f
C3538 bgr_11_0.1st_Vout_2.t14 GNDA_2 0.011681f
C3539 bgr_11_0.1st_Vout_2.n6 GNDA_2 0.010675f
C3540 bgr_11_0.1st_Vout_2.n7 GNDA_2 0.115898f
C3541 bgr_11_0.1st_Vout_2.n8 GNDA_2 0.0146f
C3542 bgr_11_0.1st_Vout_2.t15 GNDA_2 0.011528f
C3543 bgr_11_0.1st_Vout_2.t29 GNDA_2 0.194725f
C3544 bgr_11_0.1st_Vout_2.t32 GNDA_2 0.198042f
C3545 bgr_11_0.1st_Vout_2.t27 GNDA_2 0.194725f
C3546 bgr_11_0.1st_Vout_2.t20 GNDA_2 0.194725f
C3547 bgr_11_0.1st_Vout_2.t12 GNDA_2 0.198042f
C3548 bgr_11_0.1st_Vout_2.t13 GNDA_2 0.198042f
C3549 bgr_11_0.1st_Vout_2.t31 GNDA_2 0.194725f
C3550 bgr_11_0.1st_Vout_2.t25 GNDA_2 0.194725f
C3551 bgr_11_0.1st_Vout_2.t19 GNDA_2 0.198042f
C3552 bgr_11_0.1st_Vout_2.t30 GNDA_2 0.198042f
C3553 bgr_11_0.1st_Vout_2.t24 GNDA_2 0.194725f
C3554 bgr_11_0.1st_Vout_2.t18 GNDA_2 0.194725f
C3555 bgr_11_0.1st_Vout_2.t11 GNDA_2 0.198042f
C3556 bgr_11_0.1st_Vout_2.t23 GNDA_2 0.198042f
C3557 bgr_11_0.1st_Vout_2.t17 GNDA_2 0.194725f
C3558 bgr_11_0.1st_Vout_2.t10 GNDA_2 0.194725f
C3559 bgr_11_0.1st_Vout_2.t28 GNDA_2 0.198042f
C3560 bgr_11_0.1st_Vout_2.t8 GNDA_2 0.198042f
C3561 bgr_11_0.1st_Vout_2.t16 GNDA_2 0.194725f
C3562 bgr_11_0.1st_Vout_2.t22 GNDA_2 0.194725f
C3563 bgr_11_0.1st_Vout_2.n9 GNDA_2 0.641071f
C3564 bgr_11_0.1st_Vout_2.n10 GNDA_2 0.010675f
C3565 bgr_11_0.1st_Vout_2.n11 GNDA_2 0.0146f
C3566 bgr_11_0.1st_Vout_2.n12 GNDA_2 0.14235f
C3567 bgr_11_0.1st_Vout_2.t6 GNDA_2 0.044569f
.ends

