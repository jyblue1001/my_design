* NGSPICE file created from pfdpfd.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

.subckt pfdpfd A B VGND VNB VPB VPWR Y
Xsky130_fd_sc_hd__nor2_1_0 sky130_fd_sc_hd__nor2_1_0/A sky130_fd_sc_hd__nor2_1_0/B
+ sky130_fd_sc_hd__nor2_1_0/VGND VNB VPB sky130_fd_sc_hd__nor2_1_0/VPWR sky130_fd_sc_hd__nor2_1_0/Y
+ sky130_fd_sc_hd__nor2_1
.ends

