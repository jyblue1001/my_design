magic
tech sky130A
timestamp 1738187251
<< nwell >>
rect -2400 460 -2160 545
rect -3070 220 -1755 460
rect -500 225 200 1065
<< pwell >>
rect -2565 120 -2550 125
rect -3070 -45 -1755 115
rect -3070 -70 -1815 -45
rect -1760 -70 -1755 -45
rect -3070 -90 -1755 -70
rect -2100 -165 -2080 -90
<< nmos >>
rect -3000 10 -2985 110
rect -2855 10 -2840 110
rect -2710 10 -2695 110
rect -2565 10 -2550 110
rect -2420 10 -2405 110
rect -2275 10 -2260 110
rect -2130 10 -2115 110
rect -1985 10 -1970 110
rect -1840 10 -1825 110
rect -930 -255 -870 145
rect -430 -255 -370 145
rect 70 -255 130 145
<< pmos >>
rect -3000 240 -2985 440
rect -2855 240 -2840 440
rect -2710 240 -2695 440
rect -2565 240 -2550 440
rect -2420 240 -2405 440
rect -2275 240 -2260 440
rect -2130 240 -2115 440
rect -1985 240 -1970 440
rect -1840 240 -1825 440
rect -430 245 -370 1045
rect 70 245 130 1045
<< ndiff >>
rect -3050 95 -3000 110
rect -3050 25 -3035 95
rect -3015 25 -3000 95
rect -3050 10 -3000 25
rect -2985 95 -2935 110
rect -2985 25 -2970 95
rect -2950 25 -2935 95
rect -2985 10 -2935 25
rect -2905 95 -2855 110
rect -2905 25 -2890 95
rect -2870 25 -2855 95
rect -2905 10 -2855 25
rect -2840 95 -2790 110
rect -2840 25 -2825 95
rect -2805 25 -2790 95
rect -2840 10 -2790 25
rect -2760 95 -2710 110
rect -2760 25 -2745 95
rect -2725 25 -2710 95
rect -2760 10 -2710 25
rect -2695 95 -2645 110
rect -2695 25 -2680 95
rect -2660 25 -2645 95
rect -2695 10 -2645 25
rect -2615 95 -2565 110
rect -2615 25 -2600 95
rect -2580 25 -2565 95
rect -2615 10 -2565 25
rect -2550 95 -2500 110
rect -2550 25 -2535 95
rect -2515 25 -2500 95
rect -2550 10 -2500 25
rect -2470 95 -2420 110
rect -2470 25 -2455 95
rect -2435 25 -2420 95
rect -2470 10 -2420 25
rect -2405 95 -2355 110
rect -2405 25 -2390 95
rect -2370 25 -2355 95
rect -2405 10 -2355 25
rect -2325 95 -2275 110
rect -2325 25 -2310 95
rect -2290 25 -2275 95
rect -2325 10 -2275 25
rect -2260 95 -2210 110
rect -2260 25 -2245 95
rect -2225 25 -2210 95
rect -2260 10 -2210 25
rect -2180 95 -2130 110
rect -2180 25 -2165 95
rect -2145 25 -2130 95
rect -2180 10 -2130 25
rect -2115 95 -2065 110
rect -2115 25 -2100 95
rect -2080 25 -2065 95
rect -2115 10 -2065 25
rect -2035 95 -1985 110
rect -2035 25 -2020 95
rect -2000 25 -1985 95
rect -2035 10 -1985 25
rect -1970 95 -1920 110
rect -1970 25 -1955 95
rect -1935 25 -1920 95
rect -1970 10 -1920 25
rect -1890 95 -1840 110
rect -1890 25 -1875 95
rect -1855 25 -1840 95
rect -1890 10 -1840 25
rect -1825 95 -1775 110
rect -1825 25 -1810 95
rect -1790 25 -1775 95
rect -1825 10 -1775 25
rect -980 130 -930 145
rect -980 -240 -965 130
rect -945 -240 -930 130
rect -980 -255 -930 -240
rect -870 130 -820 145
rect -870 -240 -855 130
rect -835 -240 -820 130
rect -870 -255 -820 -240
rect -480 130 -430 145
rect -480 -240 -465 130
rect -445 -240 -430 130
rect -480 -255 -430 -240
rect -370 130 -320 145
rect -370 -240 -355 130
rect -335 -240 -320 130
rect -370 -255 -320 -240
rect 20 130 70 145
rect 20 -240 35 130
rect 55 -240 70 130
rect 20 -255 70 -240
rect 130 130 180 145
rect 130 -240 145 130
rect 165 -240 180 130
rect 130 -255 180 -240
<< pdiff >>
rect -480 1030 -430 1045
rect -3050 425 -3000 440
rect -3050 255 -3035 425
rect -3015 255 -3000 425
rect -3050 240 -3000 255
rect -2985 425 -2935 440
rect -2985 255 -2970 425
rect -2950 255 -2935 425
rect -2985 240 -2935 255
rect -2905 425 -2855 440
rect -2905 255 -2890 425
rect -2870 255 -2855 425
rect -2905 240 -2855 255
rect -2840 425 -2790 440
rect -2840 255 -2825 425
rect -2805 255 -2790 425
rect -2840 240 -2790 255
rect -2760 425 -2710 440
rect -2760 255 -2745 425
rect -2725 255 -2710 425
rect -2760 240 -2710 255
rect -2695 425 -2645 440
rect -2695 255 -2680 425
rect -2660 255 -2645 425
rect -2695 240 -2645 255
rect -2615 425 -2565 440
rect -2615 255 -2600 425
rect -2580 255 -2565 425
rect -2615 240 -2565 255
rect -2550 425 -2500 440
rect -2550 255 -2535 425
rect -2515 255 -2500 425
rect -2550 240 -2500 255
rect -2470 425 -2420 440
rect -2470 255 -2455 425
rect -2435 255 -2420 425
rect -2470 240 -2420 255
rect -2405 425 -2355 440
rect -2405 255 -2390 425
rect -2370 255 -2355 425
rect -2405 240 -2355 255
rect -2325 425 -2275 440
rect -2325 255 -2310 425
rect -2290 255 -2275 425
rect -2325 240 -2275 255
rect -2260 425 -2210 440
rect -2260 255 -2245 425
rect -2225 255 -2210 425
rect -2260 240 -2210 255
rect -2180 425 -2130 440
rect -2180 255 -2165 425
rect -2145 255 -2130 425
rect -2180 240 -2130 255
rect -2115 425 -2065 440
rect -2115 255 -2100 425
rect -2080 255 -2065 425
rect -2115 240 -2065 255
rect -2035 425 -1985 440
rect -2035 255 -2020 425
rect -2000 255 -1985 425
rect -2035 240 -1985 255
rect -1970 425 -1920 440
rect -1970 255 -1955 425
rect -1935 255 -1920 425
rect -1970 240 -1920 255
rect -1890 425 -1840 440
rect -1890 255 -1875 425
rect -1855 255 -1840 425
rect -1890 240 -1840 255
rect -1825 425 -1775 440
rect -1825 255 -1810 425
rect -1790 255 -1775 425
rect -1825 240 -1775 255
rect -480 260 -465 1030
rect -445 260 -430 1030
rect -480 245 -430 260
rect -370 1030 -320 1045
rect -370 260 -355 1030
rect -335 260 -320 1030
rect -370 245 -320 260
rect 20 1030 70 1045
rect 20 260 35 1030
rect 55 260 70 1030
rect 20 245 70 260
rect 130 1030 180 1045
rect 130 260 145 1030
rect 165 260 180 1030
rect 130 245 180 260
<< ndiffc >>
rect -3035 25 -3015 95
rect -2970 25 -2950 95
rect -2890 25 -2870 95
rect -2825 25 -2805 95
rect -2745 25 -2725 95
rect -2680 25 -2660 95
rect -2600 25 -2580 95
rect -2535 25 -2515 95
rect -2455 25 -2435 95
rect -2390 25 -2370 95
rect -2310 25 -2290 95
rect -2245 25 -2225 95
rect -2165 25 -2145 95
rect -2100 25 -2080 95
rect -2020 25 -2000 95
rect -1955 25 -1935 95
rect -1875 25 -1855 95
rect -1810 25 -1790 95
rect -965 -240 -945 130
rect -855 -240 -835 130
rect -465 -240 -445 130
rect -355 -240 -335 130
rect 35 -240 55 130
rect 145 -240 165 130
<< pdiffc >>
rect -3035 255 -3015 425
rect -2970 255 -2950 425
rect -2890 255 -2870 425
rect -2825 255 -2805 425
rect -2745 255 -2725 425
rect -2680 255 -2660 425
rect -2600 255 -2580 425
rect -2535 255 -2515 425
rect -2455 255 -2435 425
rect -2390 255 -2370 425
rect -2310 255 -2290 425
rect -2245 255 -2225 425
rect -2165 255 -2145 425
rect -2100 255 -2080 425
rect -2020 255 -2000 425
rect -1955 255 -1935 425
rect -1875 255 -1855 425
rect -1810 255 -1790 425
rect -465 260 -445 1030
rect -355 260 -335 1030
rect 35 260 55 1030
rect 145 260 165 1030
<< psubdiff >>
rect -2590 -40 -2490 -25
rect -2590 -60 -2575 -40
rect -2505 -60 -2490 -40
rect -2590 -75 -2490 -60
rect -820 130 -770 145
rect -820 -240 -805 130
rect -785 -240 -770 130
rect -820 -255 -770 -240
rect -320 130 -270 145
rect -320 -240 -305 130
rect -285 -240 -270 130
rect -320 -255 -270 -240
rect -30 130 20 145
rect -30 -240 -15 130
rect 5 -240 20 130
rect -30 -255 20 -240
<< nsubdiff >>
rect -2380 510 -2180 525
rect -2380 490 -2365 510
rect -2195 490 -2180 510
rect -2380 475 -2180 490
rect -320 1030 -270 1045
rect -320 260 -305 1030
rect -285 260 -270 1030
rect -320 245 -270 260
rect -30 1030 20 1045
rect -30 260 -15 1030
rect 5 260 20 1030
rect -30 245 20 260
<< psubdiffcont >>
rect -2575 -60 -2505 -40
rect -805 -240 -785 130
rect -305 -240 -285 130
rect -15 -240 5 130
<< nsubdiffcont >>
rect -2365 490 -2195 510
rect -305 260 -285 1030
rect -15 260 5 1030
<< poly >>
rect -1365 1245 395 1260
rect -1365 885 -1350 1245
rect -1485 875 -1350 885
rect -2670 870 -1350 875
rect -1255 1120 85 1135
rect -2670 860 -1470 870
rect -2670 700 -2655 860
rect -1620 715 -1580 725
rect -1620 700 -1610 715
rect -2690 690 -2650 700
rect -2690 670 -2680 690
rect -2660 670 -2650 690
rect -2690 660 -2650 670
rect -2610 695 -1610 700
rect -1590 695 -1580 715
rect -2610 690 -1580 695
rect -2610 670 -2600 690
rect -2580 685 -1580 690
rect -2580 670 -2570 685
rect -2610 660 -2570 670
rect -1255 660 -1240 1120
rect 70 1060 85 1120
rect -430 1045 -370 1060
rect 70 1045 130 1060
rect -2530 650 -1240 660
rect -2530 630 -2520 650
rect -2500 645 -1800 650
rect -2500 630 -2490 645
rect -2530 620 -2490 630
rect -1810 630 -1800 645
rect -1780 645 -1240 650
rect -1780 630 -1770 645
rect -1810 620 -1770 630
rect -2710 580 -1825 595
rect -3000 440 -2985 455
rect -2855 440 -2840 455
rect -2710 440 -2695 580
rect -2565 440 -2550 455
rect -2420 440 -2405 455
rect -2275 440 -2260 455
rect -2130 440 -2115 455
rect -1985 440 -1970 455
rect -1840 440 -1825 580
rect -1620 585 -1580 595
rect -1620 565 -1610 585
rect -1590 565 -1580 585
rect -1620 555 -1580 565
rect -1620 250 -1605 555
rect -3000 185 -2985 240
rect -2855 200 -2840 240
rect -2710 200 -2695 240
rect -2565 225 -2550 240
rect -3065 170 -2985 185
rect -3000 110 -2985 170
rect -2880 190 -2840 200
rect -2880 170 -2870 190
rect -2850 170 -2840 190
rect -2880 160 -2840 170
rect -2735 190 -2695 200
rect -2735 170 -2725 190
rect -2705 170 -2695 190
rect -2670 215 -2550 225
rect -2670 195 -2660 215
rect -2640 210 -2550 215
rect -2640 195 -2630 210
rect -2670 185 -2630 195
rect -2735 160 -2695 170
rect -2855 110 -2840 160
rect -2710 135 -2695 160
rect -2710 120 -2550 135
rect -2710 110 -2695 120
rect -2565 110 -2550 120
rect -2420 110 -2405 240
rect -2275 230 -2260 240
rect -2355 215 -2260 230
rect -2235 215 -2195 225
rect -2130 215 -2115 240
rect -1985 215 -1970 240
rect -1840 225 -1825 240
rect -1620 235 -805 250
rect 380 875 395 1245
rect 435 875 475 885
rect 380 860 445 875
rect 435 855 445 860
rect 465 855 475 875
rect 435 845 475 855
rect 435 245 475 255
rect -430 235 -370 245
rect -830 220 -370 235
rect 70 235 130 245
rect 435 240 445 245
rect 290 235 445 240
rect 70 225 445 235
rect 465 225 475 245
rect 70 220 475 225
rect 435 215 475 220
rect -2355 165 -2340 215
rect -2235 195 -2225 215
rect -2205 200 -1860 215
rect -2205 195 -2195 200
rect -2235 190 -2195 195
rect -2380 155 -2340 165
rect -2195 160 -2155 165
rect -2380 135 -2370 155
rect -2350 135 -2340 155
rect -2380 125 -2340 135
rect -2275 155 -2155 160
rect -2275 145 -2185 155
rect -2275 110 -2260 145
rect -2195 135 -2185 145
rect -2165 135 -2155 155
rect -2195 125 -2155 135
rect -2130 110 -2115 200
rect -1875 165 -1860 200
rect -975 190 -935 200
rect -975 175 -965 190
rect -1755 170 -965 175
rect -945 175 -935 190
rect -945 170 -370 175
rect -2090 150 -2050 160
rect -1875 150 -1825 165
rect -2090 130 -2080 150
rect -2060 135 -2050 150
rect -2060 130 -1970 135
rect -2090 120 -1970 130
rect -1985 110 -1970 120
rect -1840 110 -1825 150
rect -1755 160 -370 170
rect -3000 -5 -2985 10
rect -2855 -5 -2840 10
rect -2710 -5 -2695 10
rect -2565 -5 -2550 10
rect -2420 -120 -2405 10
rect -2275 -5 -2260 10
rect -2130 -5 -2115 10
rect -1985 -5 -1970 10
rect -1840 -5 -1825 10
rect -1945 -15 -1905 -5
rect -1945 -35 -1935 -15
rect -1915 -30 -1905 -15
rect -1755 -30 -1740 160
rect -930 155 -370 160
rect -930 145 -870 155
rect -430 145 -370 155
rect 70 155 295 170
rect 70 145 130 155
rect -1915 -35 -1740 -30
rect -1945 -45 -1740 -35
rect -2040 -80 -1470 -70
rect -2040 -100 -2030 -80
rect -2010 -85 -1810 -80
rect -2010 -100 -2000 -85
rect -2040 -110 -2000 -100
rect -1820 -100 -1810 -85
rect -1790 -85 -1470 -80
rect -1790 -100 -1780 -85
rect -1820 -110 -1780 -100
rect -3065 -135 -2405 -120
rect -2120 -135 -2080 -125
rect -2120 -155 -2110 -135
rect -2090 -150 -2080 -135
rect -1485 -150 -1470 -85
rect -2090 -155 -1600 -150
rect -2120 -165 -1600 -155
rect -1485 -165 -1350 -150
rect -1615 -350 -1600 -165
rect -1615 -360 -1575 -350
rect -1615 -380 -1605 -360
rect -1585 -380 -1575 -360
rect -1615 -390 -1575 -380
rect -1365 -465 -1350 -165
rect 280 125 295 155
rect 435 125 475 135
rect 280 110 445 125
rect 435 105 445 110
rect 465 105 475 125
rect 435 95 475 105
rect 435 -155 475 -145
rect 435 -160 445 -155
rect 385 -175 445 -160
rect 465 -175 475 -155
rect -930 -270 -870 -255
rect -430 -270 -370 -255
rect 70 -270 130 -255
rect -1275 -370 -1235 -360
rect -1275 -390 -1265 -370
rect -1245 -375 -1235 -370
rect 70 -375 85 -270
rect -1245 -390 85 -375
rect -1275 -400 -1235 -390
rect 385 -465 400 -175
rect 435 -185 475 -175
rect -1365 -480 400 -465
<< polycont >>
rect -2680 670 -2660 690
rect -1610 695 -1590 715
rect -2600 670 -2580 690
rect -2520 630 -2500 650
rect -1800 630 -1780 650
rect -1610 565 -1590 585
rect -2870 170 -2850 190
rect -2725 170 -2705 190
rect -2660 195 -2640 215
rect 445 855 465 875
rect 445 225 465 245
rect -2225 195 -2205 215
rect -2370 135 -2350 155
rect -2185 135 -2165 155
rect -965 170 -945 190
rect -2080 130 -2060 150
rect -1935 -35 -1915 -15
rect -2030 -100 -2010 -80
rect -1810 -100 -1790 -80
rect -2110 -155 -2090 -135
rect -1605 -380 -1585 -360
rect 445 105 465 125
rect 445 -175 465 -155
rect -1265 -390 -1245 -370
<< locali >>
rect -475 1030 -435 1040
rect -1620 715 -1580 725
rect -2690 690 -2650 700
rect -2690 670 -2680 690
rect -2660 670 -2650 690
rect -2690 660 -2650 670
rect -2670 435 -2650 660
rect -3045 425 -3005 435
rect -3045 255 -3035 425
rect -3015 255 -3005 425
rect -3045 245 -3005 255
rect -2980 425 -2940 435
rect -2980 255 -2970 425
rect -2950 255 -2940 425
rect -2980 245 -2940 255
rect -2900 425 -2860 435
rect -2900 255 -2890 425
rect -2870 255 -2860 425
rect -2900 245 -2860 255
rect -2835 425 -2795 435
rect -2835 255 -2825 425
rect -2805 255 -2795 425
rect -2835 245 -2795 255
rect -2755 425 -2715 435
rect -2755 255 -2745 425
rect -2725 255 -2715 425
rect -2755 245 -2715 255
rect -2690 425 -2650 435
rect -2690 255 -2680 425
rect -2660 255 -2650 425
rect -2690 245 -2650 255
rect -2610 690 -2570 700
rect -2610 670 -2600 690
rect -2580 670 -2570 690
rect -2610 660 -2570 670
rect -1620 695 -1610 715
rect -1590 695 -1580 715
rect -1620 685 -1580 695
rect -2610 435 -2590 660
rect -2530 650 -2490 660
rect -2530 630 -2520 650
rect -2500 630 -2490 650
rect -2530 620 -2490 630
rect -1810 650 -1770 660
rect -1810 630 -1800 650
rect -1780 630 -1770 650
rect -1810 620 -1770 630
rect -2530 435 -2510 620
rect -1810 530 -1790 620
rect -1620 595 -1600 685
rect -1620 585 -1580 595
rect -1620 565 -1610 585
rect -1590 565 -1580 585
rect -1620 555 -1580 565
rect -2375 510 -2185 520
rect -2375 490 -2365 510
rect -2195 490 -2185 510
rect -2375 480 -2185 490
rect -1810 435 -1790 510
rect -2610 425 -2570 435
rect -2610 255 -2600 425
rect -2580 255 -2570 425
rect -2610 245 -2570 255
rect -2545 425 -2505 435
rect -2545 255 -2535 425
rect -2515 255 -2505 425
rect -2545 245 -2505 255
rect -2465 425 -2425 435
rect -2465 255 -2455 425
rect -2435 255 -2425 425
rect -2465 245 -2425 255
rect -2400 425 -2360 435
rect -2400 255 -2390 425
rect -2370 275 -2360 425
rect -2320 425 -2280 435
rect -2370 255 -2355 275
rect -2400 245 -2355 255
rect -2320 255 -2310 425
rect -2290 255 -2280 425
rect -2320 245 -2280 255
rect -2255 425 -2215 435
rect -2255 255 -2245 425
rect -2225 255 -2215 425
rect -2255 245 -2215 255
rect -2175 425 -2135 435
rect -2175 255 -2165 425
rect -2145 255 -2135 425
rect -2175 245 -2135 255
rect -2110 425 -2070 435
rect -2110 255 -2100 425
rect -2080 255 -2070 425
rect -2110 245 -2070 255
rect -2030 425 -1990 435
rect -2030 255 -2020 425
rect -2000 255 -1990 425
rect -2030 245 -1990 255
rect -1965 425 -1925 435
rect -1965 255 -1955 425
rect -1935 255 -1925 425
rect -1965 245 -1925 255
rect -1885 425 -1845 435
rect -1885 255 -1875 425
rect -1855 255 -1845 425
rect -1885 245 -1845 255
rect -1820 425 -1780 435
rect -1820 255 -1810 425
rect -1790 255 -1780 425
rect -1820 245 -1780 255
rect -475 260 -465 1030
rect -445 260 -435 1030
rect -475 250 -435 260
rect -365 1030 -275 1040
rect -365 260 -355 1030
rect -335 260 -305 1030
rect -285 260 -275 1030
rect -365 250 -275 260
rect -25 1030 65 1040
rect -25 260 -15 1030
rect 5 260 35 1030
rect 55 260 65 1030
rect -25 250 65 260
rect 135 1030 175 1040
rect 135 260 145 1030
rect 165 260 175 1030
rect 515 890 570 900
rect 435 875 475 885
rect 515 875 525 890
rect 435 855 445 875
rect 465 855 525 875
rect 560 855 570 890
rect 435 845 475 855
rect 515 845 570 855
rect 135 250 175 260
rect 515 295 570 305
rect 515 260 525 295
rect 560 260 570 295
rect 435 250 475 255
rect 515 250 570 260
rect -2960 190 -2940 245
rect -2880 190 -2840 200
rect -2960 170 -2870 190
rect -2850 170 -2840 190
rect -2960 105 -2940 170
rect -2880 160 -2840 170
rect -2815 190 -2795 245
rect -2670 225 -2650 245
rect -2670 215 -2630 225
rect -2735 190 -2695 200
rect -2815 170 -2725 190
rect -2705 170 -2695 190
rect -2815 105 -2795 170
rect -2735 160 -2695 170
rect -2670 195 -2660 215
rect -2640 195 -2630 215
rect -2670 185 -2630 195
rect -2670 105 -2650 185
rect -2600 105 -2580 245
rect -2545 105 -2525 245
rect -2445 225 -2425 245
rect -2310 225 -2290 245
rect -2445 205 -2290 225
rect -2445 105 -2425 205
rect -2380 155 -2340 165
rect -2380 135 -2370 155
rect -2350 135 -2340 155
rect -2380 125 -2340 135
rect -2380 105 -2360 125
rect -2310 105 -2290 205
rect -2245 225 -2225 245
rect -2245 215 -2195 225
rect -2245 195 -2225 215
rect -2205 195 -2195 215
rect -2245 190 -2195 195
rect -2245 105 -2225 190
rect -2170 165 -2150 245
rect -2195 155 -2150 165
rect -2195 135 -2185 155
rect -2165 135 -2150 155
rect -2195 125 -2150 135
rect -2090 160 -2070 245
rect -2090 150 -2050 160
rect -2090 130 -2080 150
rect -2060 130 -2050 150
rect -2090 120 -2050 130
rect -2090 105 -2070 120
rect -2020 105 -2000 245
rect -1955 105 -1935 245
rect -975 190 -935 200
rect -975 170 -965 190
rect -945 170 -935 190
rect -975 160 -935 170
rect -965 140 -945 160
rect -465 140 -445 250
rect 145 195 165 250
rect 435 245 540 250
rect 435 225 445 245
rect 465 230 540 245
rect 465 225 475 230
rect 435 215 475 225
rect 145 185 420 195
rect 145 175 1250 185
rect 145 140 165 175
rect 385 165 1250 175
rect -975 130 -935 140
rect -3045 95 -3005 105
rect -3045 25 -3035 95
rect -3015 25 -3005 95
rect -3045 15 -3005 25
rect -2980 95 -2940 105
rect -2980 25 -2970 95
rect -2950 25 -2940 95
rect -2980 15 -2940 25
rect -2900 95 -2860 105
rect -2900 25 -2890 95
rect -2870 25 -2860 95
rect -2900 15 -2860 25
rect -2835 95 -2795 105
rect -2835 25 -2825 95
rect -2805 25 -2795 95
rect -2835 15 -2795 25
rect -2755 95 -2715 105
rect -2755 25 -2745 95
rect -2725 25 -2715 95
rect -2755 15 -2715 25
rect -2690 95 -2650 105
rect -2690 25 -2680 95
rect -2660 25 -2650 95
rect -2690 15 -2650 25
rect -2610 95 -2570 105
rect -2610 25 -2600 95
rect -2580 25 -2570 95
rect -2610 15 -2570 25
rect -2545 95 -2505 105
rect -2545 25 -2535 95
rect -2515 25 -2505 95
rect -2545 15 -2505 25
rect -2465 95 -2425 105
rect -2465 25 -2455 95
rect -2435 25 -2425 95
rect -2465 15 -2425 25
rect -2400 95 -2360 105
rect -2400 25 -2390 95
rect -2370 25 -2360 95
rect -2400 15 -2360 25
rect -2320 95 -2280 105
rect -2320 25 -2310 95
rect -2290 25 -2280 95
rect -2320 15 -2280 25
rect -2255 95 -2215 105
rect -2255 25 -2245 95
rect -2225 25 -2215 95
rect -2255 15 -2215 25
rect -2175 95 -2135 105
rect -2175 25 -2165 95
rect -2145 25 -2135 95
rect -2175 15 -2135 25
rect -2110 95 -2070 105
rect -2110 25 -2100 95
rect -2080 25 -2070 95
rect -2110 15 -2070 25
rect -2030 95 -1990 105
rect -2030 25 -2020 95
rect -2000 25 -1990 95
rect -2030 15 -1990 25
rect -1965 95 -1920 105
rect -1965 25 -1955 95
rect -1935 25 -1920 95
rect -1965 15 -1920 25
rect -1885 95 -1845 105
rect -1885 25 -1875 95
rect -1855 25 -1845 95
rect -1885 15 -1845 25
rect -1820 95 -1780 105
rect -1820 25 -1810 95
rect -1790 25 -1780 95
rect -1820 15 -1780 25
rect -2585 -40 -2495 -30
rect -2585 -60 -2575 -40
rect -2505 -60 -2495 -40
rect -2585 -70 -2495 -60
rect -2100 -125 -2080 15
rect -2020 -70 -2000 15
rect -1945 -5 -1925 15
rect -1945 -15 -1905 -5
rect -1945 -35 -1935 -15
rect -1915 -35 -1905 -15
rect -1945 -45 -1905 -35
rect -1810 -45 -1790 15
rect -2040 -80 -2000 -70
rect -2040 -100 -2030 -80
rect -2010 -100 -2000 -80
rect -2040 -110 -2000 -100
rect -1820 -80 -1780 -70
rect -1820 -100 -1810 -80
rect -1790 -100 -1780 -80
rect -1820 -110 -1780 -100
rect -2120 -135 -2080 -125
rect -2120 -155 -2110 -135
rect -2090 -155 -2080 -135
rect -2120 -165 -2080 -155
rect -975 -200 -965 130
rect -1500 -210 -965 -200
rect -3065 -220 -965 -210
rect -3065 -230 -1470 -220
rect -975 -240 -965 -220
rect -945 -240 -935 130
rect -975 -250 -935 -240
rect -865 130 -775 140
rect -865 -240 -855 130
rect -835 -240 -805 130
rect -785 -240 -775 130
rect -865 -250 -775 -240
rect -475 130 -435 140
rect -475 -240 -465 130
rect -445 -240 -435 130
rect -475 -250 -435 -240
rect -365 130 -275 140
rect -365 -240 -355 130
rect -335 -240 -305 130
rect -285 -240 -275 130
rect -365 -250 -275 -240
rect -25 130 65 140
rect -25 -240 -15 130
rect 5 -240 35 130
rect 55 -240 65 130
rect -25 -250 65 -240
rect 135 130 175 140
rect 135 -240 145 130
rect 165 -240 175 130
rect 435 125 475 135
rect 435 105 445 125
rect 465 120 475 125
rect 465 105 550 120
rect 435 100 550 105
rect 435 95 475 100
rect 515 90 570 100
rect 515 55 525 90
rect 560 55 570 90
rect 515 45 570 55
rect 515 -130 570 -120
rect 435 -155 475 -145
rect 515 -155 525 -130
rect 435 -175 445 -155
rect 465 -165 525 -155
rect 560 -165 570 -130
rect 465 -175 570 -165
rect 435 -185 475 -175
rect 135 -250 175 -240
rect -1615 -360 -1575 -350
rect -1615 -380 -1605 -360
rect -1585 -370 -1575 -360
rect -1275 -370 -1235 -360
rect -1585 -380 -1265 -370
rect -1615 -390 -1265 -380
rect -1245 -390 -1235 -370
rect -1275 -400 -1235 -390
<< viali >>
rect -3035 255 -3015 425
rect -2890 255 -2870 425
rect -2745 255 -2725 425
rect -2365 490 -2195 510
rect -2390 255 -2370 425
rect -2165 255 -2145 425
rect -1875 255 -1855 425
rect -355 260 -335 1030
rect -305 260 -285 1030
rect -15 260 5 1030
rect 35 260 55 1030
rect 525 855 560 890
rect 525 260 560 295
rect -3035 25 -3015 95
rect -2890 25 -2870 95
rect -2745 25 -2725 95
rect -2390 25 -2370 95
rect -2165 25 -2145 95
rect -1875 25 -1855 95
rect -2575 -60 -2505 -40
rect -855 -240 -835 130
rect -805 -240 -785 130
rect -355 -240 -335 130
rect -305 -240 -285 130
rect -15 -240 5 130
rect 35 -240 55 130
rect 525 55 560 90
rect 525 -165 560 -130
<< metal1 >>
rect -1355 1030 180 1045
rect -2380 510 -2180 525
rect -2380 490 -2365 510
rect -2195 490 -2180 510
rect -2380 440 -2180 490
rect -1355 450 -355 1030
rect -1485 440 -355 450
rect -3100 425 -355 440
rect -3100 255 -3035 425
rect -3015 255 -2890 425
rect -2870 255 -2745 425
rect -2725 255 -2390 425
rect -2370 255 -2165 425
rect -2145 255 -1875 425
rect -1855 260 -355 425
rect -335 260 -305 1030
rect -285 260 -15 1030
rect 5 260 35 1030
rect 55 260 180 1030
rect 515 890 570 900
rect 515 855 525 890
rect 560 855 570 890
rect 515 845 570 855
rect -1855 255 180 260
rect -3100 250 180 255
rect 515 295 570 305
rect 515 260 525 295
rect 560 260 570 295
rect 515 250 570 260
rect -3100 240 -1415 250
rect -1360 245 180 250
rect -1350 130 180 145
rect -1350 120 -855 130
rect -1645 110 -855 120
rect -3100 95 -855 110
rect -3100 25 -3035 95
rect -3015 25 -2890 95
rect -2870 25 -2745 95
rect -2725 25 -2390 95
rect -2370 25 -2165 95
rect -2145 25 -1875 95
rect -1855 25 -855 95
rect -3100 10 -855 25
rect -3100 0 -1465 10
rect -2590 -40 -2485 0
rect -2590 -60 -2575 -40
rect -2505 -60 -2485 -40
rect -2590 -75 -2485 -60
rect -1350 -240 -855 10
rect -835 -240 -805 130
rect -785 -240 -355 130
rect -335 -240 -305 130
rect -285 -240 -15 130
rect 5 -240 35 130
rect 55 -240 180 130
rect 515 90 570 100
rect 515 55 525 90
rect 560 55 570 90
rect 515 45 570 55
rect 515 -130 570 -120
rect 515 -165 525 -130
rect 560 -165 570 -130
rect 515 -175 570 -165
rect -1350 -255 180 -240
<< via1 >>
rect 525 855 560 890
rect 525 260 560 295
rect 525 55 560 90
rect 525 -165 560 -130
<< metal2 >>
rect 515 890 570 900
rect 515 855 525 890
rect 560 855 570 890
rect 515 845 570 855
rect 515 295 570 305
rect 515 260 525 295
rect 560 260 570 295
rect 515 250 570 260
rect 515 90 570 100
rect 515 55 525 90
rect 560 55 570 90
rect 515 45 570 55
rect 515 -130 570 -120
rect 515 -165 525 -130
rect 560 -165 570 -130
rect 515 -175 570 -165
<< via2 >>
rect 525 855 560 890
rect 525 260 560 295
rect 525 55 560 90
rect 525 -165 560 -130
<< metal3 >>
rect 690 900 1140 925
rect 515 890 1140 900
rect 515 855 525 890
rect 560 855 1140 890
rect 515 845 1140 855
rect 690 305 1140 845
rect 515 295 1140 305
rect 515 260 525 295
rect 560 260 1140 295
rect 515 250 1140 260
rect 690 235 1140 250
rect 690 100 980 115
rect 515 90 980 100
rect 515 55 525 90
rect 560 55 980 90
rect 515 45 980 55
rect 690 -120 980 45
rect 515 -130 980 -120
rect 515 -165 525 -130
rect 560 -165 980 -130
rect 515 -175 980 -165
<< via3 >>
rect 525 260 560 295
rect 525 55 560 90
<< mimcap >>
rect 705 295 1125 910
rect 705 260 715 295
rect 750 260 1125 295
rect 705 250 1125 260
rect 705 90 965 100
rect 705 55 715 90
rect 750 55 965 90
rect 705 -160 965 55
<< mimcapcontact >>
rect 715 260 750 295
rect 715 55 750 90
<< metal4 >>
rect 515 295 760 305
rect 515 260 525 295
rect 560 260 715 295
rect 750 260 760 295
rect 515 250 760 260
rect 515 90 760 100
rect 515 55 525 90
rect 560 55 715 90
rect 750 55 760 90
rect 515 45 760 55
<< labels >>
flabel locali -3065 -220 -3065 -220 7 FreeSans 400 0 -200 0 I_IN
flabel poly -3065 -125 -3065 -125 7 FreeSans 400 0 -200 0 DOWN_PFD
flabel poly -3065 175 -3065 175 7 FreeSans 400 0 -200 0 UP_PFD
flabel metal1 -3100 340 -3100 340 7 FreeSans 400 0 -200 0 VDDA
flabel metal1 -3100 60 -3100 60 7 FreeSans 400 0 -200 0 GNDA
flabel locali 1250 175 1250 175 3 FreeSans 400 0 80 0 VOUT
flabel poly -2130 -5 -2130 -5 7 FreeSans 400 0 -200 -200 DOWN_b
flabel poly -2670 820 -2670 820 7 FreeSans 400 0 -200 0 UP_b
flabel poly -2120 -165 -2120 -165 7 FreeSans 400 0 -200 -200 DOWN
flabel poly -2710 595 -2710 595 7 FreeSans 400 0 -200 0 UP
<< end >>
