* PEX produced on Mon Feb 24 09:52:34 AM CET 2025 using /foss/tools/osic-multitool/iic-pex.sh with m=3 and s=1
* NGSPICE file created from pfd_cp_lf_magic_2.ext - technology: sky130A

.subckt pfd_cp_lf_magic V_OUT VDDA GNDA F_REF F_VCO I_IN
X0 GNDA.t86 a_6200_5250.t2 a_6200_5250.t3 GNDA.t85 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X1 a_5970_4630.t7 opamp_cell_4_0.VIN- a_6200_5250.t5 VDDA.t88 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X2 pfd_8_0.DOWN_b.t1 VDDA.t130 pfd_8_0.DOWN_PFD_b.t3 GNDA.t55 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X3 a_870_1400.t0 pfd_8_0.QA_b.t3 VDDA.t128 VDDA.t39 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X4 pfd_8_0.DOWN.t1 pfd_8_0.DOWN_b.t2 VDDA.t13 VDDA.t12 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X5 GNDA.t128 GNDA.t126 GNDA.t128 GNDA.t127 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0 ps=0 w=2 l=0.6
X6 VDDA.t26 pfd_8_0.UP_input.t13 opamp_cell_4_0.VIN+.t4 VDDA.t25 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X7 opamp_cell_4_0.n_right.t1 opamp_cell_4_0.VIN+.t6 a_6320_5840.t0 GNDA.t70 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X8 opamp_cell_4_0.n_right.t4 opamp_cell_4_0.n_left.t6 VDDA.t53 VDDA.t52 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X9 pfd_8_0.UP_input.t10 opamp_cell_4_0.n_right.t5 VDDA.t84 VDDA.t83 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X10 pfd_8_0.UP_input.t7 a_6490_4630.t5 GNDA.t69 GNDA.t68 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X11 a_2350_1400.t0 pfd_8_0.before_Reset.t3 GNDA.t72 GNDA.t71 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X12 pfd_8_0.DOWN.t0 pfd_8_0.DOWN_b.t3 GNDA.t48 GNDA.t47 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X13 VDDA.t74 opamp_cell_4_0.p_bias.t7 opamp_cell_4_0.p_bias.t8 VDDA.t73 sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X14 a_n30_1400.t0 F_REF.t0 VDDA.t6 VDDA.t5 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X15 GNDA.t31 pfd_8_0.QA.t3 pfd_8_0.QA_b.t1 GNDA.t30 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X16 a_6200_5250.t1 a_6200_5250.t0 GNDA.t84 GNDA.t83 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X17 a_6200_5250.t4 opamp_cell_4_0.VIN- a_5970_4630.t6 VDDA.t87 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X18 VDDA.t47 opamp_cell_4_0.p_bias.t9 a_5970_4630.t2 VDDA.t46 sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X19 VDDA.t125 VDDA.t122 VDDA.t124 VDDA.t123 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=0 ps=0 w=2 l=0.6
X20 pfd_8_0.DOWN_input.t1 pfd_8_0.DOWN_b.t4 I_IN.t5 VDDA.t7 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X21 VDDA.t121 VDDA.t119 VDDA.t121 VDDA.t120 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0 ps=0 w=2 l=0.6
X22 VDDA.t11 pfd_8_0.UP_input.t14 V_OUT.t5 VDDA.t10 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X23 a_1910_2020.t1 pfd_8_0.QB.t3 GNDA.t33 GNDA.t32 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X24 a_6220_5810.t8 a_6220_5810.t7 GNDA.t40 GNDA.t39 sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0.3125 ps=1.75 w=1.25 l=0.5
X25 GNDA.t138 pfd_8_0.DOWN_input.t3 V_OUT.t1 GNDA.t137 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X26 pfd_8_0.UP.t1 pfd_8_0.UP_PFD_b.t2 VDDA.t86 VDDA.t85 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X27 a_6320_5840.t9 a_6220_5810.t9 GNDA.t140 GNDA.t139 sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0.3125 ps=1.75 w=1.25 l=0.5
X28 pfd_8_0.UP_input.t12 pfd_8_0.UP.t2 pfd_8_0.UP_input.t11 GNDA.t76 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0 ps=0 w=1 l=0.15
X29 pfd_8_0.QA.t1 pfd_8_0.QA_b.t4 GNDA.t1 GNDA.t0 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X30 a_5970_4630.t5 opamp_cell_4_0.p_bias.t10 VDDA.t68 VDDA.t67 sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X31 pfd_8_0.DOWN_input.t0 pfd_8_0.DOWN.t2 I_IN.t4 GNDA.t73 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X32 GNDA.t134 I_IN.t6 opamp_cell_4_0.VIN+.t5 GNDA.t133 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X33 a_1390_1400.t0 pfd_8_0.E.t3 pfd_8_0.E_b.t0 VDDA.t22 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X34 a_870_640.t1 pfd_8_0.QB_b.t3 VDDA.t40 VDDA.t39 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X35 VDDA.t118 VDDA.t115 VDDA.t117 VDDA.t116 sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0 ps=0 w=1 l=0.15
X36 V_OUT.t6 loop_filter_2_0.R1_C1.t0 GNDA.t36 sky130_fd_pr__res_xhigh_po_0p35 l=7.52
X37 VDDA.t17 a_2530_190.t2 a_2200_190.t1 VDDA.t16 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=0.15
X38 GNDA.t125 GNDA.t123 GNDA.t125 GNDA.t124 sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0 ps=0 w=1.25 l=0.5
X39 GNDA.t122 GNDA.t119 GNDA.t121 GNDA.t120 sky130_fd_pr__nfet_01v8 ad=0.25 pd=2 as=0 ps=0 w=0.5 l=0.15
X40 opamp_cell_4_0.p_bias.t6 opamp_cell_4_0.p_bias.t5 VDDA.t76 VDDA.t75 sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X41 VDDA.t114 VDDA.t112 VDDA.t114 VDDA.t113 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0 ps=0 w=2 l=0.6
X42 V_OUT.t4 pfd_8_0.UP_input.t15 VDDA.t72 VDDA.t71 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X43 pfd_8_0.DOWN_input.t2 pfd_8_0.DOWN_b.t5 GNDA.t13 GNDA.t12 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X44 GNDA.t17 a_2530_190.t3 a_2200_190.t0 GNDA.t16 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X45 pfd_8_0.F.t2 pfd_8_0.QB_b.t4 GNDA.t50 GNDA.t49 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X46 GNDA.t118 GNDA.t115 GNDA.t117 GNDA.t116 sky130_fd_pr__nfet_01v8 ad=0.625 pd=3.5 as=0 ps=0 w=1.25 l=0.5
X47 pfd_8_0.UP_input.t16 a_9360_6440.t0 sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X48 V_OUT.t0 pfd_8_0.DOWN_input.t4 GNDA.t136 GNDA.t135 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X49 pfd_8_0.UP_b.t0 pfd_8_0.UP.t3 GNDA.t153 GNDA.t152 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X50 GNDA.t147 pfd_8_0.E_b.t3 pfd_8_0.E.t1 GNDA.t146 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X51 GNDA.t145 a_6220_5810.t10 a_6320_5840.t11 GNDA.t144 sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0.3125 ps=1.75 w=1.25 l=0.5
X52 a_1390_640.t0 pfd_8_0.F.t3 pfd_8_0.F_b.t1 VDDA.t22 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X53 a_2350_1400.t1 pfd_8_0.before_Reset.t4 VDDA.t66 VDDA.t65 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=0.15
X54 opamp_cell_4_0.VIN+.t0 I_IN.t7 GNDA.t25 GNDA.t24 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X55 GNDA.t44 a_6220_5810.t5 a_6220_5810.t6 GNDA.t43 sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0.3125 ps=1.75 w=1.25 l=0.5
X56 GNDA.t114 GNDA.t112 GNDA.t114 GNDA.t113 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0 ps=0 w=0.5 l=0.15
X57 a_5970_4630.t12 a_5970_4630.t11 a_5970_4630.t12 VDDA.t90 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0 ps=0 w=1 l=0.15
X58 pfd_8_0.F_b.t2 pfd_8_0.F.t4 GNDA.t19 GNDA.t18 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X59 VDDA.t9 pfd_8_0.UP_input.t17 V_OUT.t3 VDDA.t8 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X60 GNDA.t156 loop_filter_2_0.R1_C1.t1 sky130_fd_pr__cap_mim_m3_1 l=60 w=69.8
X61 VDDA.t36 pfd_8_0.F.t5 a_490_640.t1 VDDA.t35 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X62 VDDA.t111 VDDA.t109 VDDA.t111 VDDA.t110 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0 ps=0 w=1 l=0.15
X63 GNDA.t111 GNDA.t109 GNDA.t111 GNDA.t110 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0 ps=0 w=2 l=0.6
X64 pfd_8_0.QA_b.t2 pfd_8_0.QA.t4 a_n30_1400.t1 VDDA.t4 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X65 GNDA.t108 GNDA.t106 GNDA.t108 GNDA.t107 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0 ps=0 w=0.5 l=0.15
X66 pfd_8_0.UP_input.t18 charge_pump_cell_6_0.UP_b.t1 sky130_fd_pr__cap_mim_m3_1 l=16 w=13.9
X67 GNDA.t54 pfd_8_0.F.t6 pfd_8_0.QB.t0 GNDA.t53 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X68 GNDA.t105 GNDA.t103 GNDA.t105 GNDA.t104 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0 ps=0 w=2 l=0.6
X69 pfd_8_0.before_Reset.t1 pfd_8_0.QB.t4 VDDA.t24 VDDA.t23 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.805 ps=5 w=2 l=0.15
X70 GNDA.t67 a_6490_4630.t6 pfd_8_0.UP_input.t6 GNDA.t66 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X71 VDDA.t28 opamp_cell_4_0.n_right.t6 pfd_8_0.UP_input.t1 VDDA.t27 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X72 opamp_cell_4_0.VIN+.t3 pfd_8_0.UP_input.t19 VDDA.t55 VDDA.t54 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X73 pfd_8_0.UP_input.t9 pfd_8_0.UP_b.t2 pfd_8_0.UP_input.t8 VDDA.t7 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=0 ps=0 w=2 l=0.15
X74 a_490_1400.t1 pfd_8_0.QA_b.t5 pfd_8_0.QA.t0 VDDA.t58 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X75 V_OUT.t2 pfd_8_0.UP_input.t20 VDDA.t1 VDDA.t0 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X76 GNDA.t42 pfd_8_0.Reset.t2 pfd_8_0.E_b.t2 GNDA.t41 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X77 a_2530_190.t0 a_2350_1400.t2 GNDA.t61 GNDA.t60 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X78 VDDA.t82 opamp_cell_4_0.n_left.t2 opamp_cell_4_0.n_left.t3 VDDA.t81 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X79 a_6320_5840.t7 opamp_cell_4_0.VIN- opamp_cell_4_0.n_left.t5 GNDA.t130 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X80 GNDA.t7 I_IN.t2 I_IN.t3 GNDA.t6 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X81 pfd_8_0.E.t2 pfd_8_0.E_b.t4 a_870_1400.t1 VDDA.t19 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X82 pfd_8_0.UP_b.t1 pfd_8_0.UP.t4 VDDA.t129 VDDA.t12 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X83 a_5970_4630.t10 a_5970_4630.t8 a_5970_4630.t9 VDDA.t89 sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0 ps=0 w=1 l=0.15
X84 GNDA.t102 GNDA.t99 GNDA.t101 GNDA.t100 sky130_fd_pr__nfet_01v8 ad=0.25 pd=2 as=0 ps=0 w=0.5 l=0.15
X85 pfd_8_0.DOWN_input.t5 charge_pump_cell_6_0.DOWN.t0 sky130_fd_pr__cap_mim_m3_1 l=2.6 w=3.8
X86 VDDA.t60 a_1870_190.t2 pfd_8_0.Reset.t1 VDDA.t59 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=0.15
X87 pfd_8_0.UP_input.t5 a_6490_4630.t7 GNDA.t65 GNDA.t64 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X88 pfd_8_0.UP_input.t0 opamp_cell_4_0.n_right.t7 VDDA.t21 VDDA.t20 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X89 GNDA.t21 a_1870_190.t3 pfd_8_0.Reset.t0 GNDA.t20 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X90 VDDA.t108 VDDA.t105 VDDA.t107 VDDA.t106 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=0 ps=0 w=2 l=0.6
X91 opamp_cell_4_0.p_bias.t4 opamp_cell_4_0.p_bias.t3 VDDA.t78 VDDA.t77 sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X92 I_IN.t1 I_IN.t0 GNDA.t38 GNDA.t37 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X93 opamp_cell_4_0.p_bias.t0 a_6220_5810.t0 GNDA.t35 sky130_fd_pr__res_xhigh_po_5p73 l=1
X94 opamp_cell_4_0.n_left.t1 opamp_cell_4_0.n_left.t0 VDDA.t57 VDDA.t56 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X95 GNDA.t157 V_OUT.t7 sky130_fd_pr__cap_mim_m3_1 l=60 w=13.8
X96 opamp_cell_4_0.n_left.t4 opamp_cell_4_0.VIN- a_6320_5840.t8 GNDA.t129 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X97 a_5970_4630.t4 opamp_cell_4_0.p_bias.t11 VDDA.t64 VDDA.t63 sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X98 pfd_8_0.before_Reset.t0 pfd_8_0.QA.t5 a_1910_2020.t0 GNDA.t15 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X99 pfd_8_0.UP_PFD_b.t0 pfd_8_0.QA.t6 GNDA.t9 GNDA.t8 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X100 GNDA.t98 GNDA.t95 GNDA.t97 GNDA.t96 sky130_fd_pr__nfet_01v8 ad=1 pd=5 as=0 ps=0 w=2 l=0.6
X101 GNDA.t155 pfd_8_0.E.t4 pfd_8_0.QA.t2 GNDA.t154 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X102 a_9360_6440.t1 a_6490_4630.t2 GNDA.t34 sky130_fd_pr__res_xhigh_po_0p35 l=0.86
X103 pfd_8_0.F.t1 pfd_8_0.F_b.t3 a_870_640.t0 VDDA.t19 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X104 VDDA.t34 pfd_8_0.Reset.t3 a_1390_1400.t1 VDDA.t33 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X105 VDDA.t104 VDDA.t102 VDDA.t104 VDDA.t103 sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0 ps=0 w=2.5 l=0.5
X106 GNDA.t94 GNDA.t91 GNDA.t93 GNDA.t92 sky130_fd_pr__nfet_01v8 ad=1 pd=5 as=0 ps=0 w=2 l=0.6
X107 a_2530_190.t1 a_2350_1400.t3 VDDA.t42 VDDA.t41 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=0.15
X108 GNDA.t57 a_6220_5810.t3 a_6220_5810.t4 GNDA.t56 sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0.3125 ps=1.75 w=1.25 l=0.5
X109 GNDA.t63 a_6490_4630.t8 pfd_8_0.UP_input.t4 GNDA.t62 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X110 VDDA.t30 opamp_cell_4_0.n_right.t8 pfd_8_0.UP_input.t2 VDDA.t29 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X111 VDDA.t101 VDDA.t98 VDDA.t100 VDDA.t99 sky130_fd_pr__pfet_01v8 ad=1.25 pd=6 as=0 ps=0 w=2.5 l=0.5
X112 GNDA.t5 pfd_8_0.F_b.t4 pfd_8_0.F.t0 GNDA.t4 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X113 GNDA.t90 GNDA.t87 GNDA.t89 GNDA.t88 sky130_fd_pr__nfet_01v8 ad=1 pd=5 as=0 ps=0 w=2 l=0.6
X114 GNDA.t143 a_6220_5810.t11 a_6320_5840.t10 GNDA.t142 sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0.3125 ps=1.75 w=1.25 l=0.5
X115 pfd_8_0.QB_b.t1 pfd_8_0.QB.t5 a_n30_640.t1 VDDA.t4 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X116 GNDA.t82 a_6200_5250.t6 a_6490_4630.t4 GNDA.t81 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X117 a_5970_4630.t0 opamp_cell_4_0.VIN+.t7 a_6490_4630.t1 VDDA.t14 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X118 VDDA.t62 opamp_cell_4_0.p_bias.t12 a_5970_4630.t3 VDDA.t61 sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X119 VDDA.t127 pfd_8_0.Reset.t4 a_1390_640.t1 VDDA.t33 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X120 VDDA.t80 opamp_cell_4_0.p_bias.t1 opamp_cell_4_0.p_bias.t2 VDDA.t79 sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X121 pfd_8_0.UP_input.t3 pfd_8_0.UP.t5 VDDA.t38 VDDA.t37 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X122 opamp_cell_4_0.n_right.t2 charge_pump_cell_6_0.UP_b.t0 GNDA.t22 sky130_fd_pr__res_xhigh_po_0p35 l=1.14
X123 VDDA.t97 VDDA.t94 VDDA.t96 VDDA.t95 sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0 ps=0 w=1 l=0.15
X124 a_6320_5840.t6 a_6320_5840.t4 a_6320_5840.t5 GNDA.t141 sky130_fd_pr__nfet_01v8 ad=0.25 pd=2 as=0 ps=0 w=0.5 l=0.15
X125 GNDA.t3 pfd_8_0.QB.t6 pfd_8_0.QB_b.t2 GNDA.t2 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X126 a_6320_5840.t12 a_6220_5810.t12 GNDA.t151 GNDA.t150 sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0.3125 ps=1.75 w=1.25 l=0.5
X127 GNDA.t29 pfd_8_0.Reset.t5 pfd_8_0.F_b.t0 GNDA.t28 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X128 a_6320_5840.t3 a_6320_5840.t2 a_6320_5840.t3 GNDA.t23 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0 ps=0 w=0.5 l=0.15
X129 VDDA.t93 VDDA.t91 VDDA.t93 VDDA.t92 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0 ps=0 w=1 l=0.15
X130 a_6220_5810.t2 a_6220_5810.t1 GNDA.t59 GNDA.t58 sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0.3125 ps=1.75 w=1.25 l=0.5
X131 pfd_8_0.E.t0 pfd_8_0.QA_b.t6 GNDA.t11 GNDA.t10 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X132 VDDA.t45 pfd_8_0.QA.t7 pfd_8_0.before_Reset.t2 VDDA.t44 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X133 a_n30_640.t0 F_VCO.t0 VDDA.t18 VDDA.t5 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X134 pfd_8_0.UP_PFD_b.t1 pfd_8_0.QA.t8 VDDA.t15 VDDA.t2 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X135 a_6490_4630.t3 a_6200_5250.t7 GNDA.t80 GNDA.t79 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X136 a_6490_4630.t0 opamp_cell_4_0.VIN+.t8 a_5970_4630.t1 VDDA.t43 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X137 VDDA.t126 pfd_8_0.E.t5 a_490_1400.t0 VDDA.t35 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X138 VDDA.t32 a_2200_190.t2 a_1870_190.t1 VDDA.t31 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=0.15
X139 pfd_8_0.QA_b.t0 F_REF.t1 GNDA.t27 GNDA.t26 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X140 pfd_8_0.QB_b.t0 F_VCO.t1 GNDA.t52 GNDA.t51 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X141 a_490_640.t0 pfd_8_0.QB_b.t5 pfd_8_0.QB.t1 VDDA.t58 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X142 VDDA.t49 pfd_8_0.UP_input.t21 opamp_cell_4_0.VIN+.t2 VDDA.t48 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X143 GNDA.t75 a_2200_190.t3 a_1870_190.t0 GNDA.t74 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X144 a_6320_5840.t1 opamp_cell_4_0.VIN+.t9 opamp_cell_4_0.n_right.t0 GNDA.t14 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X145 VDDA.t51 opamp_cell_4_0.n_left.t7 opamp_cell_4_0.n_right.t3 VDDA.t50 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X146 pfd_8_0.QB.t2 pfd_8_0.QB_b.t6 GNDA.t149 GNDA.t148 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X147 pfd_8_0.DOWN_PFD_b.t0 pfd_8_0.QB.t7 VDDA.t3 VDDA.t2 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X148 pfd_8_0.UP.t0 pfd_8_0.UP_PFD_b.t3 GNDA.t78 GNDA.t77 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X149 pfd_8_0.DOWN_PFD_b.t2 pfd_8_0.QB.t8 GNDA.t132 GNDA.t131 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X150 pfd_8_0.E_b.t1 pfd_8_0.E.t6 GNDA.t46 GNDA.t45 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X151 opamp_cell_4_0.VIN+.t1 pfd_8_0.UP_input.t22 VDDA.t70 VDDA.t69 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X152 pfd_8_0.DOWN_b.t0 GNDA.t158 pfd_8_0.DOWN_PFD_b.t1 VDDA.t85 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
R0 a_6200_5250.n5 a_6200_5250.n4 427.647
R1 a_6200_5250.n1 a_6200_5250.t6 321.334
R2 a_6200_5250.n4 a_6200_5250.n0 210.601
R3 a_6200_5250.n2 a_6200_5250.n1 208.868
R4 a_6200_5250.n3 a_6200_5250.t0 174.056
R5 a_6200_5250.n4 a_6200_5250.n3 152
R6 a_6200_5250.n1 a_6200_5250.t7 112.468
R7 a_6200_5250.n2 a_6200_5250.t2 112.468
R8 a_6200_5250.n3 a_6200_5250.n2 61.5894
R9 a_6200_5250.n0 a_6200_5250.t3 60.0005
R10 a_6200_5250.n0 a_6200_5250.t1 60.0005
R11 a_6200_5250.n5 a_6200_5250.t5 49.2505
R12 a_6200_5250.t4 a_6200_5250.n5 49.2505
R13 GNDA.n396 GNDA.n395 348175
R14 GNDA.n395 GNDA.n394 292776
R15 GNDA.n269 GNDA.t76 25257.7
R16 GNDA.n275 GNDA.n269 15376.3
R17 GNDA.n394 GNDA.t12 2083.03
R18 GNDA.t18 GNDA.t4 1939.79
R19 GNDA.t148 GNDA.t2 1939.79
R20 GNDA.n213 GNDA.n24 1860.65
R21 GNDA.t55 GNDA.t131 1845.16
R22 GNDA.t47 GNDA.t73 1372.04
R23 GNDA.t20 GNDA.n399 1253.76
R24 GNDA.n402 GNDA.n23 1230.11
R25 GNDA.n259 GNDA.n258 1186
R26 GNDA.n212 GNDA.n211 1186
R27 GNDA.n205 GNDA.n204 1186
R28 GNDA.n266 GNDA.n265 1186
R29 GNDA.n268 GNDA.n267 1170
R30 GNDA.n393 GNDA.t73 1064.52
R31 GNDA.n356 GNDA.t55 1064.52
R32 GNDA.n394 GNDA.n26 1052.76
R33 GNDA.t16 GNDA.n401 922.582
R34 GNDA.t74 GNDA.n400 922.582
R35 GNDA.n106 GNDA.t26 783.001
R36 GNDA.t12 GNDA.n393 780.645
R37 GNDA.n356 GNDA.t47 780.645
R38 GNDA.t131 GNDA.n23 780.645
R39 GNDA.n328 GNDA.n327 669.307
R40 GNDA.n330 GNDA.n46 669.307
R41 GNDA.n323 GNDA.n322 669.307
R42 GNDA.n320 GNDA.n50 669.307
R43 GNDA.n274 GNDA.n273 669.307
R44 GNDA.n277 GNDA.n276 669.307
R45 GNDA.n402 GNDA.t16 638.711
R46 GNDA.n401 GNDA.t74 638.711
R47 GNDA.n400 GNDA.t20 638.711
R48 GNDA.n399 GNDA.t28 638.711
R49 GNDA.t49 GNDA.n398 638.711
R50 GNDA.n398 GNDA.t53 638.711
R51 GNDA.t51 GNDA.n396 638.711
R52 GNDA.t146 GNDA.t45 601.333
R53 GNDA.t30 GNDA.t0 601.333
R54 GNDA.t127 GNDA.t137 593.865
R55 GNDA.t137 GNDA.t135 593.865
R56 GNDA.t135 GNDA.t96 593.865
R57 GNDA.t133 GNDA.t110 593.865
R58 GNDA.t24 GNDA.t133 593.865
R59 GNDA.t92 GNDA.t24 593.865
R60 GNDA.t104 GNDA.t6 593.865
R61 GNDA.t6 GNDA.t37 593.865
R62 GNDA.t37 GNDA.t88 593.865
R63 GNDA.n105 GNDA.n104 585.003
R64 GNDA.n398 GNDA.n397 585.003
R65 GNDA.n102 GNDA.n101 585.001
R66 GNDA.n100 GNDA.n86 585.001
R67 GNDA.n99 GNDA.n83 585.001
R68 GNDA.n80 GNDA.n25 585.001
R69 GNDA.n257 GNDA.n256 585.001
R70 GNDA.n214 GNDA.n213 585.001
R71 GNDA.n175 GNDA.n174 585.001
R72 GNDA.n75 GNDA.n72 585.001
R73 GNDA.n77 GNDA.n76 585.001
R74 GNDA.n393 GNDA.n392 585.001
R75 GNDA.n357 GNDA.n356 585.001
R76 GNDA.n362 GNDA.n23 585.001
R77 GNDA.n403 GNDA.n402 585.001
R78 GNDA.n401 GNDA.n19 585.001
R79 GNDA.n400 GNDA.n16 585.001
R80 GNDA.n399 GNDA.n13 585.001
R81 GNDA.n396 GNDA.n2 585.001
R82 GNDA.n272 GNDA.n270 585
R83 GNDA.n68 GNDA.n66 585
R84 GNDA.n54 GNDA.n51 585
R85 GNDA.n57 GNDA.n56 585
R86 GNDA.n49 GNDA.n48 585
R87 GNDA.n332 GNDA.n331 585
R88 GNDA.n31 GNDA.n30 585
R89 GNDA.n30 GNDA.n26 585
R90 GNDA.n34 GNDA.n33 585
R91 GNDA.n36 GNDA.n28 585
R92 GNDA.n38 GNDA.n37 585
R93 GNDA.n37 GNDA.n26 585
R94 GNDA.n375 GNDA.t158 566.966
R95 GNDA.n275 GNDA.t127 566.871
R96 GNDA.n324 GNDA.t96 566.871
R97 GNDA.t110 GNDA.n324 566.871
R98 GNDA.n329 GNDA.t92 566.871
R99 GNDA.n329 GNDA.t104 566.871
R100 GNDA.t88 GNDA.n26 566.871
R101 GNDA.t34 GNDA.n266 564.696
R102 GNDA.n269 GNDA.t22 534.24
R103 GNDA.t28 GNDA.t18 520.431
R104 GNDA.t4 GNDA.t49 520.431
R105 GNDA.t53 GNDA.t148 520.431
R106 GNDA.t2 GNDA.t51 520.431
R107 GNDA.t22 GNDA.t34 509.197
R108 GNDA.t76 GNDA.t152 425.334
R109 GNDA.n76 GNDA.t60 418
R110 GNDA.n175 GNDA.t77 344.668
R111 GNDA.t8 GNDA.n75 344.668
R112 GNDA.n325 GNDA.t103 336.329
R113 GNDA.n325 GNDA.t91 336.329
R114 GNDA.n52 GNDA.t109 336.329
R115 GNDA.n52 GNDA.t95 336.329
R116 GNDA.n39 GNDA.t87 320.7
R117 GNDA.n278 GNDA.t126 320.7
R118 GNDA.n269 GNDA.n268 309.736
R119 GNDA.n176 GNDA.t106 304.634
R120 GNDA.n260 GNDA.t119 304.634
R121 GNDA.n210 GNDA.t99 304.634
R122 GNDA.n206 GNDA.t112 304.634
R123 GNDA.n255 GNDA.t123 292.584
R124 GNDA.n215 GNDA.t115 292.584
R125 GNDA.t71 GNDA.n25 286
R126 GNDA.t15 GNDA.n99 286
R127 GNDA.n275 GNDA.n274 250.349
R128 GNDA.n276 GNDA.n275 250.349
R129 GNDA.n324 GNDA.n323 250.349
R130 GNDA.n324 GNDA.n50 250.349
R131 GNDA.n329 GNDA.n328 250.349
R132 GNDA.n330 GNDA.n329 250.349
R133 GNDA.n35 GNDA.n26 250.349
R134 GNDA.n265 GNDA.t108 245
R135 GNDA.n259 GNDA.t122 245
R136 GNDA.n211 GNDA.t102 245
R137 GNDA.n205 GNDA.t114 245
R138 GNDA.t152 GNDA.n175 227.333
R139 GNDA.n75 GNDA.t77 227.333
R140 GNDA.n76 GNDA.t8 227.333
R141 GNDA.n102 GNDA.n100 205.333
R142 GNDA.n262 GNDA.n178 204.201
R143 GNDA.n208 GNDA.n202 204.201
R144 GNDA.n209 GNDA.n201 204.201
R145 GNDA.n207 GNDA.n203 204.201
R146 GNDA.n261 GNDA.n179 204.201
R147 GNDA.n264 GNDA.n263 204.201
R148 GNDA.n3 GNDA.t3 198.058
R149 GNDA.n444 GNDA.t149 198.058
R150 GNDA.n432 GNDA.t5 198.058
R151 GNDA.n11 GNDA.t19 198.058
R152 GNDA.n131 GNDA.t46 198.058
R153 GNDA.n126 GNDA.t147 198.058
R154 GNDA.n96 GNDA.t1 198.058
R155 GNDA.n112 GNDA.t31 198.058
R156 GNDA.n99 GNDA.t71 198
R157 GNDA.n100 GNDA.t32 198
R158 GNDA.t41 GNDA.n102 198
R159 GNDA.n105 GNDA.t10 198
R160 GNDA.t154 GNDA.n105 198
R161 GNDA.n331 GNDA.n49 197
R162 GNDA.n56 GNDA.n51 197
R163 GNDA.n270 GNDA.n68 197
R164 GNDA.n34 GNDA.n30 197
R165 GNDA.n37 GNDA.n36 197
R166 GNDA.n327 GNDA.n326 185
R167 GNDA.n326 GNDA.n46 185
R168 GNDA.n322 GNDA.n321 185
R169 GNDA.n321 GNDA.n320 185
R170 GNDA.n273 GNDA.n67 185
R171 GNDA.n277 GNDA.n67 185
R172 GNDA.n31 GNDA.n29 185
R173 GNDA.n38 GNDA.n29 185
R174 GNDA.n327 GNDA.n325 166.63
R175 GNDA.n322 GNDA.n52 166.63
R176 GNDA.t32 GNDA.t15 161.333
R177 GNDA.t45 GNDA.t41 161.333
R178 GNDA.t10 GNDA.t146 161.333
R179 GNDA.t0 GNDA.t154 161.333
R180 GNDA.t26 GNDA.t30 161.333
R181 GNDA.n256 GNDA.t125 134.501
R182 GNDA.n214 GNDA.t118 134.501
R183 GNDA.n7 GNDA.t54 130.713
R184 GNDA.n106 GNDA.t27 130.001
R185 GNDA.n101 GNDA.t42 130.001
R186 GNDA.n86 GNDA.t33 130.001
R187 GNDA.n83 GNDA.t72 130.001
R188 GNDA.n80 GNDA.t61 130.001
R189 GNDA.n2 GNDA.t52 130.001
R190 GNDA.n13 GNDA.t29 130.001
R191 GNDA.n16 GNDA.t21 130.001
R192 GNDA.n19 GNDA.t75 130.001
R193 GNDA.n403 GNDA.t17 130.001
R194 GNDA.n103 GNDA.t11 130.001
R195 GNDA.n95 GNDA.t155 130.001
R196 GNDA.n8 GNDA.t50 130.001
R197 GNDA.n77 GNDA.t9 122.501
R198 GNDA.n72 GNDA.t78 122.501
R199 GNDA.n174 GNDA.t153 122.501
R200 GNDA.n362 GNDA.t132 122.501
R201 GNDA.n357 GNDA.t48 122.501
R202 GNDA.n392 GNDA.t13 122.501
R203 GNDA.n257 GNDA.t23 112.157
R204 GNDA.n183 GNDA.n182 97.8707
R205 GNDA.n187 GNDA.n186 97.8707
R206 GNDA.n191 GNDA.n190 97.8707
R207 GNDA.n195 GNDA.n194 97.8707
R208 GNDA.n200 GNDA.n199 97.8707
R209 GNDA.n204 GNDA.t39 97.7783
R210 GNDA.n266 GNDA.t107 94.9025
R211 GNDA.n258 GNDA.t120 94.9025
R212 GNDA.n287 GNDA.n62 92.2612
R213 GNDA.n280 GNDA.n65 92.2612
R214 GNDA.n314 GNDA.n293 92.2612
R215 GNDA.n308 GNDA.n296 92.2612
R216 GNDA.n336 GNDA.n335 92.2612
R217 GNDA.n343 GNDA.n342 92.2612
R218 GNDA.n326 GNDA.n47 91.3721
R219 GNDA.n334 GNDA.n45 91.3721
R220 GNDA.n334 GNDA.n333 91.3721
R221 GNDA.n321 GNDA.n55 91.3721
R222 GNDA.n292 GNDA.n53 91.3721
R223 GNDA.n292 GNDA.n58 91.3721
R224 GNDA.n271 GNDA.n67 90.7567
R225 GNDA.n32 GNDA.n29 90.7567
R226 GNDA.t39 GNDA.t141 89.1508
R227 GNDA.n212 GNDA.t116 86.275
R228 GNDA.n274 GNDA.n270 84.306
R229 GNDA.n276 GNDA.n68 84.306
R230 GNDA.n323 GNDA.n51 84.306
R231 GNDA.n56 GNDA.n50 84.306
R232 GNDA.n328 GNDA.n49 84.306
R233 GNDA.n331 GNDA.n330 84.306
R234 GNDA.n35 GNDA.n34 84.306
R235 GNDA.n36 GNDA.n35 84.306
R236 GNDA.n267 GNDA.t157 84.2543
R237 GNDA.n208 GNDA.n207 83.2005
R238 GNDA.n209 GNDA.n208 83.2005
R239 GNDA.n267 GNDA.t156 81.0543
R240 GNDA.n395 GNDA.n24 80.6672
R241 GNDA.t43 GNDA.t113 77.6476
R242 GNDA.t66 GNDA.t107 74.7717
R243 GNDA.t64 GNDA.t66 74.7717
R244 GNDA.t62 GNDA.t64 74.7717
R245 GNDA.t68 GNDA.t62 74.7717
R246 GNDA.t120 GNDA.t68 74.7717
R247 GNDA.n258 GNDA.n257 74.7717
R248 GNDA.t130 GNDA.t70 74.7717
R249 GNDA.t81 GNDA.t79 74.7717
R250 GNDA.t83 GNDA.t100 74.7717
R251 GNDA.n395 GNDA.n25 73.3338
R252 GNDA.t14 GNDA.t124 71.8959
R253 GNDA.t144 GNDA.t85 71.8959
R254 GNDA.n263 GNDA.n262 66.5605
R255 GNDA.n262 GNDA.n261 66.5605
R256 GNDA.t129 GNDA.t139 66.1443
R257 GNDA.n262 GNDA.n177 65.9634
R258 GNDA.n107 GNDA.n106 60.29
R259 GNDA.n101 GNDA.n89 60.29
R260 GNDA.n139 GNDA.n86 60.29
R261 GNDA.n146 GNDA.n83 60.29
R262 GNDA.n152 GNDA.n80 60.29
R263 GNDA.n404 GNDA.n403 60.29
R264 GNDA.n411 GNDA.n19 60.29
R265 GNDA.n417 GNDA.n16 60.29
R266 GNDA.n424 GNDA.n13 60.29
R267 GNDA.n452 GNDA.n2 60.29
R268 GNDA.n178 GNDA.t65 60.0005
R269 GNDA.n178 GNDA.t63 60.0005
R270 GNDA.n202 GNDA.t80 60.0005
R271 GNDA.n202 GNDA.t86 60.0005
R272 GNDA.n201 GNDA.t84 60.0005
R273 GNDA.n201 GNDA.t101 60.0005
R274 GNDA.t114 GNDA.n203 60.0005
R275 GNDA.n203 GNDA.t82 60.0005
R276 GNDA.n179 GNDA.t69 60.0005
R277 GNDA.n179 GNDA.t121 60.0005
R278 GNDA.t108 GNDA.n264 60.0005
R279 GNDA.n264 GNDA.t67 60.0005
R280 GNDA.n160 GNDA.n77 59.5478
R281 GNDA.n167 GNDA.n72 59.5478
R282 GNDA.n174 GNDA.n173 59.5478
R283 GNDA.n380 GNDA.n357 58.9809
R284 GNDA.n363 GNDA.n362 58.9809
R285 GNDA.n392 GNDA.n391 58.9809
R286 GNDA.n268 GNDA.t36 56.0165
R287 GNDA.n120 GNDA.n95 54.4005
R288 GNDA.n103 GNDA.n94 54.4005
R289 GNDA.n437 GNDA.n8 54.4005
R290 GNDA.n439 GNDA.n7 54.4005
R291 GNDA.t56 GNDA.t129 48.8894
R292 GNDA.t60 GNDA.n24 44.0005
R293 GNDA.t142 GNDA.t14 43.1378
R294 GNDA.t85 GNDA.t150 43.1378
R295 GNDA.n208 GNDA.n197 41.6005
R296 GNDA.n349 GNDA.n348 41.3005
R297 GNDA.n252 GNDA.n177 39.4985
R298 GNDA.t113 GNDA.t58 37.3861
R299 GNDA.t58 GNDA.t81 37.3861
R300 GNDA.n107 GNDA.n0 33.0991
R301 GNDA.n453 GNDA.n452 33.0991
R302 GNDA.n288 GNDA.n287 32.0005
R303 GNDA.n288 GNDA.n59 32.0005
R304 GNDA.n282 GNDA.n281 32.0005
R305 GNDA.n282 GNDA.n63 32.0005
R306 GNDA.n286 GNDA.n63 32.0005
R307 GNDA.n315 GNDA.n60 32.0005
R308 GNDA.n313 GNDA.n294 32.0005
R309 GNDA.n309 GNDA.n294 32.0005
R310 GNDA.n309 GNDA.n308 32.0005
R311 GNDA.n307 GNDA.n297 32.0005
R312 GNDA.n303 GNDA.n297 32.0005
R313 GNDA.n302 GNDA.n301 32.0005
R314 GNDA.n301 GNDA.n44 32.0005
R315 GNDA.n337 GNDA.n42 32.0005
R316 GNDA.n341 GNDA.n42 32.0005
R317 GNDA.n344 GNDA.n40 32.0005
R318 GNDA.n173 GNDA.n172 32.0005
R319 GNDA.n172 GNDA.n70 32.0005
R320 GNDA.n168 GNDA.n70 32.0005
R321 GNDA.n166 GNDA.n165 32.0005
R322 GNDA.n165 GNDA.n73 32.0005
R323 GNDA.n161 GNDA.n73 32.0005
R324 GNDA.n159 GNDA.n158 32.0005
R325 GNDA.n158 GNDA.n78 32.0005
R326 GNDA.n154 GNDA.n78 32.0005
R327 GNDA.n154 GNDA.n153 32.0005
R328 GNDA.n151 GNDA.n81 32.0005
R329 GNDA.n147 GNDA.n81 32.0005
R330 GNDA.n145 GNDA.n144 32.0005
R331 GNDA.n144 GNDA.n84 32.0005
R332 GNDA.n140 GNDA.n84 32.0005
R333 GNDA.n138 GNDA.n137 32.0005
R334 GNDA.n137 GNDA.n87 32.0005
R335 GNDA.n133 GNDA.n132 32.0005
R336 GNDA.n132 GNDA.n131 32.0005
R337 GNDA.n131 GNDA.n90 32.0005
R338 GNDA.n127 GNDA.n90 32.0005
R339 GNDA.n127 GNDA.n126 32.0005
R340 GNDA.n126 GNDA.n125 32.0005
R341 GNDA.n125 GNDA.n92 32.0005
R342 GNDA.n119 GNDA.n118 32.0005
R343 GNDA.n118 GNDA.n96 32.0005
R344 GNDA.n114 GNDA.n96 32.0005
R345 GNDA.n114 GNDA.n113 32.0005
R346 GNDA.n113 GNDA.n112 32.0005
R347 GNDA.n112 GNDA.n98 32.0005
R348 GNDA.n108 GNDA.n98 32.0005
R349 GNDA.n252 GNDA.n251 32.0005
R350 GNDA.n251 GNDA.n250 32.0005
R351 GNDA.n250 GNDA.n181 32.0005
R352 GNDA.n246 GNDA.n181 32.0005
R353 GNDA.n246 GNDA.n245 32.0005
R354 GNDA.n245 GNDA.n244 32.0005
R355 GNDA.n244 GNDA.n185 32.0005
R356 GNDA.n240 GNDA.n185 32.0005
R357 GNDA.n240 GNDA.n239 32.0005
R358 GNDA.n239 GNDA.n238 32.0005
R359 GNDA.n238 GNDA.n189 32.0005
R360 GNDA.n234 GNDA.n189 32.0005
R361 GNDA.n234 GNDA.n233 32.0005
R362 GNDA.n233 GNDA.n232 32.0005
R363 GNDA.n232 GNDA.n193 32.0005
R364 GNDA.n228 GNDA.n227 32.0005
R365 GNDA.n227 GNDA.n226 32.0005
R366 GNDA.n226 GNDA.n198 32.0005
R367 GNDA.n221 GNDA.n198 32.0005
R368 GNDA.n221 GNDA.n220 32.0005
R369 GNDA.n220 GNDA.n219 32.0005
R370 GNDA.n390 GNDA.n352 32.0005
R371 GNDA.n386 GNDA.n352 32.0005
R372 GNDA.n386 GNDA.n385 32.0005
R373 GNDA.n385 GNDA.n384 32.0005
R374 GNDA.n384 GNDA.n354 32.0005
R375 GNDA.n380 GNDA.n354 32.0005
R376 GNDA.n380 GNDA.n379 32.0005
R377 GNDA.n379 GNDA.n378 32.0005
R378 GNDA.n378 GNDA.n358 32.0005
R379 GNDA.n373 GNDA.n358 32.0005
R380 GNDA.n373 GNDA.n372 32.0005
R381 GNDA.n372 GNDA.n371 32.0005
R382 GNDA.n371 GNDA.n360 32.0005
R383 GNDA.n367 GNDA.n366 32.0005
R384 GNDA.n366 GNDA.n365 32.0005
R385 GNDA.n365 GNDA.n22 32.0005
R386 GNDA.n405 GNDA.n22 32.0005
R387 GNDA.n409 GNDA.n20 32.0005
R388 GNDA.n410 GNDA.n409 32.0005
R389 GNDA.n412 GNDA.n17 32.0005
R390 GNDA.n416 GNDA.n17 32.0005
R391 GNDA.n419 GNDA.n418 32.0005
R392 GNDA.n419 GNDA.n14 32.0005
R393 GNDA.n423 GNDA.n14 32.0005
R394 GNDA.n426 GNDA.n425 32.0005
R395 GNDA.n426 GNDA.n11 32.0005
R396 GNDA.n430 GNDA.n11 32.0005
R397 GNDA.n431 GNDA.n430 32.0005
R398 GNDA.n432 GNDA.n431 32.0005
R399 GNDA.n432 GNDA.n9 32.0005
R400 GNDA.n436 GNDA.n9 32.0005
R401 GNDA.n440 GNDA.n5 32.0005
R402 GNDA.n444 GNDA.n5 32.0005
R403 GNDA.n445 GNDA.n444 32.0005
R404 GNDA.n446 GNDA.n445 32.0005
R405 GNDA.n446 GNDA.n3 32.0005
R406 GNDA.n450 GNDA.n3 32.0005
R407 GNDA.n451 GNDA.n450 32.0005
R408 GNDA.t70 GNDA.t142 31.6345
R409 GNDA.n302 GNDA.n46 29.0291
R410 GNDA.n320 GNDA.n319 29.0291
R411 GNDA.n168 GNDA.n167 28.8005
R412 GNDA.n152 GNDA.n151 28.8005
R413 GNDA.n213 GNDA.n212 28.7587
R414 GNDA.n260 GNDA.n259 27.2005
R415 GNDA.n265 GNDA.n176 27.2005
R416 GNDA.t141 GNDA.t56 25.8829
R417 GNDA.n319 GNDA.n60 25.6005
R418 GNDA.n337 GNDA.n336 25.6005
R419 GNDA.n343 GNDA.n341 25.6005
R420 GNDA.n161 GNDA.n160 25.6005
R421 GNDA.n140 GNDA.n139 25.6005
R422 GNDA.n89 GNDA.n87 25.6005
R423 GNDA.n121 GNDA.n94 25.6005
R424 GNDA.n121 GNDA.n120 25.6005
R425 GNDA.n211 GNDA.n210 25.6005
R426 GNDA.n206 GNDA.n205 25.6005
R427 GNDA.n228 GNDA.n197 25.6005
R428 GNDA.n219 GNDA 25.6005
R429 GNDA.n391 GNDA.n390 25.6005
R430 GNDA.n363 GNDA.n360 25.6005
R431 GNDA.n404 GNDA.n20 25.6005
R432 GNDA.n417 GNDA.n416 25.6005
R433 GNDA.n424 GNDA.n423 25.6005
R434 GNDA.n438 GNDA.n437 25.6005
R435 GNDA.n256 GNDA.n255 24.8279
R436 GNDA.n215 GNDA.n214 24.8279
R437 GNDA.n182 GNDA.t125 24.0005
R438 GNDA.n182 GNDA.t143 24.0005
R439 GNDA.n186 GNDA.t140 24.0005
R440 GNDA.n186 GNDA.t57 24.0005
R441 GNDA.n190 GNDA.t40 24.0005
R442 GNDA.n190 GNDA.t44 24.0005
R443 GNDA.n194 GNDA.t59 24.0005
R444 GNDA.n194 GNDA.t145 24.0005
R445 GNDA.n199 GNDA.t151 24.0005
R446 GNDA.n199 GNDA.t117 24.0005
R447 GNDA.n439 GNDA.n438 22.4005
R448 GNDA.n279 GNDA.n278 20.9665
R449 GNDA.n315 GNDA.n314 19.2005
R450 GNDA.n314 GNDA.n313 19.2005
R451 GNDA.n146 GNDA.n145 19.2005
R452 GNDA.t35 GNDA.t83 17.8306
R453 GNDA.n204 GNDA.t43 17.2554
R454 GNDA.n411 GNDA.n410 16.0005
R455 GNDA.n412 GNDA.n411 16.0005
R456 GNDA.n217 GNDA 15.7005
R457 GNDA.n278 GNDA.n277 15.6449
R458 GNDA.n39 GNDA.n38 15.6449
R459 GNDA.n62 GNDA.t136 15.0005
R460 GNDA.n62 GNDA.t97 15.0005
R461 GNDA.t128 GNDA.n65 15.0005
R462 GNDA.n65 GNDA.t138 15.0005
R463 GNDA.n293 GNDA.t111 15.0005
R464 GNDA.n293 GNDA.t134 15.0005
R465 GNDA.n296 GNDA.t25 15.0005
R466 GNDA.n296 GNDA.t93 15.0005
R467 GNDA.n335 GNDA.t105 15.0005
R468 GNDA.n335 GNDA.t7 15.0005
R469 GNDA.n342 GNDA.t38 15.0005
R470 GNDA.n342 GNDA.t89 15.0005
R471 GNDA.t105 GNDA.n334 15.0005
R472 GNDA.n326 GNDA.t94 15.0005
R473 GNDA.t111 GNDA.n292 15.0005
R474 GNDA.n321 GNDA.t98 15.0005
R475 GNDA.n67 GNDA.t128 15.0005
R476 GNDA.n29 GNDA.t90 15.0005
R477 GNDA.n40 GNDA.n39 14.4005
R478 GNDA.n261 GNDA.n260 14.0805
R479 GNDA.n263 GNDA.n176 14.0805
R480 GNDA.n391 GNDA.n351 13.9181
R481 GNDA.t150 GNDA.t35 13.8044
R482 GNDA.n217 GNDA.n27 13.1958
R483 GNDA.n69 GNDA.n27 12.8163
R484 GNDA.n319 GNDA.n59 12.8005
R485 GNDA.n281 GNDA.n280 12.8005
R486 GNDA.n336 GNDA.n44 12.8005
R487 GNDA.n344 GNDA.n343 12.8005
R488 GNDA.n147 GNDA.n146 12.8005
R489 GNDA.n210 GNDA.n209 12.8005
R490 GNDA.n207 GNDA.n206 12.8005
R491 GNDA GNDA.n0 12.7806
R492 GNDA GNDA.n453 11.8829
R493 GNDA.n351 GNDA.n350 11.8528
R494 GNDA.n350 GNDA.n349 11.6542
R495 GNDA.n440 GNDA.n439 9.6005
R496 GNDA.n255 GNDA.n254 9.58175
R497 GNDA.n223 GNDA.n215 9.58175
R498 GNDA.n122 GNDA.n121 9.3005
R499 GNDA.n109 GNDA.n108 9.3005
R500 GNDA.n110 GNDA.n98 9.3005
R501 GNDA.n112 GNDA.n111 9.3005
R502 GNDA.n113 GNDA.n97 9.3005
R503 GNDA.n115 GNDA.n114 9.3005
R504 GNDA.n116 GNDA.n96 9.3005
R505 GNDA.n118 GNDA.n117 9.3005
R506 GNDA.n119 GNDA.n93 9.3005
R507 GNDA.n123 GNDA.n92 9.3005
R508 GNDA.n125 GNDA.n124 9.3005
R509 GNDA.n126 GNDA.n91 9.3005
R510 GNDA.n128 GNDA.n127 9.3005
R511 GNDA.n129 GNDA.n90 9.3005
R512 GNDA.n131 GNDA.n130 9.3005
R513 GNDA.n132 GNDA.n88 9.3005
R514 GNDA.n134 GNDA.n133 9.3005
R515 GNDA.n135 GNDA.n87 9.3005
R516 GNDA.n137 GNDA.n136 9.3005
R517 GNDA.n138 GNDA.n85 9.3005
R518 GNDA.n141 GNDA.n140 9.3005
R519 GNDA.n142 GNDA.n84 9.3005
R520 GNDA.n144 GNDA.n143 9.3005
R521 GNDA.n145 GNDA.n82 9.3005
R522 GNDA.n148 GNDA.n147 9.3005
R523 GNDA.n149 GNDA.n81 9.3005
R524 GNDA.n151 GNDA.n150 9.3005
R525 GNDA.n153 GNDA.n79 9.3005
R526 GNDA.n155 GNDA.n154 9.3005
R527 GNDA.n156 GNDA.n78 9.3005
R528 GNDA.n158 GNDA.n157 9.3005
R529 GNDA.n159 GNDA.n74 9.3005
R530 GNDA.n162 GNDA.n161 9.3005
R531 GNDA.n163 GNDA.n73 9.3005
R532 GNDA.n165 GNDA.n164 9.3005
R533 GNDA.n166 GNDA.n71 9.3005
R534 GNDA.n169 GNDA.n168 9.3005
R535 GNDA.n170 GNDA.n70 9.3005
R536 GNDA.n172 GNDA.n171 9.3005
R537 GNDA.n253 GNDA.n252 9.3005
R538 GNDA.n251 GNDA.n180 9.3005
R539 GNDA.n250 GNDA.n249 9.3005
R540 GNDA.n248 GNDA.n181 9.3005
R541 GNDA.n247 GNDA.n246 9.3005
R542 GNDA.n245 GNDA.n184 9.3005
R543 GNDA.n244 GNDA.n243 9.3005
R544 GNDA.n242 GNDA.n185 9.3005
R545 GNDA.n241 GNDA.n240 9.3005
R546 GNDA.n239 GNDA.n188 9.3005
R547 GNDA.n238 GNDA.n237 9.3005
R548 GNDA.n236 GNDA.n189 9.3005
R549 GNDA.n235 GNDA.n234 9.3005
R550 GNDA.n233 GNDA.n192 9.3005
R551 GNDA.n232 GNDA.n231 9.3005
R552 GNDA.n230 GNDA.n193 9.3005
R553 GNDA.n229 GNDA.n228 9.3005
R554 GNDA.n227 GNDA.n196 9.3005
R555 GNDA.n226 GNDA.n225 9.3005
R556 GNDA.n224 GNDA.n198 9.3005
R557 GNDA.n222 GNDA.n221 9.3005
R558 GNDA.n220 GNDA.n216 9.3005
R559 GNDA.n219 GNDA.n218 9.3005
R560 GNDA.n348 GNDA.n347 9.3005
R561 GNDA.n346 GNDA.n40 9.3005
R562 GNDA.n345 GNDA.n344 9.3005
R563 GNDA.n343 GNDA.n41 9.3005
R564 GNDA.n341 GNDA.n340 9.3005
R565 GNDA.n339 GNDA.n42 9.3005
R566 GNDA.n338 GNDA.n337 9.3005
R567 GNDA.n336 GNDA.n43 9.3005
R568 GNDA.n299 GNDA.n44 9.3005
R569 GNDA.n301 GNDA.n300 9.3005
R570 GNDA.n302 GNDA.n298 9.3005
R571 GNDA.n281 GNDA.n64 9.3005
R572 GNDA.n283 GNDA.n282 9.3005
R573 GNDA.n284 GNDA.n63 9.3005
R574 GNDA.n286 GNDA.n285 9.3005
R575 GNDA.n287 GNDA.n61 9.3005
R576 GNDA.n289 GNDA.n288 9.3005
R577 GNDA.n290 GNDA.n59 9.3005
R578 GNDA.n319 GNDA.n318 9.3005
R579 GNDA.n317 GNDA.n60 9.3005
R580 GNDA.n316 GNDA.n315 9.3005
R581 GNDA.n314 GNDA.n291 9.3005
R582 GNDA.n313 GNDA.n312 9.3005
R583 GNDA.n311 GNDA.n294 9.3005
R584 GNDA.n310 GNDA.n309 9.3005
R585 GNDA.n308 GNDA.n295 9.3005
R586 GNDA.n307 GNDA.n306 9.3005
R587 GNDA.n305 GNDA.n297 9.3005
R588 GNDA.n304 GNDA.n303 9.3005
R589 GNDA.n390 GNDA.n389 9.3005
R590 GNDA.n388 GNDA.n352 9.3005
R591 GNDA.n387 GNDA.n386 9.3005
R592 GNDA.n385 GNDA.n353 9.3005
R593 GNDA.n384 GNDA.n383 9.3005
R594 GNDA.n382 GNDA.n354 9.3005
R595 GNDA.n381 GNDA.n380 9.3005
R596 GNDA.n379 GNDA.n355 9.3005
R597 GNDA.n378 GNDA.n377 9.3005
R598 GNDA.n376 GNDA.n358 9.3005
R599 GNDA.n374 GNDA.n373 9.3005
R600 GNDA.n372 GNDA.n359 9.3005
R601 GNDA.n371 GNDA.n370 9.3005
R602 GNDA.n369 GNDA.n360 9.3005
R603 GNDA.n368 GNDA.n367 9.3005
R604 GNDA.n366 GNDA.n361 9.3005
R605 GNDA.n365 GNDA.n364 9.3005
R606 GNDA.n22 GNDA.n21 9.3005
R607 GNDA.n406 GNDA.n405 9.3005
R608 GNDA.n407 GNDA.n20 9.3005
R609 GNDA.n409 GNDA.n408 9.3005
R610 GNDA.n410 GNDA.n18 9.3005
R611 GNDA.n413 GNDA.n412 9.3005
R612 GNDA.n414 GNDA.n17 9.3005
R613 GNDA.n416 GNDA.n415 9.3005
R614 GNDA.n418 GNDA.n15 9.3005
R615 GNDA.n420 GNDA.n419 9.3005
R616 GNDA.n421 GNDA.n14 9.3005
R617 GNDA.n423 GNDA.n422 9.3005
R618 GNDA.n425 GNDA.n12 9.3005
R619 GNDA.n427 GNDA.n426 9.3005
R620 GNDA.n428 GNDA.n11 9.3005
R621 GNDA.n430 GNDA.n429 9.3005
R622 GNDA.n431 GNDA.n10 9.3005
R623 GNDA.n433 GNDA.n432 9.3005
R624 GNDA.n434 GNDA.n9 9.3005
R625 GNDA.n436 GNDA.n435 9.3005
R626 GNDA.n438 GNDA.n6 9.3005
R627 GNDA.n441 GNDA.n440 9.3005
R628 GNDA.n442 GNDA.n5 9.3005
R629 GNDA.n444 GNDA.n443 9.3005
R630 GNDA.n445 GNDA.n4 9.3005
R631 GNDA.n447 GNDA.n446 9.3005
R632 GNDA.n448 GNDA.n3 9.3005
R633 GNDA.n450 GNDA.n449 9.3005
R634 GNDA.n451 GNDA.n1 9.3005
R635 GNDA.t139 GNDA.t130 8.62795
R636 GNDA.t100 GNDA.t116 8.62795
R637 GNDA.n173 GNDA.n69 7.49888
R638 GNDA.n273 GNDA.n272 7.11161
R639 GNDA.n277 GNDA.n66 7.11161
R640 GNDA.n33 GNDA.n31 7.11161
R641 GNDA.n38 GNDA.n28 7.11161
R642 GNDA.n280 GNDA.n279 6.69883
R643 GNDA.n287 GNDA.n286 6.4005
R644 GNDA.n308 GNDA.n307 6.4005
R645 GNDA.n303 GNDA.n302 6.4005
R646 GNDA.n160 GNDA.n159 6.4005
R647 GNDA.n139 GNDA.n138 6.4005
R648 GNDA.n133 GNDA.n89 6.4005
R649 GNDA.n94 GNDA.n92 6.4005
R650 GNDA.n120 GNDA.n119 6.4005
R651 GNDA.n108 GNDA.n107 6.4005
R652 GNDA.n197 GNDA.n193 6.4005
R653 GNDA.n367 GNDA.n363 6.4005
R654 GNDA.n405 GNDA.n404 6.4005
R655 GNDA.n418 GNDA.n417 6.4005
R656 GNDA.n425 GNDA.n424 6.4005
R657 GNDA.n437 GNDA.n436 6.4005
R658 GNDA.n452 GNDA.n451 6.4005
R659 GNDA.n348 GNDA.n40 6.4005
R660 GNDA.n104 GNDA.n103 5.68939
R661 GNDA.n104 GNDA.n95 5.68939
R662 GNDA.n397 GNDA.n8 5.68939
R663 GNDA.n397 GNDA.n7 4.97828
R664 GNDA.n272 GNDA.n271 3.48951
R665 GNDA.n271 GNDA.n66 3.48951
R666 GNDA.n33 GNDA.n32 3.48951
R667 GNDA.n32 GNDA.n28 3.48951
R668 GNDA.n167 GNDA.n166 3.2005
R669 GNDA.n153 GNDA.n152 3.2005
R670 GNDA.t124 GNDA.t23 2.87632
R671 GNDA.t79 GNDA.t144 2.87632
R672 GNDA.n48 GNDA.n45 2.25882
R673 GNDA.n48 GNDA.n47 2.25882
R674 GNDA.n333 GNDA.n46 2.25882
R675 GNDA.n332 GNDA.n47 2.25882
R676 GNDA.n327 GNDA.n45 2.25882
R677 GNDA.n333 GNDA.n332 2.25882
R678 GNDA.n54 GNDA.n53 2.25882
R679 GNDA.n55 GNDA.n54 2.25882
R680 GNDA.n320 GNDA.n58 2.25882
R681 GNDA.n57 GNDA.n55 2.25882
R682 GNDA.n322 GNDA.n53 2.25882
R683 GNDA.n58 GNDA.n57 2.25882
R684 GNDA.n350 GNDA.n27 0.9875
R685 GNDA.n279 GNDA.n64 0.703977
R686 GNDA.n171 GNDA.n69 0.193977
R687 GNDA.n109 GNDA.n0 0.193881
R688 GNDA.n453 GNDA.n1 0.193881
R689 GNDA.n389 GNDA.n351 0.193695
R690 GNDA.n218 GNDA.n217 0.188
R691 GNDA.n171 GNDA.n170 0.15675
R692 GNDA.n170 GNDA.n169 0.15675
R693 GNDA.n169 GNDA.n71 0.15675
R694 GNDA.n164 GNDA.n71 0.15675
R695 GNDA.n164 GNDA.n163 0.15675
R696 GNDA.n163 GNDA.n162 0.15675
R697 GNDA.n162 GNDA.n74 0.15675
R698 GNDA.n157 GNDA.n74 0.15675
R699 GNDA.n157 GNDA.n156 0.15675
R700 GNDA.n156 GNDA.n155 0.15675
R701 GNDA.n155 GNDA.n79 0.15675
R702 GNDA.n150 GNDA.n79 0.15675
R703 GNDA.n150 GNDA.n149 0.15675
R704 GNDA.n149 GNDA.n148 0.15675
R705 GNDA.n148 GNDA.n82 0.15675
R706 GNDA.n143 GNDA.n82 0.15675
R707 GNDA.n143 GNDA.n142 0.15675
R708 GNDA.n142 GNDA.n141 0.15675
R709 GNDA.n141 GNDA.n85 0.15675
R710 GNDA.n136 GNDA.n85 0.15675
R711 GNDA.n136 GNDA.n135 0.15675
R712 GNDA.n135 GNDA.n134 0.15675
R713 GNDA.n134 GNDA.n88 0.15675
R714 GNDA.n130 GNDA.n88 0.15675
R715 GNDA.n130 GNDA.n129 0.15675
R716 GNDA.n129 GNDA.n128 0.15675
R717 GNDA.n128 GNDA.n91 0.15675
R718 GNDA.n124 GNDA.n91 0.15675
R719 GNDA.n124 GNDA.n123 0.15675
R720 GNDA.n123 GNDA.n122 0.15675
R721 GNDA.n122 GNDA.n93 0.15675
R722 GNDA.n117 GNDA.n93 0.15675
R723 GNDA.n117 GNDA.n116 0.15675
R724 GNDA.n116 GNDA.n115 0.15675
R725 GNDA.n115 GNDA.n97 0.15675
R726 GNDA.n111 GNDA.n97 0.15675
R727 GNDA.n111 GNDA.n110 0.15675
R728 GNDA.n110 GNDA.n109 0.15675
R729 GNDA.n253 GNDA.n180 0.15675
R730 GNDA.n249 GNDA.n248 0.15675
R731 GNDA.n248 GNDA.n247 0.15675
R732 GNDA.n247 GNDA.n184 0.15675
R733 GNDA.n243 GNDA.n242 0.15675
R734 GNDA.n242 GNDA.n241 0.15675
R735 GNDA.n241 GNDA.n188 0.15675
R736 GNDA.n237 GNDA.n236 0.15675
R737 GNDA.n236 GNDA.n235 0.15675
R738 GNDA.n235 GNDA.n192 0.15675
R739 GNDA.n231 GNDA.n230 0.15675
R740 GNDA.n230 GNDA.n229 0.15675
R741 GNDA.n229 GNDA.n196 0.15675
R742 GNDA.n225 GNDA.n224 0.15675
R743 GNDA.n222 GNDA.n216 0.15675
R744 GNDA.n218 GNDA.n216 0.15675
R745 GNDA.n283 GNDA.n64 0.15675
R746 GNDA.n284 GNDA.n283 0.15675
R747 GNDA.n285 GNDA.n284 0.15675
R748 GNDA.n285 GNDA.n61 0.15675
R749 GNDA.n289 GNDA.n61 0.15675
R750 GNDA.n290 GNDA.n289 0.15675
R751 GNDA.n318 GNDA.n290 0.15675
R752 GNDA.n318 GNDA.n317 0.15675
R753 GNDA.n317 GNDA.n316 0.15675
R754 GNDA.n316 GNDA.n291 0.15675
R755 GNDA.n312 GNDA.n291 0.15675
R756 GNDA.n312 GNDA.n311 0.15675
R757 GNDA.n311 GNDA.n310 0.15675
R758 GNDA.n310 GNDA.n295 0.15675
R759 GNDA.n306 GNDA.n295 0.15675
R760 GNDA.n306 GNDA.n305 0.15675
R761 GNDA.n305 GNDA.n304 0.15675
R762 GNDA.n304 GNDA.n298 0.15675
R763 GNDA.n300 GNDA.n298 0.15675
R764 GNDA.n300 GNDA.n299 0.15675
R765 GNDA.n299 GNDA.n43 0.15675
R766 GNDA.n338 GNDA.n43 0.15675
R767 GNDA.n339 GNDA.n338 0.15675
R768 GNDA.n340 GNDA.n339 0.15675
R769 GNDA.n340 GNDA.n41 0.15675
R770 GNDA.n345 GNDA.n41 0.15675
R771 GNDA.n346 GNDA.n345 0.15675
R772 GNDA.n347 GNDA.n346 0.15675
R773 GNDA.n389 GNDA.n388 0.15675
R774 GNDA.n388 GNDA.n387 0.15675
R775 GNDA.n387 GNDA.n353 0.15675
R776 GNDA.n383 GNDA.n353 0.15675
R777 GNDA.n383 GNDA.n382 0.15675
R778 GNDA.n382 GNDA.n381 0.15675
R779 GNDA.n381 GNDA.n355 0.15675
R780 GNDA.n377 GNDA.n355 0.15675
R781 GNDA.n377 GNDA.n376 0.15675
R782 GNDA.n374 GNDA.n359 0.15675
R783 GNDA.n370 GNDA.n359 0.15675
R784 GNDA.n370 GNDA.n369 0.15675
R785 GNDA.n369 GNDA.n368 0.15675
R786 GNDA.n368 GNDA.n361 0.15675
R787 GNDA.n364 GNDA.n361 0.15675
R788 GNDA.n364 GNDA.n21 0.15675
R789 GNDA.n406 GNDA.n21 0.15675
R790 GNDA.n407 GNDA.n406 0.15675
R791 GNDA.n408 GNDA.n407 0.15675
R792 GNDA.n408 GNDA.n18 0.15675
R793 GNDA.n413 GNDA.n18 0.15675
R794 GNDA.n414 GNDA.n413 0.15675
R795 GNDA.n415 GNDA.n414 0.15675
R796 GNDA.n415 GNDA.n15 0.15675
R797 GNDA.n420 GNDA.n15 0.15675
R798 GNDA.n421 GNDA.n420 0.15675
R799 GNDA.n422 GNDA.n421 0.15675
R800 GNDA.n422 GNDA.n12 0.15675
R801 GNDA.n427 GNDA.n12 0.15675
R802 GNDA.n428 GNDA.n427 0.15675
R803 GNDA.n429 GNDA.n428 0.15675
R804 GNDA.n429 GNDA.n10 0.15675
R805 GNDA.n433 GNDA.n10 0.15675
R806 GNDA.n434 GNDA.n433 0.15675
R807 GNDA.n435 GNDA.n434 0.15675
R808 GNDA.n435 GNDA.n6 0.15675
R809 GNDA.n441 GNDA.n6 0.15675
R810 GNDA.n442 GNDA.n441 0.15675
R811 GNDA.n443 GNDA.n442 0.15675
R812 GNDA.n443 GNDA.n4 0.15675
R813 GNDA.n447 GNDA.n4 0.15675
R814 GNDA.n448 GNDA.n447 0.15675
R815 GNDA.n449 GNDA.n448 0.15675
R816 GNDA.n449 GNDA.n1 0.15675
R817 GNDA.n254 GNDA.n177 0.131895
R818 GNDA.n347 GNDA 0.1255
R819 GNDA.n376 GNDA.n375 0.109875
R820 GNDA.n183 GNDA.n180 0.09425
R821 GNDA.n187 GNDA.n184 0.09425
R822 GNDA.n191 GNDA.n188 0.09425
R823 GNDA.n195 GNDA.n192 0.09425
R824 GNDA.n200 GNDA.n196 0.09425
R825 GNDA.n224 GNDA.n223 0.09425
R826 GNDA.n254 GNDA.n253 0.063
R827 GNDA.n249 GNDA.n183 0.063
R828 GNDA.n243 GNDA.n187 0.063
R829 GNDA.n237 GNDA.n191 0.063
R830 GNDA.n231 GNDA.n195 0.063
R831 GNDA.n225 GNDA.n200 0.063
R832 GNDA.n223 GNDA.n222 0.063
R833 GNDA.n349 GNDA 0.063
R834 GNDA.n375 GNDA.n374 0.047375
R835 a_5970_4630.n8 a_5970_4630.n6 522.322
R836 a_5970_4630.n3 a_5970_4630.t8 384.967
R837 a_5970_4630.n0 a_5970_4630.t11 384.967
R838 a_5970_4630.n3 a_5970_4630.t10 379.166
R839 a_5970_4630.t12 a_5970_4630.n0 376.56
R840 a_5970_4630.n5 a_5970_4630.n1 315.647
R841 a_5970_4630.n4 a_5970_4630.n2 315.647
R842 a_5970_4630.n11 a_5970_4630.n10 314.502
R843 a_5970_4630.n8 a_5970_4630.n7 160.721
R844 a_5970_4630.n5 a_5970_4630.n4 83.2005
R845 a_5970_4630.n1 a_5970_4630.t1 49.2505
R846 a_5970_4630.n1 a_5970_4630.t7 49.2505
R847 a_5970_4630.n2 a_5970_4630.t6 49.2505
R848 a_5970_4630.n2 a_5970_4630.t9 49.2505
R849 a_5970_4630.t12 a_5970_4630.n11 49.2505
R850 a_5970_4630.n11 a_5970_4630.t0 49.2505
R851 a_5970_4630.n10 a_5970_4630.n9 42.6672
R852 a_5970_4630.n9 a_5970_4630.n8 37.763
R853 a_5970_4630.n9 a_5970_4630.n5 23.4672
R854 a_5970_4630.n6 a_5970_4630.t2 19.7005
R855 a_5970_4630.n6 a_5970_4630.t4 19.7005
R856 a_5970_4630.n7 a_5970_4630.t3 19.7005
R857 a_5970_4630.n7 a_5970_4630.t5 19.7005
R858 a_5970_4630.n4 a_5970_4630.n3 16.0005
R859 a_5970_4630.n10 a_5970_4630.n0 16.0005
R860 VDDA.n468 VDDA.n460 831.25
R861 VDDA.n463 VDDA.n462 831.25
R862 VDDA.n457 VDDA.n449 831.25
R863 VDDA.n452 VDDA.n451 831.25
R864 VDDA.n461 VDDA.n460 585
R865 VDDA.n465 VDDA.n463 585
R866 VDDA.n361 VDDA.n355 585
R867 VDDA.n356 VDDA.n355 585
R868 VDDA.n367 VDDA.n44 585
R869 VDDA.n371 VDDA.n44 585
R870 VDDA.n312 VDDA.n50 585
R871 VDDA.n307 VDDA.n50 585
R872 VDDA.n288 VDDA.n283 585
R873 VDDA.n292 VDDA.n283 585
R874 VDDA.n450 VDDA.n449 585
R875 VDDA.n454 VDDA.n452 585
R876 VDDA.n352 VDDA.n346 585
R877 VDDA.n347 VDDA.n346 585
R878 VDDA.n58 VDDA.n51 585
R879 VDDA.n53 VDDA.n51 585
R880 VDDA.n123 VDDA.n116 585
R881 VDDA.n105 VDDA.n97 585
R882 VDDA.n271 VDDA.n175 585
R883 VDDA.n264 VDDA.n175 585
R884 VDDA.n261 VDDA.n260 585
R885 VDDA.n260 VDDA.n259 585
R886 VDDA.n230 VDDA.n229 585
R887 VDDA.n230 VDDA.n219 585
R888 VDDA.n467 VDDA.t128 465.079
R889 VDDA.t128 VDDA.n466 465.079
R890 VDDA.n456 VDDA.t40 465.079
R891 VDDA.t40 VDDA.n455 465.079
R892 VDDA.t17 VDDA.n336 464.281
R893 VDDA.n338 VDDA.t17 464.281
R894 VDDA.n444 VDDA.t6 464.281
R895 VDDA.t6 VDDA.n443 464.281
R896 VDDA.n481 VDDA.t34 464.281
R897 VDDA.t34 VDDA.n480 464.281
R898 VDDA.n425 VDDA.t24 464.281
R899 VDDA.t24 VDDA.n424 464.281
R900 VDDA.n403 VDDA.t66 464.281
R901 VDDA.t66 VDDA.n402 464.281
R902 VDDA.n333 VDDA.t42 464.281
R903 VDDA.t42 VDDA.n332 464.281
R904 VDDA.t18 VDDA.n433 464.281
R905 VDDA.n434 VDDA.t18 464.281
R906 VDDA.t127 VDDA.n17 464.281
R907 VDDA.n471 VDDA.t127 464.281
R908 VDDA.t60 VDDA.n25 464.281
R909 VDDA.n406 VDDA.t60 464.281
R910 VDDA.t32 VDDA.n321 464.281
R911 VDDA.n322 VDDA.t32 464.281
R912 VDDA.n41 VDDA.t130 415.336
R913 VDDA.n86 VDDA.t109 384.967
R914 VDDA.n128 VDDA.t115 384.967
R915 VDDA.n91 VDDA.t94 384.967
R916 VDDA.n111 VDDA.t91 384.967
R917 VDDA.n123 VDDA.t102 374.878
R918 VDDA.t113 VDDA.t8 360.346
R919 VDDA.t8 VDDA.t0 360.346
R920 VDDA.t0 VDDA.t10 360.346
R921 VDDA.t10 VDDA.t71 360.346
R922 VDDA.t71 VDDA.t106 360.346
R923 VDDA.t48 VDDA.t120 360.346
R924 VDDA.t69 VDDA.t48 360.346
R925 VDDA.t25 VDDA.t69 360.346
R926 VDDA.t54 VDDA.t25 360.346
R927 VDDA.t123 VDDA.t54 360.346
R928 VDDA.n96 VDDA.t98 352.834
R929 VDDA.n225 VDDA.t113 343.966
R930 VDDA.n263 VDDA.t106 343.966
R931 VDDA.t120 VDDA.n263 343.966
R932 VDDA.n269 VDDA.t123 343.966
R933 VDDA.n112 VDDA.t93 341.752
R934 VDDA.n127 VDDA.t118 341.752
R935 VDDA.n87 VDDA.t111 341.752
R936 VDDA.n92 VDDA.t97 341.752
R937 VDDA.n258 VDDA.t119 336.329
R938 VDDA.n258 VDDA.t105 336.329
R939 VDDA.n220 VDDA.t112 320.7
R940 VDDA.n272 VDDA.t122 320.7
R941 VDDA.n85 VDDA.n83 315.647
R942 VDDA.n79 VDDA.n78 315.647
R943 VDDA.n110 VDDA.n109 315.647
R944 VDDA.n90 VDDA.n89 315.647
R945 VDDA.n130 VDDA.n82 315.647
R946 VDDA.n129 VDDA.n84 315.647
R947 VDDA.n24 VDDA.t45 315.25
R948 VDDA.t22 VDDA.t19 314.113
R949 VDDA.t58 VDDA.t4 314.113
R950 VDDA.t110 VDDA.n87 304.659
R951 VDDA.n260 VDDA.n183 291.363
R952 VDDA.n256 VDDA.n181 291.363
R953 VDDA.n257 VDDA.n256 291.363
R954 VDDA.n359 VDDA.n355 290.733
R955 VDDA.n365 VDDA.n44 290.733
R956 VDDA.n310 VDDA.n50 290.733
R957 VDDA.n286 VDDA.n283 290.733
R958 VDDA.n350 VDDA.n346 290.733
R959 VDDA.n52 VDDA.n51 290.733
R960 VDDA.n121 VDDA.n116 290.733
R961 VDDA.n117 VDDA.n116 290.733
R962 VDDA.n103 VDDA.n97 290.733
R963 VDDA.n98 VDDA.n97 290.733
R964 VDDA.n265 VDDA.n175 290.733
R965 VDDA.n230 VDDA.n218 290.733
R966 VDDA.n445 VDDA.n444 243.698
R967 VDDA.n482 VDDA.n481 243.698
R968 VDDA.n426 VDDA.n425 243.698
R969 VDDA.n404 VDDA.n403 243.698
R970 VDDA.n334 VDDA.n333 243.698
R971 VDDA.n434 VDDA.n431 243.698
R972 VDDA.n475 VDDA.n471 243.698
R973 VDDA.n410 VDDA.n406 243.698
R974 VDDA.n322 VDDA.n319 243.698
R975 VDDA.n430 VDDA.n1 238.367
R976 VDDA.n469 VDDA.n468 238.367
R977 VDDA.n462 VDDA.n429 238.367
R978 VDDA.n428 VDDA.n16 238.367
R979 VDDA.n421 VDDA.n19 238.367
R980 VDDA.n399 VDDA.n27 238.367
R981 VDDA.n318 VDDA.n35 238.367
R982 VDDA.n438 VDDA.n2 238.367
R983 VDDA.n458 VDDA.n457 238.367
R984 VDDA.n485 VDDA.n484 238.367
R985 VDDA.n413 VDDA.n412 238.367
R986 VDDA.n326 VDDA.n31 238.367
R987 VDDA.n451 VDDA.n447 238.367
R988 VDDA.n117 VDDA.n88 233.841
R989 VDDA.n98 VDDA.n94 233.841
R990 VDDA.n362 VDDA.n361 230.308
R991 VDDA.n356 VDDA.n315 230.308
R992 VDDA.n368 VDDA.n367 230.308
R993 VDDA.n371 VDDA.n370 230.308
R994 VDDA.n313 VDDA.n312 230.308
R995 VDDA.n307 VDDA.n46 230.308
R996 VDDA.n289 VDDA.n288 230.308
R997 VDDA.n292 VDDA.n291 230.308
R998 VDDA.n353 VDDA.n352 230.308
R999 VDDA.n58 VDDA.n48 230.308
R1000 VDDA.n53 VDDA.n47 230.308
R1001 VDDA.n347 VDDA.n344 230.308
R1002 VDDA.n124 VDDA.n123 230.308
R1003 VDDA.n271 VDDA.n270 230.308
R1004 VDDA.n268 VDDA.n264 230.308
R1005 VDDA.n262 VDDA.n261 230.308
R1006 VDDA.n259 VDDA.n178 230.308
R1007 VDDA.t7 VDDA.t12 222.178
R1008 VDDA.n363 VDDA.n343 199.195
R1009 VDDA.n192 VDDA.n191 196.502
R1010 VDDA.n189 VDDA.n188 196.502
R1011 VDDA.n255 VDDA.n254 196.502
R1012 VDDA.n246 VDDA.n211 196.502
R1013 VDDA.n239 VDDA.n214 196.502
R1014 VDDA.n232 VDDA.n231 196.502
R1015 VDDA.n338 VDDA.n317 190.333
R1016 VDDA.n127 VDDA.n126 185.001
R1017 VDDA.n113 VDDA.n112 185.001
R1018 VDDA.n108 VDDA.n92 185.001
R1019 VDDA.n57 VDDA.n56 185
R1020 VDDA.n55 VDDA.n54 185
R1021 VDDA.n351 VDDA.n345 185
R1022 VDDA.n349 VDDA.n348 185
R1023 VDDA.n325 VDDA.n324 185
R1024 VDDA.n323 VDDA.n320 185
R1025 VDDA.n407 VDDA.n26 185
R1026 VDDA.n409 VDDA.n408 185
R1027 VDDA.n472 VDDA.n18 185
R1028 VDDA.n474 VDDA.n473 185
R1029 VDDA.n450 VDDA.n448 185
R1030 VDDA.n454 VDDA.n453 185
R1031 VDDA.n437 VDDA.n436 185
R1032 VDDA.n435 VDDA.n432 185
R1033 VDDA.n287 VDDA.n285 185
R1034 VDDA.n284 VDDA.n282 185
R1035 VDDA.n311 VDDA.n49 185
R1036 VDDA.n309 VDDA.n308 185
R1037 VDDA.n366 VDDA.n364 185
R1038 VDDA.n45 VDDA.n43 185
R1039 VDDA.n360 VDDA.n354 185
R1040 VDDA.n358 VDDA.n357 185
R1041 VDDA.n329 VDDA.n328 185
R1042 VDDA.n331 VDDA.n330 185
R1043 VDDA.n29 VDDA.n28 185
R1044 VDDA.n401 VDDA.n400 185
R1045 VDDA.n21 VDDA.n20 185
R1046 VDDA.n423 VDDA.n422 185
R1047 VDDA.n477 VDDA.n476 185
R1048 VDDA.n479 VDDA.n478 185
R1049 VDDA.n461 VDDA.n459 185
R1050 VDDA.n465 VDDA.n464 185
R1051 VDDA.n440 VDDA.n439 185
R1052 VDDA.n442 VDDA.n441 185
R1053 VDDA.n342 VDDA.n34 185
R1054 VDDA.n343 VDDA.n342 185
R1055 VDDA.n341 VDDA.n340 185
R1056 VDDA.n339 VDDA.n337 185
R1057 VDDA.n343 VDDA.n317 185
R1058 VDDA.n122 VDDA.n115 185
R1059 VDDA.n120 VDDA.n114 185
R1060 VDDA.n125 VDDA.n114 185
R1061 VDDA.n119 VDDA.n118 185
R1062 VDDA.n106 VDDA.n105 185
R1063 VDDA.n107 VDDA.n106 185
R1064 VDDA.n104 VDDA.n95 185
R1065 VDDA.n102 VDDA.n101 185
R1066 VDDA.n100 VDDA.n99 185
R1067 VDDA.n182 VDDA.n179 185
R1068 VDDA.n185 VDDA.n184 185
R1069 VDDA.n177 VDDA.n176 185
R1070 VDDA.n267 VDDA.n266 185
R1071 VDDA.n229 VDDA.n221 185
R1072 VDDA.n225 VDDA.n221 185
R1073 VDDA.n228 VDDA.n227 185
R1074 VDDA.n223 VDDA.n222 185
R1075 VDDA.n224 VDDA.n219 185
R1076 VDDA.n225 VDDA.n224 185
R1077 VDDA.n290 VDDA.t7 172.38
R1078 VDDA.t85 VDDA.n314 172.38
R1079 VDDA.n369 VDDA.t2 172.38
R1080 VDDA.n259 VDDA.n258 166.63
R1081 VDDA.n441 VDDA.n439 150
R1082 VDDA.n464 VDDA.n459 150
R1083 VDDA.n478 VDDA.n476 150
R1084 VDDA.n422 VDDA.n20 150
R1085 VDDA.n400 VDDA.n28 150
R1086 VDDA.n330 VDDA.n328 150
R1087 VDDA.n437 VDDA.n432 150
R1088 VDDA.n453 VDDA.n448 150
R1089 VDDA.n474 VDDA.n18 150
R1090 VDDA.n409 VDDA.n26 150
R1091 VDDA.n325 VDDA.n320 150
R1092 VDDA.n342 VDDA.n341 150
R1093 VDDA.n337 VDDA.n317 150
R1094 VDDA.t79 VDDA.t75 145.038
R1095 VDDA.n335 VDDA.n327 137.904
R1096 VDDA.n411 VDDA.n405 137.904
R1097 VDDA.n290 VDDA.t37 126.412
R1098 VDDA.n314 VDDA.t12 126.412
R1099 VDDA.n369 VDDA.t85 126.412
R1100 VDDA.t2 VDDA.n363 126.412
R1101 VDDA.t126 VDDA.n460 123.126
R1102 VDDA.n463 VDDA.t126 123.126
R1103 VDDA.t36 VDDA.n449 123.126
R1104 VDDA.n452 VDDA.t36 123.126
R1105 VDDA.n357 VDDA.n354 120.001
R1106 VDDA.n364 VDDA.n45 120.001
R1107 VDDA.n308 VDDA.n49 120.001
R1108 VDDA.n285 VDDA.n284 120.001
R1109 VDDA.n348 VDDA.n345 120.001
R1110 VDDA.n56 VDDA.n55 120.001
R1111 VDDA.n115 VDDA.n114 120.001
R1112 VDDA.n118 VDDA.n114 120.001
R1113 VDDA.n106 VDDA.n95 120.001
R1114 VDDA.n101 VDDA.n100 120.001
R1115 VDDA.n267 VDDA.n177 120.001
R1116 VDDA.n184 VDDA.n179 120.001
R1117 VDDA.n227 VDDA.n221 120.001
R1118 VDDA.n224 VDDA.n223 120.001
R1119 VDDA.n161 VDDA.n67 119.737
R1120 VDDA.n154 VDDA.n70 119.737
R1121 VDDA.n147 VDDA.n73 119.737
R1122 VDDA.n140 VDDA.n76 119.737
R1123 VDDA.n132 VDDA.n81 119.737
R1124 VDDA.n126 VDDA.t116 119.656
R1125 VDDA.n125 VDDA.n113 108.779
R1126 VDDA.n483 VDDA.n427 107.258
R1127 VDDA.n483 VDDA.t33 103.427
R1128 VDDA.t39 VDDA.n470 103.427
R1129 VDDA.n470 VDDA.t35 103.427
R1130 VDDA.t5 VDDA.n446 103.427
R1131 VDDA.n427 VDDA.t59 95.7666
R1132 VDDA.t27 VDDA.t110 94.2753
R1133 VDDA.t20 VDDA.t27 94.2753
R1134 VDDA.t29 VDDA.t20 94.2753
R1135 VDDA.t83 VDDA.t29 94.2753
R1136 VDDA.t116 VDDA.t83 94.2753
R1137 VDDA.t50 VDDA.t52 94.2753
R1138 VDDA.t56 VDDA.t95 94.2753
R1139 VDDA.t77 VDDA.n108 94.2753
R1140 VDDA.t90 VDDA.t14 94.2753
R1141 VDDA.t88 VDDA.t87 94.2753
R1142 VDDA.t41 VDDA.t16 91.936
R1143 VDDA.t65 VDDA.t31 91.936
R1144 VDDA.t44 VDDA.t23 84.2747
R1145 VDDA.t33 VDDA.t22 84.2747
R1146 VDDA.t19 VDDA.t39 84.2747
R1147 VDDA.t35 VDDA.t58 84.2747
R1148 VDDA.t4 VDDA.t5 84.2747
R1149 VDDA.t103 VDDA.t92 83.3974
R1150 VDDA.t61 VDDA.t43 83.3974
R1151 VDDA.n110 VDDA.n79 83.2005
R1152 VDDA.n90 VDDA.n79 83.2005
R1153 VDDA.n130 VDDA.n83 83.2005
R1154 VDDA.n130 VDDA.n129 83.2005
R1155 VDDA.t63 VDDA.t81 76.1455
R1156 VDDA.t99 VDDA.t89 76.1455
R1157 VDDA.n314 VDDA.n48 69.8479
R1158 VDDA.n314 VDDA.n47 69.8479
R1159 VDDA.n363 VDDA.n353 69.8479
R1160 VDDA.n363 VDDA.n344 69.8479
R1161 VDDA.n290 VDDA.n289 69.8479
R1162 VDDA.n291 VDDA.n290 69.8479
R1163 VDDA.n314 VDDA.n313 69.8479
R1164 VDDA.n314 VDDA.n46 69.8479
R1165 VDDA.n369 VDDA.n368 69.8479
R1166 VDDA.n370 VDDA.n369 69.8479
R1167 VDDA.n363 VDDA.n362 69.8479
R1168 VDDA.n363 VDDA.n315 69.8479
R1169 VDDA.n125 VDDA.n124 69.8479
R1170 VDDA.n125 VDDA.n88 69.8479
R1171 VDDA.n107 VDDA.n93 69.8479
R1172 VDDA.n107 VDDA.n94 69.8479
R1173 VDDA.n263 VDDA.n262 69.8479
R1174 VDDA.n263 VDDA.n178 69.8479
R1175 VDDA.n270 VDDA.n269 69.8479
R1176 VDDA.n269 VDDA.n268 69.8479
R1177 VDDA.n226 VDDA.n225 69.8479
R1178 VDDA.n131 VDDA.n130 69.3203
R1179 VDDA.t81 VDDA.t73 68.8936
R1180 VDDA.t89 VDDA.n107 68.8936
R1181 VDDA.n327 VDDA.n326 65.8183
R1182 VDDA.n327 VDDA.n319 65.8183
R1183 VDDA.n412 VDDA.n411 65.8183
R1184 VDDA.n411 VDDA.n410 65.8183
R1185 VDDA.n484 VDDA.n483 65.8183
R1186 VDDA.n483 VDDA.n475 65.8183
R1187 VDDA.n470 VDDA.n458 65.8183
R1188 VDDA.n470 VDDA.n447 65.8183
R1189 VDDA.n446 VDDA.n438 65.8183
R1190 VDDA.n446 VDDA.n431 65.8183
R1191 VDDA.n335 VDDA.n334 65.8183
R1192 VDDA.n335 VDDA.n318 65.8183
R1193 VDDA.n405 VDDA.n404 65.8183
R1194 VDDA.n405 VDDA.n27 65.8183
R1195 VDDA.n427 VDDA.n426 65.8183
R1196 VDDA.n427 VDDA.n19 65.8183
R1197 VDDA.n483 VDDA.n482 65.8183
R1198 VDDA.n483 VDDA.n428 65.8183
R1199 VDDA.n470 VDDA.n469 65.8183
R1200 VDDA.n470 VDDA.n429 65.8183
R1201 VDDA.n446 VDDA.n445 65.8183
R1202 VDDA.n446 VDDA.n430 65.8183
R1203 VDDA.n343 VDDA.n316 65.8183
R1204 VDDA.t92 VDDA.t46 61.6417
R1205 VDDA.t43 VDDA.t67 61.6417
R1206 VDDA.n516 VDDA.n1 58.0576
R1207 VDDA.n486 VDDA.n16 58.0576
R1208 VDDA.n421 VDDA.n420 58.0576
R1209 VDDA.n399 VDDA.n398 58.0576
R1210 VDDA.n389 VDDA.n35 58.0576
R1211 VDDA.n516 VDDA.n2 58.0576
R1212 VDDA.n486 VDDA.n485 58.0576
R1213 VDDA.n414 VDDA.n413 58.0576
R1214 VDDA.n397 VDDA.n31 58.0576
R1215 VDDA.n390 VDDA.n34 58.0576
R1216 VDDA.n356 VDDA.n38 57.2449
R1217 VDDA.n372 VDDA.n371 57.2449
R1218 VDDA.n307 VDDA.n306 57.2449
R1219 VDDA.n293 VDDA.n292 57.2449
R1220 VDDA.n352 VDDA.n38 57.2449
R1221 VDDA.n306 VDDA.n58 57.2449
R1222 VDDA.n503 VDDA.n7 54.4005
R1223 VDDA.n9 VDDA.n7 54.4005
R1224 VDDA.n9 VDDA.n8 54.4005
R1225 VDDA.n503 VDDA.n8 54.4005
R1226 VDDA.n432 VDDA.n431 53.3664
R1227 VDDA.n453 VDDA.n447 53.3664
R1228 VDDA.n475 VDDA.n474 53.3664
R1229 VDDA.n326 VDDA.n325 53.3664
R1230 VDDA.n320 VDDA.n319 53.3664
R1231 VDDA.n412 VDDA.n26 53.3664
R1232 VDDA.n410 VDDA.n409 53.3664
R1233 VDDA.n484 VDDA.n18 53.3664
R1234 VDDA.n458 VDDA.n448 53.3664
R1235 VDDA.n438 VDDA.n437 53.3664
R1236 VDDA.n334 VDDA.n328 53.3664
R1237 VDDA.n330 VDDA.n318 53.3664
R1238 VDDA.n404 VDDA.n28 53.3664
R1239 VDDA.n400 VDDA.n27 53.3664
R1240 VDDA.n426 VDDA.n20 53.3664
R1241 VDDA.n422 VDDA.n19 53.3664
R1242 VDDA.n482 VDDA.n476 53.3664
R1243 VDDA.n478 VDDA.n428 53.3664
R1244 VDDA.n469 VDDA.n459 53.3664
R1245 VDDA.n464 VDDA.n429 53.3664
R1246 VDDA.n445 VDDA.n439 53.3664
R1247 VDDA.n441 VDDA.n430 53.3664
R1248 VDDA.n341 VDDA.n316 53.3664
R1249 VDDA.n337 VDDA.n316 53.3664
R1250 VDDA.n108 VDDA.t79 50.7639
R1251 VDDA.t111 VDDA.n85 49.2505
R1252 VDDA.n85 VDDA.t28 49.2505
R1253 VDDA.n78 VDDA.t53 49.2505
R1254 VDDA.n78 VDDA.t82 49.2505
R1255 VDDA.n109 VDDA.t93 49.2505
R1256 VDDA.n109 VDDA.t51 49.2505
R1257 VDDA.n89 VDDA.t57 49.2505
R1258 VDDA.n89 VDDA.t96 49.2505
R1259 VDDA.n82 VDDA.t21 49.2505
R1260 VDDA.n82 VDDA.t30 49.2505
R1261 VDDA.n84 VDDA.t84 49.2505
R1262 VDDA.n84 VDDA.t117 49.2505
R1263 VDDA VDDA.n517 47.763
R1264 VDDA.n348 VDDA.n344 45.3071
R1265 VDDA.n55 VDDA.n47 45.3071
R1266 VDDA.n56 VDDA.n48 45.3071
R1267 VDDA.n353 VDDA.n345 45.3071
R1268 VDDA.n289 VDDA.n285 45.3071
R1269 VDDA.n291 VDDA.n284 45.3071
R1270 VDDA.n313 VDDA.n49 45.3071
R1271 VDDA.n308 VDDA.n46 45.3071
R1272 VDDA.n368 VDDA.n364 45.3071
R1273 VDDA.n370 VDDA.n45 45.3071
R1274 VDDA.n362 VDDA.n354 45.3071
R1275 VDDA.n357 VDDA.n315 45.3071
R1276 VDDA.n118 VDDA.n88 45.3071
R1277 VDDA.n124 VDDA.n115 45.3071
R1278 VDDA.n95 VDDA.n93 45.3071
R1279 VDDA.n100 VDDA.n94 45.3071
R1280 VDDA.n101 VDDA.n93 45.3071
R1281 VDDA.n262 VDDA.n179 45.3071
R1282 VDDA.n184 VDDA.n178 45.3071
R1283 VDDA.n270 VDDA.n177 45.3071
R1284 VDDA.n268 VDDA.n267 45.3071
R1285 VDDA.n227 VDDA.n226 45.3071
R1286 VDDA.n226 VDDA.n223 45.3071
R1287 VDDA.n137 VDDA.n79 41.6005
R1288 VDDA.t75 VDDA.t90 39.886
R1289 VDDA.n131 VDDA.n80 39.4988
R1290 VDDA.n279 VDDA.n278 38.1005
R1291 VDDA.n113 VDDA.t103 36.26
R1292 VDDA.t46 VDDA.t50 32.6341
R1293 VDDA.t67 VDDA.t88 32.6341
R1294 VDDA.n261 VDDA.n180 32.2291
R1295 VDDA.n294 VDDA.n62 32.0005
R1296 VDDA.n298 VDDA.n62 32.0005
R1297 VDDA.n299 VDDA.n298 32.0005
R1298 VDDA.n300 VDDA.n299 32.0005
R1299 VDDA.n300 VDDA.n59 32.0005
R1300 VDDA.n306 VDDA.n59 32.0005
R1301 VDDA.n306 VDDA.n60 32.0005
R1302 VDDA.n60 VDDA.n42 32.0005
R1303 VDDA.n373 VDDA.n42 32.0005
R1304 VDDA.n377 VDDA.n40 32.0005
R1305 VDDA.n378 VDDA.n377 32.0005
R1306 VDDA.n379 VDDA.n378 32.0005
R1307 VDDA.n383 VDDA.n382 32.0005
R1308 VDDA.n384 VDDA.n383 32.0005
R1309 VDDA.n384 VDDA.n36 32.0005
R1310 VDDA.n388 VDDA.n36 32.0005
R1311 VDDA.n392 VDDA.n391 32.0005
R1312 VDDA.n392 VDDA.n30 32.0005
R1313 VDDA.n396 VDDA.n32 32.0005
R1314 VDDA.n419 VDDA.n22 32.0005
R1315 VDDA.n487 VDDA.n15 32.0005
R1316 VDDA.n491 VDDA.n13 32.0005
R1317 VDDA.n492 VDDA.n491 32.0005
R1318 VDDA.n493 VDDA.n492 32.0005
R1319 VDDA.n493 VDDA.n11 32.0005
R1320 VDDA.n497 VDDA.n11 32.0005
R1321 VDDA.n498 VDDA.n497 32.0005
R1322 VDDA.n499 VDDA.n498 32.0005
R1323 VDDA.n505 VDDA.n504 32.0005
R1324 VDDA.n505 VDDA.n5 32.0005
R1325 VDDA.n509 VDDA.n5 32.0005
R1326 VDDA.n510 VDDA.n509 32.0005
R1327 VDDA.n511 VDDA.n510 32.0005
R1328 VDDA.n511 VDDA.n3 32.0005
R1329 VDDA.n515 VDDA.n3 32.0005
R1330 VDDA.n135 VDDA.n80 32.0005
R1331 VDDA.n136 VDDA.n135 32.0005
R1332 VDDA.n138 VDDA.n75 32.0005
R1333 VDDA.n143 VDDA.n75 32.0005
R1334 VDDA.n144 VDDA.n143 32.0005
R1335 VDDA.n145 VDDA.n144 32.0005
R1336 VDDA.n145 VDDA.n72 32.0005
R1337 VDDA.n150 VDDA.n72 32.0005
R1338 VDDA.n151 VDDA.n150 32.0005
R1339 VDDA.n152 VDDA.n151 32.0005
R1340 VDDA.n152 VDDA.n69 32.0005
R1341 VDDA.n157 VDDA.n69 32.0005
R1342 VDDA.n158 VDDA.n157 32.0005
R1343 VDDA.n159 VDDA.n158 32.0005
R1344 VDDA.n159 VDDA.n66 32.0005
R1345 VDDA.n164 VDDA.n66 32.0005
R1346 VDDA.n165 VDDA.n164 32.0005
R1347 VDDA.n165 VDDA.n64 32.0005
R1348 VDDA.n169 VDDA.n64 32.0005
R1349 VDDA.n170 VDDA.n169 32.0005
R1350 VDDA.n274 VDDA.n172 32.0005
R1351 VDDA.n278 VDDA.n172 32.0005
R1352 VDDA.n198 VDDA.n197 32.0005
R1353 VDDA.n197 VDDA.n196 32.0005
R1354 VDDA.n204 VDDA.n186 32.0005
R1355 VDDA.n204 VDDA.n203 32.0005
R1356 VDDA.n203 VDDA.n202 32.0005
R1357 VDDA.n253 VDDA.n208 32.0005
R1358 VDDA.n248 VDDA.n247 32.0005
R1359 VDDA.n241 VDDA.n240 32.0005
R1360 VDDA.n241 VDDA.n212 32.0005
R1361 VDDA.n245 VDDA.n212 32.0005
R1362 VDDA.n234 VDDA.n233 32.0005
R1363 VDDA.n234 VDDA.n215 32.0005
R1364 VDDA.n238 VDDA.n215 32.0005
R1365 VDDA.n128 VDDA.n127 30.754
R1366 VDDA.n92 VDDA.n91 30.754
R1367 VDDA.n112 VDDA.n111 30.186
R1368 VDDA.n87 VDDA.n86 30.186
R1369 VDDA.n373 VDDA.n372 28.8005
R1370 VDDA.n273 VDDA.n174 28.8005
R1371 VDDA.n198 VDDA.n189 28.8005
R1372 VDDA.n254 VDDA.n253 28.8005
R1373 VDDA.n294 VDDA.n293 25.6005
R1374 VDDA.n379 VDDA.n38 25.6005
R1375 VDDA.n391 VDDA.n390 25.6005
R1376 VDDA.n415 VDDA.n414 25.6005
R1377 VDDA.n420 VDDA.n15 25.6005
R1378 VDDA.n487 VDDA.n486 25.6005
R1379 VDDA.n502 VDDA.n9 25.6005
R1380 VDDA.n503 VDDA.n502 25.6005
R1381 VDDA.n517 VDDA.n516 25.6005
R1382 VDDA.n137 VDDA.n136 25.6005
R1383 VDDA VDDA.n170 25.6005
R1384 VDDA.t73 VDDA.t56 25.3822
R1385 VDDA.t95 VDDA.t77 25.3822
R1386 VDDA.n355 VDDA.t15 24.6255
R1387 VDDA.n44 VDDA.t86 24.6255
R1388 VDDA.n50 VDDA.t129 24.6255
R1389 VDDA.n283 VDDA.t38 24.6255
R1390 VDDA.n346 VDDA.t3 24.6255
R1391 VDDA.n51 VDDA.t13 24.6255
R1392 VDDA.n191 VDDA.t55 24.6255
R1393 VDDA.n191 VDDA.t124 24.6255
R1394 VDDA.n188 VDDA.t70 24.6255
R1395 VDDA.n188 VDDA.t26 24.6255
R1396 VDDA.t121 VDDA.n255 24.6255
R1397 VDDA.n255 VDDA.t49 24.6255
R1398 VDDA.n211 VDDA.t72 24.6255
R1399 VDDA.n211 VDDA.t107 24.6255
R1400 VDDA.n214 VDDA.t1 24.6255
R1401 VDDA.n214 VDDA.t11 24.6255
R1402 VDDA.n231 VDDA.t114 24.6255
R1403 VDDA.n231 VDDA.t9 24.6255
R1404 VDDA.t114 VDDA.n230 24.6255
R1405 VDDA.n175 VDDA.t125 24.6255
R1406 VDDA.n256 VDDA.t121 24.6255
R1407 VDDA.n260 VDDA.t108 24.6255
R1408 VDDA.n220 VDDA.n217 24.361
R1409 VDDA.n196 VDDA.n192 22.4005
R1410 VDDA.n247 VDDA.n246 22.4005
R1411 VDDA.n248 VDDA.n180 22.4005
R1412 VDDA.n105 VDDA.n96 22.0449
R1413 VDDA.n116 VDDA.t104 19.7005
R1414 VDDA.n97 VDDA.t101 19.7005
R1415 VDDA.n67 VDDA.t68 19.7005
R1416 VDDA.n67 VDDA.t100 19.7005
R1417 VDDA.n70 VDDA.t76 19.7005
R1418 VDDA.n70 VDDA.t62 19.7005
R1419 VDDA.n73 VDDA.t78 19.7005
R1420 VDDA.n73 VDDA.t80 19.7005
R1421 VDDA.n76 VDDA.t64 19.7005
R1422 VDDA.n76 VDDA.t74 19.7005
R1423 VDDA.t104 VDDA.n81 19.7005
R1424 VDDA.n81 VDDA.t47 19.7005
R1425 VDDA.n32 VDDA.n24 19.2005
R1426 VDDA.t52 VDDA.t63 18.1303
R1427 VDDA.t87 VDDA.t99 18.1303
R1428 VDDA.n273 VDDA.n272 17.6005
R1429 VDDA.n397 VDDA.n396 16.0005
R1430 VDDA.n129 VDDA.n128 16.0005
R1431 VDDA.n91 VDDA.n90 16.0005
R1432 VDDA.n111 VDDA.n110 16.0005
R1433 VDDA.n86 VDDA.n83 16.0005
R1434 VDDA.n192 VDDA.n174 16.0005
R1435 VDDA.n208 VDDA.n180 16.0005
R1436 VDDA.n246 VDDA.n245 16.0005
R1437 VDDA.n233 VDDA.n232 16.0005
R1438 VDDA.n171 VDDA 15.7005
R1439 VDDA.n272 VDDA.n271 15.6449
R1440 VDDA.n229 VDDA.n220 15.6449
R1441 VDDA.n293 VDDA.n281 13.8989
R1442 VDDA.n398 VDDA.n30 12.8005
R1443 VDDA.n415 VDDA.n24 12.8005
R1444 VDDA.n280 VDDA.n171 12.7493
R1445 VDDA.n281 VDDA.n280 12.3383
R1446 VDDA.n280 VDDA.n279 11.579
R1447 VDDA.n343 VDDA.t41 11.4924
R1448 VDDA.t16 VDDA.n335 11.4924
R1449 VDDA.n327 VDDA.t65 11.4924
R1450 VDDA.n405 VDDA.t31 11.4924
R1451 VDDA.n411 VDDA.t44 11.4924
R1452 VDDA.t14 VDDA.t61 10.8784
R1453 VDDA.n96 VDDA.n65 9.613
R1454 VDDA.n274 VDDA.n273 9.6005
R1455 VDDA.n254 VDDA.n186 9.6005
R1456 VDDA.n202 VDDA.n189 9.6005
R1457 VDDA.n170 VDDA.n63 9.3005
R1458 VDDA.n169 VDDA.n168 9.3005
R1459 VDDA.n167 VDDA.n64 9.3005
R1460 VDDA.n166 VDDA.n165 9.3005
R1461 VDDA.n164 VDDA.n163 9.3005
R1462 VDDA.n162 VDDA.n66 9.3005
R1463 VDDA.n160 VDDA.n159 9.3005
R1464 VDDA.n158 VDDA.n68 9.3005
R1465 VDDA.n157 VDDA.n156 9.3005
R1466 VDDA.n155 VDDA.n69 9.3005
R1467 VDDA.n153 VDDA.n152 9.3005
R1468 VDDA.n151 VDDA.n71 9.3005
R1469 VDDA.n150 VDDA.n149 9.3005
R1470 VDDA.n148 VDDA.n72 9.3005
R1471 VDDA.n146 VDDA.n145 9.3005
R1472 VDDA.n144 VDDA.n74 9.3005
R1473 VDDA.n143 VDDA.n142 9.3005
R1474 VDDA.n141 VDDA.n75 9.3005
R1475 VDDA.n139 VDDA.n138 9.3005
R1476 VDDA.n133 VDDA.n80 9.3005
R1477 VDDA.n135 VDDA.n134 9.3005
R1478 VDDA.n136 VDDA.n77 9.3005
R1479 VDDA.n233 VDDA.n216 9.3005
R1480 VDDA.n235 VDDA.n234 9.3005
R1481 VDDA.n236 VDDA.n215 9.3005
R1482 VDDA.n238 VDDA.n237 9.3005
R1483 VDDA.n240 VDDA.n213 9.3005
R1484 VDDA.n242 VDDA.n241 9.3005
R1485 VDDA.n243 VDDA.n212 9.3005
R1486 VDDA.n245 VDDA.n244 9.3005
R1487 VDDA.n246 VDDA.n210 9.3005
R1488 VDDA.n247 VDDA.n209 9.3005
R1489 VDDA.n249 VDDA.n248 9.3005
R1490 VDDA.n250 VDDA.n180 9.3005
R1491 VDDA.n251 VDDA.n208 9.3005
R1492 VDDA.n253 VDDA.n252 9.3005
R1493 VDDA.n254 VDDA.n207 9.3005
R1494 VDDA.n206 VDDA.n186 9.3005
R1495 VDDA.n205 VDDA.n204 9.3005
R1496 VDDA.n203 VDDA.n187 9.3005
R1497 VDDA.n202 VDDA.n201 9.3005
R1498 VDDA.n200 VDDA.n189 9.3005
R1499 VDDA.n199 VDDA.n198 9.3005
R1500 VDDA.n197 VDDA.n190 9.3005
R1501 VDDA.n196 VDDA.n195 9.3005
R1502 VDDA.n194 VDDA.n192 9.3005
R1503 VDDA.n193 VDDA.n174 9.3005
R1504 VDDA.n273 VDDA.n173 9.3005
R1505 VDDA.n275 VDDA.n274 9.3005
R1506 VDDA.n276 VDDA.n172 9.3005
R1507 VDDA.n278 VDDA.n277 9.3005
R1508 VDDA.n517 VDDA.n0 9.3005
R1509 VDDA.n295 VDDA.n294 9.3005
R1510 VDDA.n296 VDDA.n62 9.3005
R1511 VDDA.n298 VDDA.n297 9.3005
R1512 VDDA.n299 VDDA.n61 9.3005
R1513 VDDA.n301 VDDA.n300 9.3005
R1514 VDDA.n302 VDDA.n59 9.3005
R1515 VDDA.n306 VDDA.n305 9.3005
R1516 VDDA.n304 VDDA.n60 9.3005
R1517 VDDA.n303 VDDA.n42 9.3005
R1518 VDDA.n374 VDDA.n373 9.3005
R1519 VDDA.n375 VDDA.n40 9.3005
R1520 VDDA.n377 VDDA.n376 9.3005
R1521 VDDA.n378 VDDA.n39 9.3005
R1522 VDDA.n380 VDDA.n379 9.3005
R1523 VDDA.n382 VDDA.n381 9.3005
R1524 VDDA.n383 VDDA.n37 9.3005
R1525 VDDA.n385 VDDA.n384 9.3005
R1526 VDDA.n386 VDDA.n36 9.3005
R1527 VDDA.n388 VDDA.n387 9.3005
R1528 VDDA.n391 VDDA.n33 9.3005
R1529 VDDA.n393 VDDA.n392 9.3005
R1530 VDDA.n394 VDDA.n30 9.3005
R1531 VDDA.n396 VDDA.n395 9.3005
R1532 VDDA.n32 VDDA.n23 9.3005
R1533 VDDA.n416 VDDA.n415 9.3005
R1534 VDDA.n417 VDDA.n22 9.3005
R1535 VDDA.n419 VDDA.n418 9.3005
R1536 VDDA.n15 VDDA.n14 9.3005
R1537 VDDA.n488 VDDA.n487 9.3005
R1538 VDDA.n489 VDDA.n13 9.3005
R1539 VDDA.n491 VDDA.n490 9.3005
R1540 VDDA.n492 VDDA.n12 9.3005
R1541 VDDA.n494 VDDA.n493 9.3005
R1542 VDDA.n495 VDDA.n11 9.3005
R1543 VDDA.n497 VDDA.n496 9.3005
R1544 VDDA.n498 VDDA.n10 9.3005
R1545 VDDA.n500 VDDA.n499 9.3005
R1546 VDDA.n502 VDDA.n501 9.3005
R1547 VDDA.n504 VDDA.n6 9.3005
R1548 VDDA.n506 VDDA.n505 9.3005
R1549 VDDA.n507 VDDA.n5 9.3005
R1550 VDDA.n509 VDDA.n508 9.3005
R1551 VDDA.n510 VDDA.n4 9.3005
R1552 VDDA.n512 VDDA.n511 9.3005
R1553 VDDA.n513 VDDA.n3 9.3005
R1554 VDDA.n515 VDDA.n514 9.3005
R1555 VDDA.n442 VDDA.n440 9.14336
R1556 VDDA.n479 VDDA.n477 9.14336
R1557 VDDA.n423 VDDA.n21 9.14336
R1558 VDDA.n401 VDDA.n29 9.14336
R1559 VDDA.n331 VDDA.n329 9.14336
R1560 VDDA.n436 VDDA.n435 9.14336
R1561 VDDA.n473 VDDA.n472 9.14336
R1562 VDDA.n408 VDDA.n407 9.14336
R1563 VDDA.n324 VDDA.n323 9.14336
R1564 VDDA.n340 VDDA.n339 9.14336
R1565 VDDA.t23 VDDA.t59 7.66179
R1566 VDDA.n126 VDDA.n125 7.25241
R1567 VDDA.n361 VDDA.n360 7.11161
R1568 VDDA.n358 VDDA.n356 7.11161
R1569 VDDA.n367 VDDA.n366 7.11161
R1570 VDDA.n371 VDDA.n43 7.11161
R1571 VDDA.n312 VDDA.n311 7.11161
R1572 VDDA.n309 VDDA.n307 7.11161
R1573 VDDA.n288 VDDA.n287 7.11161
R1574 VDDA.n292 VDDA.n282 7.11161
R1575 VDDA.n352 VDDA.n351 7.11161
R1576 VDDA.n349 VDDA.n347 7.11161
R1577 VDDA.n58 VDDA.n57 7.11161
R1578 VDDA.n54 VDDA.n53 7.11161
R1579 VDDA.n123 VDDA.n122 7.11161
R1580 VDDA.n120 VDDA.n119 7.11161
R1581 VDDA.n105 VDDA.n104 7.11161
R1582 VDDA.n102 VDDA.n99 7.11161
R1583 VDDA.n271 VDDA.n176 7.11161
R1584 VDDA.n266 VDDA.n264 7.11161
R1585 VDDA.n229 VDDA.n228 7.11161
R1586 VDDA.n222 VDDA.n219 7.11161
R1587 VDDA.n232 VDDA.n217 6.54033
R1588 VDDA.n382 VDDA.n38 6.4005
R1589 VDDA.n414 VDDA.n22 6.4005
R1590 VDDA.n420 VDDA.n419 6.4005
R1591 VDDA.n486 VDDA.n13 6.4005
R1592 VDDA.n499 VDDA.n9 6.4005
R1593 VDDA.n504 VDDA.n503 6.4005
R1594 VDDA.n516 VDDA.n515 6.4005
R1595 VDDA.n138 VDDA.n137 6.4005
R1596 VDDA.n465 VDDA.n461 5.81868
R1597 VDDA.n454 VDDA.n450 5.81868
R1598 VDDA.n336 VDDA.n34 5.33286
R1599 VDDA.n443 VDDA.n1 5.33286
R1600 VDDA.n480 VDDA.n16 5.33286
R1601 VDDA.n424 VDDA.n421 5.33286
R1602 VDDA.n402 VDDA.n399 5.33286
R1603 VDDA.n332 VDDA.n35 5.33286
R1604 VDDA.n433 VDDA.n2 5.33286
R1605 VDDA.n485 VDDA.n17 5.33286
R1606 VDDA.n413 VDDA.n25 5.33286
R1607 VDDA.n321 VDDA.n31 5.33286
R1608 VDDA.n444 VDDA.n440 3.75335
R1609 VDDA.n443 VDDA.n442 3.75335
R1610 VDDA.n481 VDDA.n477 3.75335
R1611 VDDA.n480 VDDA.n479 3.75335
R1612 VDDA.n425 VDDA.n21 3.75335
R1613 VDDA.n424 VDDA.n423 3.75335
R1614 VDDA.n403 VDDA.n29 3.75335
R1615 VDDA.n402 VDDA.n401 3.75335
R1616 VDDA.n333 VDDA.n329 3.75335
R1617 VDDA.n332 VDDA.n331 3.75335
R1618 VDDA.n436 VDDA.n433 3.75335
R1619 VDDA.n435 VDDA.n434 3.75335
R1620 VDDA.n472 VDDA.n17 3.75335
R1621 VDDA.n473 VDDA.n471 3.75335
R1622 VDDA.n407 VDDA.n25 3.75335
R1623 VDDA.n408 VDDA.n406 3.75335
R1624 VDDA.n324 VDDA.n321 3.75335
R1625 VDDA.n323 VDDA.n322 3.75335
R1626 VDDA.n340 VDDA.n336 3.75335
R1627 VDDA.n339 VDDA.n338 3.75335
R1628 VDDA.n360 VDDA.n359 3.53508
R1629 VDDA.n359 VDDA.n358 3.53508
R1630 VDDA.n366 VDDA.n365 3.53508
R1631 VDDA.n365 VDDA.n43 3.53508
R1632 VDDA.n311 VDDA.n310 3.53508
R1633 VDDA.n310 VDDA.n309 3.53508
R1634 VDDA.n287 VDDA.n286 3.53508
R1635 VDDA.n286 VDDA.n282 3.53508
R1636 VDDA.n351 VDDA.n350 3.53508
R1637 VDDA.n350 VDDA.n349 3.53508
R1638 VDDA.n57 VDDA.n52 3.53508
R1639 VDDA.n54 VDDA.n52 3.53508
R1640 VDDA.n122 VDDA.n121 3.53508
R1641 VDDA.n119 VDDA.n117 3.53508
R1642 VDDA.n121 VDDA.n120 3.53508
R1643 VDDA.n104 VDDA.n103 3.53508
R1644 VDDA.n99 VDDA.n98 3.53508
R1645 VDDA.n103 VDDA.n102 3.53508
R1646 VDDA.n265 VDDA.n176 3.53508
R1647 VDDA.n266 VDDA.n265 3.53508
R1648 VDDA.n228 VDDA.n218 3.53508
R1649 VDDA.n222 VDDA.n218 3.53508
R1650 VDDA.n468 VDDA.n467 3.40194
R1651 VDDA.n466 VDDA.n462 3.40194
R1652 VDDA.n457 VDDA.n456 3.40194
R1653 VDDA.n455 VDDA.n451 3.40194
R1654 VDDA.n372 VDDA.n40 3.2005
R1655 VDDA.n389 VDDA.n388 3.2005
R1656 VDDA.n390 VDDA.n389 3.2005
R1657 VDDA.n398 VDDA.n397 3.2005
R1658 VDDA.n240 VDDA.n239 3.2005
R1659 VDDA.n239 VDDA.n238 3.2005
R1660 VDDA.n467 VDDA.n461 2.39444
R1661 VDDA.n466 VDDA.n465 2.39444
R1662 VDDA.n456 VDDA.n450 2.39444
R1663 VDDA.n455 VDDA.n454 2.39444
R1664 VDDA.n462 VDDA.n7 2.32777
R1665 VDDA.n457 VDDA.n8 2.32777
R1666 VDDA.n182 VDDA.n181 2.27782
R1667 VDDA.n183 VDDA.n182 2.27782
R1668 VDDA.n259 VDDA.n257 2.27782
R1669 VDDA.n185 VDDA.n183 2.27782
R1670 VDDA.n261 VDDA.n181 2.27782
R1671 VDDA.n257 VDDA.n185 2.27782
R1672 VDDA.n217 VDDA.n216 0.703395
R1673 VDDA.n295 VDDA.n281 0.193961
R1674 VDDA.n171 VDDA.n63 0.188
R1675 VDDA.n134 VDDA.n133 0.15675
R1676 VDDA.n134 VDDA.n77 0.15675
R1677 VDDA.n139 VDDA.n77 0.15675
R1678 VDDA.n142 VDDA.n141 0.15675
R1679 VDDA.n142 VDDA.n74 0.15675
R1680 VDDA.n146 VDDA.n74 0.15675
R1681 VDDA.n149 VDDA.n148 0.15675
R1682 VDDA.n149 VDDA.n71 0.15675
R1683 VDDA.n153 VDDA.n71 0.15675
R1684 VDDA.n156 VDDA.n155 0.15675
R1685 VDDA.n156 VDDA.n68 0.15675
R1686 VDDA.n160 VDDA.n68 0.15675
R1687 VDDA.n163 VDDA.n162 0.15675
R1688 VDDA.n167 VDDA.n166 0.15675
R1689 VDDA.n168 VDDA.n167 0.15675
R1690 VDDA.n168 VDDA.n63 0.15675
R1691 VDDA.n235 VDDA.n216 0.15675
R1692 VDDA.n236 VDDA.n235 0.15675
R1693 VDDA.n237 VDDA.n236 0.15675
R1694 VDDA.n237 VDDA.n213 0.15675
R1695 VDDA.n242 VDDA.n213 0.15675
R1696 VDDA.n243 VDDA.n242 0.15675
R1697 VDDA.n244 VDDA.n243 0.15675
R1698 VDDA.n244 VDDA.n210 0.15675
R1699 VDDA.n210 VDDA.n209 0.15675
R1700 VDDA.n249 VDDA.n209 0.15675
R1701 VDDA.n250 VDDA.n249 0.15675
R1702 VDDA.n251 VDDA.n250 0.15675
R1703 VDDA.n252 VDDA.n251 0.15675
R1704 VDDA.n252 VDDA.n207 0.15675
R1705 VDDA.n207 VDDA.n206 0.15675
R1706 VDDA.n206 VDDA.n205 0.15675
R1707 VDDA.n205 VDDA.n187 0.15675
R1708 VDDA.n201 VDDA.n187 0.15675
R1709 VDDA.n201 VDDA.n200 0.15675
R1710 VDDA.n200 VDDA.n199 0.15675
R1711 VDDA.n199 VDDA.n190 0.15675
R1712 VDDA.n195 VDDA.n190 0.15675
R1713 VDDA.n195 VDDA.n194 0.15675
R1714 VDDA.n194 VDDA.n193 0.15675
R1715 VDDA.n193 VDDA.n173 0.15675
R1716 VDDA.n275 VDDA.n173 0.15675
R1717 VDDA.n276 VDDA.n275 0.15675
R1718 VDDA.n277 VDDA.n276 0.15675
R1719 VDDA.n296 VDDA.n295 0.15675
R1720 VDDA.n297 VDDA.n296 0.15675
R1721 VDDA.n297 VDDA.n61 0.15675
R1722 VDDA.n301 VDDA.n61 0.15675
R1723 VDDA.n302 VDDA.n301 0.15675
R1724 VDDA.n305 VDDA.n302 0.15675
R1725 VDDA.n305 VDDA.n304 0.15675
R1726 VDDA.n304 VDDA.n303 0.15675
R1727 VDDA.n375 VDDA.n374 0.15675
R1728 VDDA.n376 VDDA.n375 0.15675
R1729 VDDA.n376 VDDA.n39 0.15675
R1730 VDDA.n380 VDDA.n39 0.15675
R1731 VDDA.n381 VDDA.n380 0.15675
R1732 VDDA.n381 VDDA.n37 0.15675
R1733 VDDA.n385 VDDA.n37 0.15675
R1734 VDDA.n386 VDDA.n385 0.15675
R1735 VDDA.n387 VDDA.n386 0.15675
R1736 VDDA.n387 VDDA.n33 0.15675
R1737 VDDA.n393 VDDA.n33 0.15675
R1738 VDDA.n394 VDDA.n393 0.15675
R1739 VDDA.n395 VDDA.n394 0.15675
R1740 VDDA.n395 VDDA.n23 0.15675
R1741 VDDA.n416 VDDA.n23 0.15675
R1742 VDDA.n417 VDDA.n416 0.15675
R1743 VDDA.n418 VDDA.n417 0.15675
R1744 VDDA.n418 VDDA.n14 0.15675
R1745 VDDA.n488 VDDA.n14 0.15675
R1746 VDDA.n489 VDDA.n488 0.15675
R1747 VDDA.n490 VDDA.n489 0.15675
R1748 VDDA.n490 VDDA.n12 0.15675
R1749 VDDA.n494 VDDA.n12 0.15675
R1750 VDDA.n495 VDDA.n494 0.15675
R1751 VDDA.n496 VDDA.n495 0.15675
R1752 VDDA.n496 VDDA.n10 0.15675
R1753 VDDA.n500 VDDA.n10 0.15675
R1754 VDDA.n501 VDDA.n500 0.15675
R1755 VDDA.n501 VDDA.n6 0.15675
R1756 VDDA.n506 VDDA.n6 0.15675
R1757 VDDA.n507 VDDA.n506 0.15675
R1758 VDDA.n508 VDDA.n507 0.15675
R1759 VDDA.n508 VDDA.n4 0.15675
R1760 VDDA.n512 VDDA.n4 0.15675
R1761 VDDA.n513 VDDA.n512 0.15675
R1762 VDDA.n514 VDDA.n513 0.15675
R1763 VDDA.n514 VDDA.n0 0.15675
R1764 VDDA VDDA.n0 0.1255
R1765 VDDA.n277 VDDA 0.122375
R1766 VDDA.n132 VDDA.n131 0.100307
R1767 VDDA.n133 VDDA.n132 0.09425
R1768 VDDA.n141 VDDA.n140 0.09425
R1769 VDDA.n148 VDDA.n147 0.09425
R1770 VDDA.n155 VDDA.n154 0.09425
R1771 VDDA.n162 VDDA.n161 0.09425
R1772 VDDA.n166 VDDA.n65 0.09425
R1773 VDDA.n303 VDDA.n41 0.078625
R1774 VDDA.n374 VDDA.n41 0.078625
R1775 VDDA.n140 VDDA.n139 0.063
R1776 VDDA.n147 VDDA.n146 0.063
R1777 VDDA.n154 VDDA.n153 0.063
R1778 VDDA.n161 VDDA.n160 0.063
R1779 VDDA.n163 VDDA.n65 0.063
R1780 VDDA.n279 VDDA 0.0505
R1781 pfd_8_0.DOWN_PFD_b.t0 pfd_8_0.DOWN_PFD_b.n1 203.528
R1782 pfd_8_0.DOWN_PFD_b.n0 pfd_8_0.DOWN_PFD_b.t1 203.528
R1783 pfd_8_0.DOWN_PFD_b.n1 pfd_8_0.DOWN_PFD_b.t2 183.935
R1784 pfd_8_0.DOWN_PFD_b.n0 pfd_8_0.DOWN_PFD_b.t3 183.935
R1785 pfd_8_0.DOWN_PFD_b.n1 pfd_8_0.DOWN_PFD_b.n0 83.2005
R1786 pfd_8_0.DOWN_b.n0 pfd_8_0.DOWN_b.t5 1028.27
R1787 pfd_8_0.DOWN_b.n2 pfd_8_0.DOWN_b.n1 569.734
R1788 pfd_8_0.DOWN_b.n1 pfd_8_0.DOWN_b.n0 465.933
R1789 pfd_8_0.DOWN_b.n1 pfd_8_0.DOWN_b.t3 401.668
R1790 pfd_8_0.DOWN_b.n0 pfd_8_0.DOWN_b.t4 385.601
R1791 pfd_8_0.DOWN_b.n1 pfd_8_0.DOWN_b.t2 385.601
R1792 pfd_8_0.DOWN_b.t0 pfd_8_0.DOWN_b.n2 211.847
R1793 pfd_8_0.DOWN_b.n2 pfd_8_0.DOWN_b.t1 173.055
R1794 pfd_8_0.QA_b.t4 pfd_8_0.QA_b.t6 1188.93
R1795 pfd_8_0.QA_b pfd_8_0.QA_b.n2 837.38
R1796 pfd_8_0.QA_b.t6 pfd_8_0.QA_b.t3 835.467
R1797 pfd_8_0.QA_b.n0 pfd_8_0.QA_b.t5 562.333
R1798 pfd_8_0.QA_b pfd_8_0.QA_b.n0 482
R1799 pfd_8_0.QA_b.n2 pfd_8_0.QA_b.n1 247.917
R1800 pfd_8_0.QA_b.n0 pfd_8_0.QA_b.t4 224.934
R1801 pfd_8_0.QA_b.n2 pfd_8_0.QA_b.t2 221.411
R1802 pfd_8_0.QA_b.n1 pfd_8_0.QA_b.t1 24.0005
R1803 pfd_8_0.QA_b.n1 pfd_8_0.QA_b.t0 24.0005
R1804 a_870_1400.t0 a_870_1400.t1 39.4005
R1805 pfd_8_0.DOWN.n0 pfd_8_0.DOWN.t2 605.311
R1806 pfd_8_0.DOWN.t1 pfd_8_0.DOWN.n0 240.327
R1807 pfd_8_0.DOWN.n0 pfd_8_0.DOWN.t0 148.736
R1808 pfd_8_0.UP_input.n14 pfd_8_0.UP_input.n13 424.447
R1809 pfd_8_0.UP_input.n14 pfd_8_0.UP_input.n12 354.048
R1810 pfd_8_0.UP_input.t18 pfd_8_0.UP_input.n11 326.658
R1811 pfd_8_0.UP_input.n2 pfd_8_0.UP_input.n1 313
R1812 pfd_8_0.UP_input.n9 pfd_8_0.UP_input.t15 297.233
R1813 pfd_8_0.UP_input.t17 pfd_8_0.UP_input.n10 297.233
R1814 pfd_8_0.UP_input.n17 pfd_8_0.UP_input.t21 297.233
R1815 pfd_8_0.UP_input.n18 pfd_8_0.UP_input.t21 297.233
R1816 pfd_8_0.UP_input.t19 pfd_8_0.UP_input.n19 297.233
R1817 pfd_8_0.UP_input.n21 pfd_8_0.UP_input.t9 281.596
R1818 pfd_8_0.UP_input.n8 pfd_8_0.UP_input.n4 257.067
R1819 pfd_8_0.UP_input.n7 pfd_8_0.UP_input.n6 246.275
R1820 pfd_8_0.UP_input.n2 pfd_8_0.UP_input.n0 242.601
R1821 pfd_8_0.UP_input.n5 pfd_8_0.UP_input.t8 241.928
R1822 pfd_8_0.UP_input.n8 pfd_8_0.UP_input.n7 226.942
R1823 pfd_8_0.UP_input.n11 pfd_8_0.UP_input.n4 226.942
R1824 pfd_8_0.UP_input.n3 pfd_8_0.UP_input.n2 220.8
R1825 pfd_8_0.UP_input.n15 pfd_8_0.UP_input.n14 220.8
R1826 pfd_8_0.UP_input.n10 pfd_8_0.UP_input.n9 216.9
R1827 pfd_8_0.UP_input.n19 pfd_8_0.UP_input.n18 216.9
R1828 pfd_8_0.UP_input.n17 pfd_8_0.UP_input.n16 216.9
R1829 pfd_8_0.UP_input.n22 pfd_8_0.UP_input.n20 215.107
R1830 pfd_8_0.UP_input.n6 pfd_8_0.UP_input.t3 209.928
R1831 pfd_8_0.UP_input.n20 pfd_8_0.UP_input.n16 184.768
R1832 pfd_8_0.UP_input.n5 pfd_8_0.UP_input.t11 145.535
R1833 pfd_8_0.UP_input.n6 pfd_8_0.UP_input.n5 144
R1834 pfd_8_0.UP_input.n21 pfd_8_0.UP_input.t12 118.666
R1835 pfd_8_0.UP_input.n7 pfd_8_0.UP_input.t15 92.3838
R1836 pfd_8_0.UP_input.n11 pfd_8_0.UP_input.t17 92.3838
R1837 pfd_8_0.UP_input.n9 pfd_8_0.UP_input.t14 80.3338
R1838 pfd_8_0.UP_input.t14 pfd_8_0.UP_input.n8 80.3338
R1839 pfd_8_0.UP_input.n10 pfd_8_0.UP_input.t20 80.3338
R1840 pfd_8_0.UP_input.t20 pfd_8_0.UP_input.n4 80.3338
R1841 pfd_8_0.UP_input.n18 pfd_8_0.UP_input.t22 80.3338
R1842 pfd_8_0.UP_input.t22 pfd_8_0.UP_input.n17 80.3338
R1843 pfd_8_0.UP_input.n19 pfd_8_0.UP_input.t13 80.3338
R1844 pfd_8_0.UP_input.t13 pfd_8_0.UP_input.n16 80.3338
R1845 pfd_8_0.UP_input.n20 pfd_8_0.UP_input.t19 80.3338
R1846 pfd_8_0.UP_input.n23 pfd_8_0.UP_input.n22 78.9255
R1847 pfd_8_0.UP_input.n3 pfd_8_0.UP_input.t16 70.0829
R1848 pfd_8_0.UP_input.n15 pfd_8_0.UP_input.t18 63.6829
R1849 opamp_cell_4_0.VOUT pfd_8_0.UP_input.n3 62.4005
R1850 pfd_8_0.UP_input.n23 pfd_8_0.UP_input.n15 60.8005
R1851 pfd_8_0.UP_input.n22 pfd_8_0.UP_input.n21 60.2361
R1852 pfd_8_0.UP_input.n0 pfd_8_0.UP_input.t6 60.0005
R1853 pfd_8_0.UP_input.n0 pfd_8_0.UP_input.t5 60.0005
R1854 pfd_8_0.UP_input.n1 pfd_8_0.UP_input.t4 60.0005
R1855 pfd_8_0.UP_input.n1 pfd_8_0.UP_input.t7 60.0005
R1856 pfd_8_0.UP_input.n13 pfd_8_0.UP_input.t2 49.2505
R1857 pfd_8_0.UP_input.n13 pfd_8_0.UP_input.t10 49.2505
R1858 pfd_8_0.UP_input.n12 pfd_8_0.UP_input.t1 49.2505
R1859 pfd_8_0.UP_input.n12 pfd_8_0.UP_input.t0 49.2505
R1860 opamp_cell_4_0.VOUT pfd_8_0.UP_input.n23 1.6005
R1861 opamp_cell_4_0.VIN+.n0 opamp_cell_4_0.VIN+.t8 377.567
R1862 opamp_cell_4_0.VIN+.n1 opamp_cell_4_0.VIN+.t9 297.233
R1863 opamp_cell_4_0.VIN+.n2 opamp_cell_4_0.VIN+.n1 243.44
R1864 opamp_cell_4_0.VIN+.n2 opamp_cell_4_0.VIN+.n0 224.496
R1865 opamp_cell_4_0.VIN+.n0 opamp_cell_4_0.VIN+.t7 216.9
R1866 opamp_cell_4_0.VIN+.n5 opamp_cell_4_0.VIN+.n4 196.262
R1867 opamp_cell_4_0.VIN+.n5 opamp_cell_4_0.VIN+.n3 172.502
R1868 opamp_cell_4_0.VIN+.n7 opamp_cell_4_0.VIN+.n6 172.5
R1869 opamp_cell_4_0.VIN+.n1 opamp_cell_4_0.VIN+.t6 136.567
R1870 opamp_cell_4_0.VIN+.n7 opamp_cell_4_0.VIN+.n5 70.4005
R1871 opamp_cell_4_0.VIN+ opamp_cell_4_0.VIN+.n7 50.088
R1872 opamp_cell_4_0.VIN+.n3 opamp_cell_4_0.VIN+.t2 24.6255
R1873 opamp_cell_4_0.VIN+.n3 opamp_cell_4_0.VIN+.t1 24.6255
R1874 opamp_cell_4_0.VIN+.n6 opamp_cell_4_0.VIN+.t4 24.6255
R1875 opamp_cell_4_0.VIN+.n6 opamp_cell_4_0.VIN+.t3 24.6255
R1876 opamp_cell_4_0.VIN+.n4 opamp_cell_4_0.VIN+.t5 15.0005
R1877 opamp_cell_4_0.VIN+.n4 opamp_cell_4_0.VIN+.t0 15.0005
R1878 opamp_cell_4_0.VIN+ opamp_cell_4_0.VIN+.n2 3.138
R1879 a_6320_5840.n7 a_6320_5840.n5 482.582
R1880 a_6320_5840.n10 a_6320_5840.t4 304.634
R1881 a_6320_5840.n3 a_6320_5840.t2 304.634
R1882 a_6320_5840.t6 a_6320_5840.n10 277.914
R1883 a_6320_5840.n3 a_6320_5840.t3 276.289
R1884 a_6320_5840.n8 a_6320_5840.n1 204.201
R1885 a_6320_5840.n4 a_6320_5840.n2 204.201
R1886 a_6320_5840.n9 a_6320_5840.n0 204.201
R1887 a_6320_5840.n7 a_6320_5840.n6 120.981
R1888 a_6320_5840.n8 a_6320_5840.n4 74.6672
R1889 a_6320_5840.n9 a_6320_5840.n8 74.6672
R1890 a_6320_5840.n1 a_6320_5840.t0 60.0005
R1891 a_6320_5840.n1 a_6320_5840.t7 60.0005
R1892 a_6320_5840.t3 a_6320_5840.n2 60.0005
R1893 a_6320_5840.n2 a_6320_5840.t1 60.0005
R1894 a_6320_5840.n0 a_6320_5840.t8 60.0005
R1895 a_6320_5840.n0 a_6320_5840.t5 60.0005
R1896 a_6320_5840.n8 a_6320_5840.n7 37.763
R1897 a_6320_5840.n5 a_6320_5840.t11 24.0005
R1898 a_6320_5840.n5 a_6320_5840.t12 24.0005
R1899 a_6320_5840.n6 a_6320_5840.t10 24.0005
R1900 a_6320_5840.n6 a_6320_5840.t9 24.0005
R1901 a_6320_5840.n4 a_6320_5840.n3 16.0005
R1902 a_6320_5840.n10 a_6320_5840.n9 16.0005
R1903 opamp_cell_4_0.n_right.t2 opamp_cell_4_0.n_right.n6 1010.36
R1904 opamp_cell_4_0.n_right.n3 opamp_cell_4_0.n_right.n2 416.101
R1905 opamp_cell_4_0.n_right.n2 opamp_cell_4_0.n_right.n1 354.048
R1906 opamp_cell_4_0.n_right.n3 opamp_cell_4_0.n_right.t5 289.2
R1907 opamp_cell_4_0.n_right.n4 opamp_cell_4_0.n_right.t8 289.2
R1908 opamp_cell_4_0.n_right.n5 opamp_cell_4_0.n_right.t7 289.2
R1909 opamp_cell_4_0.n_right.n6 opamp_cell_4_0.n_right.t6 289.2
R1910 opamp_cell_4_0.n_right.n2 opamp_cell_4_0.n_right.n0 284.2
R1911 opamp_cell_4_0.n_right.n6 opamp_cell_4_0.n_right.n5 208.868
R1912 opamp_cell_4_0.n_right.n5 opamp_cell_4_0.n_right.n4 208.868
R1913 opamp_cell_4_0.n_right.n4 opamp_cell_4_0.n_right.n3 208.868
R1914 opamp_cell_4_0.n_right.n0 opamp_cell_4_0.n_right.t0 60.0005
R1915 opamp_cell_4_0.n_right.n0 opamp_cell_4_0.n_right.t1 60.0005
R1916 opamp_cell_4_0.n_right.n1 opamp_cell_4_0.n_right.t3 49.2505
R1917 opamp_cell_4_0.n_right.n1 opamp_cell_4_0.n_right.t4 49.2505
R1918 opamp_cell_4_0.n_left.n1 opamp_cell_4_0.n_left.t7 401.668
R1919 opamp_cell_4_0.n_left.n5 opamp_cell_4_0.n_left.n4 325.248
R1920 opamp_cell_4_0.n_left.n4 opamp_cell_4_0.n_left.n0 313
R1921 opamp_cell_4_0.n_left.n3 opamp_cell_4_0.n_left.t0 252.248
R1922 opamp_cell_4_0.n_left.n2 opamp_cell_4_0.n_left.n1 208.868
R1923 opamp_cell_4_0.n_left.n2 opamp_cell_4_0.n_left.t2 192.8
R1924 opamp_cell_4_0.n_left.n1 opamp_cell_4_0.n_left.t6 192.8
R1925 opamp_cell_4_0.n_left.n4 opamp_cell_4_0.n_left.n3 152
R1926 opamp_cell_4_0.n_left.n0 opamp_cell_4_0.n_left.t5 60.0005
R1927 opamp_cell_4_0.n_left.n0 opamp_cell_4_0.n_left.t4 60.0005
R1928 opamp_cell_4_0.n_left.n3 opamp_cell_4_0.n_left.n2 59.4472
R1929 opamp_cell_4_0.n_left.t3 opamp_cell_4_0.n_left.n5 49.2505
R1930 opamp_cell_4_0.n_left.n5 opamp_cell_4_0.n_left.t1 49.2505
R1931 a_6490_4630.t2 a_6490_4630.n6 1112.76
R1932 a_6490_4630.n3 a_6490_4630.n2 416.863
R1933 a_6490_4630.n2 a_6490_4630.n1 366.848
R1934 a_6490_4630.n2 a_6490_4630.n0 271.401
R1935 a_6490_4630.n3 a_6490_4630.t5 208.868
R1936 a_6490_4630.n6 a_6490_4630.t6 208.868
R1937 a_6490_4630.n5 a_6490_4630.t7 208.868
R1938 a_6490_4630.n4 a_6490_4630.t8 208.868
R1939 a_6490_4630.n6 a_6490_4630.n5 208.868
R1940 a_6490_4630.n5 a_6490_4630.n4 208.868
R1941 a_6490_4630.n4 a_6490_4630.n3 193.804
R1942 a_6490_4630.n0 a_6490_4630.t4 60.0005
R1943 a_6490_4630.n0 a_6490_4630.t3 60.0005
R1944 a_6490_4630.n1 a_6490_4630.t1 49.2505
R1945 a_6490_4630.n1 a_6490_4630.t0 49.2505
R1946 pfd_8_0.before_Reset.n1 pfd_8_0.before_Reset.n0 481.334
R1947 pfd_8_0.before_Reset.n0 pfd_8_0.before_Reset.t4 465.933
R1948 pfd_8_0.before_Reset.n0 pfd_8_0.before_Reset.t3 321.334
R1949 pfd_8_0.before_Reset.n2 pfd_8_0.before_Reset.n1 226.889
R1950 pfd_8_0.before_Reset.n1 pfd_8_0.before_Reset.t0 172.458
R1951 pfd_8_0.before_Reset.n2 pfd_8_0.before_Reset.t2 19.7005
R1952 pfd_8_0.before_Reset.t1 pfd_8_0.before_Reset.n2 19.7005
R1953 a_2350_1400.t1 a_2350_1400.n2 500.086
R1954 a_2350_1400.n1 a_2350_1400.n0 473.334
R1955 a_2350_1400.n0 a_2350_1400.t3 465.933
R1956 a_2350_1400.t1 a_2350_1400.n2 461.389
R1957 a_2350_1400.n0 a_2350_1400.t2 321.334
R1958 a_2350_1400.n1 a_2350_1400.t0 177.577
R1959 a_2350_1400.n2 a_2350_1400.n1 48.3899
R1960 opamp_cell_4_0.p_bias opamp_cell_4_0.p_bias.t0 918.318
R1961 opamp_cell_4_0.p_bias opamp_cell_4_0.p_bias.n11 540.801
R1962 opamp_cell_4_0.p_bias.n8 opamp_cell_4_0.p_bias.t10 377.567
R1963 opamp_cell_4_0.p_bias.n3 opamp_cell_4_0.p_bias.t9 377.567
R1964 opamp_cell_4_0.p_bias.n9 opamp_cell_4_0.p_bias.n8 257.067
R1965 opamp_cell_4_0.p_bias.n7 opamp_cell_4_0.p_bias.n6 257.067
R1966 opamp_cell_4_0.p_bias.n4 opamp_cell_4_0.p_bias.n3 257.067
R1967 opamp_cell_4_0.p_bias.n11 opamp_cell_4_0.p_bias.n0 154.321
R1968 opamp_cell_4_0.p_bias.n2 opamp_cell_4_0.p_bias.n1 154.321
R1969 opamp_cell_4_0.p_bias.n5 opamp_cell_4_0.p_bias.n2 152
R1970 opamp_cell_4_0.p_bias.n11 opamp_cell_4_0.p_bias.n10 152
R1971 opamp_cell_4_0.p_bias.n8 opamp_cell_4_0.p_bias.t12 120.501
R1972 opamp_cell_4_0.p_bias.n9 opamp_cell_4_0.p_bias.t5 120.501
R1973 opamp_cell_4_0.p_bias.n7 opamp_cell_4_0.p_bias.t1 120.501
R1974 opamp_cell_4_0.p_bias.n6 opamp_cell_4_0.p_bias.t3 120.501
R1975 opamp_cell_4_0.p_bias.n3 opamp_cell_4_0.p_bias.t11 120.501
R1976 opamp_cell_4_0.p_bias.n4 opamp_cell_4_0.p_bias.t7 120.501
R1977 opamp_cell_4_0.p_bias.n11 opamp_cell_4_0.p_bias.n2 115.201
R1978 opamp_cell_4_0.p_bias.n10 opamp_cell_4_0.p_bias.n9 85.6894
R1979 opamp_cell_4_0.p_bias.n10 opamp_cell_4_0.p_bias.n7 85.6894
R1980 opamp_cell_4_0.p_bias.n6 opamp_cell_4_0.p_bias.n5 85.6894
R1981 opamp_cell_4_0.p_bias.n5 opamp_cell_4_0.p_bias.n4 85.6894
R1982 opamp_cell_4_0.p_bias.n0 opamp_cell_4_0.p_bias.t2 19.7005
R1983 opamp_cell_4_0.p_bias.n0 opamp_cell_4_0.p_bias.t6 19.7005
R1984 opamp_cell_4_0.p_bias.n1 opamp_cell_4_0.p_bias.t8 19.7005
R1985 opamp_cell_4_0.p_bias.n1 opamp_cell_4_0.p_bias.t4 19.7005
R1986 F_REF.n0 F_REF.t0 514.134
R1987 F_REF.n0 F_REF.t1 273.134
R1988 F_REF F_REF.n0 216.9
R1989 a_n30_1400.t0 a_n30_1400.t1 39.4005
R1990 pfd_8_0.QA.t5 pfd_8_0.QA.t7 835.467
R1991 pfd_8_0.QA.n2 pfd_8_0.QA.t4 517.347
R1992 pfd_8_0.QA.n0 pfd_8_0.QA.t8 465.933
R1993 pfd_8_0.QA.n1 pfd_8_0.QA.n0 454.031
R1994 pfd_8_0.QA.n1 pfd_8_0.QA.t5 394.267
R1995 pfd_8_0.QA.n0 pfd_8_0.QA.t6 321.334
R1996 pfd_8_0.QA.n4 pfd_8_0.QA.n3 244.715
R1997 pfd_8_0.QA.n2 pfd_8_0.QA.t3 228.148
R1998 pfd_8_0.QA.n4 pfd_8_0.QA.t0 221.411
R1999 pfd_8_0.QA.n5 pfd_8_0.QA.n2 216
R2000 pfd_8_0.QA.n5 pfd_8_0.QA.n4 201.573
R2001 pfd_8_0.QA pfd_8_0.QA.n5 60.8005
R2002 pfd_8_0.QA pfd_8_0.QA.n1 56.1505
R2003 pfd_8_0.QA.n3 pfd_8_0.QA.t2 24.0005
R2004 pfd_8_0.QA.n3 pfd_8_0.QA.t1 24.0005
R2005 I_IN.n4 I_IN.n3 1269.42
R2006 I_IN.n4 I_IN.t0 275.325
R2007 I_IN.n6 I_IN.n5 248.4
R2008 I_IN.n1 I_IN.t4 238.892
R2009 I_IN I_IN.n6 214.4
R2010 I_IN.n1 I_IN.t5 161.371
R2011 I_IN.n3 I_IN.t6 151.792
R2012 I_IN I_IN.n1 149.153
R2013 I_IN.n5 I_IN.t2 140.583
R2014 I_IN.n5 I_IN.t0 140.583
R2015 I_IN.n2 I_IN.n0 95.4614
R2016 I_IN.t2 I_IN.n4 80.3338
R2017 I_IN.n3 I_IN.t7 44.2902
R2018 I_IN.n0 I_IN.t3 15.0005
R2019 I_IN.n0 I_IN.t1 15.0005
R2020 I_IN.n2 I_IN 11.488
R2021 I_IN.n6 I_IN.n2 3.2005
R2022 pfd_8_0.DOWN_input.t4 pfd_8_0.DOWN_input.t3 377.567
R2023 pfd_8_0.DOWN_input.n2 pfd_8_0.DOWN_input.t5 326.658
R2024 pfd_8_0.DOWN_input.n0 pfd_8_0.DOWN_input.t1 229.127
R2025 pfd_8_0.DOWN_input pfd_8_0.DOWN_input.n3 225.601
R2026 pfd_8_0.DOWN_input.n3 pfd_8_0.DOWN_input.n2 196.817
R2027 pfd_8_0.DOWN_input.n0 pfd_8_0.DOWN_input.t0 158.335
R2028 pfd_8_0.DOWN_input.n1 pfd_8_0.DOWN_input.t2 158.335
R2029 pfd_8_0.DOWN_input.n1 pfd_8_0.DOWN_input.n0 121.6
R2030 pfd_8_0.DOWN_input.t3 pfd_8_0.DOWN_input.n2 92.3838
R2031 pfd_8_0.DOWN_input.n3 pfd_8_0.DOWN_input.t4 92.3838
R2032 pfd_8_0.DOWN_input pfd_8_0.DOWN_input.n1 3.2005
R2033 V_OUT.n2 V_OUT.n1 242.903
R2034 V_OUT.n2 V_OUT.n0 172.502
R2035 V_OUT.n6 V_OUT.t6 164.118
R2036 V_OUT.n7 V_OUT.n4 118.35
R2037 V_OUT.n4 V_OUT.n3 106.662
R2038 V_OUT.n0 V_OUT.t3 24.6255
R2039 V_OUT.n0 V_OUT.t2 24.6255
R2040 V_OUT.n1 V_OUT.t5 24.6255
R2041 V_OUT.n1 V_OUT.t4 24.6255
R2042 V_OUT.n4 V_OUT.n2 19.2005
R2043 V_OUT.n3 V_OUT.t1 15.0005
R2044 V_OUT.n3 V_OUT.t0 15.0005
R2045 V_OUT.n7 V_OUT.n6 9.91717
R2046 V_OUT.n6 V_OUT.t7 8.246
R2047 V_OUT.n7 V_OUT.n5 0.0838333
R2048 V_OUT V_OUT.n7 0.063
R2049 pfd_8_0.QB.t4 pfd_8_0.QB.t3 835.467
R2050 pfd_8_0.QB.n1 pfd_8_0.QB.t4 564.496
R2051 pfd_8_0.QB.n2 pfd_8_0.QB.t5 517.347
R2052 pfd_8_0.QB.n0 pfd_8_0.QB.t7 514.134
R2053 pfd_8_0.QB.n1 pfd_8_0.QB.n0 455.219
R2054 pfd_8_0.QB.n5 pfd_8_0.QB.n2 363.2
R2055 pfd_8_0.QB.n0 pfd_8_0.QB.t8 273.134
R2056 pfd_8_0.QB.n4 pfd_8_0.QB.n3 244.716
R2057 pfd_8_0.QB.n2 pfd_8_0.QB.t6 228.148
R2058 pfd_8_0.QB.n4 pfd_8_0.QB.t1 221.411
R2059 pfd_8_0.QB.n5 pfd_8_0.QB.n4 54.3734
R2060 pfd_8_0.QB pfd_8_0.QB.n1 26.7568
R2061 pfd_8_0.QB.n3 pfd_8_0.QB.t0 24.0005
R2062 pfd_8_0.QB.n3 pfd_8_0.QB.t2 24.0005
R2063 pfd_8_0.QB pfd_8_0.QB.n5 6.4005
R2064 a_1910_2020.t0 a_1910_2020.t1 48.0005
R2065 a_6220_5810.n4 a_6220_5810.t12 317.317
R2066 a_6220_5810.n2 a_6220_5810.t11 317.317
R2067 a_6220_5810.n5 a_6220_5810.n4 257.067
R2068 a_6220_5810.n3 a_6220_5810.n2 257.067
R2069 a_6220_5810.n10 a_6220_5810.n9 257.067
R2070 a_6220_5810.t0 a_6220_5810.n12 194.478
R2071 a_6220_5810.n8 a_6220_5810.n7 152
R2072 a_6220_5810.n12 a_6220_5810.n11 152
R2073 a_6220_5810.n1 a_6220_5810.n0 120.981
R2074 a_6220_5810.n7 a_6220_5810.n6 117.781
R2075 a_6220_5810.n7 a_6220_5810.n1 108.8
R2076 a_6220_5810.n8 a_6220_5810.n5 85.6894
R2077 a_6220_5810.n11 a_6220_5810.n3 85.6894
R2078 a_6220_5810.n11 a_6220_5810.n10 85.6894
R2079 a_6220_5810.n9 a_6220_5810.n8 85.6894
R2080 a_6220_5810.n4 a_6220_5810.t10 60.2505
R2081 a_6220_5810.n5 a_6220_5810.t1 60.2505
R2082 a_6220_5810.n2 a_6220_5810.t9 60.2505
R2083 a_6220_5810.n3 a_6220_5810.t3 60.2505
R2084 a_6220_5810.n10 a_6220_5810.t7 60.2505
R2085 a_6220_5810.n9 a_6220_5810.t5 60.2505
R2086 a_6220_5810.n6 a_6220_5810.t6 24.0005
R2087 a_6220_5810.n6 a_6220_5810.t2 24.0005
R2088 a_6220_5810.n0 a_6220_5810.t4 24.0005
R2089 a_6220_5810.n0 a_6220_5810.t8 24.0005
R2090 a_6220_5810.n12 a_6220_5810.n1 3.2005
R2091 pfd_8_0.UP_PFD_b.n0 pfd_8_0.UP_PFD_b.t2 441.834
R2092 pfd_8_0.UP_PFD_b.n0 pfd_8_0.UP_PFD_b.t3 313.3
R2093 pfd_8_0.UP_PFD_b.n1 pfd_8_0.UP_PFD_b.n0 235.201
R2094 pfd_8_0.UP_PFD_b.t1 pfd_8_0.UP_PFD_b.n1 219.528
R2095 pfd_8_0.UP_PFD_b.n1 pfd_8_0.UP_PFD_b.t0 167.935
R2096 pfd_8_0.UP.n0 pfd_8_0.UP.t5 1205
R2097 pfd_8_0.UP.n2 pfd_8_0.UP.t4 522.168
R2098 pfd_8_0.UP.n1 pfd_8_0.UP.n0 441.834
R2099 pfd_8_0.UP.n3 pfd_8_0.UP.n2 235.201
R2100 pfd_8_0.UP.t1 pfd_8_0.UP.n3 229.127
R2101 pfd_8_0.UP.n1 pfd_8_0.UP.t3 217.905
R2102 pfd_8_0.UP.n0 pfd_8_0.UP.t2 208.868
R2103 pfd_8_0.UP.n3 pfd_8_0.UP.t0 158.335
R2104 pfd_8_0.UP.n2 pfd_8_0.UP.n1 15.063
R2105 pfd_8_0.E.n4 pfd_8_0.E.n0 1319.38
R2106 pfd_8_0.E.n0 pfd_8_0.E.t3 562.333
R2107 pfd_8_0.E.n2 pfd_8_0.E.t5 388.813
R2108 pfd_8_0.E.n2 pfd_8_0.E.t4 356.68
R2109 pfd_8_0.E.n3 pfd_8_0.E.n2 232
R2110 pfd_8_0.E.n0 pfd_8_0.E.t6 224.934
R2111 pfd_8_0.E.t2 pfd_8_0.E.n4 221.411
R2112 pfd_8_0.E.n3 pfd_8_0.E.n1 157.278
R2113 pfd_8_0.E.n4 pfd_8_0.E.n3 90.64
R2114 pfd_8_0.E.n1 pfd_8_0.E.t1 24.0005
R2115 pfd_8_0.E.n1 pfd_8_0.E.t0 24.0005
R2116 pfd_8_0.E_b.n0 pfd_8_0.E_b.t4 517.347
R2117 pfd_8_0.E_b.n2 pfd_8_0.E_b.n0 417.574
R2118 pfd_8_0.E_b.n2 pfd_8_0.E_b.n1 244.716
R2119 pfd_8_0.E_b.n0 pfd_8_0.E_b.t3 228.148
R2120 pfd_8_0.E_b.t0 pfd_8_0.E_b.n2 221.411
R2121 pfd_8_0.E_b.n1 pfd_8_0.E_b.t2 24.0005
R2122 pfd_8_0.E_b.n1 pfd_8_0.E_b.t1 24.0005
R2123 a_1390_1400.t0 a_1390_1400.t1 39.4005
R2124 pfd_8_0.QB_b.t6 pfd_8_0.QB_b.t4 1188.93
R2125 pfd_8_0.QB_b pfd_8_0.QB_b.n2 899.734
R2126 pfd_8_0.QB_b.t4 pfd_8_0.QB_b.t3 835.467
R2127 pfd_8_0.QB_b.n2 pfd_8_0.QB_b.t5 562.333
R2128 pfd_8_0.QB_b pfd_8_0.QB_b.n1 419.647
R2129 pfd_8_0.QB_b.n1 pfd_8_0.QB_b.n0 247.917
R2130 pfd_8_0.QB_b.n2 pfd_8_0.QB_b.t6 224.934
R2131 pfd_8_0.QB_b.n1 pfd_8_0.QB_b.t1 221.411
R2132 pfd_8_0.QB_b.n0 pfd_8_0.QB_b.t2 24.0005
R2133 pfd_8_0.QB_b.n0 pfd_8_0.QB_b.t0 24.0005
R2134 a_870_640.t0 a_870_640.t1 39.4005
R2135 loop_filter_2_0.R1_C1.t0 loop_filter_2_0.R1_C1.t1 167.429
R2136 a_2530_190.t1 a_2530_190.n2 500.086
R2137 a_2530_190.n0 a_2530_190.t2 465.933
R2138 a_2530_190.t1 a_2530_190.n2 461.389
R2139 a_2530_190.n1 a_2530_190.n0 392.623
R2140 a_2530_190.n0 a_2530_190.t3 321.334
R2141 a_2530_190.n1 a_2530_190.t0 177.577
R2142 a_2530_190.n2 a_2530_190.n1 48.3899
R2143 a_2200_190.t1 a_2200_190.n2 500.086
R2144 a_2200_190.n1 a_2200_190.n0 473.334
R2145 a_2200_190.n0 a_2200_190.t2 465.933
R2146 a_2200_190.t1 a_2200_190.n2 461.389
R2147 a_2200_190.n0 a_2200_190.t3 321.334
R2148 a_2200_190.n1 a_2200_190.t0 177.577
R2149 a_2200_190.n2 a_2200_190.n1 48.3898
R2150 pfd_8_0.F.n4 pfd_8_0.F.n0 1319.38
R2151 pfd_8_0.F.n0 pfd_8_0.F.t3 562.333
R2152 pfd_8_0.F.n2 pfd_8_0.F.t5 388.813
R2153 pfd_8_0.F.n2 pfd_8_0.F.t6 356.68
R2154 pfd_8_0.F.n3 pfd_8_0.F.n2 232
R2155 pfd_8_0.F.n0 pfd_8_0.F.t4 224.934
R2156 pfd_8_0.F.t1 pfd_8_0.F.n4 221.411
R2157 pfd_8_0.F.n3 pfd_8_0.F.n1 157.278
R2158 pfd_8_0.F.n4 pfd_8_0.F.n3 90.64
R2159 pfd_8_0.F.n1 pfd_8_0.F.t0 24.0005
R2160 pfd_8_0.F.n1 pfd_8_0.F.t2 24.0005
R2161 a_9360_6440.t1 a_9360_6440.t0 245.883
R2162 pfd_8_0.UP_b.n0 pfd_8_0.UP_b.t2 778.601
R2163 pfd_8_0.UP_b.t1 pfd_8_0.UP_b.n0 209.928
R2164 pfd_8_0.UP_b.n0 pfd_8_0.UP_b.t0 177.536
R2165 pfd_8_0.F_b.n0 pfd_8_0.F_b.t3 517.347
R2166 pfd_8_0.F_b.n2 pfd_8_0.F_b.n0 417.574
R2167 pfd_8_0.F_b.n2 pfd_8_0.F_b.n1 244.716
R2168 pfd_8_0.F_b.n0 pfd_8_0.F_b.t4 228.148
R2169 pfd_8_0.F_b.t1 pfd_8_0.F_b.n2 221.411
R2170 pfd_8_0.F_b.n1 pfd_8_0.F_b.t0 24.0005
R2171 pfd_8_0.F_b.n1 pfd_8_0.F_b.t2 24.0005
R2172 a_1390_640.t0 a_1390_640.t1 39.4005
R2173 a_490_640.t0 a_490_640.t1 39.4005
R2174 charge_pump_cell_6_0.UP_b.n0 charge_pump_cell_6_0.UP_b.t1 0.00505063
R2175 charge_pump_cell_6_0.UP_b charge_pump_cell_6_0.UP_b.n0 12.0576
R2176 charge_pump_cell_6_0.UP_b.n0 charge_pump_cell_6_0.UP_b.t0 323.788
R2177 a_490_1400.t0 a_490_1400.t1 39.4005
R2178 pfd_8_0.Reset.n1 pfd_8_0.Reset.t3 562.333
R2179 pfd_8_0.Reset.n2 pfd_8_0.Reset.n1 480.45
R2180 pfd_8_0.Reset.n0 pfd_8_0.Reset.t4 417.733
R2181 pfd_8_0.Reset.n0 pfd_8_0.Reset.t5 369.534
R2182 pfd_8_0.Reset.n3 pfd_8_0.Reset.n2 328.733
R2183 pfd_8_0.Reset.t1 pfd_8_0.Reset.n3 288.37
R2184 pfd_8_0.Reset.n1 pfd_8_0.Reset.t2 224.934
R2185 pfd_8_0.Reset.n3 pfd_8_0.Reset.t0 177.577
R2186 pfd_8_0.Reset.n2 pfd_8_0.Reset.n0 176.733
R2187 charge_pump_cell_6_0.DOWN charge_pump_cell_6_0.DOWN.t0 12.0533
R2188 a_1870_190.t1 a_1870_190.n2 500.086
R2189 a_1870_190.n1 a_1870_190.n0 473.334
R2190 a_1870_190.n0 a_1870_190.t2 465.933
R2191 a_1870_190.t1 a_1870_190.n2 461.389
R2192 a_1870_190.n0 a_1870_190.t3 321.334
R2193 a_1870_190.n1 a_1870_190.t0 177.577
R2194 a_1870_190.n2 a_1870_190.n1 48.3898
R2195 a_n30_640.t0 a_n30_640.t1 39.4005
R2196 F_VCO.n0 F_VCO.t0 514.134
R2197 F_VCO.n0 F_VCO.t1 273.134
R2198 F_VCO F_VCO.n0 216.9
C0 pfd_8_0.QB pfd_8_0.QA 0.074487f
C1 I_IN charge_pump_cell_6_0.DOWN 0.010902f
C2 opamp_cell_4_0.p_bias VDDA 2.86573f
C3 VDDA pfd_8_0.DOWN_input 0.221393f
C4 opamp_cell_4_0.p_bias opamp_cell_4_0.VIN+ 0.098414f
C5 opamp_cell_4_0.VIN+ pfd_8_0.DOWN_input 0.072856f
C6 pfd_8_0.QA_b pfd_8_0.QA 0.422694f
C7 F_REF pfd_8_0.QA 0.056f
C8 charge_pump_cell_6_0.UP_b VDDA 0.396833f
C9 charge_pump_cell_6_0.UP_b opamp_cell_4_0.VIN+ 0.011697f
C10 V_OUT opamp_cell_4_0.p_bias 0.041726f
C11 pfd_8_0.QB_b F_VCO 0.039516f
C12 V_OUT pfd_8_0.DOWN_input 0.389513f
C13 I_IN VDDA 0.591539f
C14 VDDA F_VCO 0.12889f
C15 opamp_cell_4_0.p_bias opamp_cell_4_0.VIN- 0.010861f
C16 pfd_8_0.QB F_VCO 0.058558f
C17 I_IN opamp_cell_4_0.VIN+ 0.17405f
C18 charge_pump_cell_6_0.UP_b V_OUT 0.805699f
C19 V_OUT charge_pump_cell_6_0.DOWN 0.033524f
C20 pfd_8_0.QB_b VDDA 0.511838f
C21 pfd_8_0.QB pfd_8_0.QB_b 0.388258f
C22 pfd_8_0.QB VDDA 2.7499f
C23 VDDA opamp_cell_4_0.VIN+ 0.924492f
C24 charge_pump_cell_6_0.UP_b opamp_cell_4_0.p_bias 0.041967f
C25 pfd_8_0.QA_b VDDA 0.52066f
C26 VDDA F_REF 0.098433f
C27 V_OUT VDDA 0.793021f
C28 charge_pump_cell_6_0.DOWN pfd_8_0.DOWN_input 0.200808f
C29 V_OUT opamp_cell_4_0.VIN+ 1.07111f
C30 VDDA opamp_cell_4_0.VIN- 0.171047f
C31 I_IN pfd_8_0.DOWN_input 0.943218f
C32 opamp_cell_4_0.VIN+ opamp_cell_4_0.VIN- 0.133176f
C33 charge_pump_cell_6_0.UP_b charge_pump_cell_6_0.DOWN 0.049574f
C34 pfd_8_0.QA_b F_REF 0.027208f
C35 VDDA pfd_8_0.QA 0.550605f
C36 F_VCO GNDA 0.389374f
C37 I_IN GNDA 3.03352f
C38 V_OUT GNDA 24.114231f
C39 F_REF GNDA 0.277742f
C40 VDDA GNDA 44.36703f
C41 charge_pump_cell_6_0.DOWN GNDA 2.95069f
C42 pfd_8_0.DOWN_input GNDA 3.10504f
C43 pfd_8_0.QB_b GNDA 1.05311f
C44 pfd_8_0.QB GNDA 1.307381f
C45 pfd_8_0.QA GNDA 3.10102f
C46 pfd_8_0.QA_b GNDA 1.05138f
C47 charge_pump_cell_6_0.UP_b GNDA 5.40697f
C48 opamp_cell_4_0.VIN+ GNDA 2.9096f
C49 opamp_cell_4_0.VIN- GNDA 1.24398f
C50 opamp_cell_4_0.p_bias GNDA 3.947561f
C51 loop_filter_2_0.R1_C1.t1 GNDA 2.39887f
C52 pfd_8_0.QB.t7 GNDA 0.066708f
C53 pfd_8_0.QB.t8 GNDA 0.031333f
C54 pfd_8_0.QB.n0 GNDA 0.096363f
C55 pfd_8_0.QB.t3 GNDA 0.066708f
C56 pfd_8_0.QB.t4 GNDA 0.100569f
C57 pfd_8_0.QB.n1 GNDA 1.20598f
C58 pfd_8_0.QB.t5 GNDA 0.067367f
C59 pfd_8_0.QB.t6 GNDA 0.029539f
C60 pfd_8_0.QB.n2 GNDA 0.170164f
C61 pfd_8_0.QB.t1 GNDA 0.14186f
C62 pfd_8_0.QB.t0 GNDA 0.026953f
C63 pfd_8_0.QB.t2 GNDA 0.026953f
C64 pfd_8_0.QB.n3 GNDA 0.143916f
C65 pfd_8_0.QB.n4 GNDA 0.255686f
C66 pfd_8_0.QB.n5 GNDA 0.218372f
C67 V_OUT.n2 GNDA 0.013414f
C68 V_OUT.n4 GNDA 0.010429f
C69 V_OUT.t7 GNDA 5.06829f
C70 V_OUT.n6 GNDA 0.112288f
C71 V_OUT.n7 GNDA 0.06102f
C72 opamp_cell_4_0.p_bias.t0 GNDA 1.66267f
C73 opamp_cell_4_0.p_bias.t2 GNDA 0.019693f
C74 opamp_cell_4_0.p_bias.t6 GNDA 0.019693f
C75 opamp_cell_4_0.p_bias.n0 GNDA 0.054067f
C76 opamp_cell_4_0.p_bias.t8 GNDA 0.019693f
C77 opamp_cell_4_0.p_bias.t4 GNDA 0.019693f
C78 opamp_cell_4_0.p_bias.n1 GNDA 0.054067f
C79 opamp_cell_4_0.p_bias.n2 GNDA 0.068502f
C80 opamp_cell_4_0.p_bias.t1 GNDA 0.054353f
C81 opamp_cell_4_0.p_bias.t3 GNDA 0.054353f
C82 opamp_cell_4_0.p_bias.t7 GNDA 0.054353f
C83 opamp_cell_4_0.p_bias.t11 GNDA 0.054353f
C84 opamp_cell_4_0.p_bias.t9 GNDA 0.074733f
C85 opamp_cell_4_0.p_bias.n3 GNDA 0.04185f
C86 opamp_cell_4_0.p_bias.n4 GNDA 0.029697f
C87 opamp_cell_4_0.p_bias.n5 GNDA 0.012761f
C88 opamp_cell_4_0.p_bias.n6 GNDA 0.029697f
C89 opamp_cell_4_0.p_bias.n7 GNDA 0.029697f
C90 opamp_cell_4_0.p_bias.t5 GNDA 0.054353f
C91 opamp_cell_4_0.p_bias.t12 GNDA 0.054353f
C92 opamp_cell_4_0.p_bias.t10 GNDA 0.074733f
C93 opamp_cell_4_0.p_bias.n8 GNDA 0.04185f
C94 opamp_cell_4_0.p_bias.n9 GNDA 0.029697f
C95 opamp_cell_4_0.p_bias.n10 GNDA 0.012761f
C96 opamp_cell_4_0.p_bias.n11 GNDA 0.120625f
C97 opamp_cell_4_0.VIN+.t8 GNDA 0.023149f
C98 opamp_cell_4_0.VIN+.t7 GNDA 0.016337f
C99 opamp_cell_4_0.VIN+.n0 GNDA 0.042889f
C100 opamp_cell_4_0.VIN+.t9 GNDA 0.014474f
C101 opamp_cell_4_0.VIN+.n1 GNDA 0.038113f
C102 opamp_cell_4_0.VIN+.n2 GNDA 0.297842f
C103 opamp_cell_4_0.VIN+.t2 GNDA 0.039604f
C104 opamp_cell_4_0.VIN+.t1 GNDA 0.039604f
C105 opamp_cell_4_0.VIN+.n3 GNDA 0.097602f
C106 opamp_cell_4_0.VIN+.t5 GNDA 0.039604f
C107 opamp_cell_4_0.VIN+.t0 GNDA 0.039604f
C108 opamp_cell_4_0.VIN+.n4 GNDA 0.265157f
C109 opamp_cell_4_0.VIN+.n5 GNDA 0.416646f
C110 opamp_cell_4_0.VIN+.t4 GNDA 0.039604f
C111 opamp_cell_4_0.VIN+.t3 GNDA 0.039604f
C112 opamp_cell_4_0.VIN+.n6 GNDA 0.097602f
C113 opamp_cell_4_0.VIN+.n7 GNDA 0.468809f
C114 pfd_8_0.UP_input.t16 GNDA 3.21937f
C115 pfd_8_0.UP_input.n2 GNDA 0.032389f
C116 pfd_8_0.UP_input.n3 GNDA 0.028023f
C117 pfd_8_0.UP_input.n4 GNDA 0.01708f
C118 pfd_8_0.UP_input.t20 GNDA 0.018899f
C119 pfd_8_0.UP_input.t15 GNDA 0.032499f
C120 pfd_8_0.UP_input.t11 GNDA 0.015109f
C121 pfd_8_0.UP_input.t8 GNDA 0.036635f
C122 pfd_8_0.UP_input.n5 GNDA 0.044925f
C123 pfd_8_0.UP_input.t3 GNDA 0.033269f
C124 pfd_8_0.UP_input.n6 GNDA 0.157493f
C125 pfd_8_0.UP_input.n7 GNDA 0.033703f
C126 pfd_8_0.UP_input.n8 GNDA 0.01708f
C127 pfd_8_0.UP_input.t14 GNDA 0.018899f
C128 pfd_8_0.UP_input.n9 GNDA 0.022781f
C129 pfd_8_0.UP_input.n10 GNDA 0.022781f
C130 pfd_8_0.UP_input.t17 GNDA 0.032499f
C131 pfd_8_0.UP_input.n11 GNDA 0.033125f
C132 pfd_8_0.UP_input.t18 GNDA 4.68775f
C133 pfd_8_0.UP_input.n12 GNDA 0.010188f
C134 pfd_8_0.UP_input.n13 GNDA 0.0132f
C135 pfd_8_0.UP_input.n14 GNDA 0.043547f
C136 pfd_8_0.UP_input.n15 GNDA 0.028715f
C137 pfd_8_0.UP_input.n16 GNDA 0.017667f
C138 pfd_8_0.UP_input.t13 GNDA 0.018899f
C139 pfd_8_0.UP_input.t21 GNDA 0.043264f
C140 pfd_8_0.UP_input.n17 GNDA 0.022781f
C141 pfd_8_0.UP_input.t22 GNDA 0.018899f
C142 pfd_8_0.UP_input.n18 GNDA 0.022781f
C143 pfd_8_0.UP_input.n19 GNDA 0.022781f
C144 pfd_8_0.UP_input.t19 GNDA 0.031081f
C145 pfd_8_0.UP_input.n20 GNDA 0.021568f
C146 pfd_8_0.UP_input.t9 GNDA 0.040417f
C147 pfd_8_0.UP_input.t12 GNDA 0.012763f
C148 pfd_8_0.UP_input.n21 GNDA 0.051561f
C149 pfd_8_0.UP_input.n22 GNDA 0.272518f
C150 pfd_8_0.UP_input.n23 GNDA 0.160077f
C151 VDDA.n1 GNDA 0.011281f
C152 VDDA.n2 GNDA 0.011281f
C153 VDDA.n16 GNDA 0.011281f
C154 VDDA.t59 GNDA 0.047758f
C155 VDDA.t45 GNDA 0.01732f
C156 VDDA.n24 GNDA 0.018969f
C157 VDDA.t31 GNDA 0.047758f
C158 VDDA.n31 GNDA 0.011281f
C159 VDDA.n34 GNDA 0.010259f
C160 VDDA.n35 GNDA 0.011281f
C161 VDDA.n41 GNDA 0.043944f
C162 VDDA.n43 GNDA 0.010271f
C163 VDDA.n44 GNDA 0.017118f
C164 VDDA.t12 GNDA 0.160962f
C165 VDDA.n50 GNDA 0.017118f
C166 VDDA.n51 GNDA 0.017118f
C167 VDDA.n53 GNDA 0.010366f
C168 VDDA.n54 GNDA 0.010271f
C169 VDDA.n57 GNDA 0.010271f
C170 VDDA.n58 GNDA 0.012107f
C171 VDDA.n67 GNDA 0.014937f
C172 VDDA.n70 GNDA 0.014937f
C173 VDDA.n73 GNDA 0.014937f
C174 VDDA.n76 GNDA 0.014937f
C175 VDDA.n79 GNDA 0.015944f
C176 VDDA.n81 GNDA 0.014937f
C177 VDDA.n83 GNDA 0.012338f
C178 VDDA.t118 GNDA 0.010226f
C179 VDDA.t111 GNDA 0.013084f
C180 VDDA.n87 GNDA 0.078421f
C181 VDDA.t110 GNDA 0.192072f
C182 VDDA.t27 GNDA 0.097171f
C183 VDDA.t20 GNDA 0.097171f
C184 VDDA.t29 GNDA 0.097171f
C185 VDDA.t83 GNDA 0.097171f
C186 VDDA.t116 GNDA 0.110251f
C187 VDDA.n90 GNDA 0.012338f
C188 VDDA.t97 GNDA 0.010226f
C189 VDDA.n92 GNDA 0.021462f
C190 VDDA.t98 GNDA 0.028263f
C191 VDDA.n97 GNDA 0.021397f
C192 VDDA.n98 GNDA 0.010209f
C193 VDDA.n99 GNDA 0.010271f
C194 VDDA.n102 GNDA 0.010271f
C195 VDDA.n104 GNDA 0.010271f
C196 VDDA.n107 GNDA 0.155099f
C197 VDDA.t89 GNDA 0.074747f
C198 VDDA.t99 GNDA 0.048585f
C199 VDDA.t87 GNDA 0.057929f
C200 VDDA.t88 GNDA 0.065403f
C201 VDDA.t67 GNDA 0.048585f
C202 VDDA.t43 GNDA 0.074747f
C203 VDDA.t61 GNDA 0.048585f
C204 VDDA.t14 GNDA 0.054191f
C205 VDDA.t90 GNDA 0.069141f
C206 VDDA.t75 GNDA 0.095302f
C207 VDDA.t79 GNDA 0.100908f
C208 VDDA.n108 GNDA 0.08054f
C209 VDDA.t77 GNDA 0.061666f
C210 VDDA.t95 GNDA 0.061666f
C211 VDDA.t56 GNDA 0.061666f
C212 VDDA.t73 GNDA 0.048585f
C213 VDDA.t81 GNDA 0.074747f
C214 VDDA.t63 GNDA 0.048585f
C215 VDDA.t52 GNDA 0.057929f
C216 VDDA.t50 GNDA 0.065403f
C217 VDDA.t46 GNDA 0.048585f
C218 VDDA.t92 GNDA 0.074747f
C219 VDDA.t103 GNDA 0.061666f
C220 VDDA.t93 GNDA 0.013084f
C221 VDDA.n110 GNDA 0.012338f
C222 VDDA.n112 GNDA 0.025501f
C223 VDDA.n113 GNDA 0.08055f
C224 VDDA.t102 GNDA 0.028842f
C225 VDDA.t104 GNDA 0.014265f
C226 VDDA.n116 GNDA 0.021397f
C227 VDDA.n117 GNDA 0.010209f
C228 VDDA.n119 GNDA 0.010271f
C229 VDDA.n120 GNDA 0.010271f
C230 VDDA.n122 GNDA 0.010271f
C231 VDDA.n123 GNDA 0.020153f
C232 VDDA.n125 GNDA 0.059797f
C233 VDDA.n126 GNDA 0.071197f
C234 VDDA.n127 GNDA 0.021462f
C235 VDDA.n129 GNDA 0.012338f
C236 VDDA.n130 GNDA 0.01766f
C237 VDDA.n131 GNDA 0.051309f
C238 VDDA.n132 GNDA 0.051555f
C239 VDDA.n140 GNDA 0.049996f
C240 VDDA.n147 GNDA 0.049996f
C241 VDDA.n154 GNDA 0.049996f
C242 VDDA.n161 GNDA 0.049996f
C243 VDDA.n171 GNDA 0.033572f
C244 VDDA.n175 GNDA 0.017118f
C245 VDDA.n176 GNDA 0.010271f
C246 VDDA.t106 GNDA 0.071152f
C247 VDDA.n182 GNDA 0.015976f
C248 VDDA.n185 GNDA 0.015976f
C249 VDDA.n188 GNDA 0.016498f
C250 VDDA.n189 GNDA 0.023215f
C251 VDDA.n191 GNDA 0.016498f
C252 VDDA.n192 GNDA 0.023215f
C253 VDDA.n211 GNDA 0.016498f
C254 VDDA.n214 GNDA 0.016498f
C255 VDDA.n216 GNDA 0.014676f
C256 VDDA.t112 GNDA 0.028441f
C257 VDDA.n220 GNDA 0.011186f
C258 VDDA.n222 GNDA 0.010271f
C259 VDDA.t71 GNDA 0.072807f
C260 VDDA.t10 GNDA 0.072807f
C261 VDDA.t0 GNDA 0.072807f
C262 VDDA.t8 GNDA 0.072807f
C263 VDDA.t113 GNDA 0.071152f
C264 VDDA.n225 GNDA 0.064533f
C265 VDDA.n228 GNDA 0.010271f
C266 VDDA.n229 GNDA 0.010364f
C267 VDDA.n230 GNDA 0.017118f
C268 VDDA.t114 GNDA 0.011412f
C269 VDDA.n231 GNDA 0.016498f
C270 VDDA.n232 GNDA 0.023509f
C271 VDDA.n239 GNDA 0.022074f
C272 VDDA.n246 GNDA 0.023215f
C273 VDDA.n254 GNDA 0.023215f
C274 VDDA.n255 GNDA 0.016498f
C275 VDDA.t121 GNDA 0.011412f
C276 VDDA.n256 GNDA 0.017118f
C277 VDDA.t105 GNDA 0.026837f
C278 VDDA.t119 GNDA 0.026837f
C279 VDDA.n258 GNDA 0.01209f
C280 VDDA.n259 GNDA 0.020603f
C281 VDDA.n260 GNDA 0.017118f
C282 VDDA.n261 GNDA 0.01941f
C283 VDDA.n263 GNDA 0.069497f
C284 VDDA.t120 GNDA 0.071152f
C285 VDDA.t48 GNDA 0.072807f
C286 VDDA.t69 GNDA 0.072807f
C287 VDDA.t25 GNDA 0.072807f
C288 VDDA.t54 GNDA 0.072807f
C289 VDDA.t123 GNDA 0.071152f
C290 VDDA.n264 GNDA 0.010366f
C291 VDDA.n266 GNDA 0.010271f
C292 VDDA.n269 GNDA 0.064533f
C293 VDDA.n271 GNDA 0.011486f
C294 VDDA.t122 GNDA 0.028441f
C295 VDDA.n279 GNDA 0.023362f
C296 VDDA.n280 GNDA 0.244464f
C297 VDDA.n281 GNDA 0.04381f
C298 VDDA.n282 GNDA 0.010271f
C299 VDDA.n283 GNDA 0.017118f
C300 VDDA.t37 GNDA 0.168037f
C301 VDDA.t7 GNDA 0.182188f
C302 VDDA.n287 GNDA 0.010271f
C303 VDDA.n288 GNDA 0.010366f
C304 VDDA.n290 GNDA 0.137968f
C305 VDDA.n292 GNDA 0.012107f
C306 VDDA.n307 GNDA 0.012107f
C307 VDDA.n309 GNDA 0.010271f
C308 VDDA.n311 GNDA 0.010271f
C309 VDDA.n312 GNDA 0.010366f
C310 VDDA.n314 GNDA 0.137968f
C311 VDDA.t85 GNDA 0.137968f
C312 VDDA.t65 GNDA 0.047758f
C313 VDDA.t32 GNDA 0.012035f
C314 VDDA.n322 GNDA 0.011114f
C315 VDDA.n327 GNDA 0.068984f
C316 VDDA.t42 GNDA 0.012035f
C317 VDDA.n333 GNDA 0.011114f
C318 VDDA.n335 GNDA 0.068984f
C319 VDDA.t16 GNDA 0.047758f
C320 VDDA.t41 GNDA 0.047758f
C321 VDDA.t17 GNDA 0.012035f
C322 VDDA.n338 GNDA 0.010062f
C323 VDDA.n343 GNDA 0.097285f
C324 VDDA.n346 GNDA 0.017118f
C325 VDDA.n347 GNDA 0.010366f
C326 VDDA.n349 GNDA 0.010271f
C327 VDDA.n351 GNDA 0.010271f
C328 VDDA.n352 GNDA 0.012107f
C329 VDDA.n355 GNDA 0.017118f
C330 VDDA.n356 GNDA 0.012107f
C331 VDDA.n358 GNDA 0.010271f
C332 VDDA.n360 GNDA 0.010271f
C333 VDDA.n361 GNDA 0.010366f
C334 VDDA.n363 GNDA 0.150349f
C335 VDDA.t2 GNDA 0.137968f
C336 VDDA.n366 GNDA 0.010271f
C337 VDDA.n367 GNDA 0.010366f
C338 VDDA.n369 GNDA 0.137968f
C339 VDDA.n371 GNDA 0.012107f
C340 VDDA.n399 GNDA 0.011281f
C341 VDDA.t66 GNDA 0.012035f
C342 VDDA.n403 GNDA 0.011114f
C343 VDDA.n405 GNDA 0.068984f
C344 VDDA.t60 GNDA 0.012035f
C345 VDDA.n406 GNDA 0.011114f
C346 VDDA.t23 GNDA 0.042452f
C347 VDDA.t44 GNDA 0.04422f
C348 VDDA.n411 GNDA 0.068984f
C349 VDDA.n413 GNDA 0.011281f
C350 VDDA.n421 GNDA 0.011068f
C351 VDDA.t24 GNDA 0.011976f
C352 VDDA.n425 GNDA 0.011114f
C353 VDDA.n427 GNDA 0.093747f
C354 VDDA.t18 GNDA 0.012035f
C355 VDDA.n434 GNDA 0.011114f
C356 VDDA.t6 GNDA 0.012035f
C357 VDDA.n444 GNDA 0.011114f
C358 VDDA.n446 GNDA 0.10436f
C359 VDDA.t5 GNDA 0.086672f
C360 VDDA.t4 GNDA 0.183957f
C361 VDDA.t58 GNDA 0.183957f
C362 VDDA.t35 GNDA 0.086672f
C363 VDDA.n450 GNDA 0.012553f
C364 VDDA.n451 GNDA 0.015024f
C365 VDDA.n454 GNDA 0.012553f
C366 VDDA.t40 GNDA 0.012041f
C367 VDDA.n457 GNDA 0.012514f
C368 VDDA.n461 GNDA 0.012553f
C369 VDDA.n462 GNDA 0.012514f
C370 VDDA.n465 GNDA 0.012553f
C371 VDDA.t128 GNDA 0.012041f
C372 VDDA.n468 GNDA 0.015024f
C373 VDDA.n470 GNDA 0.095516f
C374 VDDA.t39 GNDA 0.086672f
C375 VDDA.t19 GNDA 0.183957f
C376 VDDA.t22 GNDA 0.183957f
C377 VDDA.t33 GNDA 0.086672f
C378 VDDA.t127 GNDA 0.012035f
C379 VDDA.n471 GNDA 0.011114f
C380 VDDA.t34 GNDA 0.012035f
C381 VDDA.n481 GNDA 0.011114f
C382 VDDA.n483 GNDA 0.097285f
C383 VDDA.n485 GNDA 0.011281f
C384 a_5970_4630.t11 GNDA 0.030769f
C385 a_5970_4630.n0 GNDA 0.124795f
C386 a_5970_4630.t0 GNDA 0.020325f
C387 a_5970_4630.t1 GNDA 0.020325f
C388 a_5970_4630.t7 GNDA 0.020325f
C389 a_5970_4630.n1 GNDA 0.044943f
C390 a_5970_4630.t6 GNDA 0.020325f
C391 a_5970_4630.t9 GNDA 0.020325f
C392 a_5970_4630.n2 GNDA 0.044943f
C393 a_5970_4630.t10 GNDA 0.077457f
C394 a_5970_4630.t8 GNDA 0.030769f
C395 a_5970_4630.n3 GNDA 0.097952f
C396 a_5970_4630.n4 GNDA 0.087903f
C397 a_5970_4630.n5 GNDA 0.089425f
C398 a_5970_4630.t2 GNDA 0.050813f
C399 a_5970_4630.t4 GNDA 0.050813f
C400 a_5970_4630.n6 GNDA 0.295522f
C401 a_5970_4630.t3 GNDA 0.050813f
C402 a_5970_4630.t5 GNDA 0.050813f
C403 a_5970_4630.n7 GNDA 0.144587f
C404 a_5970_4630.n8 GNDA 0.360746f
C405 a_5970_4630.n9 GNDA 0.13437f
C406 a_5970_4630.n10 GNDA 0.085474f
C407 a_5970_4630.n11 GNDA 0.045257f
C408 a_5970_4630.t12 GNDA 0.100208f
.ends

