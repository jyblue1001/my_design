magic
tech sky130A
magscale 1 2
timestamp 1740116149
<< nwell >>
rect 6010 3750 9450 4140
rect 6010 1800 9290 3750
rect 4680 1220 6110 1800
rect 6530 1280 6650 1310
<< poly >>
rect 5290 5580 6010 5600
rect 5290 5540 5310 5580
rect 5350 5570 6010 5580
rect 5350 5540 5370 5570
rect 5290 5520 5370 5540
rect -260 1920 -180 1950
rect 4360 1890 4440 1910
rect 4360 1860 4380 1890
rect 4180 1850 4380 1860
rect 4420 1850 4440 1890
rect 4180 1830 4440 1850
rect 6060 1300 6140 1320
rect 6060 1260 6080 1300
rect 6120 1280 6140 1300
rect 6530 1280 6650 1310
rect 6120 1260 6650 1280
rect 6060 1240 6650 1260
rect 8050 1280 8130 1300
rect 8050 1240 8070 1280
rect 8110 1240 8130 1280
rect 8050 1220 8130 1240
rect 8490 910 8570 930
rect 8490 870 8510 910
rect 8550 870 8570 910
rect 8490 850 8570 870
rect -260 490 -180 520
rect 4150 170 4230 190
rect 4150 130 4170 170
rect 4210 130 4230 170
rect 4150 110 4230 130
<< polycont >>
rect 5310 5540 5350 5580
rect 4380 1850 4420 1890
rect 6080 1260 6120 1300
rect 8070 1240 8110 1280
rect 8510 870 8550 910
rect 4170 130 4210 170
<< locali >>
rect 5730 6090 5830 6120
rect 5730 6050 5760 6090
rect 5800 6050 5830 6090
rect 5730 6020 5830 6050
rect 5410 5620 5490 5640
rect 5290 5580 5370 5600
rect 5290 5540 5310 5580
rect 5350 5540 5370 5580
rect 5290 3150 5370 5540
rect 5290 3110 5310 3150
rect 5350 3110 5370 3150
rect 5290 3090 5370 3110
rect 5410 5580 5430 5620
rect 5470 5580 5490 5620
rect 4760 2420 4860 2440
rect 4710 2380 4780 2420
rect 4760 2360 4780 2380
rect 4840 2360 4860 2420
rect 4760 2340 4860 2360
rect 4080 2260 5360 2300
rect 4080 2210 4120 2260
rect 4360 1890 4440 1910
rect 4360 1850 4380 1890
rect 4420 1850 4440 1890
rect 4360 1830 4440 1850
rect 4600 1890 4680 1910
rect 4600 1850 4620 1890
rect 4660 1850 4680 1890
rect 4600 1830 4680 1850
rect 5320 1320 5360 2260
rect 5280 1300 5360 1320
rect 5000 1250 5100 1280
rect 5000 1240 5030 1250
rect 4740 1200 4800 1240
rect 4840 1200 4900 1240
rect 4940 1210 5030 1240
rect 5070 1210 5100 1250
rect 5280 1260 5300 1300
rect 5340 1260 5360 1300
rect 5280 1240 5360 1260
rect 4940 1200 5100 1210
rect 5000 1180 5100 1200
rect 5410 1170 5490 5580
rect 9820 5510 11900 5550
rect 5730 4900 5830 4930
rect 5730 4860 5760 4900
rect 5800 4860 5830 4900
rect 5730 4830 5830 4860
rect 11860 3250 11900 5510
rect 5570 3210 11900 3250
rect 5570 1320 5610 3210
rect 5820 1950 5920 1980
rect 5820 1910 5850 1950
rect 5890 1910 5920 1950
rect 5820 1880 5920 1910
rect 5530 1300 5610 1320
rect 5530 1260 5550 1300
rect 5590 1280 5610 1300
rect 6060 1300 6140 1320
rect 6060 1280 6080 1300
rect 5590 1260 6080 1280
rect 6120 1260 6140 1300
rect 5530 1240 6140 1260
rect 8050 1280 8130 1300
rect 6660 1170 6740 1250
rect 8050 1240 8070 1280
rect 8110 1240 8130 1280
rect 8050 1220 8130 1240
rect 4080 1080 4400 1120
rect 5410 1090 6740 1170
rect 9250 1110 9330 1130
rect 4080 1010 4120 1080
rect 4360 1040 4400 1080
rect 9250 1070 9270 1110
rect 9310 1070 9330 1110
rect 9250 1050 9330 1070
rect 4360 1000 5800 1040
rect 5300 910 5380 930
rect 5300 870 5320 910
rect 5360 870 5380 910
rect 5300 850 5380 870
rect 8490 910 8570 930
rect 8490 870 8510 910
rect 8550 870 8570 910
rect 8490 850 8570 870
rect 5300 530 5340 850
rect 4640 490 5340 530
rect 5820 270 5920 300
rect 5820 230 5850 270
rect 5890 230 5920 270
rect 5820 200 5920 230
rect 4150 170 4230 190
rect 4150 130 4170 170
rect 4210 130 4230 170
rect 4150 110 4230 130
rect 4760 80 4860 100
rect 4760 60 4780 80
rect 4710 20 4780 60
rect 4840 20 4860 80
rect 4760 0 4860 20
rect 4760 -250 4860 -230
rect 4760 -310 4780 -250
rect 4840 -270 4860 -250
rect 4840 -310 4920 -270
rect 4960 -310 5020 -270
rect 5060 -310 5120 -270
rect 5160 -310 5220 -270
rect 5260 -310 5320 -270
rect 5360 -310 5420 -270
rect 5460 -310 5520 -270
rect 5560 -310 5620 -270
rect 5660 -310 5720 -270
rect 5760 -310 5820 -270
rect 5860 -310 5920 -270
rect 5960 -310 6020 -270
rect 6060 -310 6120 -270
rect 6160 -310 6220 -270
rect 6260 -310 6320 -270
rect 6360 -310 6420 -270
rect 6460 -310 6520 -270
rect 6560 -310 6620 -270
rect 6660 -310 6720 -270
rect 6760 -310 6820 -270
rect 6860 -310 6920 -270
rect 6960 -310 7020 -270
rect 7060 -310 7120 -270
rect 7160 -310 7220 -270
rect 7260 -310 7320 -270
rect 7360 -310 7420 -270
rect 7460 -310 7520 -270
rect 7560 -310 7620 -270
rect 7660 -310 7720 -270
rect 7760 -310 7820 -270
rect 7860 -310 7920 -270
rect 7960 -310 8020 -270
rect 8060 -310 8120 -270
rect 8160 -310 8220 -270
rect 8260 -310 8320 -270
rect 8360 -310 8420 -270
rect 8460 -310 8520 -270
rect 8560 -310 8620 -270
rect 8660 -310 8720 -270
rect 8760 -310 8820 -270
rect 8860 -310 8920 -270
rect 8960 -310 9020 -270
rect 9060 -310 9120 -270
rect 9160 -310 9220 -270
rect 9260 -310 9320 -270
rect 9360 -310 9420 -270
rect 9460 -310 9520 -270
rect 9560 -310 9620 -270
rect 9660 -310 9720 -270
rect 9760 -310 9820 -270
rect 9860 -310 9920 -270
rect 9960 -310 10020 -270
rect 10060 -310 10120 -270
rect 10160 -310 10220 -270
rect 10260 -310 10320 -270
rect 10360 -310 10420 -270
rect 10460 -310 10520 -270
rect 10560 -310 10620 -270
rect 10660 -310 10720 -270
rect 10760 -310 10820 -270
rect 10860 -310 10920 -270
rect 10960 -310 11020 -270
rect 11060 -310 11120 -270
rect 11160 -310 11220 -270
rect 11260 -310 11320 -270
rect 11360 -310 11420 -270
rect 11460 -310 11520 -270
rect 11560 -310 11620 -270
rect 11660 -310 11720 -270
rect 11760 -310 11820 -270
rect 11860 -310 11920 -270
rect 11960 -310 12020 -270
rect 12060 -310 12120 -270
rect 12160 -310 12220 -270
rect 12260 -310 12320 -270
rect 12360 -310 12420 -270
rect 12460 -310 12520 -270
rect 12560 -310 12620 -270
rect 12660 -310 12720 -270
rect 12760 -310 12820 -270
rect 12860 -310 12920 -270
rect 12960 -310 13020 -270
rect 13060 -310 13120 -270
rect 13160 -310 13220 -270
rect 13260 -310 13320 -270
rect 13360 -310 13420 -270
rect 13460 -310 13520 -270
rect 13560 -310 13620 -270
rect 13660 -310 13720 -270
rect 13760 -310 13820 -270
rect 13860 -310 13920 -270
rect 13960 -310 14020 -270
rect 14060 -310 14120 -270
rect 14160 -310 14220 -270
rect 14260 -310 14320 -270
rect 14360 -310 14420 -270
rect 14460 -310 14520 -270
rect 14560 -310 14620 -270
rect 14660 -310 14720 -270
rect 14760 -310 14820 -270
rect 14860 -310 14920 -270
rect 14960 -310 15020 -270
rect 15060 -310 15120 -270
rect 15160 -310 15220 -270
rect 15260 -310 15320 -270
rect 15360 -310 15420 -270
rect 15460 -310 15520 -270
rect 15560 -310 15620 -270
rect 15660 -310 15720 -270
rect 15760 -310 15820 -270
rect 15860 -310 15920 -270
rect 15960 -310 16020 -270
rect 16060 -310 16120 -270
rect 16160 -310 16220 -270
rect 16260 -310 16320 -270
rect 16360 -310 16420 -270
rect 16460 -310 16520 -270
rect 16560 -310 16620 -270
rect 16660 -310 16720 -270
rect 16760 -310 16820 -270
rect 16860 -310 16920 -270
rect 16960 -310 17020 -270
rect 4760 -330 4860 -310
<< viali >>
rect 5760 6050 5800 6090
rect 5310 3110 5350 3150
rect 5430 5580 5470 5620
rect 4780 2360 4840 2420
rect 4380 1850 4420 1890
rect 4620 1850 4660 1890
rect 4700 1200 4740 1240
rect 4800 1200 4840 1240
rect 4900 1200 4940 1240
rect 5030 1210 5070 1250
rect 5300 1260 5340 1300
rect 5760 4860 5800 4900
rect 5850 1910 5890 1950
rect 5550 1260 5590 1300
rect 8070 1240 8110 1280
rect 9270 1070 9310 1110
rect 5320 870 5360 910
rect 8510 870 8550 910
rect 5850 230 5890 270
rect 4170 130 4210 170
rect 4780 20 4840 80
rect 4780 -310 4840 -250
rect 4920 -310 4960 -270
rect 5020 -310 5060 -270
rect 5120 -310 5160 -270
rect 5220 -310 5260 -270
rect 5320 -310 5360 -270
rect 5420 -310 5460 -270
rect 5520 -310 5560 -270
rect 5620 -310 5660 -270
rect 5720 -310 5760 -270
rect 5820 -310 5860 -270
rect 5920 -310 5960 -270
rect 6020 -310 6060 -270
rect 6120 -310 6160 -270
rect 6220 -310 6260 -270
rect 6320 -310 6360 -270
rect 6420 -310 6460 -270
rect 6520 -310 6560 -270
rect 6620 -310 6660 -270
rect 6720 -310 6760 -270
rect 6820 -310 6860 -270
rect 6920 -310 6960 -270
rect 7020 -310 7060 -270
rect 7120 -310 7160 -270
rect 7220 -310 7260 -270
rect 7320 -310 7360 -270
rect 7420 -310 7460 -270
rect 7520 -310 7560 -270
rect 7620 -310 7660 -270
rect 7720 -310 7760 -270
rect 7820 -310 7860 -270
rect 7920 -310 7960 -270
rect 8020 -310 8060 -270
rect 8120 -310 8160 -270
rect 8220 -310 8260 -270
rect 8320 -310 8360 -270
rect 8420 -310 8460 -270
rect 8520 -310 8560 -270
rect 8620 -310 8660 -270
rect 8720 -310 8760 -270
rect 8820 -310 8860 -270
rect 8920 -310 8960 -270
rect 9020 -310 9060 -270
rect 9120 -310 9160 -270
rect 9220 -310 9260 -270
rect 9320 -310 9360 -270
rect 9420 -310 9460 -270
rect 9520 -310 9560 -270
rect 9620 -310 9660 -270
rect 9720 -310 9760 -270
rect 9820 -310 9860 -270
rect 9920 -310 9960 -270
rect 10020 -310 10060 -270
rect 10120 -310 10160 -270
rect 10220 -310 10260 -270
rect 10320 -310 10360 -270
rect 10420 -310 10460 -270
rect 10520 -310 10560 -270
rect 10620 -310 10660 -270
rect 10720 -310 10760 -270
rect 10820 -310 10860 -270
rect 10920 -310 10960 -270
rect 11020 -310 11060 -270
rect 11120 -310 11160 -270
rect 11220 -310 11260 -270
rect 11320 -310 11360 -270
rect 11420 -310 11460 -270
rect 11520 -310 11560 -270
rect 11620 -310 11660 -270
rect 11720 -310 11760 -270
rect 11820 -310 11860 -270
rect 11920 -310 11960 -270
rect 12020 -310 12060 -270
rect 12120 -310 12160 -270
rect 12220 -310 12260 -270
rect 12320 -310 12360 -270
rect 12420 -310 12460 -270
rect 12520 -310 12560 -270
rect 12620 -310 12660 -270
rect 12720 -310 12760 -270
rect 12820 -310 12860 -270
rect 12920 -310 12960 -270
rect 13020 -310 13060 -270
rect 13120 -310 13160 -270
rect 13220 -310 13260 -270
rect 13320 -310 13360 -270
rect 13420 -310 13460 -270
rect 13520 -310 13560 -270
rect 13620 -310 13660 -270
rect 13720 -310 13760 -270
rect 13820 -310 13860 -270
rect 13920 -310 13960 -270
rect 14020 -310 14060 -270
rect 14120 -310 14160 -270
rect 14220 -310 14260 -270
rect 14320 -310 14360 -270
rect 14420 -310 14460 -270
rect 14520 -310 14560 -270
rect 14620 -310 14660 -270
rect 14720 -310 14760 -270
rect 14820 -310 14860 -270
rect 14920 -310 14960 -270
rect 15020 -310 15060 -270
rect 15120 -310 15160 -270
rect 15220 -310 15260 -270
rect 15320 -310 15360 -270
rect 15420 -310 15460 -270
rect 15520 -310 15560 -270
rect 15620 -310 15660 -270
rect 15720 -310 15760 -270
rect 15820 -310 15860 -270
rect 15920 -310 15960 -270
rect 16020 -310 16060 -270
rect 16120 -310 16160 -270
rect 16220 -310 16260 -270
rect 16320 -310 16360 -270
rect 16420 -310 16460 -270
rect 16520 -310 16560 -270
rect 16620 -310 16660 -270
rect 16720 -310 16760 -270
rect 16820 -310 16860 -270
rect 16920 -310 16960 -270
<< metal1 >>
rect 5730 6100 5830 6120
rect 5730 6040 5750 6100
rect 5810 6040 5830 6100
rect 5730 6020 5830 6040
rect 5410 5620 6010 5640
rect 5410 5580 5430 5620
rect 5470 5610 6010 5620
rect 5470 5580 5490 5610
rect 5410 5560 5490 5580
rect 5730 4910 5830 4930
rect 5730 4850 5750 4910
rect 5810 4850 5830 4910
rect 5730 4830 5830 4850
rect 5290 3150 11300 3170
rect 5290 3110 5310 3150
rect 5350 3110 11300 3150
rect 5290 3090 11300 3110
rect 5040 2890 5820 3000
rect 4710 2420 4860 2440
rect 4710 2360 4780 2420
rect 4840 2360 4860 2420
rect 4760 2340 4860 2360
rect 5040 2040 5130 2890
rect 4360 1960 5130 2040
rect 5820 1960 5920 1980
rect 4360 1890 4440 1960
rect 4360 1850 4380 1890
rect 4420 1850 4440 1890
rect 4360 1830 4440 1850
rect 4600 1890 4680 1910
rect 4600 1850 4620 1890
rect 4660 1870 4680 1890
rect 5820 1900 5840 1960
rect 5900 1900 5920 1960
rect 5820 1880 5920 1900
rect 4660 1850 5190 1870
rect 4600 1830 5190 1850
rect 5000 1260 5100 1280
rect -280 1180 -230 1260
rect 4710 1240 5020 1260
rect 4740 1200 4800 1240
rect 4840 1200 4900 1240
rect 4940 1200 5020 1240
rect 5080 1200 5100 1260
rect 4710 1180 5100 1200
rect 5150 1210 5190 1830
rect 5280 1300 5360 1320
rect 5280 1260 5300 1300
rect 5340 1280 5360 1300
rect 5530 1300 5610 1320
rect 5530 1280 5550 1300
rect 5340 1260 5550 1280
rect 5590 1260 5610 1300
rect 5280 1240 5610 1260
rect 8050 1280 8130 1300
rect 8050 1240 8070 1280
rect 8110 1240 8130 1280
rect 8050 1210 8130 1240
rect 5150 1170 8130 1210
rect 11220 1130 11300 3090
rect 9250 1110 11300 1130
rect 9250 1070 9270 1110
rect 9310 1070 11300 1110
rect 9250 1050 11300 1070
rect 5300 910 8570 930
rect 5300 870 5320 910
rect 5360 890 8510 910
rect 5360 870 5380 890
rect 5300 850 5380 870
rect 8490 870 8510 890
rect 8550 870 8570 910
rect 8490 850 8570 870
rect 5820 280 5920 300
rect 5820 220 5840 280
rect 5900 220 5920 280
rect 5820 200 5920 220
rect 4150 170 5550 190
rect 4150 130 4170 170
rect 4210 150 5550 170
rect 4210 130 4230 150
rect 4150 110 4230 130
rect 4760 80 4860 100
rect 4710 20 4780 80
rect 4840 20 4860 80
rect 4710 0 4860 20
rect 5470 10 5550 150
rect 5470 -100 5820 10
rect 11220 0 11300 1050
rect 11220 -80 13220 0
rect 4760 -250 4860 -230
rect 4760 -310 4780 -250
rect 4840 -270 17020 -250
rect 4840 -310 4920 -270
rect 4960 -310 5020 -270
rect 5060 -310 5120 -270
rect 5160 -310 5220 -270
rect 5260 -310 5320 -270
rect 5360 -310 5420 -270
rect 5460 -310 5520 -270
rect 5560 -310 5620 -270
rect 5660 -310 5720 -270
rect 5760 -310 5820 -270
rect 5860 -310 5920 -270
rect 5960 -310 6020 -270
rect 6060 -310 6120 -270
rect 6160 -310 6220 -270
rect 6260 -310 6320 -270
rect 6360 -310 6420 -270
rect 6460 -310 6520 -270
rect 6560 -310 6620 -270
rect 6660 -310 6720 -270
rect 6760 -310 6820 -270
rect 6860 -310 6920 -270
rect 6960 -310 7020 -270
rect 7060 -310 7120 -270
rect 7160 -310 7220 -270
rect 7260 -310 7320 -270
rect 7360 -310 7420 -270
rect 7460 -310 7520 -270
rect 7560 -310 7620 -270
rect 7660 -310 7720 -270
rect 7760 -310 7820 -270
rect 7860 -310 7920 -270
rect 7960 -310 8020 -270
rect 8060 -310 8120 -270
rect 8160 -310 8220 -270
rect 8260 -310 8320 -270
rect 8360 -310 8420 -270
rect 8460 -310 8520 -270
rect 8560 -310 8620 -270
rect 8660 -310 8720 -270
rect 8760 -310 8820 -270
rect 8860 -310 8920 -270
rect 8960 -310 9020 -270
rect 9060 -310 9120 -270
rect 9160 -310 9220 -270
rect 9260 -310 9320 -270
rect 9360 -310 9420 -270
rect 9460 -310 9520 -270
rect 9560 -310 9620 -270
rect 9660 -310 9720 -270
rect 9760 -310 9820 -270
rect 9860 -310 9920 -270
rect 9960 -310 10020 -270
rect 10060 -310 10120 -270
rect 10160 -310 10220 -270
rect 10260 -310 10320 -270
rect 10360 -310 10420 -270
rect 10460 -310 10520 -270
rect 10560 -310 10620 -270
rect 10660 -310 10720 -270
rect 10760 -310 10820 -270
rect 10860 -310 10920 -270
rect 10960 -310 11020 -270
rect 11060 -310 11120 -270
rect 11160 -310 11220 -270
rect 11260 -310 11320 -270
rect 11360 -310 11420 -270
rect 11460 -310 11520 -270
rect 11560 -310 11620 -270
rect 11660 -310 11720 -270
rect 11760 -310 11820 -270
rect 11860 -310 11920 -270
rect 11960 -310 12020 -270
rect 12060 -310 12120 -270
rect 12160 -310 12220 -270
rect 12260 -310 12320 -270
rect 12360 -310 12420 -270
rect 12460 -310 12520 -270
rect 12560 -310 12620 -270
rect 12660 -310 12720 -270
rect 12760 -310 12820 -270
rect 12860 -310 12920 -270
rect 12960 -310 13020 -270
rect 13060 -310 13120 -270
rect 13160 -310 13220 -270
rect 13260 -310 13320 -270
rect 13360 -310 13420 -270
rect 13460 -310 13520 -270
rect 13560 -310 13620 -270
rect 13660 -310 13720 -270
rect 13760 -310 13820 -270
rect 13860 -310 13920 -270
rect 13960 -310 14020 -270
rect 14060 -310 14120 -270
rect 14160 -310 14220 -270
rect 14260 -310 14320 -270
rect 14360 -310 14420 -270
rect 14460 -310 14520 -270
rect 14560 -310 14620 -270
rect 14660 -310 14720 -270
rect 14760 -310 14820 -270
rect 14860 -310 14920 -270
rect 14960 -310 15020 -270
rect 15060 -310 15120 -270
rect 15160 -310 15220 -270
rect 15260 -310 15320 -270
rect 15360 -310 15420 -270
rect 15460 -310 15520 -270
rect 15560 -310 15620 -270
rect 15660 -310 15720 -270
rect 15760 -310 15820 -270
rect 15860 -310 15920 -270
rect 15960 -310 16020 -270
rect 16060 -310 16120 -270
rect 16160 -310 16220 -270
rect 16260 -310 16320 -270
rect 16360 -310 16420 -270
rect 16460 -310 16520 -270
rect 16560 -310 16620 -270
rect 16660 -310 16720 -270
rect 16760 -310 16820 -270
rect 16860 -310 16920 -270
rect 16960 -310 17020 -270
rect 4760 -330 17020 -310
<< via1 >>
rect 5750 6090 5810 6100
rect 5750 6050 5760 6090
rect 5760 6050 5800 6090
rect 5800 6050 5810 6090
rect 5750 6040 5810 6050
rect 5750 4900 5810 4910
rect 5750 4860 5760 4900
rect 5760 4860 5800 4900
rect 5800 4860 5810 4900
rect 5750 4850 5810 4860
rect 4780 2360 4840 2420
rect 5840 1950 5900 1960
rect 5840 1910 5850 1950
rect 5850 1910 5890 1950
rect 5890 1910 5900 1950
rect 5840 1900 5900 1910
rect 5020 1250 5080 1260
rect 5020 1210 5030 1250
rect 5030 1210 5070 1250
rect 5070 1210 5080 1250
rect 5020 1200 5080 1210
rect 5840 270 5900 280
rect 5840 230 5850 270
rect 5850 230 5890 270
rect 5890 230 5900 270
rect 5840 220 5900 230
rect 4780 20 4840 80
rect 4780 -310 4840 -250
<< metal2 >>
rect 5730 6100 5830 6120
rect 5730 6040 5750 6100
rect 5810 6040 5830 6100
rect 5730 6020 5830 6040
rect 5730 4910 5830 4930
rect 5730 4850 5750 4910
rect 5810 4850 5830 4910
rect 5730 4830 5830 4850
rect 4760 2420 4860 2440
rect 4760 2360 4780 2420
rect 4840 2360 4860 2420
rect 4760 2340 4860 2360
rect 5820 1960 5920 1980
rect 5820 1900 5840 1960
rect 5900 1900 5920 1960
rect 5820 1880 5920 1900
rect 5000 1260 5100 1280
rect 5000 1200 5020 1260
rect 5080 1200 5100 1260
rect 5000 1180 5100 1200
rect 5820 280 5920 300
rect 5820 220 5840 280
rect 5900 220 5920 280
rect 5820 200 5920 220
rect 4760 80 4860 100
rect 4760 20 4780 80
rect 4840 20 4860 80
rect 4760 0 4860 20
rect 4760 -250 4860 -230
rect 4760 -310 4780 -250
rect 4840 -310 4860 -250
rect 4760 -330 4860 -310
<< via2 >>
rect 5750 6040 5810 6100
rect 5750 4850 5810 4910
rect 4780 2360 4840 2420
rect 5840 1900 5900 1960
rect 5020 1200 5080 1260
rect 5840 220 5900 280
rect 4780 20 4840 80
rect 4780 -310 4840 -250
<< metal3 >>
rect 4760 6110 5830 6120
rect 4760 6030 4770 6110
rect 4850 6100 5830 6110
rect 4850 6040 5750 6100
rect 5810 6040 5830 6100
rect 4850 6030 5830 6040
rect 4760 6020 5830 6030
rect 5000 4920 5830 4930
rect 5000 4840 5010 4920
rect 5090 4910 5830 4920
rect 5090 4850 5750 4910
rect 5810 4850 5830 4910
rect 5090 4840 5830 4850
rect 5000 4830 5830 4840
rect 4760 2430 4860 2440
rect 4760 2350 4770 2430
rect 4850 2350 4860 2430
rect 4760 2340 4860 2350
rect 5000 1970 5920 1980
rect 5000 1890 5010 1970
rect 5090 1960 5920 1970
rect 5090 1900 5840 1960
rect 5900 1900 5920 1960
rect 5090 1890 5920 1900
rect 5000 1880 5920 1890
rect 5000 1270 5100 1280
rect 5000 1190 5010 1270
rect 5090 1190 5100 1270
rect 5000 1180 5100 1190
rect 4760 290 5920 300
rect 4760 210 4770 290
rect 4850 280 5920 290
rect 4850 220 5840 280
rect 5900 220 5920 280
rect 4850 210 5920 220
rect 4760 200 5920 210
rect 4760 90 4860 100
rect 4760 10 4770 90
rect 4850 10 4860 90
rect 4760 0 4860 10
rect 4760 -240 4860 -230
rect 4760 -320 4770 -240
rect 4850 -320 4860 -240
rect 4760 -330 4860 -320
<< via3 >>
rect 4770 6030 4850 6110
rect 5010 4840 5090 4920
rect 4770 2420 4850 2430
rect 4770 2360 4780 2420
rect 4780 2360 4840 2420
rect 4840 2360 4850 2420
rect 4770 2350 4850 2360
rect 5010 1890 5090 1970
rect 5010 1260 5090 1270
rect 5010 1200 5020 1260
rect 5020 1200 5080 1260
rect 5080 1200 5090 1260
rect 5010 1190 5090 1200
rect 4770 210 4850 290
rect 4770 80 4850 90
rect 4770 20 4780 80
rect 4780 20 4840 80
rect 4840 20 4850 80
rect 4770 10 4850 20
rect 4770 -250 4850 -240
rect 4770 -310 4780 -250
rect 4780 -310 4840 -250
rect 4840 -310 4850 -250
rect 4770 -320 4850 -310
<< metal4 >>
rect 4760 6110 4860 6120
rect 4760 6030 4770 6110
rect 4850 6030 4860 6110
rect 4760 2430 4860 6030
rect 4760 2350 4770 2430
rect 4850 2350 4860 2430
rect -560 210 -460 310
rect 4760 290 4860 2350
rect 5000 4920 5100 4930
rect 5000 4840 5010 4920
rect 5090 4840 5100 4920
rect 5000 1970 5100 4840
rect 5000 1890 5010 1970
rect 5090 1890 5100 1970
rect 5000 1270 5100 1890
rect 5000 1190 5010 1270
rect 5090 1190 5100 1270
rect 5000 1180 5100 1190
rect 4760 210 4770 290
rect 4850 210 4860 290
rect 4760 90 4860 210
rect 4760 10 4770 90
rect 4850 10 4860 90
rect 4760 -240 4860 10
rect 4760 -320 4770 -240
rect 4850 -320 4860 -240
rect 4760 -330 4860 -320
use charge_pump_cell_6  charge_pump_cell_6_0
timestamp 1739811829
transform 1 0 -12390 0 1 -3210
box 18190 3110 23240 6210
use loop_filter_2  loop_filter_2_0
timestamp 1739812747
transform 1 0 10950 0 -1 580
box 2270 -11950 19440 660
use opamp_cell_4  opamp_cell_4_0
timestamp 1739772381
transform 1 0 -670 0 -1 9710
box 6220 1794 12730 6410
use pfd_8  pfd_8_0
timestamp 1739770731
transform 1 0 -1860 0 1 9310
box 1300 -9310 6580 -6870
use VCO_FD_magic  VCO_FD_magic_0
timestamp 1740073110
transform -1 0 10755 0 -1 -267
box 0 120 12940 2300
<< labels >>
flabel locali 5760 1020 5760 1020 5 FreeSans 800 0 0 -400 I_IN
port 6 s
flabel metal1 -280 1220 -280 1220 7 FreeSans 800 0 -400 0 VDDA
port 2 w
flabel metal4 -560 260 -560 260 7 FreeSans 800 0 -400 0 GNDA
port 3 w
flabel poly -260 500 -260 500 7 FreeSans 800 0 -400 0 F_VCO
port 5 w
flabel poly -260 1930 -260 1930 7 FreeSans 800 0 -400 0 F_REF
port 4 w
flabel metal1 11300 1090 11300 1090 3 FreeSans 800 0 400 0 V_OUT
port 1 e
<< end >>
