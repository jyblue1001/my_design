magic
tech sky130A
timestamp 1746683269
<< nwell >>
rect 2960 1960 4770 2820
<< pwell >>
rect -45 1685 130 1725
rect 3220 1560 4260 1660
<< nmos >>
rect 3260 1560 3320 1660
rect 3360 1560 3420 1660
rect 3460 1560 3520 1660
rect 3560 1560 3620 1660
rect 3660 1560 3720 1660
rect 3760 1560 3820 1660
rect 3860 1560 3920 1660
rect 3960 1560 4020 1660
rect 4060 1560 4120 1660
rect 4160 1560 4220 1660
rect 3280 985 3680 1385
rect 3800 985 4200 1385
rect 3230 755 4230 855
<< pmos >>
rect 3060 2400 3120 2800
rect 3160 2400 3220 2800
rect 3260 2400 3320 2800
rect 3360 2400 3420 2800
rect 3460 2400 3520 2800
rect 3560 2400 3620 2800
rect 3660 2400 3720 2800
rect 3760 2400 3820 2800
rect 3860 2400 3920 2800
rect 3960 2400 4020 2800
rect 4060 2400 4120 2800
rect 4160 2400 4220 2800
rect 4260 2400 4320 2800
rect 4360 2400 4420 2800
rect 3060 1980 3120 2180
rect 3160 1980 3220 2180
rect 3260 1980 3320 2180
rect 3360 1980 3420 2180
rect 3460 1980 3520 2180
rect 3560 1980 3620 2180
rect 3660 1980 3720 2180
rect 3760 1980 3820 2180
rect 3860 1980 3920 2180
rect 3960 1980 4020 2180
rect 4060 1980 4120 2180
rect 4160 1980 4220 2180
rect 4260 1980 4320 2180
rect 4360 1980 4420 2180
rect 4570 1980 4585 2180
rect 4695 1980 4710 2180
<< ndiff >>
rect 3220 1645 3260 1660
rect 3220 1625 3230 1645
rect 3250 1625 3260 1645
rect 3220 1595 3260 1625
rect 3220 1575 3230 1595
rect 3250 1575 3260 1595
rect 3220 1560 3260 1575
rect 3320 1645 3360 1660
rect 3320 1625 3330 1645
rect 3350 1625 3360 1645
rect 3320 1595 3360 1625
rect 3320 1575 3330 1595
rect 3350 1575 3360 1595
rect 3320 1560 3360 1575
rect 3420 1645 3460 1660
rect 3420 1625 3430 1645
rect 3450 1625 3460 1645
rect 3420 1595 3460 1625
rect 3420 1575 3430 1595
rect 3450 1575 3460 1595
rect 3420 1560 3460 1575
rect 3520 1645 3560 1660
rect 3520 1625 3530 1645
rect 3550 1625 3560 1645
rect 3520 1595 3560 1625
rect 3520 1575 3530 1595
rect 3550 1575 3560 1595
rect 3520 1560 3560 1575
rect 3620 1645 3660 1660
rect 3620 1625 3630 1645
rect 3650 1625 3660 1645
rect 3620 1595 3660 1625
rect 3620 1575 3630 1595
rect 3650 1575 3660 1595
rect 3620 1560 3660 1575
rect 3720 1645 3760 1660
rect 3720 1625 3730 1645
rect 3750 1625 3760 1645
rect 3720 1595 3760 1625
rect 3720 1575 3730 1595
rect 3750 1575 3760 1595
rect 3720 1560 3760 1575
rect 3820 1645 3860 1660
rect 3820 1625 3830 1645
rect 3850 1625 3860 1645
rect 3820 1595 3860 1625
rect 3820 1575 3830 1595
rect 3850 1575 3860 1595
rect 3820 1560 3860 1575
rect 3920 1645 3960 1660
rect 3920 1625 3930 1645
rect 3950 1625 3960 1645
rect 3920 1595 3960 1625
rect 3920 1575 3930 1595
rect 3950 1575 3960 1595
rect 3920 1560 3960 1575
rect 4020 1645 4060 1660
rect 4020 1625 4030 1645
rect 4050 1625 4060 1645
rect 4020 1595 4060 1625
rect 4020 1575 4030 1595
rect 4050 1575 4060 1595
rect 4020 1560 4060 1575
rect 4120 1645 4160 1660
rect 4120 1625 4130 1645
rect 4150 1625 4160 1645
rect 4120 1595 4160 1625
rect 4120 1575 4130 1595
rect 4150 1575 4160 1595
rect 4120 1560 4160 1575
rect 4220 1645 4260 1660
rect 4220 1625 4230 1645
rect 4250 1625 4260 1645
rect 4220 1595 4260 1625
rect 4220 1575 4230 1595
rect 4250 1575 4260 1595
rect 4220 1560 4260 1575
rect 3240 1370 3280 1385
rect 3240 1350 3250 1370
rect 3270 1350 3280 1370
rect 3240 1320 3280 1350
rect 3240 1300 3250 1320
rect 3270 1300 3280 1320
rect 3240 1270 3280 1300
rect 3240 1250 3250 1270
rect 3270 1250 3280 1270
rect 3240 1220 3280 1250
rect 3240 1200 3250 1220
rect 3270 1200 3280 1220
rect 3240 1170 3280 1200
rect 3240 1150 3250 1170
rect 3270 1150 3280 1170
rect 3240 1120 3280 1150
rect 3240 1100 3250 1120
rect 3270 1100 3280 1120
rect 3240 1070 3280 1100
rect 3240 1050 3250 1070
rect 3270 1050 3280 1070
rect 3240 1020 3280 1050
rect 3240 1000 3250 1020
rect 3270 1000 3280 1020
rect 3240 985 3280 1000
rect 3680 1370 3720 1385
rect 3760 1370 3800 1385
rect 3680 1350 3690 1370
rect 3710 1350 3720 1370
rect 3760 1350 3770 1370
rect 3790 1350 3800 1370
rect 3680 1320 3720 1350
rect 3760 1320 3800 1350
rect 3680 1300 3690 1320
rect 3710 1300 3720 1320
rect 3760 1300 3770 1320
rect 3790 1300 3800 1320
rect 3680 1270 3720 1300
rect 3760 1270 3800 1300
rect 3680 1250 3690 1270
rect 3710 1250 3720 1270
rect 3760 1250 3770 1270
rect 3790 1250 3800 1270
rect 3680 1220 3720 1250
rect 3760 1220 3800 1250
rect 3680 1200 3690 1220
rect 3710 1200 3720 1220
rect 3760 1200 3770 1220
rect 3790 1200 3800 1220
rect 3680 1170 3720 1200
rect 3760 1170 3800 1200
rect 3680 1150 3690 1170
rect 3710 1150 3720 1170
rect 3760 1150 3770 1170
rect 3790 1150 3800 1170
rect 3680 1120 3720 1150
rect 3760 1120 3800 1150
rect 3680 1100 3690 1120
rect 3710 1100 3720 1120
rect 3760 1100 3770 1120
rect 3790 1100 3800 1120
rect 3680 1070 3720 1100
rect 3760 1070 3800 1100
rect 3680 1050 3690 1070
rect 3710 1050 3720 1070
rect 3760 1050 3770 1070
rect 3790 1050 3800 1070
rect 3680 1020 3720 1050
rect 3760 1020 3800 1050
rect 3680 1000 3690 1020
rect 3710 1000 3720 1020
rect 3760 1000 3770 1020
rect 3790 1000 3800 1020
rect 3680 985 3720 1000
rect 3760 985 3800 1000
rect 4200 1370 4240 1385
rect 4200 1350 4210 1370
rect 4230 1350 4240 1370
rect 4200 1320 4240 1350
rect 4200 1300 4210 1320
rect 4230 1300 4240 1320
rect 4200 1270 4240 1300
rect 4200 1250 4210 1270
rect 4230 1250 4240 1270
rect 4200 1220 4240 1250
rect 4200 1200 4210 1220
rect 4230 1200 4240 1220
rect 4200 1170 4240 1200
rect 4200 1150 4210 1170
rect 4230 1150 4240 1170
rect 4200 1120 4240 1150
rect 4200 1100 4210 1120
rect 4230 1100 4240 1120
rect 4200 1070 4240 1100
rect 4200 1050 4210 1070
rect 4230 1050 4240 1070
rect 4200 1020 4240 1050
rect 4200 1000 4210 1020
rect 4230 1000 4240 1020
rect 4200 985 4240 1000
rect 3190 840 3230 855
rect 3190 820 3200 840
rect 3220 820 3230 840
rect 3190 790 3230 820
rect 3190 770 3200 790
rect 3220 770 3230 790
rect 3190 755 3230 770
rect 4230 840 4270 855
rect 4230 820 4240 840
rect 4260 820 4270 840
rect 4230 790 4270 820
rect 4230 770 4240 790
rect 4260 770 4270 790
rect 4230 755 4270 770
<< pdiff >>
rect 3020 2785 3060 2800
rect 3020 2765 3030 2785
rect 3050 2765 3060 2785
rect 3020 2735 3060 2765
rect 3020 2715 3030 2735
rect 3050 2715 3060 2735
rect 3020 2685 3060 2715
rect 3020 2665 3030 2685
rect 3050 2665 3060 2685
rect 3020 2635 3060 2665
rect 3020 2615 3030 2635
rect 3050 2615 3060 2635
rect 3020 2585 3060 2615
rect 3020 2565 3030 2585
rect 3050 2565 3060 2585
rect 3020 2535 3060 2565
rect 3020 2515 3030 2535
rect 3050 2515 3060 2535
rect 3020 2485 3060 2515
rect 3020 2465 3030 2485
rect 3050 2465 3060 2485
rect 3020 2435 3060 2465
rect 3020 2415 3030 2435
rect 3050 2415 3060 2435
rect 3020 2400 3060 2415
rect 3120 2785 3160 2800
rect 3120 2765 3130 2785
rect 3150 2765 3160 2785
rect 3120 2735 3160 2765
rect 3120 2715 3130 2735
rect 3150 2715 3160 2735
rect 3120 2685 3160 2715
rect 3120 2665 3130 2685
rect 3150 2665 3160 2685
rect 3120 2635 3160 2665
rect 3120 2615 3130 2635
rect 3150 2615 3160 2635
rect 3120 2585 3160 2615
rect 3120 2565 3130 2585
rect 3150 2565 3160 2585
rect 3120 2535 3160 2565
rect 3120 2515 3130 2535
rect 3150 2515 3160 2535
rect 3120 2485 3160 2515
rect 3120 2465 3130 2485
rect 3150 2465 3160 2485
rect 3120 2435 3160 2465
rect 3120 2415 3130 2435
rect 3150 2415 3160 2435
rect 3120 2400 3160 2415
rect 3220 2785 3260 2800
rect 3220 2765 3230 2785
rect 3250 2765 3260 2785
rect 3220 2735 3260 2765
rect 3220 2715 3230 2735
rect 3250 2715 3260 2735
rect 3220 2685 3260 2715
rect 3220 2665 3230 2685
rect 3250 2665 3260 2685
rect 3220 2635 3260 2665
rect 3220 2615 3230 2635
rect 3250 2615 3260 2635
rect 3220 2585 3260 2615
rect 3220 2565 3230 2585
rect 3250 2565 3260 2585
rect 3220 2535 3260 2565
rect 3220 2515 3230 2535
rect 3250 2515 3260 2535
rect 3220 2485 3260 2515
rect 3220 2465 3230 2485
rect 3250 2465 3260 2485
rect 3220 2435 3260 2465
rect 3220 2415 3230 2435
rect 3250 2415 3260 2435
rect 3220 2400 3260 2415
rect 3320 2785 3360 2800
rect 3320 2765 3330 2785
rect 3350 2765 3360 2785
rect 3320 2735 3360 2765
rect 3320 2715 3330 2735
rect 3350 2715 3360 2735
rect 3320 2685 3360 2715
rect 3320 2665 3330 2685
rect 3350 2665 3360 2685
rect 3320 2635 3360 2665
rect 3320 2615 3330 2635
rect 3350 2615 3360 2635
rect 3320 2585 3360 2615
rect 3320 2565 3330 2585
rect 3350 2565 3360 2585
rect 3320 2535 3360 2565
rect 3320 2515 3330 2535
rect 3350 2515 3360 2535
rect 3320 2485 3360 2515
rect 3320 2465 3330 2485
rect 3350 2465 3360 2485
rect 3320 2435 3360 2465
rect 3320 2415 3330 2435
rect 3350 2415 3360 2435
rect 3320 2400 3360 2415
rect 3420 2785 3460 2800
rect 3420 2765 3430 2785
rect 3450 2765 3460 2785
rect 3420 2735 3460 2765
rect 3420 2715 3430 2735
rect 3450 2715 3460 2735
rect 3420 2685 3460 2715
rect 3420 2665 3430 2685
rect 3450 2665 3460 2685
rect 3420 2635 3460 2665
rect 3420 2615 3430 2635
rect 3450 2615 3460 2635
rect 3420 2585 3460 2615
rect 3420 2565 3430 2585
rect 3450 2565 3460 2585
rect 3420 2535 3460 2565
rect 3420 2515 3430 2535
rect 3450 2515 3460 2535
rect 3420 2485 3460 2515
rect 3420 2465 3430 2485
rect 3450 2465 3460 2485
rect 3420 2435 3460 2465
rect 3420 2415 3430 2435
rect 3450 2415 3460 2435
rect 3420 2400 3460 2415
rect 3520 2785 3560 2800
rect 3520 2765 3530 2785
rect 3550 2765 3560 2785
rect 3520 2735 3560 2765
rect 3520 2715 3530 2735
rect 3550 2715 3560 2735
rect 3520 2685 3560 2715
rect 3520 2665 3530 2685
rect 3550 2665 3560 2685
rect 3520 2635 3560 2665
rect 3520 2615 3530 2635
rect 3550 2615 3560 2635
rect 3520 2585 3560 2615
rect 3520 2565 3530 2585
rect 3550 2565 3560 2585
rect 3520 2535 3560 2565
rect 3520 2515 3530 2535
rect 3550 2515 3560 2535
rect 3520 2485 3560 2515
rect 3520 2465 3530 2485
rect 3550 2465 3560 2485
rect 3520 2435 3560 2465
rect 3520 2415 3530 2435
rect 3550 2415 3560 2435
rect 3520 2400 3560 2415
rect 3620 2785 3660 2800
rect 3620 2765 3630 2785
rect 3650 2765 3660 2785
rect 3620 2735 3660 2765
rect 3620 2715 3630 2735
rect 3650 2715 3660 2735
rect 3620 2685 3660 2715
rect 3620 2665 3630 2685
rect 3650 2665 3660 2685
rect 3620 2635 3660 2665
rect 3620 2615 3630 2635
rect 3650 2615 3660 2635
rect 3620 2585 3660 2615
rect 3620 2565 3630 2585
rect 3650 2565 3660 2585
rect 3620 2535 3660 2565
rect 3620 2515 3630 2535
rect 3650 2515 3660 2535
rect 3620 2485 3660 2515
rect 3620 2465 3630 2485
rect 3650 2465 3660 2485
rect 3620 2435 3660 2465
rect 3620 2415 3630 2435
rect 3650 2415 3660 2435
rect 3620 2400 3660 2415
rect 3720 2785 3760 2800
rect 3720 2765 3730 2785
rect 3750 2765 3760 2785
rect 3720 2735 3760 2765
rect 3720 2715 3730 2735
rect 3750 2715 3760 2735
rect 3720 2685 3760 2715
rect 3720 2665 3730 2685
rect 3750 2665 3760 2685
rect 3720 2635 3760 2665
rect 3720 2615 3730 2635
rect 3750 2615 3760 2635
rect 3720 2585 3760 2615
rect 3720 2565 3730 2585
rect 3750 2565 3760 2585
rect 3720 2535 3760 2565
rect 3720 2515 3730 2535
rect 3750 2515 3760 2535
rect 3720 2485 3760 2515
rect 3720 2465 3730 2485
rect 3750 2465 3760 2485
rect 3720 2435 3760 2465
rect 3720 2415 3730 2435
rect 3750 2415 3760 2435
rect 3720 2400 3760 2415
rect 3820 2785 3860 2800
rect 3820 2765 3830 2785
rect 3850 2765 3860 2785
rect 3820 2735 3860 2765
rect 3820 2715 3830 2735
rect 3850 2715 3860 2735
rect 3820 2685 3860 2715
rect 3820 2665 3830 2685
rect 3850 2665 3860 2685
rect 3820 2635 3860 2665
rect 3820 2615 3830 2635
rect 3850 2615 3860 2635
rect 3820 2585 3860 2615
rect 3820 2565 3830 2585
rect 3850 2565 3860 2585
rect 3820 2535 3860 2565
rect 3820 2515 3830 2535
rect 3850 2515 3860 2535
rect 3820 2485 3860 2515
rect 3820 2465 3830 2485
rect 3850 2465 3860 2485
rect 3820 2435 3860 2465
rect 3820 2415 3830 2435
rect 3850 2415 3860 2435
rect 3820 2400 3860 2415
rect 3920 2785 3960 2800
rect 3920 2765 3930 2785
rect 3950 2765 3960 2785
rect 3920 2735 3960 2765
rect 3920 2715 3930 2735
rect 3950 2715 3960 2735
rect 3920 2685 3960 2715
rect 3920 2665 3930 2685
rect 3950 2665 3960 2685
rect 3920 2635 3960 2665
rect 3920 2615 3930 2635
rect 3950 2615 3960 2635
rect 3920 2585 3960 2615
rect 3920 2565 3930 2585
rect 3950 2565 3960 2585
rect 3920 2535 3960 2565
rect 3920 2515 3930 2535
rect 3950 2515 3960 2535
rect 3920 2485 3960 2515
rect 3920 2465 3930 2485
rect 3950 2465 3960 2485
rect 3920 2435 3960 2465
rect 3920 2415 3930 2435
rect 3950 2415 3960 2435
rect 3920 2400 3960 2415
rect 4020 2785 4060 2800
rect 4020 2765 4030 2785
rect 4050 2765 4060 2785
rect 4020 2735 4060 2765
rect 4020 2715 4030 2735
rect 4050 2715 4060 2735
rect 4020 2685 4060 2715
rect 4020 2665 4030 2685
rect 4050 2665 4060 2685
rect 4020 2635 4060 2665
rect 4020 2615 4030 2635
rect 4050 2615 4060 2635
rect 4020 2585 4060 2615
rect 4020 2565 4030 2585
rect 4050 2565 4060 2585
rect 4020 2535 4060 2565
rect 4020 2515 4030 2535
rect 4050 2515 4060 2535
rect 4020 2485 4060 2515
rect 4020 2465 4030 2485
rect 4050 2465 4060 2485
rect 4020 2435 4060 2465
rect 4020 2415 4030 2435
rect 4050 2415 4060 2435
rect 4020 2400 4060 2415
rect 4120 2785 4160 2800
rect 4120 2765 4130 2785
rect 4150 2765 4160 2785
rect 4120 2735 4160 2765
rect 4120 2715 4130 2735
rect 4150 2715 4160 2735
rect 4120 2685 4160 2715
rect 4120 2665 4130 2685
rect 4150 2665 4160 2685
rect 4120 2635 4160 2665
rect 4120 2615 4130 2635
rect 4150 2615 4160 2635
rect 4120 2585 4160 2615
rect 4120 2565 4130 2585
rect 4150 2565 4160 2585
rect 4120 2535 4160 2565
rect 4120 2515 4130 2535
rect 4150 2515 4160 2535
rect 4120 2485 4160 2515
rect 4120 2465 4130 2485
rect 4150 2465 4160 2485
rect 4120 2435 4160 2465
rect 4120 2415 4130 2435
rect 4150 2415 4160 2435
rect 4120 2400 4160 2415
rect 4220 2785 4260 2800
rect 4220 2765 4230 2785
rect 4250 2765 4260 2785
rect 4220 2735 4260 2765
rect 4220 2715 4230 2735
rect 4250 2715 4260 2735
rect 4220 2685 4260 2715
rect 4220 2665 4230 2685
rect 4250 2665 4260 2685
rect 4220 2635 4260 2665
rect 4220 2615 4230 2635
rect 4250 2615 4260 2635
rect 4220 2585 4260 2615
rect 4220 2565 4230 2585
rect 4250 2565 4260 2585
rect 4220 2535 4260 2565
rect 4220 2515 4230 2535
rect 4250 2515 4260 2535
rect 4220 2485 4260 2515
rect 4220 2465 4230 2485
rect 4250 2465 4260 2485
rect 4220 2435 4260 2465
rect 4220 2415 4230 2435
rect 4250 2415 4260 2435
rect 4220 2400 4260 2415
rect 4320 2785 4360 2800
rect 4320 2765 4330 2785
rect 4350 2765 4360 2785
rect 4320 2735 4360 2765
rect 4320 2715 4330 2735
rect 4350 2715 4360 2735
rect 4320 2685 4360 2715
rect 4320 2665 4330 2685
rect 4350 2665 4360 2685
rect 4320 2635 4360 2665
rect 4320 2615 4330 2635
rect 4350 2615 4360 2635
rect 4320 2585 4360 2615
rect 4320 2565 4330 2585
rect 4350 2565 4360 2585
rect 4320 2535 4360 2565
rect 4320 2515 4330 2535
rect 4350 2515 4360 2535
rect 4320 2485 4360 2515
rect 4320 2465 4330 2485
rect 4350 2465 4360 2485
rect 4320 2435 4360 2465
rect 4320 2415 4330 2435
rect 4350 2415 4360 2435
rect 4320 2400 4360 2415
rect 4420 2785 4460 2800
rect 4420 2765 4430 2785
rect 4450 2765 4460 2785
rect 4420 2735 4460 2765
rect 4420 2715 4430 2735
rect 4450 2715 4460 2735
rect 4420 2685 4460 2715
rect 4420 2665 4430 2685
rect 4450 2665 4460 2685
rect 4420 2635 4460 2665
rect 4420 2615 4430 2635
rect 4450 2615 4460 2635
rect 4420 2585 4460 2615
rect 4420 2565 4430 2585
rect 4450 2565 4460 2585
rect 4420 2535 4460 2565
rect 4420 2515 4430 2535
rect 4450 2515 4460 2535
rect 4420 2485 4460 2515
rect 4420 2465 4430 2485
rect 4450 2465 4460 2485
rect 4420 2435 4460 2465
rect 4420 2415 4430 2435
rect 4450 2415 4460 2435
rect 4420 2400 4460 2415
rect 3020 2165 3060 2180
rect 3020 2145 3030 2165
rect 3050 2145 3060 2165
rect 3020 2115 3060 2145
rect 3020 2095 3030 2115
rect 3050 2095 3060 2115
rect 3020 2065 3060 2095
rect 3020 2045 3030 2065
rect 3050 2045 3060 2065
rect 3020 2015 3060 2045
rect 3020 1995 3030 2015
rect 3050 1995 3060 2015
rect 3020 1980 3060 1995
rect 3120 2165 3160 2180
rect 3120 2145 3130 2165
rect 3150 2145 3160 2165
rect 3120 2115 3160 2145
rect 3120 2095 3130 2115
rect 3150 2095 3160 2115
rect 3120 2065 3160 2095
rect 3120 2045 3130 2065
rect 3150 2045 3160 2065
rect 3120 2015 3160 2045
rect 3120 1995 3130 2015
rect 3150 1995 3160 2015
rect 3120 1980 3160 1995
rect 3220 2165 3260 2180
rect 3220 2145 3230 2165
rect 3250 2145 3260 2165
rect 3220 2115 3260 2145
rect 3220 2095 3230 2115
rect 3250 2095 3260 2115
rect 3220 2065 3260 2095
rect 3220 2045 3230 2065
rect 3250 2045 3260 2065
rect 3220 2015 3260 2045
rect 3220 1995 3230 2015
rect 3250 1995 3260 2015
rect 3220 1980 3260 1995
rect 3320 2165 3360 2180
rect 3320 2145 3330 2165
rect 3350 2145 3360 2165
rect 3320 2115 3360 2145
rect 3320 2095 3330 2115
rect 3350 2095 3360 2115
rect 3320 2065 3360 2095
rect 3320 2045 3330 2065
rect 3350 2045 3360 2065
rect 3320 2015 3360 2045
rect 3320 1995 3330 2015
rect 3350 1995 3360 2015
rect 3320 1980 3360 1995
rect 3420 2165 3460 2180
rect 3420 2145 3430 2165
rect 3450 2145 3460 2165
rect 3420 2115 3460 2145
rect 3420 2095 3430 2115
rect 3450 2095 3460 2115
rect 3420 2065 3460 2095
rect 3420 2045 3430 2065
rect 3450 2045 3460 2065
rect 3420 2015 3460 2045
rect 3420 1995 3430 2015
rect 3450 1995 3460 2015
rect 3420 1980 3460 1995
rect 3520 2165 3560 2180
rect 3520 2145 3530 2165
rect 3550 2145 3560 2165
rect 3520 2115 3560 2145
rect 3520 2095 3530 2115
rect 3550 2095 3560 2115
rect 3520 2065 3560 2095
rect 3520 2045 3530 2065
rect 3550 2045 3560 2065
rect 3520 2015 3560 2045
rect 3520 1995 3530 2015
rect 3550 1995 3560 2015
rect 3520 1980 3560 1995
rect 3620 2165 3660 2180
rect 3620 2145 3630 2165
rect 3650 2145 3660 2165
rect 3620 2115 3660 2145
rect 3620 2095 3630 2115
rect 3650 2095 3660 2115
rect 3620 2065 3660 2095
rect 3620 2045 3630 2065
rect 3650 2045 3660 2065
rect 3620 2015 3660 2045
rect 3620 1995 3630 2015
rect 3650 1995 3660 2015
rect 3620 1980 3660 1995
rect 3720 2165 3760 2180
rect 3720 2145 3730 2165
rect 3750 2145 3760 2165
rect 3720 2115 3760 2145
rect 3720 2095 3730 2115
rect 3750 2095 3760 2115
rect 3720 2065 3760 2095
rect 3720 2045 3730 2065
rect 3750 2045 3760 2065
rect 3720 2015 3760 2045
rect 3720 1995 3730 2015
rect 3750 1995 3760 2015
rect 3720 1980 3760 1995
rect 3820 2165 3860 2180
rect 3820 2145 3830 2165
rect 3850 2145 3860 2165
rect 3820 2115 3860 2145
rect 3820 2095 3830 2115
rect 3850 2095 3860 2115
rect 3820 2065 3860 2095
rect 3820 2045 3830 2065
rect 3850 2045 3860 2065
rect 3820 2015 3860 2045
rect 3820 1995 3830 2015
rect 3850 1995 3860 2015
rect 3820 1980 3860 1995
rect 3920 2165 3960 2180
rect 3920 2145 3930 2165
rect 3950 2145 3960 2165
rect 3920 2115 3960 2145
rect 3920 2095 3930 2115
rect 3950 2095 3960 2115
rect 3920 2065 3960 2095
rect 3920 2045 3930 2065
rect 3950 2045 3960 2065
rect 3920 2015 3960 2045
rect 3920 1995 3930 2015
rect 3950 1995 3960 2015
rect 3920 1980 3960 1995
rect 4020 2165 4060 2180
rect 4020 2145 4030 2165
rect 4050 2145 4060 2165
rect 4020 2115 4060 2145
rect 4020 2095 4030 2115
rect 4050 2095 4060 2115
rect 4020 2065 4060 2095
rect 4020 2045 4030 2065
rect 4050 2045 4060 2065
rect 4020 2015 4060 2045
rect 4020 1995 4030 2015
rect 4050 1995 4060 2015
rect 4020 1980 4060 1995
rect 4120 2165 4160 2180
rect 4120 2145 4130 2165
rect 4150 2145 4160 2165
rect 4120 2115 4160 2145
rect 4120 2095 4130 2115
rect 4150 2095 4160 2115
rect 4120 2065 4160 2095
rect 4120 2045 4130 2065
rect 4150 2045 4160 2065
rect 4120 2015 4160 2045
rect 4120 1995 4130 2015
rect 4150 1995 4160 2015
rect 4120 1980 4160 1995
rect 4220 2165 4260 2180
rect 4220 2145 4230 2165
rect 4250 2145 4260 2165
rect 4220 2115 4260 2145
rect 4220 2095 4230 2115
rect 4250 2095 4260 2115
rect 4220 2065 4260 2095
rect 4220 2045 4230 2065
rect 4250 2045 4260 2065
rect 4220 2015 4260 2045
rect 4220 1995 4230 2015
rect 4250 1995 4260 2015
rect 4220 1980 4260 1995
rect 4320 2165 4360 2180
rect 4320 2145 4330 2165
rect 4350 2145 4360 2165
rect 4320 2115 4360 2145
rect 4320 2095 4330 2115
rect 4350 2095 4360 2115
rect 4320 2065 4360 2095
rect 4320 2045 4330 2065
rect 4350 2045 4360 2065
rect 4320 2015 4360 2045
rect 4320 1995 4330 2015
rect 4350 1995 4360 2015
rect 4320 1980 4360 1995
rect 4420 2165 4460 2180
rect 4420 2145 4430 2165
rect 4450 2145 4460 2165
rect 4420 2115 4460 2145
rect 4420 2095 4430 2115
rect 4450 2095 4460 2115
rect 4420 2065 4460 2095
rect 4420 2045 4430 2065
rect 4450 2045 4460 2065
rect 4420 2015 4460 2045
rect 4420 1995 4430 2015
rect 4450 1995 4460 2015
rect 4420 1980 4460 1995
rect 4530 2165 4570 2180
rect 4530 2145 4540 2165
rect 4560 2145 4570 2165
rect 4530 2115 4570 2145
rect 4530 2095 4540 2115
rect 4560 2095 4570 2115
rect 4530 2065 4570 2095
rect 4530 2045 4540 2065
rect 4560 2045 4570 2065
rect 4530 2015 4570 2045
rect 4530 1995 4540 2015
rect 4560 1995 4570 2015
rect 4530 1980 4570 1995
rect 4585 2165 4625 2180
rect 4585 2145 4595 2165
rect 4615 2145 4625 2165
rect 4585 2115 4625 2145
rect 4585 2095 4595 2115
rect 4615 2095 4625 2115
rect 4585 2065 4625 2095
rect 4585 2045 4595 2065
rect 4615 2045 4625 2065
rect 4585 2015 4625 2045
rect 4585 1995 4595 2015
rect 4615 1995 4625 2015
rect 4585 1980 4625 1995
rect 4655 2165 4695 2180
rect 4655 2145 4665 2165
rect 4685 2145 4695 2165
rect 4655 2115 4695 2145
rect 4655 2095 4665 2115
rect 4685 2095 4695 2115
rect 4655 2065 4695 2095
rect 4655 2045 4665 2065
rect 4685 2045 4695 2065
rect 4655 2015 4695 2045
rect 4655 1995 4665 2015
rect 4685 1995 4695 2015
rect 4655 1980 4695 1995
rect 4710 2165 4750 2180
rect 4710 2145 4720 2165
rect 4740 2145 4750 2165
rect 4710 2115 4750 2145
rect 4710 2095 4720 2115
rect 4740 2095 4750 2115
rect 4710 2065 4750 2095
rect 4710 2045 4720 2065
rect 4740 2045 4750 2065
rect 4710 2015 4750 2045
rect 4710 1995 4720 2015
rect 4740 1995 4750 2015
rect 4710 1980 4750 1995
<< ndiffc >>
rect 3230 1625 3250 1645
rect 3230 1575 3250 1595
rect 3330 1625 3350 1645
rect 3330 1575 3350 1595
rect 3430 1625 3450 1645
rect 3430 1575 3450 1595
rect 3530 1625 3550 1645
rect 3530 1575 3550 1595
rect 3630 1625 3650 1645
rect 3630 1575 3650 1595
rect 3730 1625 3750 1645
rect 3730 1575 3750 1595
rect 3830 1625 3850 1645
rect 3830 1575 3850 1595
rect 3930 1625 3950 1645
rect 3930 1575 3950 1595
rect 4030 1625 4050 1645
rect 4030 1575 4050 1595
rect 4130 1625 4150 1645
rect 4130 1575 4150 1595
rect 4230 1625 4250 1645
rect 4230 1575 4250 1595
rect 3250 1350 3270 1370
rect 3250 1300 3270 1320
rect 3250 1250 3270 1270
rect 3250 1200 3270 1220
rect 3250 1150 3270 1170
rect 3250 1100 3270 1120
rect 3250 1050 3270 1070
rect 3250 1000 3270 1020
rect 3690 1350 3710 1370
rect 3770 1350 3790 1370
rect 3690 1300 3710 1320
rect 3770 1300 3790 1320
rect 3690 1250 3710 1270
rect 3770 1250 3790 1270
rect 3690 1200 3710 1220
rect 3770 1200 3790 1220
rect 3690 1150 3710 1170
rect 3770 1150 3790 1170
rect 3690 1100 3710 1120
rect 3770 1100 3790 1120
rect 3690 1050 3710 1070
rect 3770 1050 3790 1070
rect 3690 1000 3710 1020
rect 3770 1000 3790 1020
rect 4210 1350 4230 1370
rect 4210 1300 4230 1320
rect 4210 1250 4230 1270
rect 4210 1200 4230 1220
rect 4210 1150 4230 1170
rect 4210 1100 4230 1120
rect 4210 1050 4230 1070
rect 4210 1000 4230 1020
rect 3200 820 3220 840
rect 3200 770 3220 790
rect 4240 820 4260 840
rect 4240 770 4260 790
<< pdiffc >>
rect 3030 2765 3050 2785
rect 3030 2715 3050 2735
rect 3030 2665 3050 2685
rect 3030 2615 3050 2635
rect 3030 2565 3050 2585
rect 3030 2515 3050 2535
rect 3030 2465 3050 2485
rect 3030 2415 3050 2435
rect 3130 2765 3150 2785
rect 3130 2715 3150 2735
rect 3130 2665 3150 2685
rect 3130 2615 3150 2635
rect 3130 2565 3150 2585
rect 3130 2515 3150 2535
rect 3130 2465 3150 2485
rect 3130 2415 3150 2435
rect 3230 2765 3250 2785
rect 3230 2715 3250 2735
rect 3230 2665 3250 2685
rect 3230 2615 3250 2635
rect 3230 2565 3250 2585
rect 3230 2515 3250 2535
rect 3230 2465 3250 2485
rect 3230 2415 3250 2435
rect 3330 2765 3350 2785
rect 3330 2715 3350 2735
rect 3330 2665 3350 2685
rect 3330 2615 3350 2635
rect 3330 2565 3350 2585
rect 3330 2515 3350 2535
rect 3330 2465 3350 2485
rect 3330 2415 3350 2435
rect 3430 2765 3450 2785
rect 3430 2715 3450 2735
rect 3430 2665 3450 2685
rect 3430 2615 3450 2635
rect 3430 2565 3450 2585
rect 3430 2515 3450 2535
rect 3430 2465 3450 2485
rect 3430 2415 3450 2435
rect 3530 2765 3550 2785
rect 3530 2715 3550 2735
rect 3530 2665 3550 2685
rect 3530 2615 3550 2635
rect 3530 2565 3550 2585
rect 3530 2515 3550 2535
rect 3530 2465 3550 2485
rect 3530 2415 3550 2435
rect 3630 2765 3650 2785
rect 3630 2715 3650 2735
rect 3630 2665 3650 2685
rect 3630 2615 3650 2635
rect 3630 2565 3650 2585
rect 3630 2515 3650 2535
rect 3630 2465 3650 2485
rect 3630 2415 3650 2435
rect 3730 2765 3750 2785
rect 3730 2715 3750 2735
rect 3730 2665 3750 2685
rect 3730 2615 3750 2635
rect 3730 2565 3750 2585
rect 3730 2515 3750 2535
rect 3730 2465 3750 2485
rect 3730 2415 3750 2435
rect 3830 2765 3850 2785
rect 3830 2715 3850 2735
rect 3830 2665 3850 2685
rect 3830 2615 3850 2635
rect 3830 2565 3850 2585
rect 3830 2515 3850 2535
rect 3830 2465 3850 2485
rect 3830 2415 3850 2435
rect 3930 2765 3950 2785
rect 3930 2715 3950 2735
rect 3930 2665 3950 2685
rect 3930 2615 3950 2635
rect 3930 2565 3950 2585
rect 3930 2515 3950 2535
rect 3930 2465 3950 2485
rect 3930 2415 3950 2435
rect 4030 2765 4050 2785
rect 4030 2715 4050 2735
rect 4030 2665 4050 2685
rect 4030 2615 4050 2635
rect 4030 2565 4050 2585
rect 4030 2515 4050 2535
rect 4030 2465 4050 2485
rect 4030 2415 4050 2435
rect 4130 2765 4150 2785
rect 4130 2715 4150 2735
rect 4130 2665 4150 2685
rect 4130 2615 4150 2635
rect 4130 2565 4150 2585
rect 4130 2515 4150 2535
rect 4130 2465 4150 2485
rect 4130 2415 4150 2435
rect 4230 2765 4250 2785
rect 4230 2715 4250 2735
rect 4230 2665 4250 2685
rect 4230 2615 4250 2635
rect 4230 2565 4250 2585
rect 4230 2515 4250 2535
rect 4230 2465 4250 2485
rect 4230 2415 4250 2435
rect 4330 2765 4350 2785
rect 4330 2715 4350 2735
rect 4330 2665 4350 2685
rect 4330 2615 4350 2635
rect 4330 2565 4350 2585
rect 4330 2515 4350 2535
rect 4330 2465 4350 2485
rect 4330 2415 4350 2435
rect 4430 2765 4450 2785
rect 4430 2715 4450 2735
rect 4430 2665 4450 2685
rect 4430 2615 4450 2635
rect 4430 2565 4450 2585
rect 4430 2515 4450 2535
rect 4430 2465 4450 2485
rect 4430 2415 4450 2435
rect 3030 2145 3050 2165
rect 3030 2095 3050 2115
rect 3030 2045 3050 2065
rect 3030 1995 3050 2015
rect 3130 2145 3150 2165
rect 3130 2095 3150 2115
rect 3130 2045 3150 2065
rect 3130 1995 3150 2015
rect 3230 2145 3250 2165
rect 3230 2095 3250 2115
rect 3230 2045 3250 2065
rect 3230 1995 3250 2015
rect 3330 2145 3350 2165
rect 3330 2095 3350 2115
rect 3330 2045 3350 2065
rect 3330 1995 3350 2015
rect 3430 2145 3450 2165
rect 3430 2095 3450 2115
rect 3430 2045 3450 2065
rect 3430 1995 3450 2015
rect 3530 2145 3550 2165
rect 3530 2095 3550 2115
rect 3530 2045 3550 2065
rect 3530 1995 3550 2015
rect 3630 2145 3650 2165
rect 3630 2095 3650 2115
rect 3630 2045 3650 2065
rect 3630 1995 3650 2015
rect 3730 2145 3750 2165
rect 3730 2095 3750 2115
rect 3730 2045 3750 2065
rect 3730 1995 3750 2015
rect 3830 2145 3850 2165
rect 3830 2095 3850 2115
rect 3830 2045 3850 2065
rect 3830 1995 3850 2015
rect 3930 2145 3950 2165
rect 3930 2095 3950 2115
rect 3930 2045 3950 2065
rect 3930 1995 3950 2015
rect 4030 2145 4050 2165
rect 4030 2095 4050 2115
rect 4030 2045 4050 2065
rect 4030 1995 4050 2015
rect 4130 2145 4150 2165
rect 4130 2095 4150 2115
rect 4130 2045 4150 2065
rect 4130 1995 4150 2015
rect 4230 2145 4250 2165
rect 4230 2095 4250 2115
rect 4230 2045 4250 2065
rect 4230 1995 4250 2015
rect 4330 2145 4350 2165
rect 4330 2095 4350 2115
rect 4330 2045 4350 2065
rect 4330 1995 4350 2015
rect 4430 2145 4450 2165
rect 4430 2095 4450 2115
rect 4430 2045 4450 2065
rect 4430 1995 4450 2015
rect 4540 2145 4560 2165
rect 4540 2095 4560 2115
rect 4540 2045 4560 2065
rect 4540 1995 4560 2015
rect 4595 2145 4615 2165
rect 4595 2095 4615 2115
rect 4595 2045 4615 2065
rect 4595 1995 4615 2015
rect 4665 2145 4685 2165
rect 4665 2095 4685 2115
rect 4665 2045 4685 2065
rect 4665 1995 4685 2015
rect 4720 2145 4740 2165
rect 4720 2095 4740 2115
rect 4720 2045 4740 2065
rect 4720 1995 4740 2015
<< psubdiff >>
rect -50 1715 100 1730
rect -50 1695 -35 1715
rect -15 1695 15 1715
rect 35 1695 65 1715
rect 85 1695 100 1715
rect -50 1680 100 1695
rect 3720 1370 3760 1385
rect 3720 1350 3730 1370
rect 3750 1350 3760 1370
rect 3720 1320 3760 1350
rect 3720 1300 3730 1320
rect 3750 1300 3760 1320
rect 3720 1270 3760 1300
rect 3720 1250 3730 1270
rect 3750 1250 3760 1270
rect 3720 1220 3760 1250
rect 3720 1200 3730 1220
rect 3750 1200 3760 1220
rect 3720 1170 3760 1200
rect 3720 1150 3730 1170
rect 3750 1150 3760 1170
rect 3720 1120 3760 1150
rect 3720 1100 3730 1120
rect 3750 1100 3760 1120
rect 3720 1070 3760 1100
rect 3720 1050 3730 1070
rect 3750 1050 3760 1070
rect 3720 1020 3760 1050
rect 3720 1000 3730 1020
rect 3750 1000 3760 1020
rect 3720 985 3760 1000
rect 4270 840 4310 855
rect 4270 820 4280 840
rect 4300 820 4310 840
rect 4270 790 4310 820
rect 4270 770 4280 790
rect 4300 770 4310 790
rect 4270 755 4310 770
<< nsubdiff >>
rect 2980 2785 3020 2800
rect 2980 2765 2990 2785
rect 3010 2765 3020 2785
rect 2980 2735 3020 2765
rect 2980 2715 2990 2735
rect 3010 2715 3020 2735
rect 2980 2685 3020 2715
rect 2980 2665 2990 2685
rect 3010 2665 3020 2685
rect 2980 2635 3020 2665
rect 2980 2615 2990 2635
rect 3010 2615 3020 2635
rect 2980 2585 3020 2615
rect 2980 2565 2990 2585
rect 3010 2565 3020 2585
rect 2980 2535 3020 2565
rect 2980 2515 2990 2535
rect 3010 2515 3020 2535
rect 2980 2485 3020 2515
rect 2980 2465 2990 2485
rect 3010 2465 3020 2485
rect 2980 2435 3020 2465
rect 2980 2415 2990 2435
rect 3010 2415 3020 2435
rect 2980 2400 3020 2415
rect 4460 2785 4500 2800
rect 4460 2765 4470 2785
rect 4490 2765 4500 2785
rect 4460 2735 4500 2765
rect 4460 2715 4470 2735
rect 4490 2715 4500 2735
rect 4460 2685 4500 2715
rect 4460 2665 4470 2685
rect 4490 2665 4500 2685
rect 4460 2635 4500 2665
rect 4460 2615 4470 2635
rect 4490 2615 4500 2635
rect 4460 2585 4500 2615
rect 4460 2565 4470 2585
rect 4490 2565 4500 2585
rect 4460 2535 4500 2565
rect 4460 2515 4470 2535
rect 4490 2515 4500 2535
rect 4460 2485 4500 2515
rect 4460 2465 4470 2485
rect 4490 2465 4500 2485
rect 4460 2435 4500 2465
rect 4460 2415 4470 2435
rect 4490 2415 4500 2435
rect 4460 2400 4500 2415
rect 2980 2165 3020 2180
rect 2980 2145 2990 2165
rect 3010 2145 3020 2165
rect 2980 2115 3020 2145
rect 2980 2095 2990 2115
rect 3010 2095 3020 2115
rect 2980 2065 3020 2095
rect 2980 2045 2990 2065
rect 3010 2045 3020 2065
rect 2980 2015 3020 2045
rect 2980 1995 2990 2015
rect 3010 1995 3020 2015
rect 2980 1980 3020 1995
rect 4460 2165 4500 2180
rect 4460 2145 4470 2165
rect 4490 2145 4500 2165
rect 4460 2115 4500 2145
rect 4460 2095 4470 2115
rect 4490 2095 4500 2115
rect 4460 2065 4500 2095
rect 4460 2045 4470 2065
rect 4490 2045 4500 2065
rect 4460 2015 4500 2045
rect 4460 1995 4470 2015
rect 4490 1995 4500 2015
rect 4460 1980 4500 1995
<< psubdiffcont >>
rect -35 1695 -15 1715
rect 15 1695 35 1715
rect 65 1695 85 1715
rect 3730 1350 3750 1370
rect 3730 1300 3750 1320
rect 3730 1250 3750 1270
rect 3730 1200 3750 1220
rect 3730 1150 3750 1170
rect 3730 1100 3750 1120
rect 3730 1050 3750 1070
rect 3730 1000 3750 1020
rect 4280 820 4300 840
rect 4280 770 4300 790
<< nsubdiffcont >>
rect 2990 2765 3010 2785
rect 2990 2715 3010 2735
rect 2990 2665 3010 2685
rect 2990 2615 3010 2635
rect 2990 2565 3010 2585
rect 2990 2515 3010 2535
rect 2990 2465 3010 2485
rect 2990 2415 3010 2435
rect 4470 2765 4490 2785
rect 4470 2715 4490 2735
rect 4470 2665 4490 2685
rect 4470 2615 4490 2635
rect 4470 2565 4490 2585
rect 4470 2515 4490 2535
rect 4470 2465 4490 2485
rect 4470 2415 4490 2435
rect 2990 2145 3010 2165
rect 2990 2095 3010 2115
rect 2990 2045 3010 2065
rect 2990 1995 3010 2015
rect 4470 2145 4490 2165
rect 4470 2095 4490 2115
rect 4470 2045 4490 2065
rect 4470 1995 4490 2015
<< poly >>
rect 3070 2845 3110 2855
rect 3070 2825 3080 2845
rect 3100 2825 3110 2845
rect 3070 2815 3110 2825
rect 4370 2845 4410 2855
rect 4370 2825 4380 2845
rect 4400 2825 4410 2845
rect 4370 2815 4410 2825
rect 3060 2800 3120 2815
rect 3160 2800 3220 2815
rect 3260 2800 3320 2815
rect 3360 2800 3420 2815
rect 3460 2800 3520 2815
rect 3560 2800 3620 2815
rect 3660 2800 3720 2815
rect 3760 2800 3820 2815
rect 3860 2800 3920 2815
rect 3960 2800 4020 2815
rect 4060 2800 4120 2815
rect 4160 2800 4220 2815
rect 4260 2800 4320 2815
rect 4360 2800 4420 2815
rect 3060 2385 3120 2400
rect 3160 2390 3220 2400
rect 3260 2390 3320 2400
rect 3360 2390 3420 2400
rect 3460 2390 3520 2400
rect 3560 2390 3620 2400
rect 3660 2390 3720 2400
rect 3760 2390 3820 2400
rect 3860 2390 3920 2400
rect 3960 2390 4020 2400
rect 4060 2390 4120 2400
rect 4160 2390 4220 2400
rect 4260 2390 4320 2400
rect 3160 2375 4320 2390
rect 4360 2385 4420 2400
rect 4270 2355 4280 2375
rect 4300 2355 4310 2375
rect 4270 2345 4310 2355
rect 4670 2265 4710 2275
rect 4670 2245 4680 2265
rect 4700 2245 4710 2265
rect 4670 2235 4710 2245
rect 3070 2225 3110 2235
rect 3070 2205 3080 2225
rect 3100 2205 3110 2225
rect 3070 2195 3110 2205
rect 4370 2225 4410 2235
rect 4370 2205 4380 2225
rect 4400 2205 4410 2225
rect 4370 2195 4410 2205
rect 3060 2180 3120 2195
rect 3160 2180 3220 2195
rect 3260 2180 3320 2195
rect 3360 2180 3420 2195
rect 3460 2180 3520 2195
rect 3560 2180 3620 2195
rect 3660 2180 3720 2195
rect 3760 2180 3820 2195
rect 3860 2180 3920 2195
rect 3960 2180 4020 2195
rect 4060 2180 4120 2195
rect 4160 2180 4220 2195
rect 4260 2180 4320 2195
rect 4360 2180 4420 2195
rect 4570 2180 4585 2195
rect 4695 2180 4710 2235
rect 3060 1965 3120 1980
rect 3160 1965 3220 1980
rect 3260 1970 3320 1980
rect 3360 1970 3420 1980
rect 3460 1970 3520 1980
rect 3560 1970 3620 1980
rect 3180 1915 3200 1965
rect 3260 1955 3620 1970
rect 3660 1970 3720 1980
rect 3760 1970 3820 1980
rect 3660 1955 3820 1970
rect 3860 1970 3920 1980
rect 3960 1970 4020 1980
rect 4060 1970 4120 1980
rect 4160 1970 4220 1980
rect 3860 1955 4220 1970
rect 4260 1965 4320 1980
rect 4360 1965 4420 1980
rect 3320 1950 3360 1955
rect 3320 1930 3330 1950
rect 3350 1930 3360 1950
rect 3320 1920 3360 1930
rect 3680 1915 3700 1955
rect 3780 1915 3800 1955
rect 4120 1950 4160 1955
rect 4120 1930 4130 1950
rect 4150 1930 4160 1950
rect 4120 1920 4160 1930
rect 4280 1915 4300 1965
rect 4570 1940 4585 1980
rect 4695 1965 4710 1980
rect 4640 1940 4680 1950
rect 4570 1920 4650 1940
rect 4670 1920 4680 1940
rect 3170 1905 3210 1915
rect 3170 1885 3180 1905
rect 3200 1885 3210 1905
rect 3170 1875 3210 1885
rect 3670 1905 3710 1915
rect 3670 1885 3680 1905
rect 3700 1885 3710 1905
rect 3670 1875 3710 1885
rect 3770 1905 3810 1915
rect 3770 1885 3780 1905
rect 3800 1885 3810 1905
rect 3770 1875 3810 1885
rect 4270 1905 4310 1915
rect 4640 1910 4680 1920
rect 4270 1885 4280 1905
rect 4300 1885 4310 1905
rect 4270 1875 4310 1885
rect 3370 1700 3410 1710
rect 3370 1680 3380 1700
rect 3400 1680 3410 1700
rect 3670 1700 3710 1710
rect 3670 1685 3680 1700
rect 3370 1675 3410 1680
rect 3660 1680 3680 1685
rect 3700 1685 3710 1700
rect 3770 1700 3810 1710
rect 3770 1685 3780 1700
rect 3700 1680 3780 1685
rect 3800 1685 3810 1700
rect 4070 1700 4110 1710
rect 3800 1680 3820 1685
rect 3260 1660 3320 1675
rect 3360 1660 3420 1675
rect 3460 1660 3520 1675
rect 3560 1660 3620 1675
rect 3660 1670 3820 1680
rect 4070 1680 4080 1700
rect 4100 1680 4110 1700
rect 4070 1675 4110 1680
rect 3660 1660 3720 1670
rect 3760 1660 3820 1670
rect 3860 1660 3920 1675
rect 3960 1660 4020 1675
rect 4060 1660 4120 1675
rect 4160 1660 4220 1675
rect 3260 1545 3320 1560
rect 3360 1545 3420 1560
rect 3460 1550 3520 1560
rect 3560 1550 3620 1560
rect 3270 1540 3310 1545
rect 3270 1520 3280 1540
rect 3300 1520 3310 1540
rect 3460 1535 3620 1550
rect 3660 1545 3720 1560
rect 3760 1545 3820 1560
rect 3860 1550 3920 1560
rect 3960 1550 4020 1560
rect 3860 1535 4020 1550
rect 4060 1545 4120 1560
rect 4160 1545 4220 1560
rect 4170 1540 4210 1545
rect 3270 1510 3310 1520
rect 3520 1515 3530 1535
rect 3550 1515 3560 1535
rect 3520 1505 3560 1515
rect 3920 1515 3930 1535
rect 3950 1515 3960 1535
rect 3920 1505 3960 1515
rect 4170 1520 4180 1540
rect 4200 1520 4210 1540
rect 4170 1510 4210 1520
rect 3280 1430 3680 1440
rect 3280 1410 3290 1430
rect 3310 1410 3330 1430
rect 3350 1410 3370 1430
rect 3390 1410 3410 1430
rect 3430 1410 3450 1430
rect 3470 1410 3490 1430
rect 3510 1410 3530 1430
rect 3550 1410 3570 1430
rect 3590 1410 3610 1430
rect 3630 1410 3650 1430
rect 3670 1410 3680 1430
rect 3280 1385 3680 1410
rect 3800 1430 4200 1440
rect 3800 1410 3810 1430
rect 3830 1410 3850 1430
rect 3870 1410 3890 1430
rect 3910 1410 3930 1430
rect 3950 1410 3970 1430
rect 3990 1410 4010 1430
rect 4030 1410 4050 1430
rect 4070 1410 4090 1430
rect 4110 1410 4130 1430
rect 4150 1410 4170 1430
rect 4190 1410 4200 1430
rect 3800 1385 4200 1410
rect 3280 970 3680 985
rect 3800 970 4200 985
rect 3230 900 3270 910
rect 3230 880 3240 900
rect 3260 880 3270 900
rect 3230 870 3270 880
rect 3310 900 3350 910
rect 3310 880 3320 900
rect 3340 880 3350 900
rect 3310 870 3350 880
rect 3390 900 3430 910
rect 3390 880 3400 900
rect 3420 880 3430 900
rect 3390 870 3430 880
rect 3470 900 3510 910
rect 3470 880 3480 900
rect 3500 880 3510 900
rect 3470 870 3510 880
rect 3550 900 3590 910
rect 3550 880 3560 900
rect 3580 880 3590 900
rect 3550 870 3590 880
rect 3630 900 3670 910
rect 3630 880 3640 900
rect 3660 880 3670 900
rect 3630 870 3670 880
rect 3710 900 3750 910
rect 3710 880 3720 900
rect 3740 880 3750 900
rect 3710 870 3750 880
rect 3790 900 3830 910
rect 3790 880 3800 900
rect 3820 880 3830 900
rect 3790 870 3830 880
rect 3870 900 3910 910
rect 3870 880 3880 900
rect 3900 880 3910 900
rect 3870 870 3910 880
rect 3950 900 3990 910
rect 3950 880 3960 900
rect 3980 880 3990 900
rect 3950 870 3990 880
rect 4030 900 4070 910
rect 4030 880 4040 900
rect 4060 880 4070 900
rect 4030 870 4070 880
rect 4110 900 4150 910
rect 4110 880 4120 900
rect 4140 880 4150 900
rect 4110 870 4150 880
rect 4190 900 4230 910
rect 4190 880 4200 900
rect 4220 880 4230 900
rect 4190 870 4230 880
rect 3230 855 4230 870
rect 3230 740 4230 755
<< polycont >>
rect 3080 2825 3100 2845
rect 4380 2825 4400 2845
rect 4280 2355 4300 2375
rect 4680 2245 4700 2265
rect 3080 2205 3100 2225
rect 4380 2205 4400 2225
rect 3330 1930 3350 1950
rect 4130 1930 4150 1950
rect 4650 1920 4670 1940
rect 3180 1885 3200 1905
rect 3680 1885 3700 1905
rect 3780 1885 3800 1905
rect 4280 1885 4300 1905
rect 3380 1680 3400 1700
rect 3680 1680 3700 1700
rect 3780 1680 3800 1700
rect 4080 1680 4100 1700
rect 3280 1520 3300 1540
rect 3530 1515 3550 1535
rect 3930 1515 3950 1535
rect 4180 1520 4200 1540
rect 3290 1410 3310 1430
rect 3330 1410 3350 1430
rect 3370 1410 3390 1430
rect 3410 1410 3430 1430
rect 3450 1410 3470 1430
rect 3490 1410 3510 1430
rect 3530 1410 3550 1430
rect 3570 1410 3590 1430
rect 3610 1410 3630 1430
rect 3650 1410 3670 1430
rect 3810 1410 3830 1430
rect 3850 1410 3870 1430
rect 3890 1410 3910 1430
rect 3930 1410 3950 1430
rect 3970 1410 3990 1430
rect 4010 1410 4030 1430
rect 4050 1410 4070 1430
rect 4090 1410 4110 1430
rect 4130 1410 4150 1430
rect 4170 1410 4190 1430
rect 3240 880 3260 900
rect 3320 880 3340 900
rect 3400 880 3420 900
rect 3480 880 3500 900
rect 3560 880 3580 900
rect 3640 880 3660 900
rect 3720 880 3740 900
rect 3800 880 3820 900
rect 3880 880 3900 900
rect 3960 880 3980 900
rect 4040 880 4060 900
rect 4120 880 4140 900
rect 4200 880 4220 900
<< xpolycontact >>
rect 1705 2565 1925 2600
rect 2469 2565 2689 2600
rect 1705 2505 1925 2540
rect 2469 2505 2689 2540
rect 1705 2445 1925 2480
rect 2469 2445 2689 2480
rect 1705 2385 1925 2420
rect 2469 2385 2689 2420
rect 1705 2325 1925 2360
rect 2469 2325 2689 2360
rect 1705 2265 1925 2300
rect 2469 2265 2689 2300
rect 1705 2205 1925 2240
rect 2469 2205 2689 2240
rect 1705 2145 1925 2180
rect 2469 2145 2689 2180
rect 1705 2085 1925 2120
rect 2469 2085 2689 2120
rect 1705 2025 1925 2060
rect 2259 2025 2479 2060
rect 1705 1965 1925 2000
rect 2469 1965 2689 2000
rect 1705 1905 1925 1940
rect 2469 1905 2689 1940
rect 1705 1845 1925 1880
rect 2469 1845 2689 1880
rect 1705 1785 1925 1820
rect 2469 1785 2689 1820
rect 1705 1725 1925 1760
rect 2469 1725 2689 1760
rect 1705 1665 1925 1700
rect 2469 1665 2689 1700
rect 1705 1605 1925 1640
rect 2469 1605 2689 1640
rect 1705 1545 1925 1580
rect 2469 1545 2689 1580
rect 1705 1485 1925 1520
rect 2469 1485 2689 1520
<< xpolyres >>
rect 1925 2565 2469 2600
rect 1925 2505 2469 2540
rect 1925 2445 2469 2480
rect 1925 2385 2469 2420
rect 1925 2325 2469 2360
rect 1925 2265 2469 2300
rect 1925 2205 2469 2240
rect 1925 2145 2469 2180
rect 1925 2085 2469 2120
rect 1925 2025 2259 2060
rect 1925 1965 2469 2000
rect 1925 1905 2469 1940
rect 1925 1845 2469 1880
rect 1925 1785 2469 1820
rect 1925 1725 2469 1760
rect 1925 1665 2469 1700
rect 1925 1605 2469 1640
rect 1925 1545 2469 1580
rect 1925 1485 2469 1520
<< locali >>
rect 3020 2845 3120 2855
rect 3020 2825 3030 2845
rect 3050 2825 3080 2845
rect 3100 2825 3120 2845
rect 3020 2815 3120 2825
rect 3220 2845 3260 2855
rect 3220 2825 3230 2845
rect 3250 2825 3260 2845
rect 3220 2815 3260 2825
rect 3420 2845 3460 2855
rect 3420 2825 3430 2845
rect 3450 2825 3460 2845
rect 3420 2815 3460 2825
rect 3620 2845 3660 2855
rect 3620 2825 3630 2845
rect 3650 2825 3660 2845
rect 3620 2815 3660 2825
rect 3720 2845 3760 2855
rect 3720 2825 3730 2845
rect 3750 2825 3760 2845
rect 3720 2815 3760 2825
rect 3820 2845 3860 2855
rect 3820 2825 3830 2845
rect 3850 2825 3860 2845
rect 3820 2815 3860 2825
rect 4020 2845 4060 2855
rect 4020 2825 4030 2845
rect 4050 2825 4060 2845
rect 4020 2815 4060 2825
rect 4220 2845 4260 2855
rect 4220 2825 4230 2845
rect 4250 2825 4260 2845
rect 4220 2815 4260 2825
rect 4360 2845 4460 2855
rect 4360 2825 4380 2845
rect 4400 2825 4430 2845
rect 4450 2825 4460 2845
rect 4360 2815 4460 2825
rect 3030 2795 3050 2815
rect 3230 2795 3250 2815
rect 3430 2795 3450 2815
rect 3630 2795 3650 2815
rect 3730 2795 3750 2815
rect 3830 2795 3850 2815
rect 4030 2795 4050 2815
rect 4230 2795 4250 2815
rect 4430 2795 4450 2815
rect 2985 2785 3055 2795
rect 2985 2765 2990 2785
rect 3010 2765 3030 2785
rect 3050 2765 3055 2785
rect 2985 2735 3055 2765
rect 2985 2715 2990 2735
rect 3010 2715 3030 2735
rect 3050 2715 3055 2735
rect 650 2055 775 2700
rect 1330 2055 1455 2700
rect 2985 2685 3055 2715
rect 2985 2665 2990 2685
rect 3010 2665 3030 2685
rect 3050 2665 3055 2685
rect 2985 2635 3055 2665
rect 2985 2615 2990 2635
rect 3010 2615 3030 2635
rect 3050 2615 3055 2635
rect 1660 2595 1705 2600
rect 1660 2570 1670 2595
rect 1695 2570 1705 2595
rect 1660 2565 1705 2570
rect 2689 2565 2769 2600
rect 1660 2535 1705 2540
rect 1660 2510 1670 2535
rect 1695 2510 1705 2535
rect 1660 2505 1705 2510
rect 2689 2505 2729 2540
rect 1660 2475 1705 2480
rect 1660 2450 1670 2475
rect 1695 2450 1705 2475
rect 1660 2445 1705 2450
rect 2654 2420 2689 2445
rect 1625 2385 1705 2420
rect 1625 2120 1645 2385
rect 2709 2360 2729 2505
rect 1665 2325 1705 2360
rect 2689 2325 2729 2360
rect 1665 2180 1685 2325
rect 2749 2300 2769 2565
rect 2985 2585 3055 2615
rect 2985 2565 2990 2585
rect 3010 2565 3030 2585
rect 3050 2565 3055 2585
rect 2985 2535 3055 2565
rect 2985 2515 2990 2535
rect 3010 2515 3030 2535
rect 3050 2515 3055 2535
rect 2985 2485 3055 2515
rect 2985 2465 2990 2485
rect 3010 2465 3030 2485
rect 3050 2465 3055 2485
rect 2985 2435 3055 2465
rect 2985 2415 2990 2435
rect 3010 2415 3030 2435
rect 3050 2415 3055 2435
rect 2985 2405 3055 2415
rect 3125 2785 3155 2795
rect 3125 2765 3130 2785
rect 3150 2765 3155 2785
rect 3125 2735 3155 2765
rect 3125 2715 3130 2735
rect 3150 2715 3155 2735
rect 3125 2685 3155 2715
rect 3125 2665 3130 2685
rect 3150 2665 3155 2685
rect 3125 2635 3155 2665
rect 3125 2615 3130 2635
rect 3150 2615 3155 2635
rect 3125 2585 3155 2615
rect 3125 2565 3130 2585
rect 3150 2565 3155 2585
rect 3125 2535 3155 2565
rect 3125 2515 3130 2535
rect 3150 2515 3155 2535
rect 3125 2485 3155 2515
rect 3125 2465 3130 2485
rect 3150 2465 3155 2485
rect 3125 2435 3155 2465
rect 3125 2415 3130 2435
rect 3150 2415 3155 2435
rect 3125 2405 3155 2415
rect 3225 2785 3255 2795
rect 3225 2765 3230 2785
rect 3250 2765 3255 2785
rect 3225 2735 3255 2765
rect 3225 2715 3230 2735
rect 3250 2715 3255 2735
rect 3225 2685 3255 2715
rect 3225 2665 3230 2685
rect 3250 2665 3255 2685
rect 3225 2635 3255 2665
rect 3225 2615 3230 2635
rect 3250 2615 3255 2635
rect 3225 2585 3255 2615
rect 3225 2565 3230 2585
rect 3250 2565 3255 2585
rect 3225 2535 3255 2565
rect 3225 2515 3230 2535
rect 3250 2515 3255 2535
rect 3225 2485 3255 2515
rect 3225 2465 3230 2485
rect 3250 2465 3255 2485
rect 3225 2435 3255 2465
rect 3225 2415 3230 2435
rect 3250 2415 3255 2435
rect 3225 2405 3255 2415
rect 3325 2785 3355 2795
rect 3325 2765 3330 2785
rect 3350 2765 3355 2785
rect 3325 2735 3355 2765
rect 3325 2715 3330 2735
rect 3350 2715 3355 2735
rect 3325 2685 3355 2715
rect 3325 2665 3330 2685
rect 3350 2665 3355 2685
rect 3325 2635 3355 2665
rect 3325 2615 3330 2635
rect 3350 2615 3355 2635
rect 3325 2585 3355 2615
rect 3325 2565 3330 2585
rect 3350 2565 3355 2585
rect 3325 2535 3355 2565
rect 3325 2515 3330 2535
rect 3350 2515 3355 2535
rect 3325 2485 3355 2515
rect 3325 2465 3330 2485
rect 3350 2465 3355 2485
rect 3325 2435 3355 2465
rect 3325 2415 3330 2435
rect 3350 2415 3355 2435
rect 3325 2405 3355 2415
rect 3425 2785 3455 2795
rect 3425 2765 3430 2785
rect 3450 2765 3455 2785
rect 3425 2735 3455 2765
rect 3425 2715 3430 2735
rect 3450 2715 3455 2735
rect 3425 2685 3455 2715
rect 3425 2665 3430 2685
rect 3450 2665 3455 2685
rect 3425 2635 3455 2665
rect 3425 2615 3430 2635
rect 3450 2615 3455 2635
rect 3425 2585 3455 2615
rect 3425 2565 3430 2585
rect 3450 2565 3455 2585
rect 3425 2535 3455 2565
rect 3425 2515 3430 2535
rect 3450 2515 3455 2535
rect 3425 2485 3455 2515
rect 3425 2465 3430 2485
rect 3450 2465 3455 2485
rect 3425 2435 3455 2465
rect 3425 2415 3430 2435
rect 3450 2415 3455 2435
rect 3425 2405 3455 2415
rect 3525 2785 3555 2795
rect 3525 2765 3530 2785
rect 3550 2765 3555 2785
rect 3525 2735 3555 2765
rect 3525 2715 3530 2735
rect 3550 2715 3555 2735
rect 3525 2685 3555 2715
rect 3525 2665 3530 2685
rect 3550 2665 3555 2685
rect 3525 2635 3555 2665
rect 3525 2615 3530 2635
rect 3550 2615 3555 2635
rect 3525 2585 3555 2615
rect 3525 2565 3530 2585
rect 3550 2565 3555 2585
rect 3525 2535 3555 2565
rect 3525 2515 3530 2535
rect 3550 2515 3555 2535
rect 3525 2485 3555 2515
rect 3525 2465 3530 2485
rect 3550 2465 3555 2485
rect 3525 2435 3555 2465
rect 3525 2415 3530 2435
rect 3550 2415 3555 2435
rect 3525 2405 3555 2415
rect 3625 2785 3655 2795
rect 3625 2765 3630 2785
rect 3650 2765 3655 2785
rect 3625 2735 3655 2765
rect 3625 2715 3630 2735
rect 3650 2715 3655 2735
rect 3625 2685 3655 2715
rect 3625 2665 3630 2685
rect 3650 2665 3655 2685
rect 3625 2635 3655 2665
rect 3625 2615 3630 2635
rect 3650 2615 3655 2635
rect 3625 2585 3655 2615
rect 3625 2565 3630 2585
rect 3650 2565 3655 2585
rect 3625 2535 3655 2565
rect 3625 2515 3630 2535
rect 3650 2515 3655 2535
rect 3625 2485 3655 2515
rect 3625 2465 3630 2485
rect 3650 2465 3655 2485
rect 3625 2435 3655 2465
rect 3625 2415 3630 2435
rect 3650 2415 3655 2435
rect 3625 2405 3655 2415
rect 3725 2785 3755 2795
rect 3725 2765 3730 2785
rect 3750 2765 3755 2785
rect 3725 2735 3755 2765
rect 3725 2715 3730 2735
rect 3750 2715 3755 2735
rect 3725 2685 3755 2715
rect 3725 2665 3730 2685
rect 3750 2665 3755 2685
rect 3725 2635 3755 2665
rect 3725 2615 3730 2635
rect 3750 2615 3755 2635
rect 3725 2585 3755 2615
rect 3725 2565 3730 2585
rect 3750 2565 3755 2585
rect 3725 2535 3755 2565
rect 3725 2515 3730 2535
rect 3750 2515 3755 2535
rect 3725 2485 3755 2515
rect 3725 2465 3730 2485
rect 3750 2465 3755 2485
rect 3725 2435 3755 2465
rect 3725 2415 3730 2435
rect 3750 2415 3755 2435
rect 3725 2405 3755 2415
rect 3825 2785 3855 2795
rect 3825 2765 3830 2785
rect 3850 2765 3855 2785
rect 3825 2735 3855 2765
rect 3825 2715 3830 2735
rect 3850 2715 3855 2735
rect 3825 2685 3855 2715
rect 3825 2665 3830 2685
rect 3850 2665 3855 2685
rect 3825 2635 3855 2665
rect 3825 2615 3830 2635
rect 3850 2615 3855 2635
rect 3825 2585 3855 2615
rect 3825 2565 3830 2585
rect 3850 2565 3855 2585
rect 3825 2535 3855 2565
rect 3825 2515 3830 2535
rect 3850 2515 3855 2535
rect 3825 2485 3855 2515
rect 3825 2465 3830 2485
rect 3850 2465 3855 2485
rect 3825 2435 3855 2465
rect 3825 2415 3830 2435
rect 3850 2415 3855 2435
rect 3825 2405 3855 2415
rect 3925 2785 3955 2795
rect 3925 2765 3930 2785
rect 3950 2765 3955 2785
rect 3925 2735 3955 2765
rect 3925 2715 3930 2735
rect 3950 2715 3955 2735
rect 3925 2685 3955 2715
rect 3925 2665 3930 2685
rect 3950 2665 3955 2685
rect 3925 2635 3955 2665
rect 3925 2615 3930 2635
rect 3950 2615 3955 2635
rect 3925 2585 3955 2615
rect 3925 2565 3930 2585
rect 3950 2565 3955 2585
rect 3925 2535 3955 2565
rect 3925 2515 3930 2535
rect 3950 2515 3955 2535
rect 3925 2485 3955 2515
rect 3925 2465 3930 2485
rect 3950 2465 3955 2485
rect 3925 2435 3955 2465
rect 3925 2415 3930 2435
rect 3950 2415 3955 2435
rect 3925 2405 3955 2415
rect 4025 2785 4055 2795
rect 4025 2765 4030 2785
rect 4050 2765 4055 2785
rect 4025 2735 4055 2765
rect 4025 2715 4030 2735
rect 4050 2715 4055 2735
rect 4025 2685 4055 2715
rect 4025 2665 4030 2685
rect 4050 2665 4055 2685
rect 4025 2635 4055 2665
rect 4025 2615 4030 2635
rect 4050 2615 4055 2635
rect 4025 2585 4055 2615
rect 4025 2565 4030 2585
rect 4050 2565 4055 2585
rect 4025 2535 4055 2565
rect 4025 2515 4030 2535
rect 4050 2515 4055 2535
rect 4025 2485 4055 2515
rect 4025 2465 4030 2485
rect 4050 2465 4055 2485
rect 4025 2435 4055 2465
rect 4025 2415 4030 2435
rect 4050 2415 4055 2435
rect 4025 2405 4055 2415
rect 4125 2785 4155 2795
rect 4125 2765 4130 2785
rect 4150 2765 4155 2785
rect 4125 2735 4155 2765
rect 4125 2715 4130 2735
rect 4150 2715 4155 2735
rect 4125 2685 4155 2715
rect 4125 2665 4130 2685
rect 4150 2665 4155 2685
rect 4125 2635 4155 2665
rect 4125 2615 4130 2635
rect 4150 2615 4155 2635
rect 4125 2585 4155 2615
rect 4125 2565 4130 2585
rect 4150 2565 4155 2585
rect 4125 2535 4155 2565
rect 4125 2515 4130 2535
rect 4150 2515 4155 2535
rect 4125 2485 4155 2515
rect 4125 2465 4130 2485
rect 4150 2465 4155 2485
rect 4125 2435 4155 2465
rect 4125 2415 4130 2435
rect 4150 2415 4155 2435
rect 4125 2405 4155 2415
rect 4225 2785 4255 2795
rect 4225 2765 4230 2785
rect 4250 2765 4255 2785
rect 4225 2735 4255 2765
rect 4225 2715 4230 2735
rect 4250 2715 4255 2735
rect 4225 2685 4255 2715
rect 4225 2665 4230 2685
rect 4250 2665 4255 2685
rect 4225 2635 4255 2665
rect 4225 2615 4230 2635
rect 4250 2615 4255 2635
rect 4225 2585 4255 2615
rect 4225 2565 4230 2585
rect 4250 2565 4255 2585
rect 4225 2535 4255 2565
rect 4225 2515 4230 2535
rect 4250 2515 4255 2535
rect 4225 2485 4255 2515
rect 4225 2465 4230 2485
rect 4250 2465 4255 2485
rect 4225 2435 4255 2465
rect 4225 2415 4230 2435
rect 4250 2415 4255 2435
rect 4225 2405 4255 2415
rect 4325 2785 4355 2795
rect 4325 2765 4330 2785
rect 4350 2765 4355 2785
rect 4325 2735 4355 2765
rect 4325 2715 4330 2735
rect 4350 2715 4355 2735
rect 4325 2685 4355 2715
rect 4325 2665 4330 2685
rect 4350 2665 4355 2685
rect 4325 2635 4355 2665
rect 4325 2615 4330 2635
rect 4350 2615 4355 2635
rect 4325 2585 4355 2615
rect 4325 2565 4330 2585
rect 4350 2565 4355 2585
rect 4325 2535 4355 2565
rect 4325 2515 4330 2535
rect 4350 2515 4355 2535
rect 4325 2485 4355 2515
rect 4325 2465 4330 2485
rect 4350 2465 4355 2485
rect 4325 2435 4355 2465
rect 4325 2415 4330 2435
rect 4350 2415 4355 2435
rect 4325 2405 4355 2415
rect 4425 2785 4495 2795
rect 4425 2765 4430 2785
rect 4450 2765 4470 2785
rect 4490 2765 4495 2785
rect 4425 2735 4495 2765
rect 4425 2715 4430 2735
rect 4450 2715 4470 2735
rect 4490 2715 4495 2735
rect 4425 2685 4495 2715
rect 4425 2665 4430 2685
rect 4450 2665 4470 2685
rect 4490 2665 4495 2685
rect 4425 2635 4495 2665
rect 4425 2615 4430 2635
rect 4450 2615 4470 2635
rect 4490 2615 4495 2635
rect 4425 2585 4495 2615
rect 4425 2565 4430 2585
rect 4450 2565 4470 2585
rect 4490 2565 4495 2585
rect 4425 2535 4495 2565
rect 4425 2515 4430 2535
rect 4450 2515 4470 2535
rect 4490 2515 4495 2535
rect 4425 2485 4495 2515
rect 4425 2465 4430 2485
rect 4450 2465 4470 2485
rect 4490 2465 4495 2485
rect 4425 2435 4495 2465
rect 4425 2415 4430 2435
rect 4450 2415 4470 2435
rect 4490 2415 4495 2435
rect 4425 2405 4495 2415
rect 2689 2265 2769 2300
rect 3130 2295 3150 2405
rect 3330 2340 3350 2405
rect 3530 2385 3550 2405
rect 3520 2375 3560 2385
rect 3520 2355 3530 2375
rect 3550 2355 3560 2375
rect 3520 2345 3560 2355
rect 3330 2330 3370 2340
rect 3330 2310 3340 2330
rect 3360 2310 3370 2330
rect 3330 2300 3370 2310
rect 3730 2295 3750 2405
rect 3930 2385 3950 2405
rect 3920 2375 3960 2385
rect 3920 2355 3930 2375
rect 3950 2355 3960 2375
rect 3920 2345 3960 2355
rect 4130 2340 4150 2405
rect 4270 2375 4310 2385
rect 4270 2355 4280 2375
rect 4300 2355 4310 2375
rect 4270 2345 4310 2355
rect 4110 2330 4150 2340
rect 4110 2310 4120 2330
rect 4140 2310 4150 2330
rect 4110 2300 4150 2310
rect 4330 2295 4350 2405
rect 3120 2285 3160 2295
rect 3120 2265 3130 2285
rect 3150 2265 3160 2285
rect 1705 2240 1740 2265
rect 3120 2255 3160 2265
rect 3720 2285 3760 2295
rect 3720 2265 3730 2285
rect 3750 2265 3760 2285
rect 3720 2255 3760 2265
rect 4320 2285 4360 2295
rect 4320 2265 4330 2285
rect 4350 2265 4360 2285
rect 4320 2255 4360 2265
rect 4530 2275 4570 2285
rect 4530 2255 4540 2275
rect 4560 2265 4710 2275
rect 4560 2255 4680 2265
rect 4530 2245 4570 2255
rect 4670 2245 4680 2255
rect 4700 2245 4710 2265
rect 2689 2205 2769 2240
rect 1665 2145 1705 2180
rect 2689 2145 2729 2180
rect 1625 2085 1705 2120
rect 125 2015 1455 2055
rect 1520 2055 1565 2060
rect 1520 2030 1530 2055
rect 1555 2030 1565 2055
rect 1520 2025 1565 2030
rect 1660 2055 1705 2060
rect 1660 2030 1670 2055
rect 1695 2030 1705 2055
rect 1660 2025 1705 2030
rect 2479 2055 2524 2060
rect 2479 2030 2489 2055
rect 2514 2030 2524 2055
rect 2479 2025 2524 2030
rect -45 1715 130 1725
rect -45 1695 -35 1715
rect -15 1695 15 1715
rect 35 1695 65 1715
rect 85 1695 130 1715
rect -45 1685 130 1695
rect 650 1375 775 2015
rect 1330 1375 1455 2015
rect 2654 2000 2689 2085
rect 1625 1965 1705 2000
rect 1625 1700 1645 1965
rect 2709 1940 2729 2145
rect 1665 1905 1705 1940
rect 2689 1905 2729 1940
rect 1665 1760 1685 1905
rect 2749 1880 2769 2205
rect 3020 2225 3120 2235
rect 3020 2205 3030 2225
rect 3050 2205 3080 2225
rect 3100 2205 3120 2225
rect 3020 2195 3120 2205
rect 3220 2225 3260 2235
rect 3220 2205 3230 2225
rect 3250 2205 3260 2225
rect 3220 2195 3260 2205
rect 3420 2225 3460 2235
rect 3420 2205 3430 2225
rect 3450 2205 3460 2225
rect 3420 2195 3460 2205
rect 3620 2225 3660 2235
rect 3620 2205 3630 2225
rect 3650 2205 3660 2225
rect 3620 2195 3660 2205
rect 3820 2225 3860 2235
rect 3820 2205 3830 2225
rect 3850 2205 3860 2225
rect 3820 2195 3860 2205
rect 4020 2225 4060 2235
rect 4020 2205 4030 2225
rect 4050 2205 4060 2225
rect 4020 2195 4060 2205
rect 4220 2225 4260 2235
rect 4220 2205 4230 2225
rect 4250 2205 4260 2225
rect 4220 2195 4260 2205
rect 4370 2225 4460 2235
rect 4370 2205 4380 2225
rect 4400 2205 4430 2225
rect 4450 2205 4460 2225
rect 4370 2195 4460 2205
rect 3030 2175 3050 2195
rect 3230 2175 3250 2195
rect 3430 2175 3450 2195
rect 3630 2175 3650 2195
rect 3830 2175 3850 2195
rect 4030 2175 4050 2195
rect 4230 2175 4250 2195
rect 4430 2175 4450 2195
rect 4540 2175 4560 2245
rect 4670 2235 4710 2245
rect 4740 2225 4780 2235
rect 4740 2205 4750 2225
rect 4770 2205 4780 2225
rect 4740 2195 4780 2205
rect 4750 2175 4770 2195
rect 2985 2165 3055 2175
rect 2985 2145 2990 2165
rect 3010 2145 3030 2165
rect 3050 2145 3055 2165
rect 2985 2115 3055 2145
rect 2985 2095 2990 2115
rect 3010 2095 3030 2115
rect 3050 2095 3055 2115
rect 2985 2065 3055 2095
rect 2985 2045 2990 2065
rect 3010 2045 3030 2065
rect 3050 2045 3055 2065
rect 2985 2015 3055 2045
rect 2985 1995 2990 2015
rect 3010 1995 3030 2015
rect 3050 1995 3055 2015
rect 2985 1985 3055 1995
rect 3125 2165 3155 2175
rect 3125 2145 3130 2165
rect 3150 2145 3155 2165
rect 3125 2115 3155 2145
rect 3125 2095 3130 2115
rect 3150 2095 3155 2115
rect 3125 2065 3155 2095
rect 3125 2045 3130 2065
rect 3150 2045 3155 2065
rect 3125 2015 3155 2045
rect 3125 1995 3130 2015
rect 3150 1995 3155 2015
rect 3125 1985 3155 1995
rect 3225 2165 3255 2175
rect 3225 2145 3230 2165
rect 3250 2145 3255 2165
rect 3225 2115 3255 2145
rect 3225 2095 3230 2115
rect 3250 2095 3255 2115
rect 3225 2065 3255 2095
rect 3225 2045 3230 2065
rect 3250 2045 3255 2065
rect 3225 2015 3255 2045
rect 3225 1995 3230 2015
rect 3250 1995 3255 2015
rect 3225 1985 3255 1995
rect 3325 2165 3355 2175
rect 3325 2145 3330 2165
rect 3350 2145 3355 2165
rect 3325 2115 3355 2145
rect 3325 2095 3330 2115
rect 3350 2095 3355 2115
rect 3325 2065 3355 2095
rect 3325 2045 3330 2065
rect 3350 2045 3355 2065
rect 3325 2015 3355 2045
rect 3325 1995 3330 2015
rect 3350 1995 3355 2015
rect 3325 1985 3355 1995
rect 3425 2165 3455 2175
rect 3425 2145 3430 2165
rect 3450 2145 3455 2165
rect 3425 2115 3455 2145
rect 3425 2095 3430 2115
rect 3450 2095 3455 2115
rect 3425 2065 3455 2095
rect 3425 2045 3430 2065
rect 3450 2045 3455 2065
rect 3425 2015 3455 2045
rect 3425 1995 3430 2015
rect 3450 1995 3455 2015
rect 3425 1985 3455 1995
rect 3525 2165 3555 2175
rect 3525 2145 3530 2165
rect 3550 2145 3555 2165
rect 3525 2115 3555 2145
rect 3525 2095 3530 2115
rect 3550 2095 3555 2115
rect 3525 2065 3555 2095
rect 3525 2045 3530 2065
rect 3550 2045 3555 2065
rect 3525 2015 3555 2045
rect 3525 1995 3530 2015
rect 3550 1995 3555 2015
rect 3525 1985 3555 1995
rect 3625 2165 3655 2175
rect 3625 2145 3630 2165
rect 3650 2145 3655 2165
rect 3625 2115 3655 2145
rect 3625 2095 3630 2115
rect 3650 2095 3655 2115
rect 3625 2065 3655 2095
rect 3625 2045 3630 2065
rect 3650 2045 3655 2065
rect 3625 2015 3655 2045
rect 3625 1995 3630 2015
rect 3650 1995 3655 2015
rect 3625 1985 3655 1995
rect 3725 2165 3755 2175
rect 3725 2145 3730 2165
rect 3750 2145 3755 2165
rect 3725 2115 3755 2145
rect 3725 2095 3730 2115
rect 3750 2095 3755 2115
rect 3725 2065 3755 2095
rect 3725 2045 3730 2065
rect 3750 2045 3755 2065
rect 3725 2015 3755 2045
rect 3725 1995 3730 2015
rect 3750 1995 3755 2015
rect 3725 1985 3755 1995
rect 3825 2165 3855 2175
rect 3825 2145 3830 2165
rect 3850 2145 3855 2165
rect 3825 2115 3855 2145
rect 3825 2095 3830 2115
rect 3850 2095 3855 2115
rect 3825 2065 3855 2095
rect 3825 2045 3830 2065
rect 3850 2045 3855 2065
rect 3825 2015 3855 2045
rect 3825 1995 3830 2015
rect 3850 1995 3855 2015
rect 3825 1985 3855 1995
rect 3925 2165 3955 2175
rect 3925 2145 3930 2165
rect 3950 2145 3955 2165
rect 3925 2115 3955 2145
rect 3925 2095 3930 2115
rect 3950 2095 3955 2115
rect 3925 2065 3955 2095
rect 3925 2045 3930 2065
rect 3950 2045 3955 2065
rect 3925 2015 3955 2045
rect 3925 1995 3930 2015
rect 3950 1995 3955 2015
rect 3925 1985 3955 1995
rect 4025 2165 4055 2175
rect 4025 2145 4030 2165
rect 4050 2145 4055 2165
rect 4025 2115 4055 2145
rect 4025 2095 4030 2115
rect 4050 2095 4055 2115
rect 4025 2065 4055 2095
rect 4025 2045 4030 2065
rect 4050 2045 4055 2065
rect 4025 2015 4055 2045
rect 4025 1995 4030 2015
rect 4050 1995 4055 2015
rect 4025 1985 4055 1995
rect 4125 2165 4155 2175
rect 4125 2145 4130 2165
rect 4150 2145 4155 2165
rect 4125 2115 4155 2145
rect 4125 2095 4130 2115
rect 4150 2095 4155 2115
rect 4125 2065 4155 2095
rect 4125 2045 4130 2065
rect 4150 2045 4155 2065
rect 4125 2015 4155 2045
rect 4125 1995 4130 2015
rect 4150 1995 4155 2015
rect 4125 1985 4155 1995
rect 4225 2165 4255 2175
rect 4225 2145 4230 2165
rect 4250 2145 4255 2165
rect 4225 2115 4255 2145
rect 4225 2095 4230 2115
rect 4250 2095 4255 2115
rect 4225 2065 4255 2095
rect 4225 2045 4230 2065
rect 4250 2045 4255 2065
rect 4225 2015 4255 2045
rect 4225 1995 4230 2015
rect 4250 1995 4255 2015
rect 4225 1985 4255 1995
rect 4325 2165 4355 2175
rect 4325 2145 4330 2165
rect 4350 2145 4355 2165
rect 4325 2115 4355 2145
rect 4325 2095 4330 2115
rect 4350 2095 4355 2115
rect 4325 2065 4355 2095
rect 4325 2045 4330 2065
rect 4350 2045 4355 2065
rect 4325 2015 4355 2045
rect 4325 1995 4330 2015
rect 4350 1995 4355 2015
rect 4325 1985 4355 1995
rect 4425 2165 4495 2175
rect 4425 2145 4430 2165
rect 4450 2145 4470 2165
rect 4490 2145 4495 2165
rect 4425 2115 4495 2145
rect 4425 2095 4430 2115
rect 4450 2095 4470 2115
rect 4490 2095 4495 2115
rect 4425 2065 4495 2095
rect 4425 2045 4430 2065
rect 4450 2045 4470 2065
rect 4490 2045 4495 2065
rect 4425 2015 4495 2045
rect 4425 1995 4430 2015
rect 4450 1995 4470 2015
rect 4490 1995 4495 2015
rect 4425 1985 4495 1995
rect 4535 2165 4565 2175
rect 4535 2145 4540 2165
rect 4560 2145 4565 2165
rect 4535 2115 4565 2145
rect 4535 2095 4540 2115
rect 4560 2095 4565 2115
rect 4535 2065 4565 2095
rect 4535 2045 4540 2065
rect 4560 2045 4565 2065
rect 4535 2015 4565 2045
rect 4535 1995 4540 2015
rect 4560 1995 4565 2015
rect 4535 1985 4565 1995
rect 4590 2165 4620 2175
rect 4590 2145 4595 2165
rect 4615 2145 4620 2165
rect 4590 2115 4620 2145
rect 4590 2095 4595 2115
rect 4615 2095 4620 2115
rect 4590 2065 4620 2095
rect 4590 2045 4595 2065
rect 4615 2045 4620 2065
rect 4590 2015 4620 2045
rect 4590 1995 4595 2015
rect 4615 1995 4620 2015
rect 4590 1985 4620 1995
rect 4660 2165 4690 2175
rect 4660 2145 4665 2165
rect 4685 2145 4690 2165
rect 4660 2115 4690 2145
rect 4660 2095 4665 2115
rect 4685 2095 4690 2115
rect 4660 2065 4690 2095
rect 4660 2045 4665 2065
rect 4685 2045 4690 2065
rect 4660 2015 4690 2045
rect 4660 1995 4665 2015
rect 4685 1995 4690 2015
rect 4660 1985 4690 1995
rect 4715 2165 4770 2175
rect 4715 2145 4720 2165
rect 4740 2145 4770 2165
rect 4715 2115 4750 2145
rect 4715 2095 4720 2115
rect 4740 2095 4750 2115
rect 4715 2065 4750 2095
rect 4715 2045 4720 2065
rect 4740 2045 4750 2065
rect 4715 2015 4750 2045
rect 4715 1995 4720 2015
rect 4740 1995 4750 2015
rect 4715 1985 4750 1995
rect 2689 1845 2769 1880
rect 3130 1860 3150 1985
rect 3330 1960 3350 1985
rect 3320 1950 3360 1960
rect 3320 1930 3330 1950
rect 3350 1930 3360 1950
rect 3320 1920 3360 1930
rect 3530 1915 3550 1985
rect 3170 1905 3210 1915
rect 3170 1885 3180 1905
rect 3200 1885 3210 1905
rect 3170 1875 3210 1885
rect 3520 1905 3560 1915
rect 3520 1885 3530 1905
rect 3550 1885 3560 1905
rect 3520 1875 3560 1885
rect 3670 1905 3710 1915
rect 3670 1885 3680 1905
rect 3700 1885 3710 1905
rect 3670 1875 3710 1885
rect 3730 1860 3750 1985
rect 3930 1915 3950 1985
rect 4130 1960 4150 1985
rect 4120 1950 4160 1960
rect 4120 1930 4130 1950
rect 4150 1930 4160 1950
rect 4120 1920 4160 1930
rect 3770 1905 3810 1915
rect 3770 1885 3780 1905
rect 3800 1885 3810 1905
rect 3770 1875 3810 1885
rect 3920 1905 3960 1915
rect 3920 1885 3930 1905
rect 3950 1885 3960 1905
rect 3920 1875 3960 1885
rect 4270 1905 4310 1915
rect 4270 1885 4280 1905
rect 4300 1885 4310 1905
rect 4270 1875 4310 1885
rect 4330 1860 4350 1985
rect 4530 1975 4570 1985
rect 4530 1955 4540 1975
rect 4560 1955 4570 1975
rect 4530 1945 4570 1955
rect 3120 1850 3160 1860
rect 1705 1820 1740 1845
rect 3120 1830 3130 1850
rect 3150 1830 3160 1850
rect 3120 1820 3160 1830
rect 3720 1850 3760 1860
rect 3720 1830 3730 1850
rect 3750 1830 3760 1850
rect 3720 1820 3760 1830
rect 4320 1850 4360 1860
rect 4320 1830 4330 1850
rect 4350 1830 4360 1850
rect 4320 1820 4360 1830
rect 2689 1785 2769 1820
rect 1665 1725 1705 1760
rect 2689 1725 2729 1760
rect 1625 1665 1705 1700
rect 2654 1640 2689 1665
rect 1660 1635 1705 1640
rect 1660 1610 1670 1635
rect 1695 1610 1705 1635
rect 1660 1605 1705 1610
rect 2709 1580 2729 1725
rect 1660 1575 1705 1580
rect 1660 1550 1670 1575
rect 1695 1550 1705 1575
rect 1660 1545 1705 1550
rect 2689 1545 2729 1580
rect 1660 1515 1705 1525
rect 2749 1520 2769 1785
rect 3320 1790 3360 1800
rect 3320 1770 3330 1790
rect 3350 1770 3360 1790
rect 3320 1760 3360 1770
rect 3720 1790 3760 1800
rect 3720 1770 3730 1790
rect 3750 1770 3760 1790
rect 3720 1760 3760 1770
rect 4120 1790 4160 1800
rect 4120 1770 4130 1790
rect 4150 1770 4160 1790
rect 4120 1760 4160 1770
rect 3330 1655 3350 1760
rect 3520 1745 3560 1755
rect 3520 1725 3530 1745
rect 3550 1725 3560 1745
rect 3520 1715 3560 1725
rect 3370 1700 3410 1710
rect 3370 1680 3380 1700
rect 3400 1680 3410 1700
rect 3370 1670 3410 1680
rect 3530 1655 3550 1715
rect 3670 1700 3710 1710
rect 3670 1680 3680 1700
rect 3700 1680 3710 1700
rect 3670 1670 3710 1680
rect 3730 1655 3750 1760
rect 3920 1745 3960 1755
rect 3920 1725 3930 1745
rect 3950 1725 3960 1745
rect 3920 1715 3960 1725
rect 3770 1700 3810 1710
rect 3770 1680 3780 1700
rect 3800 1680 3810 1700
rect 3770 1670 3810 1680
rect 3930 1655 3950 1715
rect 4070 1700 4110 1710
rect 4070 1680 4080 1700
rect 4100 1680 4110 1700
rect 4070 1670 4110 1680
rect 4130 1655 4150 1760
rect 4595 1710 4615 1985
rect 4660 1950 4680 1985
rect 4640 1940 4680 1950
rect 4640 1920 4650 1940
rect 4670 1920 4680 1940
rect 4640 1910 4680 1920
rect 4585 1700 4625 1710
rect 4585 1680 4595 1700
rect 4615 1680 4625 1700
rect 4585 1670 4625 1680
rect 3225 1645 3255 1655
rect 3225 1630 3230 1645
rect 3185 1625 3230 1630
rect 3250 1625 3255 1645
rect 3185 1620 3255 1625
rect 3185 1600 3195 1620
rect 3215 1600 3255 1620
rect 3185 1595 3255 1600
rect 3185 1590 3230 1595
rect 3225 1575 3230 1590
rect 3250 1575 3255 1595
rect 3225 1565 3255 1575
rect 3325 1645 3355 1655
rect 3325 1625 3330 1645
rect 3350 1625 3355 1645
rect 3325 1595 3355 1625
rect 3325 1575 3330 1595
rect 3350 1575 3355 1595
rect 3325 1565 3355 1575
rect 3425 1645 3455 1655
rect 3425 1625 3430 1645
rect 3450 1625 3455 1645
rect 3425 1595 3455 1625
rect 3425 1575 3430 1595
rect 3450 1575 3455 1595
rect 3425 1565 3455 1575
rect 3525 1645 3555 1655
rect 3525 1625 3530 1645
rect 3550 1625 3555 1645
rect 3525 1595 3555 1625
rect 3525 1575 3530 1595
rect 3550 1575 3555 1595
rect 3525 1565 3555 1575
rect 3625 1645 3655 1655
rect 3625 1625 3630 1645
rect 3650 1625 3655 1645
rect 3625 1595 3655 1625
rect 3625 1575 3630 1595
rect 3650 1575 3655 1595
rect 3625 1565 3655 1575
rect 3725 1645 3755 1655
rect 3725 1625 3730 1645
rect 3750 1625 3755 1645
rect 3725 1595 3755 1625
rect 3725 1575 3730 1595
rect 3750 1575 3755 1595
rect 3725 1565 3755 1575
rect 3825 1645 3855 1655
rect 3825 1625 3830 1645
rect 3850 1625 3855 1645
rect 3825 1595 3855 1625
rect 3825 1575 3830 1595
rect 3850 1575 3855 1595
rect 3825 1565 3855 1575
rect 3925 1645 3955 1655
rect 3925 1625 3930 1645
rect 3950 1625 3955 1645
rect 3925 1595 3955 1625
rect 3925 1575 3930 1595
rect 3950 1575 3955 1595
rect 3925 1565 3955 1575
rect 4025 1645 4055 1655
rect 4025 1625 4030 1645
rect 4050 1625 4055 1645
rect 4025 1595 4055 1625
rect 4025 1575 4030 1595
rect 4050 1575 4055 1595
rect 4025 1565 4055 1575
rect 4125 1645 4155 1655
rect 4125 1625 4130 1645
rect 4150 1625 4155 1645
rect 4125 1595 4155 1625
rect 4125 1575 4130 1595
rect 4150 1575 4155 1595
rect 4125 1565 4155 1575
rect 4225 1645 4255 1655
rect 4225 1625 4230 1645
rect 4250 1625 4255 1645
rect 4225 1595 4255 1625
rect 4225 1575 4230 1595
rect 4250 1575 4255 1595
rect 4225 1565 4255 1575
rect 3230 1540 3250 1565
rect 3270 1540 3310 1550
rect 3230 1520 3280 1540
rect 3300 1520 3310 1540
rect 1660 1490 1670 1515
rect 1695 1490 1705 1515
rect 1660 1480 1705 1490
rect 2689 1485 2769 1520
rect 3270 1510 3310 1520
rect 3430 1500 3450 1565
rect 3520 1535 3560 1545
rect 3520 1515 3530 1535
rect 3550 1515 3560 1535
rect 3520 1505 3560 1515
rect 3630 1500 3650 1565
rect 3830 1500 3850 1565
rect 3920 1535 3960 1545
rect 3920 1515 3930 1535
rect 3950 1515 3960 1535
rect 3920 1505 3960 1515
rect 4030 1500 4050 1565
rect 4170 1540 4210 1550
rect 4230 1540 4250 1565
rect 4170 1520 4180 1540
rect 4200 1520 4250 1540
rect 4170 1510 4210 1520
rect 3420 1490 3460 1500
rect 3420 1470 3430 1490
rect 3450 1470 3460 1490
rect 3420 1460 3460 1470
rect 3620 1490 3660 1500
rect 3620 1470 3630 1490
rect 3650 1470 3660 1490
rect 3620 1460 3660 1470
rect 3820 1490 3860 1500
rect 3820 1470 3830 1490
rect 3850 1470 3860 1490
rect 3820 1460 3860 1470
rect 4020 1490 4060 1500
rect 4020 1470 4030 1490
rect 4050 1470 4060 1490
rect 4020 1460 4060 1470
rect 3430 1440 3450 1460
rect 3630 1440 3650 1460
rect 3245 1430 3680 1440
rect 3245 1410 3290 1430
rect 3310 1410 3330 1430
rect 3350 1410 3370 1430
rect 3390 1410 3410 1430
rect 3430 1410 3450 1430
rect 3470 1410 3490 1430
rect 3510 1410 3530 1430
rect 3550 1410 3570 1430
rect 3590 1410 3610 1430
rect 3630 1410 3650 1430
rect 3670 1410 3680 1430
rect 3245 1400 3680 1410
rect 3800 1430 4240 1440
rect 3800 1410 3810 1430
rect 3830 1410 3850 1430
rect 3870 1410 3890 1430
rect 3910 1410 3930 1430
rect 3950 1410 3970 1430
rect 3990 1410 4010 1430
rect 4030 1410 4050 1430
rect 4070 1410 4090 1430
rect 4110 1410 4130 1430
rect 4150 1410 4170 1430
rect 4190 1410 4210 1430
rect 4230 1410 4240 1430
rect 3800 1400 4240 1410
rect 125 1335 2185 1375
rect 650 690 775 1335
rect 1330 690 1455 1335
rect 2060 695 2185 1335
rect 3245 1370 3275 1400
rect 3245 1350 3250 1370
rect 3270 1350 3275 1370
rect 3245 1320 3275 1350
rect 3245 1300 3250 1320
rect 3270 1300 3275 1320
rect 3245 1270 3275 1300
rect 3245 1250 3250 1270
rect 3270 1250 3275 1270
rect 3245 1220 3275 1250
rect 3245 1200 3250 1220
rect 3270 1200 3275 1220
rect 3245 1170 3275 1200
rect 3245 1150 3250 1170
rect 3270 1150 3275 1170
rect 3245 1120 3275 1150
rect 3245 1100 3250 1120
rect 3270 1100 3275 1120
rect 3245 1070 3275 1100
rect 3245 1050 3250 1070
rect 3270 1050 3275 1070
rect 3245 1020 3275 1050
rect 3245 1000 3250 1020
rect 3270 1000 3275 1020
rect 3245 990 3275 1000
rect 3685 1370 3795 1380
rect 3685 1350 3690 1370
rect 3710 1350 3730 1370
rect 3750 1350 3770 1370
rect 3790 1350 3795 1370
rect 3685 1320 3795 1350
rect 3685 1300 3690 1320
rect 3710 1300 3730 1320
rect 3750 1300 3770 1320
rect 3790 1300 3795 1320
rect 3685 1270 3795 1300
rect 3685 1250 3690 1270
rect 3710 1250 3730 1270
rect 3750 1250 3770 1270
rect 3790 1250 3795 1270
rect 3685 1220 3795 1250
rect 3685 1200 3690 1220
rect 3710 1200 3730 1220
rect 3750 1200 3770 1220
rect 3790 1200 3795 1220
rect 3685 1170 3795 1200
rect 3685 1150 3690 1170
rect 3710 1150 3730 1170
rect 3750 1150 3770 1170
rect 3790 1150 3795 1170
rect 3685 1120 3795 1150
rect 3685 1100 3690 1120
rect 3710 1100 3730 1120
rect 3750 1100 3770 1120
rect 3790 1100 3795 1120
rect 3685 1070 3795 1100
rect 3685 1050 3690 1070
rect 3710 1050 3730 1070
rect 3750 1050 3770 1070
rect 3790 1050 3795 1070
rect 3685 1020 3795 1050
rect 3685 1000 3690 1020
rect 3710 1000 3730 1020
rect 3750 1000 3770 1020
rect 3790 1000 3795 1020
rect 3685 990 3795 1000
rect 4205 1370 4235 1400
rect 4205 1350 4210 1370
rect 4230 1350 4235 1370
rect 4205 1320 4235 1350
rect 4205 1300 4210 1320
rect 4230 1300 4235 1320
rect 4205 1270 4235 1300
rect 4205 1250 4210 1270
rect 4230 1250 4235 1270
rect 4205 1220 4235 1250
rect 4205 1200 4210 1220
rect 4230 1200 4235 1220
rect 4205 1170 4235 1200
rect 4205 1150 4210 1170
rect 4230 1150 4235 1170
rect 4205 1120 4235 1150
rect 4205 1100 4210 1120
rect 4230 1100 4235 1120
rect 4205 1070 4235 1100
rect 4205 1050 4210 1070
rect 4230 1050 4235 1070
rect 4205 1020 4235 1050
rect 4205 1000 4210 1020
rect 4230 1000 4235 1020
rect 4205 990 4235 1000
rect 3690 970 3710 990
rect 3730 970 3750 990
rect 3770 970 3790 990
rect 3680 960 3800 970
rect 3680 940 3690 960
rect 3710 940 3730 960
rect 3750 940 3770 960
rect 3790 940 3800 960
rect 3680 930 3800 940
rect 3200 900 4270 910
rect 3200 880 3240 900
rect 3260 880 3320 900
rect 3340 880 3400 900
rect 3420 880 3480 900
rect 3500 880 3560 900
rect 3580 880 3640 900
rect 3660 880 3720 900
rect 3740 880 3800 900
rect 3820 880 3880 900
rect 3900 880 3960 900
rect 3980 880 4040 900
rect 4060 880 4120 900
rect 4140 880 4200 900
rect 4220 880 4240 900
rect 4260 880 4270 900
rect 3200 870 4270 880
rect 3200 850 3220 870
rect 3195 840 3225 850
rect 3195 820 3200 840
rect 3220 820 3225 840
rect 3195 790 3225 820
rect 3195 770 3200 790
rect 3220 770 3225 790
rect 3195 760 3225 770
rect 4235 840 4305 850
rect 4235 820 4240 840
rect 4260 820 4280 840
rect 4300 825 4305 840
rect 4300 820 4345 825
rect 4235 815 4345 820
rect 4235 795 4315 815
rect 4335 795 4345 815
rect 4235 790 4345 795
rect 4235 770 4240 790
rect 4260 770 4280 790
rect 4300 785 4345 790
rect 4300 770 4305 785
rect 4235 760 4305 770
<< viali >>
rect 3030 2825 3050 2845
rect 3230 2825 3250 2845
rect 3430 2825 3450 2845
rect 3630 2825 3650 2845
rect 3730 2825 3750 2845
rect 3830 2825 3850 2845
rect 4030 2825 4050 2845
rect 4230 2825 4250 2845
rect 4430 2825 4450 2845
rect 1670 2570 1695 2595
rect 1670 2510 1695 2535
rect 1670 2450 1695 2475
rect 3530 2355 3550 2375
rect 3340 2310 3360 2330
rect 3930 2355 3950 2375
rect 4280 2355 4300 2375
rect 4120 2310 4140 2330
rect 3130 2265 3150 2285
rect 3730 2265 3750 2285
rect 4330 2265 4350 2285
rect 4540 2255 4560 2275
rect 1530 2030 1555 2055
rect 1670 2030 1695 2055
rect 2489 2030 2514 2055
rect -35 1695 -15 1715
rect 3030 2205 3050 2225
rect 3230 2205 3250 2225
rect 3430 2205 3450 2225
rect 3630 2205 3650 2225
rect 3830 2205 3850 2225
rect 4030 2205 4050 2225
rect 4230 2205 4250 2225
rect 4430 2205 4450 2225
rect 4750 2205 4770 2225
rect 3330 1930 3350 1950
rect 3180 1885 3200 1905
rect 3530 1885 3550 1905
rect 3680 1885 3700 1905
rect 4130 1930 4150 1950
rect 3780 1885 3800 1905
rect 3930 1885 3950 1905
rect 4280 1885 4300 1905
rect 4540 1955 4560 1975
rect 3130 1830 3150 1850
rect 3730 1830 3750 1850
rect 4330 1830 4350 1850
rect 1670 1610 1695 1635
rect 1670 1550 1695 1575
rect 3330 1770 3350 1790
rect 3730 1770 3750 1790
rect 4130 1770 4150 1790
rect 3530 1725 3550 1745
rect 3380 1680 3400 1700
rect 3680 1680 3700 1700
rect 3930 1725 3950 1745
rect 3780 1680 3800 1700
rect 4080 1680 4100 1700
rect 4650 1920 4670 1940
rect 4595 1680 4615 1700
rect 3195 1600 3215 1620
rect 1670 1490 1695 1515
rect 3530 1515 3550 1535
rect 3930 1515 3950 1535
rect 4180 1520 4200 1540
rect 3430 1470 3450 1490
rect 3630 1470 3650 1490
rect 3830 1470 3850 1490
rect 4030 1470 4050 1490
rect 4210 1410 4230 1430
rect 3690 940 3710 960
rect 3730 940 3750 960
rect 3770 940 3790 960
rect 4240 880 4260 900
rect 4315 795 4335 815
<< metal1 >>
rect 1555 2900 1705 2910
rect 1555 2870 1565 2900
rect 1595 2870 1615 2900
rect 1645 2870 1665 2900
rect 1695 2870 1705 2900
rect 1555 2860 1705 2870
rect 275 2200 1520 2550
rect 1570 2480 1590 2860
rect 1620 2540 1640 2860
rect 1670 2600 1690 2860
rect 3730 2855 3750 3175
rect 3020 2850 3060 2855
rect 3020 2820 3025 2850
rect 3055 2820 3060 2850
rect 3020 2815 3060 2820
rect 3220 2850 3260 2855
rect 3220 2820 3225 2850
rect 3255 2820 3260 2850
rect 3220 2815 3260 2820
rect 3420 2850 3460 2855
rect 3420 2820 3425 2850
rect 3455 2820 3460 2850
rect 3420 2815 3460 2820
rect 3620 2850 3660 2855
rect 3620 2820 3625 2850
rect 3655 2820 3660 2850
rect 3620 2815 3660 2820
rect 3720 2845 3760 2855
rect 3720 2825 3730 2845
rect 3750 2825 3760 2845
rect 3720 2815 3760 2825
rect 3820 2850 3860 2855
rect 3820 2820 3825 2850
rect 3855 2820 3860 2850
rect 3820 2815 3860 2820
rect 4020 2850 4060 2855
rect 4020 2820 4025 2850
rect 4055 2820 4060 2850
rect 4020 2815 4060 2820
rect 4220 2850 4260 2855
rect 4220 2820 4225 2850
rect 4255 2820 4260 2850
rect 4220 2815 4260 2820
rect 4420 2850 4460 2855
rect 4420 2820 4425 2850
rect 4455 2820 4460 2850
rect 4420 2815 4460 2820
rect 1660 2565 1665 2600
rect 1700 2565 1705 2600
rect 1610 2535 1645 2540
rect 1610 2505 1615 2535
rect 1660 2505 1665 2540
rect 1700 2505 1705 2540
rect 1610 2500 1645 2505
rect 1560 2475 1600 2480
rect 1560 2445 1565 2475
rect 1595 2445 1600 2475
rect 1660 2445 1665 2480
rect 1700 2445 1705 2480
rect 1560 2440 1600 2445
rect 2855 2380 2895 2385
rect 2855 2350 2860 2380
rect 2890 2350 2895 2380
rect 2855 2345 2895 2350
rect 3520 2380 3560 2385
rect 3520 2350 3525 2380
rect 3555 2350 3560 2380
rect 3520 2345 3560 2350
rect 3920 2380 3960 2385
rect 3920 2350 3925 2380
rect 3955 2350 3960 2380
rect 3920 2345 3960 2350
rect 4270 2380 4310 2385
rect 4270 2350 4275 2380
rect 4305 2350 4310 2380
rect 4270 2345 4310 2350
rect 4530 2380 4570 2385
rect 4530 2350 4535 2380
rect 4565 2350 4570 2380
rect 4530 2345 4570 2350
rect 2800 2290 2840 2295
rect 2800 2260 2805 2290
rect 2835 2260 2840 2290
rect 2800 2255 2840 2260
rect 1485 2060 1520 2200
rect 1485 2025 1525 2060
rect 1560 2025 1565 2060
rect 1660 2025 1665 2060
rect 1700 2025 1705 2060
rect 2479 2025 2484 2060
rect 2519 2025 2524 2060
rect 1485 1870 1520 2025
rect -110 1720 -70 1725
rect -110 1690 -105 1720
rect -75 1715 -70 1720
rect -45 1720 -5 1725
rect -45 1715 -40 1720
rect -75 1695 -40 1715
rect -75 1690 -70 1695
rect -110 1685 -70 1690
rect -45 1690 -40 1695
rect -10 1690 -5 1720
rect -45 1685 -5 1690
rect 275 1520 1520 1870
rect 1550 1635 1590 1640
rect 1550 1605 1555 1635
rect 1585 1605 1590 1635
rect 1660 1605 1665 1640
rect 1700 1605 1705 1640
rect 1550 1600 1590 1605
rect 1485 1190 1520 1520
rect 1560 1400 1580 1600
rect 1605 1575 1645 1580
rect 1605 1545 1610 1575
rect 1640 1545 1645 1575
rect 1660 1545 1665 1580
rect 1700 1545 1705 1580
rect 1605 1540 1645 1545
rect 1615 1445 1635 1540
rect 1660 1520 1705 1525
rect 1660 1485 1665 1520
rect 1700 1485 1705 1520
rect 2810 1490 2830 2255
rect 2865 1710 2885 2345
rect 2910 2335 2950 2340
rect 2910 2305 2915 2335
rect 2945 2305 2950 2335
rect 2910 2300 2950 2305
rect 3330 2335 3370 2340
rect 3330 2305 3335 2335
rect 3365 2305 3370 2335
rect 3330 2300 3370 2305
rect 4110 2335 4150 2340
rect 4110 2305 4115 2335
rect 4145 2305 4150 2335
rect 4110 2300 4150 2305
rect 2920 2060 2940 2300
rect 3120 2290 3160 2295
rect 3120 2260 3125 2290
rect 3155 2260 3160 2290
rect 3120 2255 3160 2260
rect 3720 2290 3760 2295
rect 3720 2260 3725 2290
rect 3755 2260 3760 2290
rect 3720 2255 3760 2260
rect 4320 2290 4360 2295
rect 4320 2260 4325 2290
rect 4355 2260 4360 2290
rect 4540 2285 4560 2345
rect 4320 2255 4360 2260
rect 4530 2275 4570 2285
rect 4530 2255 4540 2275
rect 4560 2255 4570 2275
rect 4530 2245 4570 2255
rect 3020 2230 3060 2235
rect 3020 2200 3025 2230
rect 3055 2200 3060 2230
rect 3020 2195 3060 2200
rect 3220 2230 3260 2235
rect 3220 2200 3225 2230
rect 3255 2200 3260 2230
rect 3220 2195 3260 2200
rect 3420 2230 3460 2235
rect 3420 2200 3425 2230
rect 3455 2200 3460 2230
rect 3420 2195 3460 2200
rect 3620 2230 3660 2235
rect 3620 2200 3625 2230
rect 3655 2200 3660 2230
rect 3620 2195 3660 2200
rect 3820 2230 3860 2235
rect 3820 2200 3825 2230
rect 3855 2200 3860 2230
rect 3820 2195 3860 2200
rect 4020 2230 4060 2235
rect 4020 2200 4025 2230
rect 4055 2200 4060 2230
rect 4020 2195 4060 2200
rect 4220 2230 4260 2235
rect 4220 2200 4225 2230
rect 4255 2200 4260 2230
rect 4220 2195 4260 2200
rect 4420 2230 4460 2235
rect 4420 2200 4425 2230
rect 4455 2200 4460 2230
rect 4420 2195 4460 2200
rect 4740 2230 4780 2235
rect 4740 2200 4745 2230
rect 4775 2200 4780 2230
rect 4740 2195 4780 2200
rect 2910 2055 2950 2060
rect 2910 2025 2915 2055
rect 2945 2025 2950 2055
rect 2910 2020 2950 2025
rect 2855 1705 2895 1710
rect 2855 1675 2860 1705
rect 2890 1675 2895 1705
rect 2855 1670 2895 1675
rect 1660 1480 1705 1485
rect 2800 1485 2840 1490
rect 2800 1455 2805 1485
rect 2835 1455 2840 1485
rect 2800 1450 2840 1455
rect 2865 1445 2885 1670
rect 2920 1545 2940 2020
rect 4530 1980 4570 1985
rect 3320 1955 3360 1960
rect 3320 1925 3325 1955
rect 3355 1925 3360 1955
rect 3320 1920 3360 1925
rect 4120 1955 4160 1960
rect 4120 1925 4125 1955
rect 4155 1925 4160 1955
rect 4530 1950 4535 1980
rect 4565 1950 4570 1980
rect 4530 1945 4570 1950
rect 4120 1920 4160 1925
rect 3170 1910 3210 1915
rect 3170 1880 3175 1910
rect 3205 1880 3210 1910
rect 3170 1875 3210 1880
rect 3120 1855 3160 1860
rect 3120 1825 3125 1855
rect 3155 1825 3160 1855
rect 3120 1820 3160 1825
rect 3330 1800 3350 1920
rect 3520 1910 3560 1915
rect 3520 1880 3525 1910
rect 3555 1880 3560 1910
rect 3520 1875 3560 1880
rect 3670 1910 3710 1915
rect 3670 1880 3675 1910
rect 3705 1880 3710 1910
rect 3670 1875 3710 1880
rect 3770 1910 3810 1915
rect 3770 1880 3775 1910
rect 3805 1880 3810 1910
rect 3770 1875 3810 1880
rect 3920 1910 3960 1915
rect 3920 1880 3925 1910
rect 3955 1880 3960 1910
rect 3920 1875 3960 1880
rect 4270 1910 4310 1915
rect 4270 1880 4275 1910
rect 4305 1880 4310 1910
rect 4270 1875 4310 1880
rect 3720 1855 3760 1860
rect 3720 1825 3725 1855
rect 3755 1825 3760 1855
rect 3720 1820 3760 1825
rect 3320 1795 3360 1800
rect 3320 1765 3325 1795
rect 3355 1765 3360 1795
rect 3320 1760 3360 1765
rect 3720 1795 3760 1800
rect 3720 1765 3725 1795
rect 3755 1765 3760 1795
rect 3720 1760 3760 1765
rect 3930 1755 3950 1875
rect 4540 1860 4560 1945
rect 4640 1940 4680 1950
rect 4640 1920 4650 1940
rect 4670 1920 4680 1940
rect 4640 1910 4680 1920
rect 4320 1855 4360 1860
rect 4320 1825 4325 1855
rect 4355 1825 4360 1855
rect 4320 1820 4360 1825
rect 4530 1855 4570 1860
rect 4530 1825 4535 1855
rect 4565 1825 4570 1855
rect 4530 1820 4570 1825
rect 4120 1795 4160 1800
rect 4120 1765 4125 1795
rect 4155 1765 4160 1795
rect 4120 1760 4160 1765
rect 3520 1750 3560 1755
rect 3520 1720 3525 1750
rect 3555 1720 3560 1750
rect 3520 1715 3560 1720
rect 3920 1750 3960 1755
rect 3920 1720 3925 1750
rect 3955 1720 3960 1750
rect 3920 1715 3960 1720
rect 3370 1705 3410 1710
rect 3370 1675 3375 1705
rect 3405 1675 3410 1705
rect 3370 1670 3410 1675
rect 3670 1705 3710 1710
rect 3670 1675 3675 1705
rect 3705 1675 3710 1705
rect 3670 1670 3710 1675
rect 3770 1705 3810 1710
rect 3770 1675 3775 1705
rect 3805 1675 3810 1705
rect 3770 1670 3810 1675
rect 4070 1705 4110 1710
rect 4070 1675 4075 1705
rect 4105 1675 4110 1705
rect 4070 1670 4110 1675
rect 3105 1625 3145 1630
rect 3105 1595 3110 1625
rect 3140 1595 3145 1625
rect 3105 1590 3145 1595
rect 3185 1625 3225 1630
rect 3185 1595 3190 1625
rect 3220 1595 3225 1625
rect 3185 1590 3225 1595
rect 2910 1540 2950 1545
rect 2910 1510 2915 1540
rect 2945 1510 2950 1540
rect 2910 1505 2950 1510
rect 1605 1440 1645 1445
rect 1605 1410 1610 1440
rect 1640 1410 1645 1440
rect 1605 1405 1645 1410
rect 2855 1440 2895 1445
rect 2855 1410 2860 1440
rect 2890 1410 2895 1440
rect 2855 1405 2895 1410
rect 1550 1395 1590 1400
rect 1550 1365 1555 1395
rect 1585 1365 1590 1395
rect 1550 1360 1590 1365
rect 275 840 1520 1190
rect 1685 1035 2225 1190
rect 2865 1035 2885 1405
rect 2920 1400 2940 1505
rect 2910 1395 2950 1400
rect 2910 1365 2915 1395
rect 2945 1365 2950 1395
rect 2910 1360 2950 1365
rect 1685 1030 2265 1035
rect 1685 1000 2230 1030
rect 2260 1000 2265 1030
rect 1685 995 2265 1000
rect 2855 1030 2895 1035
rect 2855 1000 2860 1030
rect 2890 1000 2895 1030
rect 2855 995 2895 1000
rect 1685 840 2225 995
rect 3115 640 3135 1590
rect 4170 1545 4210 1550
rect 3520 1540 3560 1545
rect 3520 1510 3525 1540
rect 3555 1510 3560 1540
rect 3520 1505 3560 1510
rect 3920 1540 3960 1545
rect 3920 1510 3925 1540
rect 3955 1510 3960 1540
rect 4170 1515 4175 1545
rect 4205 1515 4210 1545
rect 4170 1510 4210 1515
rect 3920 1505 3960 1510
rect 3420 1495 3460 1500
rect 3420 1465 3425 1495
rect 3455 1465 3460 1495
rect 3420 1460 3460 1465
rect 3620 1495 3660 1500
rect 3620 1465 3625 1495
rect 3655 1465 3660 1495
rect 3620 1460 3660 1465
rect 3820 1495 3860 1500
rect 3820 1465 3825 1495
rect 3855 1465 3860 1495
rect 3820 1460 3860 1465
rect 4020 1495 4060 1500
rect 4020 1465 4025 1495
rect 4055 1465 4060 1495
rect 4020 1460 4060 1465
rect 4330 1440 4350 1820
rect 4585 1705 4625 1710
rect 4585 1675 4590 1705
rect 4620 1675 4625 1705
rect 4585 1670 4625 1675
rect 4200 1435 4240 1440
rect 4200 1405 4205 1435
rect 4235 1405 4240 1435
rect 4200 1400 4240 1405
rect 4320 1435 4360 1440
rect 4320 1405 4325 1435
rect 4355 1405 4360 1435
rect 4320 1400 4360 1405
rect 3680 965 3800 970
rect 3680 935 3685 965
rect 3715 935 3725 965
rect 3755 935 3765 965
rect 3795 935 3800 965
rect 3680 930 3800 935
rect 4660 910 4680 1910
rect 4230 905 4270 910
rect 4230 875 4235 905
rect 4265 875 4270 905
rect 4230 870 4270 875
rect 4650 905 4690 910
rect 4650 875 4655 905
rect 4685 875 4690 905
rect 4650 870 4690 875
rect 4305 820 4345 825
rect 4305 790 4310 820
rect 4340 790 4345 820
rect 4305 785 4345 790
rect 3100 630 3150 640
rect 3100 600 3110 630
rect 3140 600 3150 630
rect 3100 590 3150 600
<< via1 >>
rect 1565 2870 1595 2900
rect 1615 2870 1645 2900
rect 1665 2870 1695 2900
rect 3025 2845 3055 2850
rect 3025 2825 3030 2845
rect 3030 2825 3050 2845
rect 3050 2825 3055 2845
rect 3025 2820 3055 2825
rect 3225 2845 3255 2850
rect 3225 2825 3230 2845
rect 3230 2825 3250 2845
rect 3250 2825 3255 2845
rect 3225 2820 3255 2825
rect 3425 2845 3455 2850
rect 3425 2825 3430 2845
rect 3430 2825 3450 2845
rect 3450 2825 3455 2845
rect 3425 2820 3455 2825
rect 3625 2845 3655 2850
rect 3625 2825 3630 2845
rect 3630 2825 3650 2845
rect 3650 2825 3655 2845
rect 3625 2820 3655 2825
rect 3825 2845 3855 2850
rect 3825 2825 3830 2845
rect 3830 2825 3850 2845
rect 3850 2825 3855 2845
rect 3825 2820 3855 2825
rect 4025 2845 4055 2850
rect 4025 2825 4030 2845
rect 4030 2825 4050 2845
rect 4050 2825 4055 2845
rect 4025 2820 4055 2825
rect 4225 2845 4255 2850
rect 4225 2825 4230 2845
rect 4230 2825 4250 2845
rect 4250 2825 4255 2845
rect 4225 2820 4255 2825
rect 4425 2845 4455 2850
rect 4425 2825 4430 2845
rect 4430 2825 4450 2845
rect 4450 2825 4455 2845
rect 4425 2820 4455 2825
rect 1665 2595 1700 2600
rect 1665 2570 1670 2595
rect 1670 2570 1695 2595
rect 1695 2570 1700 2595
rect 1665 2565 1700 2570
rect 1615 2505 1645 2535
rect 1665 2535 1700 2540
rect 1665 2510 1670 2535
rect 1670 2510 1695 2535
rect 1695 2510 1700 2535
rect 1665 2505 1700 2510
rect 1565 2445 1595 2475
rect 1665 2475 1700 2480
rect 1665 2450 1670 2475
rect 1670 2450 1695 2475
rect 1695 2450 1700 2475
rect 1665 2445 1700 2450
rect 2860 2350 2890 2380
rect 3525 2375 3555 2380
rect 3525 2355 3530 2375
rect 3530 2355 3550 2375
rect 3550 2355 3555 2375
rect 3525 2350 3555 2355
rect 3925 2375 3955 2380
rect 3925 2355 3930 2375
rect 3930 2355 3950 2375
rect 3950 2355 3955 2375
rect 3925 2350 3955 2355
rect 4275 2375 4305 2380
rect 4275 2355 4280 2375
rect 4280 2355 4300 2375
rect 4300 2355 4305 2375
rect 4275 2350 4305 2355
rect 4535 2350 4565 2380
rect 2805 2260 2835 2290
rect 1525 2055 1560 2060
rect 1525 2030 1530 2055
rect 1530 2030 1555 2055
rect 1555 2030 1560 2055
rect 1525 2025 1560 2030
rect 1665 2055 1700 2060
rect 1665 2030 1670 2055
rect 1670 2030 1695 2055
rect 1695 2030 1700 2055
rect 1665 2025 1700 2030
rect 2484 2055 2519 2060
rect 2484 2030 2489 2055
rect 2489 2030 2514 2055
rect 2514 2030 2519 2055
rect 2484 2025 2519 2030
rect -105 1690 -75 1720
rect -40 1715 -10 1720
rect -40 1695 -35 1715
rect -35 1695 -15 1715
rect -15 1695 -10 1715
rect -40 1690 -10 1695
rect 1555 1605 1585 1635
rect 1665 1635 1700 1640
rect 1665 1610 1670 1635
rect 1670 1610 1695 1635
rect 1695 1610 1700 1635
rect 1665 1605 1700 1610
rect 1610 1545 1640 1575
rect 1665 1575 1700 1580
rect 1665 1550 1670 1575
rect 1670 1550 1695 1575
rect 1695 1550 1700 1575
rect 1665 1545 1700 1550
rect 1665 1515 1700 1520
rect 1665 1490 1670 1515
rect 1670 1490 1695 1515
rect 1695 1490 1700 1515
rect 1665 1485 1700 1490
rect 2915 2305 2945 2335
rect 3335 2330 3365 2335
rect 3335 2310 3340 2330
rect 3340 2310 3360 2330
rect 3360 2310 3365 2330
rect 3335 2305 3365 2310
rect 4115 2330 4145 2335
rect 4115 2310 4120 2330
rect 4120 2310 4140 2330
rect 4140 2310 4145 2330
rect 4115 2305 4145 2310
rect 3125 2285 3155 2290
rect 3125 2265 3130 2285
rect 3130 2265 3150 2285
rect 3150 2265 3155 2285
rect 3125 2260 3155 2265
rect 3725 2285 3755 2290
rect 3725 2265 3730 2285
rect 3730 2265 3750 2285
rect 3750 2265 3755 2285
rect 3725 2260 3755 2265
rect 4325 2285 4355 2290
rect 4325 2265 4330 2285
rect 4330 2265 4350 2285
rect 4350 2265 4355 2285
rect 4325 2260 4355 2265
rect 3025 2225 3055 2230
rect 3025 2205 3030 2225
rect 3030 2205 3050 2225
rect 3050 2205 3055 2225
rect 3025 2200 3055 2205
rect 3225 2225 3255 2230
rect 3225 2205 3230 2225
rect 3230 2205 3250 2225
rect 3250 2205 3255 2225
rect 3225 2200 3255 2205
rect 3425 2225 3455 2230
rect 3425 2205 3430 2225
rect 3430 2205 3450 2225
rect 3450 2205 3455 2225
rect 3425 2200 3455 2205
rect 3625 2225 3655 2230
rect 3625 2205 3630 2225
rect 3630 2205 3650 2225
rect 3650 2205 3655 2225
rect 3625 2200 3655 2205
rect 3825 2225 3855 2230
rect 3825 2205 3830 2225
rect 3830 2205 3850 2225
rect 3850 2205 3855 2225
rect 3825 2200 3855 2205
rect 4025 2225 4055 2230
rect 4025 2205 4030 2225
rect 4030 2205 4050 2225
rect 4050 2205 4055 2225
rect 4025 2200 4055 2205
rect 4225 2225 4255 2230
rect 4225 2205 4230 2225
rect 4230 2205 4250 2225
rect 4250 2205 4255 2225
rect 4225 2200 4255 2205
rect 4425 2225 4455 2230
rect 4425 2205 4430 2225
rect 4430 2205 4450 2225
rect 4450 2205 4455 2225
rect 4425 2200 4455 2205
rect 4745 2225 4775 2230
rect 4745 2205 4750 2225
rect 4750 2205 4770 2225
rect 4770 2205 4775 2225
rect 4745 2200 4775 2205
rect 2915 2025 2945 2055
rect 2860 1675 2890 1705
rect 2805 1455 2835 1485
rect 3325 1950 3355 1955
rect 3325 1930 3330 1950
rect 3330 1930 3350 1950
rect 3350 1930 3355 1950
rect 3325 1925 3355 1930
rect 4125 1950 4155 1955
rect 4125 1930 4130 1950
rect 4130 1930 4150 1950
rect 4150 1930 4155 1950
rect 4125 1925 4155 1930
rect 4535 1975 4565 1980
rect 4535 1955 4540 1975
rect 4540 1955 4560 1975
rect 4560 1955 4565 1975
rect 4535 1950 4565 1955
rect 3175 1905 3205 1910
rect 3175 1885 3180 1905
rect 3180 1885 3200 1905
rect 3200 1885 3205 1905
rect 3175 1880 3205 1885
rect 3125 1850 3155 1855
rect 3125 1830 3130 1850
rect 3130 1830 3150 1850
rect 3150 1830 3155 1850
rect 3125 1825 3155 1830
rect 3525 1905 3555 1910
rect 3525 1885 3530 1905
rect 3530 1885 3550 1905
rect 3550 1885 3555 1905
rect 3525 1880 3555 1885
rect 3675 1905 3705 1910
rect 3675 1885 3680 1905
rect 3680 1885 3700 1905
rect 3700 1885 3705 1905
rect 3675 1880 3705 1885
rect 3775 1905 3805 1910
rect 3775 1885 3780 1905
rect 3780 1885 3800 1905
rect 3800 1885 3805 1905
rect 3775 1880 3805 1885
rect 3925 1905 3955 1910
rect 3925 1885 3930 1905
rect 3930 1885 3950 1905
rect 3950 1885 3955 1905
rect 3925 1880 3955 1885
rect 4275 1905 4305 1910
rect 4275 1885 4280 1905
rect 4280 1885 4300 1905
rect 4300 1885 4305 1905
rect 4275 1880 4305 1885
rect 3725 1850 3755 1855
rect 3725 1830 3730 1850
rect 3730 1830 3750 1850
rect 3750 1830 3755 1850
rect 3725 1825 3755 1830
rect 3325 1790 3355 1795
rect 3325 1770 3330 1790
rect 3330 1770 3350 1790
rect 3350 1770 3355 1790
rect 3325 1765 3355 1770
rect 3725 1790 3755 1795
rect 3725 1770 3730 1790
rect 3730 1770 3750 1790
rect 3750 1770 3755 1790
rect 3725 1765 3755 1770
rect 4325 1850 4355 1855
rect 4325 1830 4330 1850
rect 4330 1830 4350 1850
rect 4350 1830 4355 1850
rect 4325 1825 4355 1830
rect 4535 1825 4565 1855
rect 4125 1790 4155 1795
rect 4125 1770 4130 1790
rect 4130 1770 4150 1790
rect 4150 1770 4155 1790
rect 4125 1765 4155 1770
rect 3525 1745 3555 1750
rect 3525 1725 3530 1745
rect 3530 1725 3550 1745
rect 3550 1725 3555 1745
rect 3525 1720 3555 1725
rect 3925 1745 3955 1750
rect 3925 1725 3930 1745
rect 3930 1725 3950 1745
rect 3950 1725 3955 1745
rect 3925 1720 3955 1725
rect 3375 1700 3405 1705
rect 3375 1680 3380 1700
rect 3380 1680 3400 1700
rect 3400 1680 3405 1700
rect 3375 1675 3405 1680
rect 3675 1700 3705 1705
rect 3675 1680 3680 1700
rect 3680 1680 3700 1700
rect 3700 1680 3705 1700
rect 3675 1675 3705 1680
rect 3775 1700 3805 1705
rect 3775 1680 3780 1700
rect 3780 1680 3800 1700
rect 3800 1680 3805 1700
rect 3775 1675 3805 1680
rect 4075 1700 4105 1705
rect 4075 1680 4080 1700
rect 4080 1680 4100 1700
rect 4100 1680 4105 1700
rect 4075 1675 4105 1680
rect 3110 1595 3140 1625
rect 3190 1620 3220 1625
rect 3190 1600 3195 1620
rect 3195 1600 3215 1620
rect 3215 1600 3220 1620
rect 3190 1595 3220 1600
rect 2915 1510 2945 1540
rect 1610 1410 1640 1440
rect 2860 1410 2890 1440
rect 1555 1365 1585 1395
rect 2915 1365 2945 1395
rect 2230 1000 2260 1030
rect 2860 1000 2890 1030
rect 3525 1535 3555 1540
rect 3525 1515 3530 1535
rect 3530 1515 3550 1535
rect 3550 1515 3555 1535
rect 3525 1510 3555 1515
rect 3925 1535 3955 1540
rect 3925 1515 3930 1535
rect 3930 1515 3950 1535
rect 3950 1515 3955 1535
rect 3925 1510 3955 1515
rect 4175 1540 4205 1545
rect 4175 1520 4180 1540
rect 4180 1520 4200 1540
rect 4200 1520 4205 1540
rect 4175 1515 4205 1520
rect 3425 1490 3455 1495
rect 3425 1470 3430 1490
rect 3430 1470 3450 1490
rect 3450 1470 3455 1490
rect 3425 1465 3455 1470
rect 3625 1490 3655 1495
rect 3625 1470 3630 1490
rect 3630 1470 3650 1490
rect 3650 1470 3655 1490
rect 3625 1465 3655 1470
rect 3825 1490 3855 1495
rect 3825 1470 3830 1490
rect 3830 1470 3850 1490
rect 3850 1470 3855 1490
rect 3825 1465 3855 1470
rect 4025 1490 4055 1495
rect 4025 1470 4030 1490
rect 4030 1470 4050 1490
rect 4050 1470 4055 1490
rect 4025 1465 4055 1470
rect 4590 1700 4620 1705
rect 4590 1680 4595 1700
rect 4595 1680 4615 1700
rect 4615 1680 4620 1700
rect 4590 1675 4620 1680
rect 4205 1430 4235 1435
rect 4205 1410 4210 1430
rect 4210 1410 4230 1430
rect 4230 1410 4235 1430
rect 4205 1405 4235 1410
rect 4325 1405 4355 1435
rect 3685 960 3715 965
rect 3685 940 3690 960
rect 3690 940 3710 960
rect 3710 940 3715 960
rect 3685 935 3715 940
rect 3725 960 3755 965
rect 3725 940 3730 960
rect 3730 940 3750 960
rect 3750 940 3755 960
rect 3725 935 3755 940
rect 3765 960 3795 965
rect 3765 940 3770 960
rect 3770 940 3790 960
rect 3790 940 3795 960
rect 3765 935 3795 940
rect 4235 900 4265 905
rect 4235 880 4240 900
rect 4240 880 4260 900
rect 4260 880 4265 900
rect 4235 875 4265 880
rect 4655 875 4685 905
rect 4310 815 4340 820
rect 4310 795 4315 815
rect 4315 795 4335 815
rect 4335 795 4340 815
rect 4310 790 4340 795
rect 3110 600 3140 630
<< metal2 >>
rect -195 2985 -155 2990
rect -195 2955 -190 2985
rect -160 2955 -155 2985
rect -195 2950 -155 2955
rect 4875 2985 4915 2990
rect 4875 2955 4880 2985
rect 4910 2955 4915 2985
rect 4875 2950 4915 2955
rect 1555 2900 1705 2910
rect 1555 2870 1565 2900
rect 1595 2870 1615 2900
rect 1645 2870 1665 2900
rect 1695 2870 1705 2900
rect 1555 2860 1705 2870
rect -195 2850 -155 2855
rect -195 2820 -190 2850
rect -160 2845 -155 2850
rect 3020 2850 3060 2855
rect 3020 2845 3025 2850
rect -160 2825 3025 2845
rect -160 2820 -155 2825
rect -195 2815 -155 2820
rect 3020 2820 3025 2825
rect 3055 2845 3060 2850
rect 3220 2850 3260 2855
rect 3220 2845 3225 2850
rect 3055 2825 3225 2845
rect 3055 2820 3060 2825
rect 3020 2815 3060 2820
rect 3220 2820 3225 2825
rect 3255 2845 3260 2850
rect 3420 2850 3460 2855
rect 3420 2845 3425 2850
rect 3255 2825 3425 2845
rect 3255 2820 3260 2825
rect 3220 2815 3260 2820
rect 3420 2820 3425 2825
rect 3455 2845 3460 2850
rect 3620 2850 3660 2855
rect 3620 2845 3625 2850
rect 3455 2825 3625 2845
rect 3455 2820 3460 2825
rect 3420 2815 3460 2820
rect 3620 2820 3625 2825
rect 3655 2845 3660 2850
rect 3820 2850 3860 2855
rect 3820 2845 3825 2850
rect 3655 2825 3825 2845
rect 3655 2820 3660 2825
rect 3620 2815 3660 2820
rect 3820 2820 3825 2825
rect 3855 2845 3860 2850
rect 4020 2850 4060 2855
rect 4020 2845 4025 2850
rect 3855 2825 4025 2845
rect 3855 2820 3860 2825
rect 3820 2815 3860 2820
rect 4020 2820 4025 2825
rect 4055 2845 4060 2850
rect 4220 2850 4260 2855
rect 4220 2845 4225 2850
rect 4055 2825 4225 2845
rect 4055 2820 4060 2825
rect 4020 2815 4060 2820
rect 4220 2820 4225 2825
rect 4255 2845 4260 2850
rect 4420 2850 4460 2855
rect 4420 2845 4425 2850
rect 4255 2825 4425 2845
rect 4255 2820 4260 2825
rect 4220 2815 4260 2820
rect 4420 2820 4425 2825
rect 4455 2845 4460 2850
rect 4875 2850 4915 2855
rect 4875 2845 4880 2850
rect 4455 2825 4880 2845
rect 4455 2820 4460 2825
rect 4420 2815 4460 2820
rect 4875 2820 4880 2825
rect 4910 2820 4915 2850
rect 4875 2815 4915 2820
rect 1660 2565 1665 2600
rect 1700 2565 1705 2600
rect 1610 2535 1645 2540
rect 1660 2535 1665 2540
rect 1610 2505 1615 2535
rect 1645 2510 1665 2535
rect 1660 2505 1665 2510
rect 1700 2505 1705 2540
rect 1610 2500 1645 2505
rect 1560 2475 1600 2480
rect 1660 2475 1665 2480
rect 1560 2445 1565 2475
rect 1595 2450 1665 2475
rect 1595 2445 1600 2450
rect 1660 2445 1665 2450
rect 1700 2445 1705 2480
rect 1560 2440 1600 2445
rect 2855 2380 2895 2385
rect 2855 2350 2860 2380
rect 2890 2375 2895 2380
rect 3520 2380 3560 2385
rect 3520 2375 3525 2380
rect 2890 2355 3525 2375
rect 2890 2350 2895 2355
rect 2855 2345 2895 2350
rect 3520 2350 3525 2355
rect 3555 2375 3560 2380
rect 3920 2380 3960 2385
rect 3920 2375 3925 2380
rect 3555 2355 3925 2375
rect 3555 2350 3560 2355
rect 3520 2345 3560 2350
rect 3920 2350 3925 2355
rect 3955 2350 3960 2380
rect 3920 2345 3960 2350
rect 4270 2380 4310 2385
rect 4270 2350 4275 2380
rect 4305 2375 4310 2380
rect 4530 2380 4570 2385
rect 4530 2375 4535 2380
rect 4305 2355 4535 2375
rect 4305 2350 4310 2355
rect 4270 2345 4310 2350
rect 4530 2350 4535 2355
rect 4565 2350 4570 2380
rect 4530 2345 4570 2350
rect 2910 2335 2950 2340
rect 2910 2305 2915 2335
rect 2945 2330 2950 2335
rect 3330 2335 3370 2340
rect 3330 2330 3335 2335
rect 2945 2310 3335 2330
rect 2945 2305 2950 2310
rect 2910 2300 2950 2305
rect 3330 2305 3335 2310
rect 3365 2330 3370 2335
rect 4110 2335 4150 2340
rect 4110 2330 4115 2335
rect 3365 2310 4115 2330
rect 3365 2305 3370 2310
rect 3330 2300 3370 2305
rect 4110 2305 4115 2310
rect 4145 2305 4150 2335
rect 4110 2300 4150 2305
rect 2800 2290 2840 2295
rect 2800 2260 2805 2290
rect 2835 2285 2840 2290
rect 3120 2290 3160 2295
rect 3120 2285 3125 2290
rect 2835 2265 3125 2285
rect 2835 2260 2840 2265
rect 2800 2255 2840 2260
rect 3120 2260 3125 2265
rect 3155 2285 3160 2290
rect 3720 2290 3760 2295
rect 3720 2285 3725 2290
rect 3155 2265 3725 2285
rect 3155 2260 3160 2265
rect 3120 2255 3160 2260
rect 3720 2260 3725 2265
rect 3755 2285 3760 2290
rect 4320 2290 4360 2295
rect 4320 2285 4325 2290
rect 3755 2265 4325 2285
rect 3755 2260 3760 2265
rect 3720 2255 3760 2260
rect 4320 2260 4325 2265
rect 4355 2260 4360 2290
rect 4320 2255 4360 2260
rect 3020 2230 3060 2235
rect 3020 2200 3025 2230
rect 3055 2225 3060 2230
rect 3220 2230 3260 2235
rect 3220 2225 3225 2230
rect 3055 2205 3225 2225
rect 3055 2200 3060 2205
rect 3020 2195 3060 2200
rect 3220 2200 3225 2205
rect 3255 2225 3260 2230
rect 3420 2230 3460 2235
rect 3420 2225 3425 2230
rect 3255 2205 3425 2225
rect 3255 2200 3260 2205
rect 3220 2195 3260 2200
rect 3420 2200 3425 2205
rect 3455 2225 3460 2230
rect 3620 2230 3660 2235
rect 3620 2225 3625 2230
rect 3455 2205 3625 2225
rect 3455 2200 3460 2205
rect 3420 2195 3460 2200
rect 3620 2200 3625 2205
rect 3655 2225 3660 2230
rect 3820 2230 3860 2235
rect 3820 2225 3825 2230
rect 3655 2205 3825 2225
rect 3655 2200 3660 2205
rect 3620 2195 3660 2200
rect 3820 2200 3825 2205
rect 3855 2225 3860 2230
rect 4020 2230 4060 2235
rect 4020 2225 4025 2230
rect 3855 2205 4025 2225
rect 3855 2200 3860 2205
rect 3820 2195 3860 2200
rect 4020 2200 4025 2205
rect 4055 2225 4060 2230
rect 4220 2230 4260 2235
rect 4220 2225 4225 2230
rect 4055 2205 4225 2225
rect 4055 2200 4060 2205
rect 4020 2195 4060 2200
rect 4220 2200 4225 2205
rect 4255 2225 4260 2230
rect 4420 2230 4460 2235
rect 4420 2225 4425 2230
rect 4255 2205 4425 2225
rect 4255 2200 4260 2205
rect 4220 2195 4260 2200
rect 4420 2200 4425 2205
rect 4455 2200 4460 2230
rect 4420 2195 4460 2200
rect 4740 2230 4780 2235
rect 4740 2200 4745 2230
rect 4775 2225 4780 2230
rect 4875 2230 4915 2235
rect 4875 2225 4880 2230
rect 4775 2205 4880 2225
rect 4775 2200 4780 2205
rect 4740 2195 4780 2200
rect 4875 2200 4880 2205
rect 4910 2200 4915 2230
rect 4875 2195 4915 2200
rect 1520 2025 1525 2060
rect 1560 2055 1565 2060
rect 1660 2055 1665 2060
rect 1560 2030 1665 2055
rect 1560 2025 1565 2030
rect 1660 2025 1665 2030
rect 1700 2025 1705 2060
rect 2479 2025 2484 2060
rect 2519 2055 2524 2060
rect 2910 2055 2950 2060
rect 2519 2030 2915 2055
rect 2519 2025 2524 2030
rect 2910 2025 2915 2030
rect 2945 2025 2950 2055
rect 2910 2020 2950 2025
rect 4530 1980 4570 1985
rect 3320 1955 3360 1960
rect 3320 1925 3325 1955
rect 3355 1950 3360 1955
rect 4120 1955 4160 1960
rect 4120 1950 4125 1955
rect 3355 1930 4125 1950
rect 3355 1925 3360 1930
rect 3320 1920 3360 1925
rect 4120 1925 4125 1930
rect 4155 1925 4160 1955
rect 4530 1950 4535 1980
rect 4565 1950 4570 1980
rect 4530 1945 4570 1950
rect 4120 1920 4160 1925
rect 3170 1910 3210 1915
rect 3170 1880 3175 1910
rect 3205 1905 3210 1910
rect 3520 1910 3560 1915
rect 3520 1905 3525 1910
rect 3205 1885 3525 1905
rect 3205 1880 3210 1885
rect 3170 1875 3210 1880
rect 3520 1880 3525 1885
rect 3555 1905 3560 1910
rect 3670 1910 3710 1915
rect 3670 1905 3675 1910
rect 3555 1885 3675 1905
rect 3555 1880 3560 1885
rect 3520 1875 3560 1880
rect 3670 1880 3675 1885
rect 3705 1905 3710 1910
rect 3770 1910 3810 1915
rect 3770 1905 3775 1910
rect 3705 1885 3775 1905
rect 3705 1880 3710 1885
rect 3670 1875 3710 1880
rect 3770 1880 3775 1885
rect 3805 1905 3810 1910
rect 3920 1910 3960 1915
rect 3920 1905 3925 1910
rect 3805 1885 3925 1905
rect 3805 1880 3810 1885
rect 3770 1875 3810 1880
rect 3920 1880 3925 1885
rect 3955 1905 3960 1910
rect 4270 1910 4310 1915
rect 4270 1905 4275 1910
rect 3955 1885 4275 1905
rect 3955 1880 3960 1885
rect 3920 1875 3960 1880
rect 4270 1880 4275 1885
rect 4305 1880 4310 1910
rect 4270 1875 4310 1880
rect 3120 1855 3160 1860
rect 3120 1825 3125 1855
rect 3155 1850 3160 1855
rect 3720 1855 3760 1860
rect 3720 1850 3725 1855
rect 3155 1830 3725 1850
rect 3155 1825 3160 1830
rect 3120 1820 3160 1825
rect 3720 1825 3725 1830
rect 3755 1850 3760 1855
rect 4320 1855 4360 1860
rect 4320 1850 4325 1855
rect 3755 1830 4325 1850
rect 3755 1825 3760 1830
rect 3720 1820 3760 1825
rect 4320 1825 4325 1830
rect 4355 1850 4360 1855
rect 4530 1855 4570 1860
rect 4530 1850 4535 1855
rect 4355 1830 4535 1850
rect 4355 1825 4360 1830
rect 4320 1820 4360 1825
rect 4530 1825 4535 1830
rect 4565 1825 4570 1855
rect 4530 1820 4570 1825
rect 3320 1795 3360 1800
rect 3320 1765 3325 1795
rect 3355 1790 3360 1795
rect 3720 1795 3760 1800
rect 3720 1790 3725 1795
rect 3355 1770 3725 1790
rect 3355 1765 3360 1770
rect 3320 1760 3360 1765
rect 3720 1765 3725 1770
rect 3755 1790 3760 1795
rect 4120 1795 4160 1800
rect 4120 1790 4125 1795
rect 3755 1770 4125 1790
rect 3755 1765 3760 1770
rect 3720 1760 3760 1765
rect 4120 1765 4125 1770
rect 4155 1765 4160 1795
rect 4120 1760 4160 1765
rect 3520 1750 3560 1755
rect -110 1720 -70 1725
rect -110 1690 -105 1720
rect -75 1690 -70 1720
rect -110 1685 -70 1690
rect -45 1720 -5 1725
rect -45 1690 -40 1720
rect -10 1690 -5 1720
rect 3520 1720 3525 1750
rect 3555 1745 3560 1750
rect 3920 1750 3960 1755
rect 3920 1745 3925 1750
rect 3555 1725 3925 1745
rect 3555 1720 3560 1725
rect 3520 1715 3560 1720
rect 3920 1720 3925 1725
rect 3955 1720 3960 1750
rect 3920 1715 3960 1720
rect -45 1685 -5 1690
rect 2855 1705 2895 1710
rect 2855 1675 2860 1705
rect 2890 1700 2895 1705
rect 3370 1705 3410 1710
rect 3370 1700 3375 1705
rect 2890 1680 3375 1700
rect 2890 1675 2895 1680
rect 2855 1670 2895 1675
rect 3370 1675 3375 1680
rect 3405 1700 3410 1705
rect 3670 1705 3710 1710
rect 3670 1700 3675 1705
rect 3405 1680 3675 1700
rect 3405 1675 3410 1680
rect 3370 1670 3410 1675
rect 3670 1675 3675 1680
rect 3705 1700 3710 1705
rect 3770 1705 3810 1710
rect 3770 1700 3775 1705
rect 3705 1680 3775 1700
rect 3705 1675 3710 1680
rect 3670 1670 3710 1675
rect 3770 1675 3775 1680
rect 3805 1700 3810 1705
rect 4070 1705 4110 1710
rect 4070 1700 4075 1705
rect 3805 1680 4075 1700
rect 3805 1675 3810 1680
rect 3770 1670 3810 1675
rect 4070 1675 4075 1680
rect 4105 1700 4110 1705
rect 4585 1705 4625 1710
rect 4585 1700 4590 1705
rect 4105 1680 4590 1700
rect 4105 1675 4110 1680
rect 4070 1670 4110 1675
rect 4585 1675 4590 1680
rect 4620 1675 4625 1705
rect 4585 1670 4625 1675
rect 1550 1635 1590 1640
rect 1660 1635 1665 1640
rect 1550 1605 1555 1635
rect 1585 1610 1665 1635
rect 1585 1605 1590 1610
rect 1660 1605 1665 1610
rect 1700 1605 1705 1640
rect 3105 1625 3145 1630
rect 1550 1600 1590 1605
rect 3105 1595 3110 1625
rect 3140 1620 3145 1625
rect 3185 1625 3225 1630
rect 3185 1620 3190 1625
rect 3140 1600 3190 1620
rect 3140 1595 3145 1600
rect 3105 1590 3145 1595
rect 3185 1595 3190 1600
rect 3220 1595 3225 1625
rect 3185 1590 3225 1595
rect 1605 1575 1645 1580
rect 1660 1575 1665 1580
rect 1605 1545 1610 1575
rect 1640 1550 1665 1575
rect 1640 1545 1645 1550
rect 1660 1545 1665 1550
rect 1700 1545 1705 1580
rect 4170 1545 4210 1550
rect 1605 1540 1645 1545
rect 2910 1540 2950 1545
rect 1660 1520 1705 1525
rect 1660 1485 1665 1520
rect 1700 1485 1705 1520
rect 2910 1510 2915 1540
rect 2945 1535 2950 1540
rect 3520 1540 3560 1545
rect 3520 1535 3525 1540
rect 2945 1515 3525 1535
rect 2945 1510 2950 1515
rect 2910 1505 2950 1510
rect 3520 1510 3525 1515
rect 3555 1535 3560 1540
rect 3920 1540 3960 1545
rect 3920 1535 3925 1540
rect 3555 1515 3925 1535
rect 3555 1510 3560 1515
rect 3520 1505 3560 1510
rect 3920 1510 3925 1515
rect 3955 1510 3960 1540
rect 4170 1515 4175 1545
rect 4205 1540 4210 1545
rect 4790 1545 4830 1550
rect 4790 1540 4795 1545
rect 4205 1520 4795 1540
rect 4205 1515 4210 1520
rect 4170 1510 4210 1515
rect 4790 1515 4795 1520
rect 4825 1515 4830 1545
rect 4790 1510 4830 1515
rect 3920 1505 3960 1510
rect 3420 1495 3460 1500
rect 1660 1480 1705 1485
rect 2800 1485 2840 1490
rect 2800 1480 2805 1485
rect 1660 1460 2805 1480
rect 2800 1455 2805 1460
rect 2835 1455 2840 1485
rect 3420 1465 3425 1495
rect 3455 1490 3460 1495
rect 3620 1495 3660 1500
rect 3620 1490 3625 1495
rect 3455 1470 3625 1490
rect 3455 1465 3460 1470
rect 3420 1460 3460 1465
rect 3620 1465 3625 1470
rect 3655 1490 3660 1495
rect 3820 1495 3860 1500
rect 3820 1490 3825 1495
rect 3655 1470 3825 1490
rect 3655 1465 3660 1470
rect 3620 1460 3660 1465
rect 3820 1465 3825 1470
rect 3855 1490 3860 1495
rect 4020 1495 4060 1500
rect 4020 1490 4025 1495
rect 3855 1470 4025 1490
rect 3855 1465 3860 1470
rect 3820 1460 3860 1465
rect 4020 1465 4025 1470
rect 4055 1465 4060 1495
rect 4020 1460 4060 1465
rect 2800 1450 2840 1455
rect 1605 1440 1645 1445
rect 1605 1410 1610 1440
rect 1640 1435 1645 1440
rect 2855 1440 2895 1445
rect 2855 1435 2860 1440
rect 1640 1415 2860 1435
rect 1640 1410 1645 1415
rect 1605 1405 1645 1410
rect 2855 1410 2860 1415
rect 2890 1410 2895 1440
rect 2855 1405 2895 1410
rect 4200 1435 4240 1440
rect 4200 1405 4205 1435
rect 4235 1430 4240 1435
rect 4320 1435 4360 1440
rect 4320 1430 4325 1435
rect 4235 1410 4325 1430
rect 4235 1405 4240 1410
rect 4200 1400 4240 1405
rect 4320 1405 4325 1410
rect 4355 1405 4360 1435
rect 4320 1400 4360 1405
rect 1550 1395 1590 1400
rect 1550 1365 1555 1395
rect 1585 1390 1590 1395
rect 2910 1395 2950 1400
rect 2910 1390 2915 1395
rect 1585 1370 2915 1390
rect 1585 1365 1590 1370
rect 1550 1360 1590 1365
rect 2910 1365 2915 1370
rect 2945 1365 2950 1395
rect 2910 1360 2950 1365
rect 2225 1030 2265 1035
rect 2225 1000 2230 1030
rect 2260 1025 2265 1030
rect 2855 1030 2895 1035
rect 2855 1025 2860 1030
rect 2260 1005 2860 1025
rect 2260 1000 2265 1005
rect 2225 995 2265 1000
rect 2855 1000 2860 1005
rect 2890 1000 2895 1030
rect 2855 995 2895 1000
rect 3680 965 3800 970
rect 3680 935 3685 965
rect 3715 935 3725 965
rect 3755 935 3765 965
rect 3795 960 3800 965
rect 4790 965 4830 970
rect 4790 960 4795 965
rect 3795 940 4795 960
rect 3795 935 3800 940
rect 3680 930 3800 935
rect 4790 935 4795 940
rect 4825 935 4830 965
rect 4790 930 4830 935
rect 4230 905 4270 910
rect 4230 875 4235 905
rect 4265 900 4270 905
rect 4650 905 4690 910
rect 4650 900 4655 905
rect 4265 880 4655 900
rect 4265 875 4270 880
rect 4230 870 4270 875
rect 4650 875 4655 880
rect 4685 875 4690 905
rect 4650 870 4690 875
rect 4305 820 4345 825
rect 4305 790 4310 820
rect 4340 815 4345 820
rect 4790 820 4830 825
rect 4790 815 4795 820
rect 4340 795 4795 815
rect 4340 790 4345 795
rect 4305 785 4345 790
rect 4790 790 4795 795
rect 4825 790 4830 820
rect 4790 785 4830 790
rect 3100 630 3150 640
rect 3100 600 3110 630
rect 3140 600 3150 630
rect 3100 590 3150 600
rect -195 550 -155 555
rect -195 520 -190 550
rect -160 520 -155 550
rect -195 515 -155 520
<< via2 >>
rect -190 2955 -160 2985
rect 4880 2955 4910 2985
rect 1565 2870 1595 2900
rect 1615 2870 1645 2900
rect 1665 2870 1695 2900
rect -190 2820 -160 2850
rect 4880 2820 4910 2850
rect 4880 2200 4910 2230
rect -105 1690 -75 1720
rect 4795 1515 4825 1545
rect 4795 935 4825 965
rect 4795 790 4825 820
rect 3110 600 3140 630
rect -190 520 -160 550
<< metal3 >>
rect -200 2990 -150 2995
rect -200 2950 -195 2990
rect -155 2950 -150 2990
rect -200 2945 -150 2950
rect 4870 2990 4920 2995
rect 4870 2950 4875 2990
rect 4915 2950 4920 2990
rect 4870 2945 4920 2950
rect -195 2850 -155 2945
rect -115 2905 -65 2910
rect -115 2865 -110 2905
rect -70 2865 -65 2905
rect -115 2860 -65 2865
rect 1555 2905 1705 2910
rect 1555 2865 1560 2905
rect 1600 2865 1610 2905
rect 1650 2865 1660 2905
rect 1700 2865 1705 2905
rect 1555 2860 1705 2865
rect 4785 2905 4835 2910
rect 4785 2865 4790 2905
rect 4830 2865 4835 2905
rect 4785 2860 4835 2865
rect -195 2820 -190 2850
rect -160 2820 -155 2850
rect -195 560 -155 2820
rect -110 1720 -70 2860
rect -110 1690 -105 1720
rect -75 1690 -70 1720
rect -110 640 -70 1690
rect 4790 1545 4830 2860
rect 4790 1515 4795 1545
rect 4825 1515 4830 1545
rect 4790 965 4830 1515
rect 4790 935 4795 965
rect 4825 935 4830 965
rect 4790 820 4830 935
rect 4790 790 4795 820
rect 4825 790 4830 820
rect 4790 640 4830 790
rect 4875 2850 4915 2945
rect 4875 2820 4880 2850
rect 4910 2820 4915 2850
rect 4875 2230 4915 2820
rect 4875 2200 4880 2230
rect 4910 2200 4915 2230
rect -115 635 -65 640
rect -115 595 -110 635
rect -70 595 -65 635
rect -115 590 -65 595
rect 3100 635 3150 640
rect 3100 595 3105 635
rect 3145 595 3150 635
rect 3100 590 3150 595
rect 4785 635 4835 640
rect 4785 595 4790 635
rect 4830 595 4835 635
rect 4785 590 4835 595
rect 4875 560 4915 2200
rect -200 555 -150 560
rect -200 515 -195 555
rect -155 515 -150 555
rect -200 510 -150 515
rect 4870 555 4920 560
rect 4870 515 4875 555
rect 4915 515 4920 555
rect 4870 510 4920 515
<< via3 >>
rect -195 2985 -155 2990
rect -195 2955 -190 2985
rect -190 2955 -160 2985
rect -160 2955 -155 2985
rect -195 2950 -155 2955
rect 4875 2985 4915 2990
rect 4875 2955 4880 2985
rect 4880 2955 4910 2985
rect 4910 2955 4915 2985
rect 4875 2950 4915 2955
rect -110 2865 -70 2905
rect 1560 2900 1600 2905
rect 1560 2870 1565 2900
rect 1565 2870 1595 2900
rect 1595 2870 1600 2900
rect 1560 2865 1600 2870
rect 1610 2900 1650 2905
rect 1610 2870 1615 2900
rect 1615 2870 1645 2900
rect 1645 2870 1650 2900
rect 1610 2865 1650 2870
rect 1660 2900 1700 2905
rect 1660 2870 1665 2900
rect 1665 2870 1695 2900
rect 1695 2870 1700 2900
rect 1660 2865 1700 2870
rect 4790 2865 4830 2905
rect -110 595 -70 635
rect 3105 630 3145 635
rect 3105 600 3110 630
rect 3110 600 3140 630
rect 3140 600 3145 630
rect 3105 595 3145 600
rect 4790 595 4830 635
rect -195 550 -155 555
rect -195 520 -190 550
rect -190 520 -160 550
rect -160 520 -155 550
rect -195 515 -155 520
rect 4875 515 4915 555
<< metal4 >>
rect -200 2990 4920 2995
rect -200 2950 -195 2990
rect -155 2950 4875 2990
rect 4915 2950 4920 2990
rect -200 2945 4920 2950
rect -115 2905 4835 2910
rect -115 2865 -110 2905
rect -70 2865 1560 2905
rect 1600 2865 1610 2905
rect 1650 2865 1660 2905
rect 1700 2865 4790 2905
rect 4830 2865 4835 2905
rect -115 2860 4835 2865
rect -115 635 4835 640
rect -115 595 -110 635
rect -70 595 3105 635
rect 3145 595 4790 635
rect 4830 595 4835 635
rect -115 590 4835 595
rect -200 555 4920 560
rect -200 515 -195 555
rect -155 515 4875 555
rect 4915 515 4920 555
rect -200 510 4920 515
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0 $PDKPATH/libs.ref/sky130_fd_pr/mag
timestamp 1723858470
transform 1 0 795 0 1 1360
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_1
timestamp 1723858470
transform 1 0 795 0 1 2040
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_2
timestamp 1723858470
transform 1 0 795 0 1 680
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_3
timestamp 1723858470
transform 1 0 115 0 1 2040
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_4
timestamp 1723858470
transform 1 0 115 0 1 1360
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5
timestamp 1723858470
transform 1 0 115 0 1 680
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_6
timestamp 1723858470
transform 1 0 1525 0 1 680
box 0 0 670 670
<< labels >>
flabel metal3 4830 1175 4830 1175 3 FreeSans 800 0 80 0 GNDA
port 6 e
flabel metal1 4680 1615 4680 1615 3 FreeSans 400 0 80 0 start_up
flabel metal1 4570 2365 4570 2365 3 FreeSans 400 0 80 0 V_TOP
flabel locali 3430 1450 3430 1450 7 FreeSans 400 0 -80 0 V_p
flabel metal2 2980 1680 2980 1680 5 FreeSans 400 0 0 -80 Vin-
flabel metal2 2980 1515 2980 1515 5 FreeSans 400 0 0 -80 Vin+
flabel metal3 4915 1400 4915 1400 3 FreeSans 800 0 80 0 VDDA
port 1 e
flabel metal2 3320 1780 3320 1780 7 FreeSans 400 0 -80 0 V_mirror
flabel metal1 3950 1810 3950 1810 3 FreeSans 400 0 80 0 1st_Vout
flabel metal1 3740 3175 3740 3175 1 FreeSans 800 0 0 400 V_OUT
port 2 n
<< end >>
