magic
tech sky130A
timestamp 1750847378
<< metal1 >>
rect 425 5135 465 5140
rect 425 5105 430 5135
rect 460 5105 465 5135
rect 425 5100 465 5105
rect 4145 5135 4185 5140
rect 4145 5105 4150 5135
rect 4180 5105 4185 5135
rect 4145 5100 4185 5105
rect 370 5090 410 5095
rect 370 5060 375 5090
rect 405 5060 410 5090
rect 370 5055 410 5060
rect 265 4515 305 4520
rect 265 4485 270 4515
rect 300 4485 305 4515
rect 265 4480 305 4485
rect 115 4390 155 4395
rect 115 4360 120 4390
rect 150 4360 155 4390
rect 115 4355 155 4360
rect -2990 1985 -2950 1990
rect -2990 1955 -2985 1985
rect -2955 1955 -2950 1985
rect -2990 1950 -2950 1955
rect -1555 1940 -1515 1945
rect -1555 1910 -1550 1940
rect -1520 1910 -1515 1940
rect -1555 1905 -1515 1910
rect -1735 1895 -1695 1900
rect -1735 1865 -1730 1895
rect -1700 1865 -1695 1895
rect -1735 1860 -1695 1865
rect 125 1855 145 4355
rect 275 4350 295 4480
rect 325 4435 365 4440
rect 325 4405 330 4435
rect 360 4405 365 4435
rect 325 4400 365 4405
rect 265 4345 305 4350
rect 265 4315 270 4345
rect 300 4315 305 4345
rect 265 4310 305 4315
rect 265 4195 305 4200
rect 265 4165 270 4195
rect 300 4165 305 4195
rect 265 4160 305 4165
rect -1915 1850 -1875 1855
rect -1915 1820 -1910 1850
rect -1880 1820 -1875 1850
rect -1915 1815 -1875 1820
rect 115 1850 155 1855
rect 115 1820 120 1850
rect 150 1820 155 1850
rect 115 1815 155 1820
rect -470 865 -450 1750
rect 275 1290 295 4160
rect 335 3450 355 4400
rect 325 3445 365 3450
rect 325 3415 330 3445
rect 360 3415 365 3445
rect 325 3410 365 3415
rect 380 1900 400 5055
rect 435 1945 455 5100
rect 2935 5035 2975 5040
rect 2935 5005 2940 5035
rect 2970 5005 2975 5035
rect 2935 5000 2975 5005
rect 2945 3045 2965 5000
rect 7120 4760 7160 4765
rect 7120 4730 7125 4760
rect 7155 4730 7160 4760
rect 7120 4725 7160 4730
rect 4075 4455 4115 4460
rect 4075 4425 4080 4455
rect 4110 4425 4115 4455
rect 4075 4420 4115 4425
rect 4075 4345 4115 4350
rect 4075 4315 4080 4345
rect 4110 4315 4115 4345
rect 4075 4310 4115 4315
rect 2990 2430 3010 2445
rect 2735 2425 2775 2430
rect 2735 2395 2740 2425
rect 2770 2395 2775 2425
rect 2735 2390 2775 2395
rect 2980 2425 3020 2430
rect 2980 2395 2985 2425
rect 3015 2395 3020 2425
rect 4085 2410 4105 4310
rect 7130 3045 7150 4725
rect 7085 2430 7105 2445
rect 7075 2425 7115 2430
rect 2980 2390 3020 2395
rect 4075 2405 4115 2410
rect 2460 2225 2500 2265
rect 2745 1990 2765 2390
rect 4075 2375 4080 2405
rect 4110 2375 4115 2405
rect 7075 2395 7080 2425
rect 7110 2395 7115 2425
rect 7075 2390 7115 2395
rect 7315 2425 7355 2430
rect 7315 2395 7320 2425
rect 7350 2395 7355 2425
rect 7315 2390 7355 2395
rect 4075 2370 4115 2375
rect 2735 1985 2775 1990
rect 2735 1955 2740 1985
rect 2770 1955 2775 1985
rect 2735 1950 2775 1955
rect 425 1940 465 1945
rect 425 1910 430 1940
rect 460 1910 465 1940
rect 425 1905 465 1910
rect 370 1895 410 1900
rect 370 1865 375 1895
rect 405 1865 410 1895
rect 370 1860 410 1865
rect 265 1285 305 1290
rect 265 1255 270 1285
rect 300 1255 305 1285
rect 265 1250 305 1255
rect 7325 865 7345 2390
rect 7590 2225 7630 2265
rect -480 860 -440 865
rect -480 830 -475 860
rect -445 830 -440 860
rect -480 825 -440 830
rect 7315 860 7355 865
rect 7315 830 7320 860
rect 7350 830 7355 860
rect 7315 825 7355 830
<< via1 >>
rect 430 5105 460 5135
rect 4150 5105 4180 5135
rect 375 5060 405 5090
rect 270 4485 300 4515
rect 120 4360 150 4390
rect -2985 1955 -2955 1985
rect -1550 1910 -1520 1940
rect -1730 1865 -1700 1895
rect 330 4405 360 4435
rect 270 4315 300 4345
rect 270 4165 300 4195
rect -1910 1820 -1880 1850
rect 120 1820 150 1850
rect 330 3415 360 3445
rect 2940 5005 2970 5035
rect 7125 4730 7155 4760
rect 4080 4425 4110 4455
rect 4080 4315 4110 4345
rect 2740 2395 2770 2425
rect 2985 2395 3015 2425
rect 4080 2375 4110 2405
rect 7080 2395 7110 2425
rect 7320 2395 7350 2425
rect 2740 1955 2770 1985
rect 430 1910 460 1940
rect 375 1865 405 1895
rect 270 1255 300 1285
rect -475 830 -445 860
rect 7320 830 7350 860
<< metal2 >>
rect 425 5135 465 5140
rect 425 5105 430 5135
rect 460 5130 465 5135
rect 4145 5135 4185 5140
rect 4145 5130 4150 5135
rect 460 5110 4150 5130
rect 460 5105 465 5110
rect 425 5100 465 5105
rect 4145 5105 4150 5110
rect 4180 5105 4185 5135
rect 4145 5100 4185 5105
rect 370 5090 410 5095
rect 370 5060 375 5090
rect 405 5085 410 5090
rect 405 5065 4200 5085
rect 405 5060 410 5065
rect 370 5055 410 5060
rect 2935 5035 2975 5040
rect 2935 5030 2940 5035
rect 305 5010 2940 5030
rect 2935 5005 2940 5010
rect 2970 5005 2975 5035
rect 2935 5000 2975 5005
rect 7120 4760 7160 4765
rect 7120 4755 7125 4760
rect 305 4735 7125 4755
rect 7120 4730 7125 4735
rect 7155 4730 7160 4760
rect 7120 4725 7160 4730
rect 265 4515 305 4520
rect 265 4485 270 4515
rect 300 4485 305 4515
rect 265 4480 305 4485
rect 4075 4455 4115 4460
rect 325 4435 365 4440
rect 325 4405 330 4435
rect 360 4430 365 4435
rect 4075 4430 4080 4455
rect 360 4425 4080 4430
rect 4110 4425 4115 4455
rect 360 4410 4115 4425
rect 360 4405 365 4410
rect 325 4400 365 4405
rect 115 4390 155 4395
rect 115 4360 120 4390
rect 150 4385 155 4390
rect 150 4365 4440 4385
rect 150 4360 155 4365
rect 115 4355 155 4360
rect 265 4345 305 4350
rect 265 4315 270 4345
rect 300 4340 305 4345
rect 4075 4345 4115 4350
rect 4075 4340 4080 4345
rect 300 4320 4080 4340
rect 300 4315 305 4320
rect 265 4310 305 4315
rect 4075 4315 4080 4320
rect 4110 4315 4115 4345
rect 4075 4310 4115 4315
rect 265 4195 305 4200
rect 265 4165 270 4195
rect 300 4165 305 4195
rect 265 4160 305 4165
rect 325 3445 365 3450
rect 325 3440 330 3445
rect 305 3420 330 3440
rect 325 3415 330 3420
rect 360 3415 365 3445
rect 325 3410 365 3415
rect 2735 2425 2775 2430
rect 2735 2395 2740 2425
rect 2770 2420 2775 2425
rect 2980 2425 3020 2430
rect 2980 2420 2985 2425
rect 2770 2400 2985 2420
rect 2770 2395 2775 2400
rect 2735 2390 2775 2395
rect 2980 2395 2985 2400
rect 3015 2395 3020 2425
rect 7075 2425 7115 2430
rect 2980 2390 3020 2395
rect 4075 2405 4115 2410
rect 4075 2375 4080 2405
rect 4110 2400 4115 2405
rect 4110 2380 4965 2400
rect 7075 2395 7080 2425
rect 7110 2420 7115 2425
rect 7315 2425 7355 2430
rect 7315 2420 7320 2425
rect 7110 2400 7320 2420
rect 7110 2395 7115 2400
rect 7075 2390 7115 2395
rect 7315 2395 7320 2400
rect 7350 2395 7355 2425
rect 7315 2390 7355 2395
rect 4110 2375 4115 2380
rect 4075 2370 4115 2375
rect 4065 2290 4080 2310
rect 2460 2225 2500 2265
rect 7590 2225 7630 2265
rect 4065 2070 4080 2090
rect -2990 1985 -2950 1990
rect -2990 1955 -2985 1985
rect -2955 1980 -2950 1985
rect 2735 1985 2775 1990
rect 2735 1980 2740 1985
rect -2955 1960 2740 1980
rect -2955 1955 -2950 1960
rect -2990 1950 -2950 1955
rect 2735 1955 2740 1960
rect 2770 1955 2775 1985
rect 2735 1950 2775 1955
rect -1555 1940 -1515 1945
rect -1555 1910 -1550 1940
rect -1520 1935 -1515 1940
rect 425 1940 465 1945
rect 425 1935 430 1940
rect -1520 1915 430 1935
rect -1520 1910 -1515 1915
rect -1555 1905 -1515 1910
rect 425 1910 430 1915
rect 460 1910 465 1940
rect 425 1905 465 1910
rect -1735 1895 -1695 1900
rect -1735 1865 -1730 1895
rect -1700 1890 -1695 1895
rect 370 1895 410 1900
rect 370 1890 375 1895
rect -1700 1870 375 1890
rect -1700 1865 -1695 1870
rect -1735 1860 -1695 1865
rect 370 1865 375 1870
rect 405 1865 410 1895
rect 370 1860 410 1865
rect -1915 1850 -1875 1855
rect -1915 1820 -1910 1850
rect -1880 1845 -1875 1850
rect 115 1850 155 1855
rect 115 1845 120 1850
rect -1880 1825 120 1845
rect -1880 1820 -1875 1825
rect -1915 1815 -1875 1820
rect 115 1820 120 1825
rect 150 1820 155 1850
rect 115 1815 155 1820
rect 265 1285 305 1290
rect 265 1255 270 1285
rect 300 1280 305 1285
rect 300 1260 3975 1280
rect 300 1255 305 1260
rect 265 1250 305 1255
rect -480 860 -440 865
rect -480 830 -475 860
rect -445 855 -440 860
rect 7315 860 7355 865
rect 7315 855 7320 860
rect -445 835 7320 855
rect -445 830 -440 835
rect -480 825 -440 830
rect 7315 830 7320 835
rect 7350 830 7355 860
rect 7315 825 7355 830
<< metal3 >>
rect -130 50 -90 2015
rect -130 45 -80 50
rect -130 5 -125 45
rect -85 5 -80 45
rect -130 0 -80 5
<< via3 >>
rect -125 5 -85 45
<< metal4 >>
rect 940 6700 990 6750
rect -130 45 0 50
rect -130 5 -125 45
rect -85 5 0 45
rect -130 0 0 5
rect 975 0 1025 50
use bgr  bgr_0
timestamp 1750847327
transform 1 0 -5795 0 1 1400
box -200 350 6100 5350
use two_stage_opamp_dummy_magic  two_stage_opamp_dummy_magic_0
timestamp 1750645408
transform 1 0 -26855 0 1 555
box 26855 -555 36545 6195
<< labels >>
flabel metal4 965 6750 965 6750 1 FreeSans 800 0 0 400 VDDA
port 1 n
flabel metal4 1000 0 1000 0 5 FreeSans 800 0 0 -400 GNDA
port 2 s
flabel metal2 7610 2225 7610 2225 5 FreeSans 400 0 0 -200 VOUT+
port 3 s
flabel metal2 2480 2225 2480 2225 5 FreeSans 400 0 0 -200 VOUT-
port 4 s
flabel metal2 4065 2080 4065 2080 7 FreeSans 400 0 -200 0 VIN+
port 5 w
flabel metal2 4065 2300 4065 2300 7 FreeSans 400 0 -200 0 VIN-
port 6 w
<< end >>
