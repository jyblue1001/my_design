magic
tech sky130A
timestamp 1748808989
<< pwell >>
rect 2945 2890 3165 2990
rect 3195 2890 5035 2990
rect 2760 2450 5140 2750
rect 2515 1900 2665 2000
rect 2695 1900 3935 2000
rect 3965 1900 5205 2000
rect -45 1685 130 1725
rect 3115 1615 3755 1665
rect 4145 1615 4785 1665
rect 2785 1210 3905 1460
rect 3995 1210 5115 1460
rect 2890 1015 5010 1115
rect 3040 810 3170 910
rect 3200 810 4950 910
<< nmos >>
rect 2985 2890 3035 2990
rect 3075 2890 3125 2990
rect 3235 2890 3285 2990
rect 3325 2890 3375 2990
rect 3415 2890 3465 2990
rect 3505 2890 3555 2990
rect 3595 2890 3645 2990
rect 3685 2890 3735 2990
rect 3775 2890 3825 2990
rect 3865 2890 3915 2990
rect 3955 2890 4005 2990
rect 4045 2890 4095 2990
rect 4135 2890 4185 2990
rect 4225 2890 4275 2990
rect 4315 2890 4365 2990
rect 4405 2890 4455 2990
rect 4495 2890 4545 2990
rect 4585 2890 4635 2990
rect 4675 2890 4725 2990
rect 4765 2890 4815 2990
rect 4855 2890 4905 2990
rect 4945 2890 4995 2990
rect 2800 2450 2850 2750
rect 2890 2450 2940 2750
rect 2980 2450 3030 2750
rect 3070 2450 3120 2750
rect 3160 2450 3210 2750
rect 3250 2450 3300 2750
rect 3340 2450 3390 2750
rect 3430 2450 3480 2750
rect 3520 2450 3570 2750
rect 3610 2450 3660 2750
rect 3700 2450 3750 2750
rect 3790 2450 3840 2750
rect 3880 2450 3930 2750
rect 3970 2450 4020 2750
rect 4060 2450 4110 2750
rect 4150 2450 4200 2750
rect 4240 2450 4290 2750
rect 4330 2450 4380 2750
rect 4420 2450 4470 2750
rect 4510 2450 4560 2750
rect 4600 2450 4650 2750
rect 4690 2450 4740 2750
rect 4780 2450 4830 2750
rect 4870 2450 4920 2750
rect 4960 2450 5010 2750
rect 5050 2450 5100 2750
rect 2555 1900 2570 2000
rect 2610 1900 2625 2000
rect 2735 1900 2755 2000
rect 2795 1900 2815 2000
rect 2855 1900 2875 2000
rect 2915 1900 2935 2000
rect 2975 1900 2995 2000
rect 3035 1900 3055 2000
rect 3095 1900 3115 2000
rect 3155 1900 3175 2000
rect 3215 1900 3235 2000
rect 3275 1900 3295 2000
rect 3335 1900 3355 2000
rect 3395 1900 3415 2000
rect 3455 1900 3475 2000
rect 3515 1900 3535 2000
rect 3575 1900 3595 2000
rect 3635 1900 3655 2000
rect 3695 1900 3715 2000
rect 3755 1900 3775 2000
rect 3815 1900 3835 2000
rect 3875 1900 3895 2000
rect 4005 1900 4025 2000
rect 4065 1900 4085 2000
rect 4125 1900 4145 2000
rect 4185 1900 4205 2000
rect 4245 1900 4265 2000
rect 4305 1900 4325 2000
rect 4365 1900 4385 2000
rect 4425 1900 4445 2000
rect 4485 1900 4505 2000
rect 4545 1900 4565 2000
rect 4605 1900 4625 2000
rect 4665 1900 4685 2000
rect 4725 1900 4745 2000
rect 4785 1900 4805 2000
rect 4845 1900 4865 2000
rect 4905 1900 4925 2000
rect 4965 1900 4985 2000
rect 5025 1900 5045 2000
rect 5085 1900 5105 2000
rect 5145 1900 5165 2000
rect 3155 1615 3175 1665
rect 3215 1615 3235 1665
rect 3275 1615 3295 1665
rect 3335 1615 3355 1665
rect 3395 1615 3415 1665
rect 3455 1615 3475 1665
rect 3515 1615 3535 1665
rect 3575 1615 3595 1665
rect 3635 1615 3655 1665
rect 3695 1615 3715 1665
rect 4185 1615 4205 1665
rect 4245 1615 4265 1665
rect 4305 1615 4325 1665
rect 4365 1615 4385 1665
rect 4425 1615 4445 1665
rect 4485 1615 4505 1665
rect 4545 1615 4565 1665
rect 4605 1615 4625 1665
rect 4665 1615 4685 1665
rect 4725 1615 4745 1665
rect 2825 1210 3325 1460
rect 3365 1210 3865 1460
rect 4035 1210 4535 1460
rect 4575 1210 5075 1460
rect 2930 1015 3930 1115
rect 3970 1015 4970 1115
rect 3080 810 3130 910
rect 3240 810 3290 910
rect 3330 810 3380 910
rect 3420 810 3470 910
rect 3510 810 3560 910
rect 3600 810 3650 910
rect 3690 810 3740 910
rect 3780 810 3830 910
rect 3870 810 3920 910
rect 3960 810 4010 910
rect 4050 810 4100 910
rect 4140 810 4190 910
rect 4230 810 4280 910
rect 4320 810 4370 910
rect 4410 810 4460 910
rect 4500 810 4550 910
rect 4590 810 4640 910
rect 4680 810 4730 910
rect 4770 810 4820 910
rect 4860 810 4910 910
<< ndiff >>
rect 2945 2975 2985 2990
rect 2945 2955 2955 2975
rect 2975 2955 2985 2975
rect 2945 2925 2985 2955
rect 2945 2905 2955 2925
rect 2975 2905 2985 2925
rect 2945 2890 2985 2905
rect 3035 2975 3075 2990
rect 3035 2955 3045 2975
rect 3065 2955 3075 2975
rect 3035 2925 3075 2955
rect 3035 2905 3045 2925
rect 3065 2905 3075 2925
rect 3035 2890 3075 2905
rect 3125 2975 3165 2990
rect 3125 2955 3135 2975
rect 3155 2955 3165 2975
rect 3125 2925 3165 2955
rect 3125 2905 3135 2925
rect 3155 2905 3165 2925
rect 3125 2890 3165 2905
rect 3195 2975 3235 2990
rect 3195 2955 3205 2975
rect 3225 2955 3235 2975
rect 3195 2925 3235 2955
rect 3195 2905 3205 2925
rect 3225 2905 3235 2925
rect 3195 2890 3235 2905
rect 3285 2975 3325 2990
rect 3285 2955 3295 2975
rect 3315 2955 3325 2975
rect 3285 2925 3325 2955
rect 3285 2905 3295 2925
rect 3315 2905 3325 2925
rect 3285 2890 3325 2905
rect 3375 2975 3415 2990
rect 3375 2955 3385 2975
rect 3405 2955 3415 2975
rect 3375 2925 3415 2955
rect 3375 2905 3385 2925
rect 3405 2905 3415 2925
rect 3375 2890 3415 2905
rect 3465 2975 3505 2990
rect 3465 2955 3475 2975
rect 3495 2955 3505 2975
rect 3465 2925 3505 2955
rect 3465 2905 3475 2925
rect 3495 2905 3505 2925
rect 3465 2890 3505 2905
rect 3555 2975 3595 2990
rect 3555 2955 3565 2975
rect 3585 2955 3595 2975
rect 3555 2925 3595 2955
rect 3555 2905 3565 2925
rect 3585 2905 3595 2925
rect 3555 2890 3595 2905
rect 3645 2975 3685 2990
rect 3645 2955 3655 2975
rect 3675 2955 3685 2975
rect 3645 2925 3685 2955
rect 3645 2905 3655 2925
rect 3675 2905 3685 2925
rect 3645 2890 3685 2905
rect 3735 2975 3775 2990
rect 3735 2955 3745 2975
rect 3765 2955 3775 2975
rect 3735 2925 3775 2955
rect 3735 2905 3745 2925
rect 3765 2905 3775 2925
rect 3735 2890 3775 2905
rect 3825 2975 3865 2990
rect 3825 2955 3835 2975
rect 3855 2955 3865 2975
rect 3825 2925 3865 2955
rect 3825 2905 3835 2925
rect 3855 2905 3865 2925
rect 3825 2890 3865 2905
rect 3915 2975 3955 2990
rect 3915 2955 3925 2975
rect 3945 2955 3955 2975
rect 3915 2925 3955 2955
rect 3915 2905 3925 2925
rect 3945 2905 3955 2925
rect 3915 2890 3955 2905
rect 4005 2975 4045 2990
rect 4005 2955 4015 2975
rect 4035 2955 4045 2975
rect 4005 2925 4045 2955
rect 4005 2905 4015 2925
rect 4035 2905 4045 2925
rect 4005 2890 4045 2905
rect 4095 2975 4135 2990
rect 4095 2955 4105 2975
rect 4125 2955 4135 2975
rect 4095 2925 4135 2955
rect 4095 2905 4105 2925
rect 4125 2905 4135 2925
rect 4095 2890 4135 2905
rect 4185 2975 4225 2990
rect 4185 2955 4195 2975
rect 4215 2955 4225 2975
rect 4185 2925 4225 2955
rect 4185 2905 4195 2925
rect 4215 2905 4225 2925
rect 4185 2890 4225 2905
rect 4275 2975 4315 2990
rect 4275 2955 4285 2975
rect 4305 2955 4315 2975
rect 4275 2925 4315 2955
rect 4275 2905 4285 2925
rect 4305 2905 4315 2925
rect 4275 2890 4315 2905
rect 4365 2975 4405 2990
rect 4365 2955 4375 2975
rect 4395 2955 4405 2975
rect 4365 2925 4405 2955
rect 4365 2905 4375 2925
rect 4395 2905 4405 2925
rect 4365 2890 4405 2905
rect 4455 2975 4495 2990
rect 4455 2955 4465 2975
rect 4485 2955 4495 2975
rect 4455 2925 4495 2955
rect 4455 2905 4465 2925
rect 4485 2905 4495 2925
rect 4455 2890 4495 2905
rect 4545 2975 4585 2990
rect 4545 2955 4555 2975
rect 4575 2955 4585 2975
rect 4545 2925 4585 2955
rect 4545 2905 4555 2925
rect 4575 2905 4585 2925
rect 4545 2890 4585 2905
rect 4635 2975 4675 2990
rect 4635 2955 4645 2975
rect 4665 2955 4675 2975
rect 4635 2925 4675 2955
rect 4635 2905 4645 2925
rect 4665 2905 4675 2925
rect 4635 2890 4675 2905
rect 4725 2975 4765 2990
rect 4725 2955 4735 2975
rect 4755 2955 4765 2975
rect 4725 2925 4765 2955
rect 4725 2905 4735 2925
rect 4755 2905 4765 2925
rect 4725 2890 4765 2905
rect 4815 2975 4855 2990
rect 4815 2955 4825 2975
rect 4845 2955 4855 2975
rect 4815 2925 4855 2955
rect 4815 2905 4825 2925
rect 4845 2905 4855 2925
rect 4815 2890 4855 2905
rect 4905 2975 4945 2990
rect 4905 2955 4915 2975
rect 4935 2955 4945 2975
rect 4905 2925 4945 2955
rect 4905 2905 4915 2925
rect 4935 2905 4945 2925
rect 4905 2890 4945 2905
rect 4995 2975 5035 2990
rect 4995 2955 5005 2975
rect 5025 2955 5035 2975
rect 4995 2925 5035 2955
rect 4995 2905 5005 2925
rect 5025 2905 5035 2925
rect 4995 2890 5035 2905
rect 2760 2735 2800 2750
rect 2760 2715 2770 2735
rect 2790 2715 2800 2735
rect 2760 2685 2800 2715
rect 2760 2665 2770 2685
rect 2790 2665 2800 2685
rect 2760 2635 2800 2665
rect 2760 2615 2770 2635
rect 2790 2615 2800 2635
rect 2760 2585 2800 2615
rect 2760 2565 2770 2585
rect 2790 2565 2800 2585
rect 2760 2535 2800 2565
rect 2760 2515 2770 2535
rect 2790 2515 2800 2535
rect 2760 2485 2800 2515
rect 2760 2465 2770 2485
rect 2790 2465 2800 2485
rect 2760 2450 2800 2465
rect 2850 2735 2890 2750
rect 2850 2715 2860 2735
rect 2880 2715 2890 2735
rect 2850 2685 2890 2715
rect 2850 2665 2860 2685
rect 2880 2665 2890 2685
rect 2850 2635 2890 2665
rect 2850 2615 2860 2635
rect 2880 2615 2890 2635
rect 2850 2585 2890 2615
rect 2850 2565 2860 2585
rect 2880 2565 2890 2585
rect 2850 2535 2890 2565
rect 2850 2515 2860 2535
rect 2880 2515 2890 2535
rect 2850 2485 2890 2515
rect 2850 2465 2860 2485
rect 2880 2465 2890 2485
rect 2850 2450 2890 2465
rect 2940 2735 2980 2750
rect 2940 2715 2950 2735
rect 2970 2715 2980 2735
rect 2940 2685 2980 2715
rect 2940 2665 2950 2685
rect 2970 2665 2980 2685
rect 2940 2635 2980 2665
rect 2940 2615 2950 2635
rect 2970 2615 2980 2635
rect 2940 2585 2980 2615
rect 2940 2565 2950 2585
rect 2970 2565 2980 2585
rect 2940 2535 2980 2565
rect 2940 2515 2950 2535
rect 2970 2515 2980 2535
rect 2940 2485 2980 2515
rect 2940 2465 2950 2485
rect 2970 2465 2980 2485
rect 2940 2450 2980 2465
rect 3030 2735 3070 2750
rect 3030 2715 3040 2735
rect 3060 2715 3070 2735
rect 3030 2685 3070 2715
rect 3030 2665 3040 2685
rect 3060 2665 3070 2685
rect 3030 2635 3070 2665
rect 3030 2615 3040 2635
rect 3060 2615 3070 2635
rect 3030 2585 3070 2615
rect 3030 2565 3040 2585
rect 3060 2565 3070 2585
rect 3030 2535 3070 2565
rect 3030 2515 3040 2535
rect 3060 2515 3070 2535
rect 3030 2485 3070 2515
rect 3030 2465 3040 2485
rect 3060 2465 3070 2485
rect 3030 2450 3070 2465
rect 3120 2735 3160 2750
rect 3120 2715 3130 2735
rect 3150 2715 3160 2735
rect 3120 2685 3160 2715
rect 3120 2665 3130 2685
rect 3150 2665 3160 2685
rect 3120 2635 3160 2665
rect 3120 2615 3130 2635
rect 3150 2615 3160 2635
rect 3120 2585 3160 2615
rect 3120 2565 3130 2585
rect 3150 2565 3160 2585
rect 3120 2535 3160 2565
rect 3120 2515 3130 2535
rect 3150 2515 3160 2535
rect 3120 2485 3160 2515
rect 3120 2465 3130 2485
rect 3150 2465 3160 2485
rect 3120 2450 3160 2465
rect 3210 2735 3250 2750
rect 3210 2715 3220 2735
rect 3240 2715 3250 2735
rect 3210 2685 3250 2715
rect 3210 2665 3220 2685
rect 3240 2665 3250 2685
rect 3210 2635 3250 2665
rect 3210 2615 3220 2635
rect 3240 2615 3250 2635
rect 3210 2585 3250 2615
rect 3210 2565 3220 2585
rect 3240 2565 3250 2585
rect 3210 2535 3250 2565
rect 3210 2515 3220 2535
rect 3240 2515 3250 2535
rect 3210 2485 3250 2515
rect 3210 2465 3220 2485
rect 3240 2465 3250 2485
rect 3210 2450 3250 2465
rect 3300 2735 3340 2750
rect 3300 2715 3310 2735
rect 3330 2715 3340 2735
rect 3300 2685 3340 2715
rect 3300 2665 3310 2685
rect 3330 2665 3340 2685
rect 3300 2635 3340 2665
rect 3300 2615 3310 2635
rect 3330 2615 3340 2635
rect 3300 2585 3340 2615
rect 3300 2565 3310 2585
rect 3330 2565 3340 2585
rect 3300 2535 3340 2565
rect 3300 2515 3310 2535
rect 3330 2515 3340 2535
rect 3300 2485 3340 2515
rect 3300 2465 3310 2485
rect 3330 2465 3340 2485
rect 3300 2450 3340 2465
rect 3390 2735 3430 2750
rect 3390 2715 3400 2735
rect 3420 2715 3430 2735
rect 3390 2685 3430 2715
rect 3390 2665 3400 2685
rect 3420 2665 3430 2685
rect 3390 2635 3430 2665
rect 3390 2615 3400 2635
rect 3420 2615 3430 2635
rect 3390 2585 3430 2615
rect 3390 2565 3400 2585
rect 3420 2565 3430 2585
rect 3390 2535 3430 2565
rect 3390 2515 3400 2535
rect 3420 2515 3430 2535
rect 3390 2485 3430 2515
rect 3390 2465 3400 2485
rect 3420 2465 3430 2485
rect 3390 2450 3430 2465
rect 3480 2735 3520 2750
rect 3480 2715 3490 2735
rect 3510 2715 3520 2735
rect 3480 2685 3520 2715
rect 3480 2665 3490 2685
rect 3510 2665 3520 2685
rect 3480 2635 3520 2665
rect 3480 2615 3490 2635
rect 3510 2615 3520 2635
rect 3480 2585 3520 2615
rect 3480 2565 3490 2585
rect 3510 2565 3520 2585
rect 3480 2535 3520 2565
rect 3480 2515 3490 2535
rect 3510 2515 3520 2535
rect 3480 2485 3520 2515
rect 3480 2465 3490 2485
rect 3510 2465 3520 2485
rect 3480 2450 3520 2465
rect 3570 2735 3610 2750
rect 3570 2715 3580 2735
rect 3600 2715 3610 2735
rect 3570 2685 3610 2715
rect 3570 2665 3580 2685
rect 3600 2665 3610 2685
rect 3570 2635 3610 2665
rect 3570 2615 3580 2635
rect 3600 2615 3610 2635
rect 3570 2585 3610 2615
rect 3570 2565 3580 2585
rect 3600 2565 3610 2585
rect 3570 2535 3610 2565
rect 3570 2515 3580 2535
rect 3600 2515 3610 2535
rect 3570 2485 3610 2515
rect 3570 2465 3580 2485
rect 3600 2465 3610 2485
rect 3570 2450 3610 2465
rect 3660 2735 3700 2750
rect 3660 2715 3670 2735
rect 3690 2715 3700 2735
rect 3660 2685 3700 2715
rect 3660 2665 3670 2685
rect 3690 2665 3700 2685
rect 3660 2635 3700 2665
rect 3660 2615 3670 2635
rect 3690 2615 3700 2635
rect 3660 2585 3700 2615
rect 3660 2565 3670 2585
rect 3690 2565 3700 2585
rect 3660 2535 3700 2565
rect 3660 2515 3670 2535
rect 3690 2515 3700 2535
rect 3660 2485 3700 2515
rect 3660 2465 3670 2485
rect 3690 2465 3700 2485
rect 3660 2450 3700 2465
rect 3750 2735 3790 2750
rect 3750 2715 3760 2735
rect 3780 2715 3790 2735
rect 3750 2685 3790 2715
rect 3750 2665 3760 2685
rect 3780 2665 3790 2685
rect 3750 2635 3790 2665
rect 3750 2615 3760 2635
rect 3780 2615 3790 2635
rect 3750 2585 3790 2615
rect 3750 2565 3760 2585
rect 3780 2565 3790 2585
rect 3750 2535 3790 2565
rect 3750 2515 3760 2535
rect 3780 2515 3790 2535
rect 3750 2485 3790 2515
rect 3750 2465 3760 2485
rect 3780 2465 3790 2485
rect 3750 2450 3790 2465
rect 3840 2735 3880 2750
rect 3840 2715 3850 2735
rect 3870 2715 3880 2735
rect 3840 2685 3880 2715
rect 3840 2665 3850 2685
rect 3870 2665 3880 2685
rect 3840 2635 3880 2665
rect 3840 2615 3850 2635
rect 3870 2615 3880 2635
rect 3840 2585 3880 2615
rect 3840 2565 3850 2585
rect 3870 2565 3880 2585
rect 3840 2535 3880 2565
rect 3840 2515 3850 2535
rect 3870 2515 3880 2535
rect 3840 2485 3880 2515
rect 3840 2465 3850 2485
rect 3870 2465 3880 2485
rect 3840 2450 3880 2465
rect 3930 2735 3970 2750
rect 3930 2715 3940 2735
rect 3960 2715 3970 2735
rect 3930 2685 3970 2715
rect 3930 2665 3940 2685
rect 3960 2665 3970 2685
rect 3930 2635 3970 2665
rect 3930 2615 3940 2635
rect 3960 2615 3970 2635
rect 3930 2585 3970 2615
rect 3930 2565 3940 2585
rect 3960 2565 3970 2585
rect 3930 2535 3970 2565
rect 3930 2515 3940 2535
rect 3960 2515 3970 2535
rect 3930 2485 3970 2515
rect 3930 2465 3940 2485
rect 3960 2465 3970 2485
rect 3930 2450 3970 2465
rect 4020 2735 4060 2750
rect 4020 2715 4030 2735
rect 4050 2715 4060 2735
rect 4020 2685 4060 2715
rect 4020 2665 4030 2685
rect 4050 2665 4060 2685
rect 4020 2635 4060 2665
rect 4020 2615 4030 2635
rect 4050 2615 4060 2635
rect 4020 2585 4060 2615
rect 4020 2565 4030 2585
rect 4050 2565 4060 2585
rect 4020 2535 4060 2565
rect 4020 2515 4030 2535
rect 4050 2515 4060 2535
rect 4020 2485 4060 2515
rect 4020 2465 4030 2485
rect 4050 2465 4060 2485
rect 4020 2450 4060 2465
rect 4110 2735 4150 2750
rect 4110 2715 4120 2735
rect 4140 2715 4150 2735
rect 4110 2685 4150 2715
rect 4110 2665 4120 2685
rect 4140 2665 4150 2685
rect 4110 2635 4150 2665
rect 4110 2615 4120 2635
rect 4140 2615 4150 2635
rect 4110 2585 4150 2615
rect 4110 2565 4120 2585
rect 4140 2565 4150 2585
rect 4110 2535 4150 2565
rect 4110 2515 4120 2535
rect 4140 2515 4150 2535
rect 4110 2485 4150 2515
rect 4110 2465 4120 2485
rect 4140 2465 4150 2485
rect 4110 2450 4150 2465
rect 4200 2735 4240 2750
rect 4200 2715 4210 2735
rect 4230 2715 4240 2735
rect 4200 2685 4240 2715
rect 4200 2665 4210 2685
rect 4230 2665 4240 2685
rect 4200 2635 4240 2665
rect 4200 2615 4210 2635
rect 4230 2615 4240 2635
rect 4200 2585 4240 2615
rect 4200 2565 4210 2585
rect 4230 2565 4240 2585
rect 4200 2535 4240 2565
rect 4200 2515 4210 2535
rect 4230 2515 4240 2535
rect 4200 2485 4240 2515
rect 4200 2465 4210 2485
rect 4230 2465 4240 2485
rect 4200 2450 4240 2465
rect 4290 2735 4330 2750
rect 4290 2715 4300 2735
rect 4320 2715 4330 2735
rect 4290 2685 4330 2715
rect 4290 2665 4300 2685
rect 4320 2665 4330 2685
rect 4290 2635 4330 2665
rect 4290 2615 4300 2635
rect 4320 2615 4330 2635
rect 4290 2585 4330 2615
rect 4290 2565 4300 2585
rect 4320 2565 4330 2585
rect 4290 2535 4330 2565
rect 4290 2515 4300 2535
rect 4320 2515 4330 2535
rect 4290 2485 4330 2515
rect 4290 2465 4300 2485
rect 4320 2465 4330 2485
rect 4290 2450 4330 2465
rect 4380 2735 4420 2750
rect 4380 2715 4390 2735
rect 4410 2715 4420 2735
rect 4380 2685 4420 2715
rect 4380 2665 4390 2685
rect 4410 2665 4420 2685
rect 4380 2635 4420 2665
rect 4380 2615 4390 2635
rect 4410 2615 4420 2635
rect 4380 2585 4420 2615
rect 4380 2565 4390 2585
rect 4410 2565 4420 2585
rect 4380 2535 4420 2565
rect 4380 2515 4390 2535
rect 4410 2515 4420 2535
rect 4380 2485 4420 2515
rect 4380 2465 4390 2485
rect 4410 2465 4420 2485
rect 4380 2450 4420 2465
rect 4470 2735 4510 2750
rect 4470 2715 4480 2735
rect 4500 2715 4510 2735
rect 4470 2685 4510 2715
rect 4470 2665 4480 2685
rect 4500 2665 4510 2685
rect 4470 2635 4510 2665
rect 4470 2615 4480 2635
rect 4500 2615 4510 2635
rect 4470 2585 4510 2615
rect 4470 2565 4480 2585
rect 4500 2565 4510 2585
rect 4470 2535 4510 2565
rect 4470 2515 4480 2535
rect 4500 2515 4510 2535
rect 4470 2485 4510 2515
rect 4470 2465 4480 2485
rect 4500 2465 4510 2485
rect 4470 2450 4510 2465
rect 4560 2735 4600 2750
rect 4560 2715 4570 2735
rect 4590 2715 4600 2735
rect 4560 2685 4600 2715
rect 4560 2665 4570 2685
rect 4590 2665 4600 2685
rect 4560 2635 4600 2665
rect 4560 2615 4570 2635
rect 4590 2615 4600 2635
rect 4560 2585 4600 2615
rect 4560 2565 4570 2585
rect 4590 2565 4600 2585
rect 4560 2535 4600 2565
rect 4560 2515 4570 2535
rect 4590 2515 4600 2535
rect 4560 2485 4600 2515
rect 4560 2465 4570 2485
rect 4590 2465 4600 2485
rect 4560 2450 4600 2465
rect 4650 2735 4690 2750
rect 4650 2715 4660 2735
rect 4680 2715 4690 2735
rect 4650 2685 4690 2715
rect 4650 2665 4660 2685
rect 4680 2665 4690 2685
rect 4650 2635 4690 2665
rect 4650 2615 4660 2635
rect 4680 2615 4690 2635
rect 4650 2585 4690 2615
rect 4650 2565 4660 2585
rect 4680 2565 4690 2585
rect 4650 2535 4690 2565
rect 4650 2515 4660 2535
rect 4680 2515 4690 2535
rect 4650 2485 4690 2515
rect 4650 2465 4660 2485
rect 4680 2465 4690 2485
rect 4650 2450 4690 2465
rect 4740 2735 4780 2750
rect 4740 2715 4750 2735
rect 4770 2715 4780 2735
rect 4740 2685 4780 2715
rect 4740 2665 4750 2685
rect 4770 2665 4780 2685
rect 4740 2635 4780 2665
rect 4740 2615 4750 2635
rect 4770 2615 4780 2635
rect 4740 2585 4780 2615
rect 4740 2565 4750 2585
rect 4770 2565 4780 2585
rect 4740 2535 4780 2565
rect 4740 2515 4750 2535
rect 4770 2515 4780 2535
rect 4740 2485 4780 2515
rect 4740 2465 4750 2485
rect 4770 2465 4780 2485
rect 4740 2450 4780 2465
rect 4830 2735 4870 2750
rect 4830 2715 4840 2735
rect 4860 2715 4870 2735
rect 4830 2685 4870 2715
rect 4830 2665 4840 2685
rect 4860 2665 4870 2685
rect 4830 2635 4870 2665
rect 4830 2615 4840 2635
rect 4860 2615 4870 2635
rect 4830 2585 4870 2615
rect 4830 2565 4840 2585
rect 4860 2565 4870 2585
rect 4830 2535 4870 2565
rect 4830 2515 4840 2535
rect 4860 2515 4870 2535
rect 4830 2485 4870 2515
rect 4830 2465 4840 2485
rect 4860 2465 4870 2485
rect 4830 2450 4870 2465
rect 4920 2735 4960 2750
rect 4920 2715 4930 2735
rect 4950 2715 4960 2735
rect 4920 2685 4960 2715
rect 4920 2665 4930 2685
rect 4950 2665 4960 2685
rect 4920 2635 4960 2665
rect 4920 2615 4930 2635
rect 4950 2615 4960 2635
rect 4920 2585 4960 2615
rect 4920 2565 4930 2585
rect 4950 2565 4960 2585
rect 4920 2535 4960 2565
rect 4920 2515 4930 2535
rect 4950 2515 4960 2535
rect 4920 2485 4960 2515
rect 4920 2465 4930 2485
rect 4950 2465 4960 2485
rect 4920 2450 4960 2465
rect 5010 2735 5050 2750
rect 5010 2715 5020 2735
rect 5040 2715 5050 2735
rect 5010 2685 5050 2715
rect 5010 2665 5020 2685
rect 5040 2665 5050 2685
rect 5010 2635 5050 2665
rect 5010 2615 5020 2635
rect 5040 2615 5050 2635
rect 5010 2585 5050 2615
rect 5010 2565 5020 2585
rect 5040 2565 5050 2585
rect 5010 2535 5050 2565
rect 5010 2515 5020 2535
rect 5040 2515 5050 2535
rect 5010 2485 5050 2515
rect 5010 2465 5020 2485
rect 5040 2465 5050 2485
rect 5010 2450 5050 2465
rect 5100 2735 5140 2750
rect 5100 2715 5110 2735
rect 5130 2715 5140 2735
rect 5100 2685 5140 2715
rect 5100 2665 5110 2685
rect 5130 2665 5140 2685
rect 5100 2635 5140 2665
rect 5100 2615 5110 2635
rect 5130 2615 5140 2635
rect 5100 2585 5140 2615
rect 5100 2565 5110 2585
rect 5130 2565 5140 2585
rect 5100 2535 5140 2565
rect 5100 2515 5110 2535
rect 5130 2515 5140 2535
rect 5100 2485 5140 2515
rect 5100 2465 5110 2485
rect 5130 2465 5140 2485
rect 5100 2450 5140 2465
rect 2515 1985 2555 2000
rect 2515 1965 2525 1985
rect 2545 1965 2555 1985
rect 2515 1935 2555 1965
rect 2515 1915 2525 1935
rect 2545 1915 2555 1935
rect 2515 1900 2555 1915
rect 2570 1985 2610 2000
rect 2570 1965 2580 1985
rect 2600 1965 2610 1985
rect 2570 1935 2610 1965
rect 2570 1915 2580 1935
rect 2600 1915 2610 1935
rect 2570 1900 2610 1915
rect 2625 1985 2665 2000
rect 2625 1965 2635 1985
rect 2655 1965 2665 1985
rect 2625 1935 2665 1965
rect 2625 1915 2635 1935
rect 2655 1915 2665 1935
rect 2625 1900 2665 1915
rect 2695 1985 2735 2000
rect 2695 1965 2705 1985
rect 2725 1965 2735 1985
rect 2695 1935 2735 1965
rect 2695 1915 2705 1935
rect 2725 1915 2735 1935
rect 2695 1900 2735 1915
rect 2755 1985 2795 2000
rect 2755 1965 2765 1985
rect 2785 1965 2795 1985
rect 2755 1935 2795 1965
rect 2755 1915 2765 1935
rect 2785 1915 2795 1935
rect 2755 1900 2795 1915
rect 2815 1985 2855 2000
rect 2815 1965 2825 1985
rect 2845 1965 2855 1985
rect 2815 1935 2855 1965
rect 2815 1915 2825 1935
rect 2845 1915 2855 1935
rect 2815 1900 2855 1915
rect 2875 1985 2915 2000
rect 2875 1965 2885 1985
rect 2905 1965 2915 1985
rect 2875 1935 2915 1965
rect 2875 1915 2885 1935
rect 2905 1915 2915 1935
rect 2875 1900 2915 1915
rect 2935 1985 2975 2000
rect 2935 1965 2945 1985
rect 2965 1965 2975 1985
rect 2935 1935 2975 1965
rect 2935 1915 2945 1935
rect 2965 1915 2975 1935
rect 2935 1900 2975 1915
rect 2995 1985 3035 2000
rect 2995 1965 3005 1985
rect 3025 1965 3035 1985
rect 2995 1935 3035 1965
rect 2995 1915 3005 1935
rect 3025 1915 3035 1935
rect 2995 1900 3035 1915
rect 3055 1985 3095 2000
rect 3055 1965 3065 1985
rect 3085 1965 3095 1985
rect 3055 1935 3095 1965
rect 3055 1915 3065 1935
rect 3085 1915 3095 1935
rect 3055 1900 3095 1915
rect 3115 1985 3155 2000
rect 3115 1965 3125 1985
rect 3145 1965 3155 1985
rect 3115 1935 3155 1965
rect 3115 1915 3125 1935
rect 3145 1915 3155 1935
rect 3115 1900 3155 1915
rect 3175 1985 3215 2000
rect 3175 1965 3185 1985
rect 3205 1965 3215 1985
rect 3175 1935 3215 1965
rect 3175 1915 3185 1935
rect 3205 1915 3215 1935
rect 3175 1900 3215 1915
rect 3235 1985 3275 2000
rect 3235 1965 3245 1985
rect 3265 1965 3275 1985
rect 3235 1935 3275 1965
rect 3235 1915 3245 1935
rect 3265 1915 3275 1935
rect 3235 1900 3275 1915
rect 3295 1985 3335 2000
rect 3295 1965 3305 1985
rect 3325 1965 3335 1985
rect 3295 1935 3335 1965
rect 3295 1915 3305 1935
rect 3325 1915 3335 1935
rect 3295 1900 3335 1915
rect 3355 1985 3395 2000
rect 3355 1965 3365 1985
rect 3385 1965 3395 1985
rect 3355 1935 3395 1965
rect 3355 1915 3365 1935
rect 3385 1915 3395 1935
rect 3355 1900 3395 1915
rect 3415 1985 3455 2000
rect 3415 1965 3425 1985
rect 3445 1965 3455 1985
rect 3415 1935 3455 1965
rect 3415 1915 3425 1935
rect 3445 1915 3455 1935
rect 3415 1900 3455 1915
rect 3475 1985 3515 2000
rect 3475 1965 3485 1985
rect 3505 1965 3515 1985
rect 3475 1935 3515 1965
rect 3475 1915 3485 1935
rect 3505 1915 3515 1935
rect 3475 1900 3515 1915
rect 3535 1985 3575 2000
rect 3535 1965 3545 1985
rect 3565 1965 3575 1985
rect 3535 1935 3575 1965
rect 3535 1915 3545 1935
rect 3565 1915 3575 1935
rect 3535 1900 3575 1915
rect 3595 1985 3635 2000
rect 3595 1965 3605 1985
rect 3625 1965 3635 1985
rect 3595 1935 3635 1965
rect 3595 1915 3605 1935
rect 3625 1915 3635 1935
rect 3595 1900 3635 1915
rect 3655 1985 3695 2000
rect 3655 1965 3665 1985
rect 3685 1965 3695 1985
rect 3655 1935 3695 1965
rect 3655 1915 3665 1935
rect 3685 1915 3695 1935
rect 3655 1900 3695 1915
rect 3715 1985 3755 2000
rect 3715 1965 3725 1985
rect 3745 1965 3755 1985
rect 3715 1935 3755 1965
rect 3715 1915 3725 1935
rect 3745 1915 3755 1935
rect 3715 1900 3755 1915
rect 3775 1985 3815 2000
rect 3775 1965 3785 1985
rect 3805 1965 3815 1985
rect 3775 1935 3815 1965
rect 3775 1915 3785 1935
rect 3805 1915 3815 1935
rect 3775 1900 3815 1915
rect 3835 1985 3875 2000
rect 3835 1965 3845 1985
rect 3865 1965 3875 1985
rect 3835 1935 3875 1965
rect 3835 1915 3845 1935
rect 3865 1915 3875 1935
rect 3835 1900 3875 1915
rect 3895 1985 3935 2000
rect 3895 1965 3905 1985
rect 3925 1965 3935 1985
rect 3895 1935 3935 1965
rect 3895 1915 3905 1935
rect 3925 1915 3935 1935
rect 3895 1900 3935 1915
rect 3965 1985 4005 2000
rect 3965 1965 3975 1985
rect 3995 1965 4005 1985
rect 3965 1935 4005 1965
rect 3965 1915 3975 1935
rect 3995 1915 4005 1935
rect 3965 1900 4005 1915
rect 4025 1985 4065 2000
rect 4025 1965 4035 1985
rect 4055 1965 4065 1985
rect 4025 1935 4065 1965
rect 4025 1915 4035 1935
rect 4055 1915 4065 1935
rect 4025 1900 4065 1915
rect 4085 1985 4125 2000
rect 4085 1965 4095 1985
rect 4115 1965 4125 1985
rect 4085 1935 4125 1965
rect 4085 1915 4095 1935
rect 4115 1915 4125 1935
rect 4085 1900 4125 1915
rect 4145 1985 4185 2000
rect 4145 1965 4155 1985
rect 4175 1965 4185 1985
rect 4145 1935 4185 1965
rect 4145 1915 4155 1935
rect 4175 1915 4185 1935
rect 4145 1900 4185 1915
rect 4205 1985 4245 2000
rect 4205 1965 4215 1985
rect 4235 1965 4245 1985
rect 4205 1935 4245 1965
rect 4205 1915 4215 1935
rect 4235 1915 4245 1935
rect 4205 1900 4245 1915
rect 4265 1985 4305 2000
rect 4265 1965 4275 1985
rect 4295 1965 4305 1985
rect 4265 1935 4305 1965
rect 4265 1915 4275 1935
rect 4295 1915 4305 1935
rect 4265 1900 4305 1915
rect 4325 1985 4365 2000
rect 4325 1965 4335 1985
rect 4355 1965 4365 1985
rect 4325 1935 4365 1965
rect 4325 1915 4335 1935
rect 4355 1915 4365 1935
rect 4325 1900 4365 1915
rect 4385 1985 4425 2000
rect 4385 1965 4395 1985
rect 4415 1965 4425 1985
rect 4385 1935 4425 1965
rect 4385 1915 4395 1935
rect 4415 1915 4425 1935
rect 4385 1900 4425 1915
rect 4445 1985 4485 2000
rect 4445 1965 4455 1985
rect 4475 1965 4485 1985
rect 4445 1935 4485 1965
rect 4445 1915 4455 1935
rect 4475 1915 4485 1935
rect 4445 1900 4485 1915
rect 4505 1985 4545 2000
rect 4505 1965 4515 1985
rect 4535 1965 4545 1985
rect 4505 1935 4545 1965
rect 4505 1915 4515 1935
rect 4535 1915 4545 1935
rect 4505 1900 4545 1915
rect 4565 1985 4605 2000
rect 4565 1965 4575 1985
rect 4595 1965 4605 1985
rect 4565 1935 4605 1965
rect 4565 1915 4575 1935
rect 4595 1915 4605 1935
rect 4565 1900 4605 1915
rect 4625 1985 4665 2000
rect 4625 1965 4635 1985
rect 4655 1965 4665 1985
rect 4625 1935 4665 1965
rect 4625 1915 4635 1935
rect 4655 1915 4665 1935
rect 4625 1900 4665 1915
rect 4685 1985 4725 2000
rect 4685 1965 4695 1985
rect 4715 1965 4725 1985
rect 4685 1935 4725 1965
rect 4685 1915 4695 1935
rect 4715 1915 4725 1935
rect 4685 1900 4725 1915
rect 4745 1985 4785 2000
rect 4745 1965 4755 1985
rect 4775 1965 4785 1985
rect 4745 1935 4785 1965
rect 4745 1915 4755 1935
rect 4775 1915 4785 1935
rect 4745 1900 4785 1915
rect 4805 1985 4845 2000
rect 4805 1965 4815 1985
rect 4835 1965 4845 1985
rect 4805 1935 4845 1965
rect 4805 1915 4815 1935
rect 4835 1915 4845 1935
rect 4805 1900 4845 1915
rect 4865 1985 4905 2000
rect 4865 1965 4875 1985
rect 4895 1965 4905 1985
rect 4865 1935 4905 1965
rect 4865 1915 4875 1935
rect 4895 1915 4905 1935
rect 4865 1900 4905 1915
rect 4925 1985 4965 2000
rect 4925 1965 4935 1985
rect 4955 1965 4965 1985
rect 4925 1935 4965 1965
rect 4925 1915 4935 1935
rect 4955 1915 4965 1935
rect 4925 1900 4965 1915
rect 4985 1985 5025 2000
rect 4985 1965 4995 1985
rect 5015 1965 5025 1985
rect 4985 1935 5025 1965
rect 4985 1915 4995 1935
rect 5015 1915 5025 1935
rect 4985 1900 5025 1915
rect 5045 1985 5085 2000
rect 5045 1965 5055 1985
rect 5075 1965 5085 1985
rect 5045 1935 5085 1965
rect 5045 1915 5055 1935
rect 5075 1915 5085 1935
rect 5045 1900 5085 1915
rect 5105 1985 5145 2000
rect 5105 1965 5115 1985
rect 5135 1965 5145 1985
rect 5105 1935 5145 1965
rect 5105 1915 5115 1935
rect 5135 1915 5145 1935
rect 5105 1900 5145 1915
rect 5165 1985 5205 2000
rect 5165 1965 5175 1985
rect 5195 1965 5205 1985
rect 5165 1935 5205 1965
rect 5165 1915 5175 1935
rect 5195 1915 5205 1935
rect 5165 1900 5205 1915
rect 3115 1650 3155 1665
rect 3115 1630 3125 1650
rect 3145 1630 3155 1650
rect 3115 1615 3155 1630
rect 3175 1650 3215 1665
rect 3175 1630 3185 1650
rect 3205 1630 3215 1650
rect 3175 1615 3215 1630
rect 3235 1650 3275 1665
rect 3235 1630 3245 1650
rect 3265 1630 3275 1650
rect 3235 1615 3275 1630
rect 3295 1650 3335 1665
rect 3295 1630 3305 1650
rect 3325 1630 3335 1650
rect 3295 1615 3335 1630
rect 3355 1650 3395 1665
rect 3355 1630 3365 1650
rect 3385 1630 3395 1650
rect 3355 1615 3395 1630
rect 3415 1650 3455 1665
rect 3415 1630 3425 1650
rect 3445 1630 3455 1650
rect 3415 1615 3455 1630
rect 3475 1650 3515 1665
rect 3475 1630 3485 1650
rect 3505 1630 3515 1650
rect 3475 1615 3515 1630
rect 3535 1650 3575 1665
rect 3535 1630 3545 1650
rect 3565 1630 3575 1650
rect 3535 1615 3575 1630
rect 3595 1650 3635 1665
rect 3595 1630 3605 1650
rect 3625 1630 3635 1650
rect 3595 1615 3635 1630
rect 3655 1650 3695 1665
rect 3655 1630 3665 1650
rect 3685 1630 3695 1650
rect 3655 1615 3695 1630
rect 3715 1650 3755 1665
rect 3715 1630 3725 1650
rect 3745 1630 3755 1650
rect 3715 1615 3755 1630
rect 4145 1650 4185 1665
rect 4145 1630 4155 1650
rect 4175 1630 4185 1650
rect 4145 1615 4185 1630
rect 4205 1650 4245 1665
rect 4205 1630 4215 1650
rect 4235 1630 4245 1650
rect 4205 1615 4245 1630
rect 4265 1650 4305 1665
rect 4265 1630 4275 1650
rect 4295 1630 4305 1650
rect 4265 1615 4305 1630
rect 4325 1650 4365 1665
rect 4325 1630 4335 1650
rect 4355 1630 4365 1650
rect 4325 1615 4365 1630
rect 4385 1650 4425 1665
rect 4385 1630 4395 1650
rect 4415 1630 4425 1650
rect 4385 1615 4425 1630
rect 4445 1650 4485 1665
rect 4445 1630 4455 1650
rect 4475 1630 4485 1650
rect 4445 1615 4485 1630
rect 4505 1650 4545 1665
rect 4505 1630 4515 1650
rect 4535 1630 4545 1650
rect 4505 1615 4545 1630
rect 4565 1650 4605 1665
rect 4565 1630 4575 1650
rect 4595 1630 4605 1650
rect 4565 1615 4605 1630
rect 4625 1650 4665 1665
rect 4625 1630 4635 1650
rect 4655 1630 4665 1650
rect 4625 1615 4665 1630
rect 4685 1650 4725 1665
rect 4685 1630 4695 1650
rect 4715 1630 4725 1650
rect 4685 1615 4725 1630
rect 4745 1650 4785 1665
rect 4745 1630 4755 1650
rect 4775 1630 4785 1650
rect 4745 1615 4785 1630
rect 2785 1445 2825 1460
rect 2785 1425 2795 1445
rect 2815 1425 2825 1445
rect 2785 1395 2825 1425
rect 2785 1375 2795 1395
rect 2815 1375 2825 1395
rect 2785 1345 2825 1375
rect 2785 1325 2795 1345
rect 2815 1325 2825 1345
rect 2785 1295 2825 1325
rect 2785 1275 2795 1295
rect 2815 1275 2825 1295
rect 2785 1245 2825 1275
rect 2785 1225 2795 1245
rect 2815 1225 2825 1245
rect 2785 1210 2825 1225
rect 3325 1445 3365 1460
rect 3325 1425 3335 1445
rect 3355 1425 3365 1445
rect 3325 1395 3365 1425
rect 3325 1375 3335 1395
rect 3355 1375 3365 1395
rect 3325 1345 3365 1375
rect 3325 1325 3335 1345
rect 3355 1325 3365 1345
rect 3325 1295 3365 1325
rect 3325 1275 3335 1295
rect 3355 1275 3365 1295
rect 3325 1245 3365 1275
rect 3325 1225 3335 1245
rect 3355 1225 3365 1245
rect 3325 1210 3365 1225
rect 3865 1445 3905 1460
rect 3865 1425 3875 1445
rect 3895 1425 3905 1445
rect 3865 1395 3905 1425
rect 3865 1375 3875 1395
rect 3895 1375 3905 1395
rect 3865 1345 3905 1375
rect 3865 1325 3875 1345
rect 3895 1325 3905 1345
rect 3865 1295 3905 1325
rect 3865 1275 3875 1295
rect 3895 1275 3905 1295
rect 3865 1245 3905 1275
rect 3865 1225 3875 1245
rect 3895 1225 3905 1245
rect 3865 1210 3905 1225
rect 3995 1445 4035 1460
rect 3995 1425 4005 1445
rect 4025 1425 4035 1445
rect 3995 1395 4035 1425
rect 3995 1375 4005 1395
rect 4025 1375 4035 1395
rect 3995 1345 4035 1375
rect 3995 1325 4005 1345
rect 4025 1325 4035 1345
rect 3995 1295 4035 1325
rect 3995 1275 4005 1295
rect 4025 1275 4035 1295
rect 3995 1245 4035 1275
rect 3995 1225 4005 1245
rect 4025 1225 4035 1245
rect 3995 1210 4035 1225
rect 4535 1445 4575 1460
rect 4535 1425 4545 1445
rect 4565 1425 4575 1445
rect 4535 1395 4575 1425
rect 4535 1375 4545 1395
rect 4565 1375 4575 1395
rect 4535 1345 4575 1375
rect 4535 1325 4545 1345
rect 4565 1325 4575 1345
rect 4535 1295 4575 1325
rect 4535 1275 4545 1295
rect 4565 1275 4575 1295
rect 4535 1245 4575 1275
rect 4535 1225 4545 1245
rect 4565 1225 4575 1245
rect 4535 1210 4575 1225
rect 5075 1445 5115 1460
rect 5075 1425 5085 1445
rect 5105 1425 5115 1445
rect 5075 1395 5115 1425
rect 5075 1375 5085 1395
rect 5105 1375 5115 1395
rect 5075 1345 5115 1375
rect 5075 1325 5085 1345
rect 5105 1325 5115 1345
rect 5075 1295 5115 1325
rect 5075 1275 5085 1295
rect 5105 1275 5115 1295
rect 5075 1245 5115 1275
rect 5075 1225 5085 1245
rect 5105 1225 5115 1245
rect 5075 1210 5115 1225
rect 2890 1100 2930 1115
rect 2890 1080 2900 1100
rect 2920 1080 2930 1100
rect 2890 1050 2930 1080
rect 2890 1030 2900 1050
rect 2920 1030 2930 1050
rect 2890 1015 2930 1030
rect 3930 1100 3970 1115
rect 3930 1080 3940 1100
rect 3960 1080 3970 1100
rect 3930 1050 3970 1080
rect 3930 1030 3940 1050
rect 3960 1030 3970 1050
rect 3930 1015 3970 1030
rect 4970 1100 5010 1115
rect 4970 1080 4980 1100
rect 5000 1080 5010 1100
rect 4970 1050 5010 1080
rect 4970 1030 4980 1050
rect 5000 1030 5010 1050
rect 4970 1015 5010 1030
rect 3040 895 3080 910
rect 3040 875 3050 895
rect 3070 875 3080 895
rect 3040 845 3080 875
rect 3040 825 3050 845
rect 3070 825 3080 845
rect 3040 810 3080 825
rect 3130 895 3170 910
rect 3130 875 3140 895
rect 3160 875 3170 895
rect 3130 845 3170 875
rect 3130 825 3140 845
rect 3160 825 3170 845
rect 3130 810 3170 825
rect 3200 895 3240 910
rect 3200 875 3210 895
rect 3230 875 3240 895
rect 3200 845 3240 875
rect 3200 825 3210 845
rect 3230 825 3240 845
rect 3200 810 3240 825
rect 3290 895 3330 910
rect 3290 875 3300 895
rect 3320 875 3330 895
rect 3290 845 3330 875
rect 3290 825 3300 845
rect 3320 825 3330 845
rect 3290 810 3330 825
rect 3380 895 3420 910
rect 3380 875 3390 895
rect 3410 875 3420 895
rect 3380 845 3420 875
rect 3380 825 3390 845
rect 3410 825 3420 845
rect 3380 810 3420 825
rect 3470 895 3510 910
rect 3470 875 3480 895
rect 3500 875 3510 895
rect 3470 845 3510 875
rect 3470 825 3480 845
rect 3500 825 3510 845
rect 3470 810 3510 825
rect 3560 895 3600 910
rect 3560 875 3570 895
rect 3590 875 3600 895
rect 3560 845 3600 875
rect 3560 825 3570 845
rect 3590 825 3600 845
rect 3560 810 3600 825
rect 3650 895 3690 910
rect 3650 875 3660 895
rect 3680 875 3690 895
rect 3650 845 3690 875
rect 3650 825 3660 845
rect 3680 825 3690 845
rect 3650 810 3690 825
rect 3740 895 3780 910
rect 3740 875 3750 895
rect 3770 875 3780 895
rect 3740 845 3780 875
rect 3740 825 3750 845
rect 3770 825 3780 845
rect 3740 810 3780 825
rect 3830 895 3870 910
rect 3830 875 3840 895
rect 3860 875 3870 895
rect 3830 845 3870 875
rect 3830 825 3840 845
rect 3860 825 3870 845
rect 3830 810 3870 825
rect 3920 895 3960 910
rect 3920 875 3930 895
rect 3950 875 3960 895
rect 3920 845 3960 875
rect 3920 825 3930 845
rect 3950 825 3960 845
rect 3920 810 3960 825
rect 4010 895 4050 910
rect 4010 875 4020 895
rect 4040 875 4050 895
rect 4010 845 4050 875
rect 4010 825 4020 845
rect 4040 825 4050 845
rect 4010 810 4050 825
rect 4100 895 4140 910
rect 4100 875 4110 895
rect 4130 875 4140 895
rect 4100 845 4140 875
rect 4100 825 4110 845
rect 4130 825 4140 845
rect 4100 810 4140 825
rect 4190 895 4230 910
rect 4190 875 4200 895
rect 4220 875 4230 895
rect 4190 845 4230 875
rect 4190 825 4200 845
rect 4220 825 4230 845
rect 4190 810 4230 825
rect 4280 895 4320 910
rect 4280 875 4290 895
rect 4310 875 4320 895
rect 4280 845 4320 875
rect 4280 825 4290 845
rect 4310 825 4320 845
rect 4280 810 4320 825
rect 4370 895 4410 910
rect 4370 875 4380 895
rect 4400 875 4410 895
rect 4370 845 4410 875
rect 4370 825 4380 845
rect 4400 825 4410 845
rect 4370 810 4410 825
rect 4460 895 4500 910
rect 4460 875 4470 895
rect 4490 875 4500 895
rect 4460 845 4500 875
rect 4460 825 4470 845
rect 4490 825 4500 845
rect 4460 810 4500 825
rect 4550 895 4590 910
rect 4550 875 4560 895
rect 4580 875 4590 895
rect 4550 845 4590 875
rect 4550 825 4560 845
rect 4580 825 4590 845
rect 4550 810 4590 825
rect 4640 895 4680 910
rect 4640 875 4650 895
rect 4670 875 4680 895
rect 4640 845 4680 875
rect 4640 825 4650 845
rect 4670 825 4680 845
rect 4640 810 4680 825
rect 4730 895 4770 910
rect 4730 875 4740 895
rect 4760 875 4770 895
rect 4730 845 4770 875
rect 4730 825 4740 845
rect 4760 825 4770 845
rect 4730 810 4770 825
rect 4820 895 4860 910
rect 4820 875 4830 895
rect 4850 875 4860 895
rect 4820 845 4860 875
rect 4820 825 4830 845
rect 4850 825 4860 845
rect 4820 810 4860 825
rect 4910 895 4950 910
rect 4910 875 4920 895
rect 4940 875 4950 895
rect 4910 845 4950 875
rect 4910 825 4920 845
rect 4940 825 4950 845
rect 4910 810 4950 825
<< ndiffc >>
rect 2955 2955 2975 2975
rect 2955 2905 2975 2925
rect 3045 2955 3065 2975
rect 3045 2905 3065 2925
rect 3135 2955 3155 2975
rect 3135 2905 3155 2925
rect 3205 2955 3225 2975
rect 3205 2905 3225 2925
rect 3295 2955 3315 2975
rect 3295 2905 3315 2925
rect 3385 2955 3405 2975
rect 3385 2905 3405 2925
rect 3475 2955 3495 2975
rect 3475 2905 3495 2925
rect 3565 2955 3585 2975
rect 3565 2905 3585 2925
rect 3655 2955 3675 2975
rect 3655 2905 3675 2925
rect 3745 2955 3765 2975
rect 3745 2905 3765 2925
rect 3835 2955 3855 2975
rect 3835 2905 3855 2925
rect 3925 2955 3945 2975
rect 3925 2905 3945 2925
rect 4015 2955 4035 2975
rect 4015 2905 4035 2925
rect 4105 2955 4125 2975
rect 4105 2905 4125 2925
rect 4195 2955 4215 2975
rect 4195 2905 4215 2925
rect 4285 2955 4305 2975
rect 4285 2905 4305 2925
rect 4375 2955 4395 2975
rect 4375 2905 4395 2925
rect 4465 2955 4485 2975
rect 4465 2905 4485 2925
rect 4555 2955 4575 2975
rect 4555 2905 4575 2925
rect 4645 2955 4665 2975
rect 4645 2905 4665 2925
rect 4735 2955 4755 2975
rect 4735 2905 4755 2925
rect 4825 2955 4845 2975
rect 4825 2905 4845 2925
rect 4915 2955 4935 2975
rect 4915 2905 4935 2925
rect 5005 2955 5025 2975
rect 5005 2905 5025 2925
rect 2770 2715 2790 2735
rect 2770 2665 2790 2685
rect 2770 2615 2790 2635
rect 2770 2565 2790 2585
rect 2770 2515 2790 2535
rect 2770 2465 2790 2485
rect 2860 2715 2880 2735
rect 2860 2665 2880 2685
rect 2860 2615 2880 2635
rect 2860 2565 2880 2585
rect 2860 2515 2880 2535
rect 2860 2465 2880 2485
rect 2950 2715 2970 2735
rect 2950 2665 2970 2685
rect 2950 2615 2970 2635
rect 2950 2565 2970 2585
rect 2950 2515 2970 2535
rect 2950 2465 2970 2485
rect 3040 2715 3060 2735
rect 3040 2665 3060 2685
rect 3040 2615 3060 2635
rect 3040 2565 3060 2585
rect 3040 2515 3060 2535
rect 3040 2465 3060 2485
rect 3130 2715 3150 2735
rect 3130 2665 3150 2685
rect 3130 2615 3150 2635
rect 3130 2565 3150 2585
rect 3130 2515 3150 2535
rect 3130 2465 3150 2485
rect 3220 2715 3240 2735
rect 3220 2665 3240 2685
rect 3220 2615 3240 2635
rect 3220 2565 3240 2585
rect 3220 2515 3240 2535
rect 3220 2465 3240 2485
rect 3310 2715 3330 2735
rect 3310 2665 3330 2685
rect 3310 2615 3330 2635
rect 3310 2565 3330 2585
rect 3310 2515 3330 2535
rect 3310 2465 3330 2485
rect 3400 2715 3420 2735
rect 3400 2665 3420 2685
rect 3400 2615 3420 2635
rect 3400 2565 3420 2585
rect 3400 2515 3420 2535
rect 3400 2465 3420 2485
rect 3490 2715 3510 2735
rect 3490 2665 3510 2685
rect 3490 2615 3510 2635
rect 3490 2565 3510 2585
rect 3490 2515 3510 2535
rect 3490 2465 3510 2485
rect 3580 2715 3600 2735
rect 3580 2665 3600 2685
rect 3580 2615 3600 2635
rect 3580 2565 3600 2585
rect 3580 2515 3600 2535
rect 3580 2465 3600 2485
rect 3670 2715 3690 2735
rect 3670 2665 3690 2685
rect 3670 2615 3690 2635
rect 3670 2565 3690 2585
rect 3670 2515 3690 2535
rect 3670 2465 3690 2485
rect 3760 2715 3780 2735
rect 3760 2665 3780 2685
rect 3760 2615 3780 2635
rect 3760 2565 3780 2585
rect 3760 2515 3780 2535
rect 3760 2465 3780 2485
rect 3850 2715 3870 2735
rect 3850 2665 3870 2685
rect 3850 2615 3870 2635
rect 3850 2565 3870 2585
rect 3850 2515 3870 2535
rect 3850 2465 3870 2485
rect 3940 2715 3960 2735
rect 3940 2665 3960 2685
rect 3940 2615 3960 2635
rect 3940 2565 3960 2585
rect 3940 2515 3960 2535
rect 3940 2465 3960 2485
rect 4030 2715 4050 2735
rect 4030 2665 4050 2685
rect 4030 2615 4050 2635
rect 4030 2565 4050 2585
rect 4030 2515 4050 2535
rect 4030 2465 4050 2485
rect 4120 2715 4140 2735
rect 4120 2665 4140 2685
rect 4120 2615 4140 2635
rect 4120 2565 4140 2585
rect 4120 2515 4140 2535
rect 4120 2465 4140 2485
rect 4210 2715 4230 2735
rect 4210 2665 4230 2685
rect 4210 2615 4230 2635
rect 4210 2565 4230 2585
rect 4210 2515 4230 2535
rect 4210 2465 4230 2485
rect 4300 2715 4320 2735
rect 4300 2665 4320 2685
rect 4300 2615 4320 2635
rect 4300 2565 4320 2585
rect 4300 2515 4320 2535
rect 4300 2465 4320 2485
rect 4390 2715 4410 2735
rect 4390 2665 4410 2685
rect 4390 2615 4410 2635
rect 4390 2565 4410 2585
rect 4390 2515 4410 2535
rect 4390 2465 4410 2485
rect 4480 2715 4500 2735
rect 4480 2665 4500 2685
rect 4480 2615 4500 2635
rect 4480 2565 4500 2585
rect 4480 2515 4500 2535
rect 4480 2465 4500 2485
rect 4570 2715 4590 2735
rect 4570 2665 4590 2685
rect 4570 2615 4590 2635
rect 4570 2565 4590 2585
rect 4570 2515 4590 2535
rect 4570 2465 4590 2485
rect 4660 2715 4680 2735
rect 4660 2665 4680 2685
rect 4660 2615 4680 2635
rect 4660 2565 4680 2585
rect 4660 2515 4680 2535
rect 4660 2465 4680 2485
rect 4750 2715 4770 2735
rect 4750 2665 4770 2685
rect 4750 2615 4770 2635
rect 4750 2565 4770 2585
rect 4750 2515 4770 2535
rect 4750 2465 4770 2485
rect 4840 2715 4860 2735
rect 4840 2665 4860 2685
rect 4840 2615 4860 2635
rect 4840 2565 4860 2585
rect 4840 2515 4860 2535
rect 4840 2465 4860 2485
rect 4930 2715 4950 2735
rect 4930 2665 4950 2685
rect 4930 2615 4950 2635
rect 4930 2565 4950 2585
rect 4930 2515 4950 2535
rect 4930 2465 4950 2485
rect 5020 2715 5040 2735
rect 5020 2665 5040 2685
rect 5020 2615 5040 2635
rect 5020 2565 5040 2585
rect 5020 2515 5040 2535
rect 5020 2465 5040 2485
rect 5110 2715 5130 2735
rect 5110 2665 5130 2685
rect 5110 2615 5130 2635
rect 5110 2565 5130 2585
rect 5110 2515 5130 2535
rect 5110 2465 5130 2485
rect 2525 1965 2545 1985
rect 2525 1915 2545 1935
rect 2580 1965 2600 1985
rect 2580 1915 2600 1935
rect 2635 1965 2655 1985
rect 2635 1915 2655 1935
rect 2705 1965 2725 1985
rect 2705 1915 2725 1935
rect 2765 1965 2785 1985
rect 2765 1915 2785 1935
rect 2825 1965 2845 1985
rect 2825 1915 2845 1935
rect 2885 1965 2905 1985
rect 2885 1915 2905 1935
rect 2945 1965 2965 1985
rect 2945 1915 2965 1935
rect 3005 1965 3025 1985
rect 3005 1915 3025 1935
rect 3065 1965 3085 1985
rect 3065 1915 3085 1935
rect 3125 1965 3145 1985
rect 3125 1915 3145 1935
rect 3185 1965 3205 1985
rect 3185 1915 3205 1935
rect 3245 1965 3265 1985
rect 3245 1915 3265 1935
rect 3305 1965 3325 1985
rect 3305 1915 3325 1935
rect 3365 1965 3385 1985
rect 3365 1915 3385 1935
rect 3425 1965 3445 1985
rect 3425 1915 3445 1935
rect 3485 1965 3505 1985
rect 3485 1915 3505 1935
rect 3545 1965 3565 1985
rect 3545 1915 3565 1935
rect 3605 1965 3625 1985
rect 3605 1915 3625 1935
rect 3665 1965 3685 1985
rect 3665 1915 3685 1935
rect 3725 1965 3745 1985
rect 3725 1915 3745 1935
rect 3785 1965 3805 1985
rect 3785 1915 3805 1935
rect 3845 1965 3865 1985
rect 3845 1915 3865 1935
rect 3905 1965 3925 1985
rect 3905 1915 3925 1935
rect 3975 1965 3995 1985
rect 3975 1915 3995 1935
rect 4035 1965 4055 1985
rect 4035 1915 4055 1935
rect 4095 1965 4115 1985
rect 4095 1915 4115 1935
rect 4155 1965 4175 1985
rect 4155 1915 4175 1935
rect 4215 1965 4235 1985
rect 4215 1915 4235 1935
rect 4275 1965 4295 1985
rect 4275 1915 4295 1935
rect 4335 1965 4355 1985
rect 4335 1915 4355 1935
rect 4395 1965 4415 1985
rect 4395 1915 4415 1935
rect 4455 1965 4475 1985
rect 4455 1915 4475 1935
rect 4515 1965 4535 1985
rect 4515 1915 4535 1935
rect 4575 1965 4595 1985
rect 4575 1915 4595 1935
rect 4635 1965 4655 1985
rect 4635 1915 4655 1935
rect 4695 1965 4715 1985
rect 4695 1915 4715 1935
rect 4755 1965 4775 1985
rect 4755 1915 4775 1935
rect 4815 1965 4835 1985
rect 4815 1915 4835 1935
rect 4875 1965 4895 1985
rect 4875 1915 4895 1935
rect 4935 1965 4955 1985
rect 4935 1915 4955 1935
rect 4995 1965 5015 1985
rect 4995 1915 5015 1935
rect 5055 1965 5075 1985
rect 5055 1915 5075 1935
rect 5115 1965 5135 1985
rect 5115 1915 5135 1935
rect 5175 1965 5195 1985
rect 5175 1915 5195 1935
rect 3125 1630 3145 1650
rect 3185 1630 3205 1650
rect 3245 1630 3265 1650
rect 3305 1630 3325 1650
rect 3365 1630 3385 1650
rect 3425 1630 3445 1650
rect 3485 1630 3505 1650
rect 3545 1630 3565 1650
rect 3605 1630 3625 1650
rect 3665 1630 3685 1650
rect 3725 1630 3745 1650
rect 4155 1630 4175 1650
rect 4215 1630 4235 1650
rect 4275 1630 4295 1650
rect 4335 1630 4355 1650
rect 4395 1630 4415 1650
rect 4455 1630 4475 1650
rect 4515 1630 4535 1650
rect 4575 1630 4595 1650
rect 4635 1630 4655 1650
rect 4695 1630 4715 1650
rect 4755 1630 4775 1650
rect 2795 1425 2815 1445
rect 2795 1375 2815 1395
rect 2795 1325 2815 1345
rect 2795 1275 2815 1295
rect 2795 1225 2815 1245
rect 3335 1425 3355 1445
rect 3335 1375 3355 1395
rect 3335 1325 3355 1345
rect 3335 1275 3355 1295
rect 3335 1225 3355 1245
rect 3875 1425 3895 1445
rect 3875 1375 3895 1395
rect 3875 1325 3895 1345
rect 3875 1275 3895 1295
rect 3875 1225 3895 1245
rect 4005 1425 4025 1445
rect 4005 1375 4025 1395
rect 4005 1325 4025 1345
rect 4005 1275 4025 1295
rect 4005 1225 4025 1245
rect 4545 1425 4565 1445
rect 4545 1375 4565 1395
rect 4545 1325 4565 1345
rect 4545 1275 4565 1295
rect 4545 1225 4565 1245
rect 5085 1425 5105 1445
rect 5085 1375 5105 1395
rect 5085 1325 5105 1345
rect 5085 1275 5105 1295
rect 5085 1225 5105 1245
rect 2900 1080 2920 1100
rect 2900 1030 2920 1050
rect 3940 1080 3960 1100
rect 3940 1030 3960 1050
rect 4980 1080 5000 1100
rect 4980 1030 5000 1050
rect 3050 875 3070 895
rect 3050 825 3070 845
rect 3140 875 3160 895
rect 3140 825 3160 845
rect 3210 875 3230 895
rect 3210 825 3230 845
rect 3300 875 3320 895
rect 3300 825 3320 845
rect 3390 875 3410 895
rect 3390 825 3410 845
rect 3480 875 3500 895
rect 3480 825 3500 845
rect 3570 875 3590 895
rect 3570 825 3590 845
rect 3660 875 3680 895
rect 3660 825 3680 845
rect 3750 875 3770 895
rect 3750 825 3770 845
rect 3840 875 3860 895
rect 3840 825 3860 845
rect 3930 875 3950 895
rect 3930 825 3950 845
rect 4020 875 4040 895
rect 4020 825 4040 845
rect 4110 875 4130 895
rect 4110 825 4130 845
rect 4200 875 4220 895
rect 4200 825 4220 845
rect 4290 875 4310 895
rect 4290 825 4310 845
rect 4380 875 4400 895
rect 4380 825 4400 845
rect 4470 875 4490 895
rect 4470 825 4490 845
rect 4560 875 4580 895
rect 4560 825 4580 845
rect 4650 875 4670 895
rect 4650 825 4670 845
rect 4740 875 4760 895
rect 4740 825 4760 845
rect 4830 875 4850 895
rect 4830 825 4850 845
rect 4920 875 4940 895
rect 4920 825 4940 845
<< psubdiff >>
rect -50 1715 100 1730
rect -50 1695 -35 1715
rect -15 1695 15 1715
rect 35 1695 65 1715
rect 85 1695 100 1715
rect -50 1680 100 1695
<< psubdiffcont >>
rect -35 1695 -15 1715
rect 15 1695 35 1715
rect 65 1695 85 1715
<< poly >>
rect 2985 2990 3035 3005
rect 3075 2990 3125 3005
rect 3235 2990 3285 3005
rect 3325 2990 3375 3005
rect 3415 2990 3465 3005
rect 3505 2990 3555 3005
rect 3595 2990 3645 3005
rect 3685 2990 3735 3005
rect 3775 2990 3825 3005
rect 3865 2990 3915 3005
rect 3955 2990 4005 3005
rect 4045 2990 4095 3005
rect 4135 2990 4185 3005
rect 4225 2990 4275 3005
rect 4315 2990 4365 3005
rect 4405 2990 4455 3005
rect 4495 2990 4545 3005
rect 4585 2990 4635 3005
rect 4675 2990 4725 3005
rect 4765 2990 4815 3005
rect 4855 2990 4905 3005
rect 4945 2990 4995 3005
rect 2985 2875 3035 2890
rect 3075 2875 3125 2890
rect 3235 2875 3285 2890
rect 3325 2875 3375 2890
rect 3415 2875 3465 2890
rect 3505 2875 3555 2890
rect 3595 2875 3645 2890
rect 3685 2875 3735 2890
rect 3775 2875 3825 2890
rect 3865 2875 3915 2890
rect 3955 2875 4005 2890
rect 4045 2875 4095 2890
rect 4135 2875 4185 2890
rect 4225 2875 4275 2890
rect 4315 2875 4365 2890
rect 4405 2875 4455 2890
rect 4495 2875 4545 2890
rect 4585 2875 4635 2890
rect 4675 2875 4725 2890
rect 4765 2875 4815 2890
rect 4855 2875 4905 2890
rect 4945 2875 4995 2890
rect 2800 2750 2850 2765
rect 2890 2750 2940 2765
rect 2980 2750 3030 2765
rect 3070 2750 3120 2765
rect 3160 2750 3210 2765
rect 3250 2750 3300 2765
rect 3340 2750 3390 2765
rect 3430 2750 3480 2765
rect 3520 2750 3570 2765
rect 3610 2750 3660 2765
rect 3700 2750 3750 2765
rect 3790 2750 3840 2765
rect 3880 2750 3930 2765
rect 3970 2750 4020 2765
rect 4060 2750 4110 2765
rect 4150 2750 4200 2765
rect 4240 2750 4290 2765
rect 4330 2750 4380 2765
rect 4420 2750 4470 2765
rect 4510 2750 4560 2765
rect 4600 2750 4650 2765
rect 4690 2750 4740 2765
rect 4780 2750 4830 2765
rect 4870 2750 4920 2765
rect 4960 2750 5010 2765
rect 5050 2750 5100 2765
rect 2800 2440 2850 2450
rect 2760 2425 2850 2440
rect 2890 2440 2940 2450
rect 2980 2440 3030 2450
rect 3070 2440 3120 2450
rect 3160 2440 3210 2450
rect 3250 2440 3300 2450
rect 3340 2440 3390 2450
rect 3430 2440 3480 2450
rect 3520 2440 3570 2450
rect 3610 2440 3660 2450
rect 3700 2440 3750 2450
rect 3790 2440 3840 2450
rect 3880 2440 3930 2450
rect 3970 2440 4020 2450
rect 4060 2440 4110 2450
rect 4150 2440 4200 2450
rect 4240 2440 4290 2450
rect 4330 2440 4380 2450
rect 4420 2440 4470 2450
rect 4510 2440 4560 2450
rect 4600 2440 4650 2450
rect 4690 2440 4740 2450
rect 4780 2440 4830 2450
rect 4870 2440 4920 2450
rect 4960 2440 5010 2450
rect 2890 2425 5010 2440
rect 5050 2440 5100 2450
rect 5050 2425 5140 2440
rect 2760 2405 2770 2425
rect 2790 2405 2800 2425
rect 2760 2395 2800 2405
rect 2940 2420 2980 2425
rect 2940 2400 2950 2420
rect 2970 2400 2980 2420
rect 2940 2390 2980 2400
rect 3835 2405 3845 2425
rect 3865 2405 3875 2425
rect 3835 2395 3875 2405
rect 5100 2405 5110 2425
rect 5130 2405 5140 2425
rect 5100 2395 5140 2405
rect 2695 2045 2735 2055
rect 2695 2025 2705 2045
rect 2725 2030 2735 2045
rect 3895 2045 3935 2055
rect 3895 2030 3905 2045
rect 2725 2025 2755 2030
rect 2695 2015 2755 2025
rect 3875 2025 3905 2030
rect 3925 2025 3935 2045
rect 3875 2015 3935 2025
rect 3965 2045 4005 2055
rect 3965 2025 3975 2045
rect 3995 2030 4005 2045
rect 5165 2045 5205 2055
rect 5165 2030 5175 2045
rect 3995 2025 4025 2030
rect 3965 2015 4025 2025
rect 5145 2025 5175 2030
rect 5195 2025 5205 2045
rect 5145 2015 5205 2025
rect 2555 2000 2570 2015
rect 2610 2000 2625 2015
rect 2735 2000 2755 2015
rect 2795 2000 2815 2015
rect 2855 2000 2875 2015
rect 2915 2000 2935 2015
rect 2975 2000 2995 2015
rect 3035 2000 3055 2015
rect 3095 2000 3115 2015
rect 3155 2000 3175 2015
rect 3215 2000 3235 2015
rect 3275 2000 3295 2015
rect 3335 2000 3355 2015
rect 3395 2000 3415 2015
rect 3455 2000 3475 2015
rect 3515 2000 3535 2015
rect 3575 2000 3595 2015
rect 3635 2000 3655 2015
rect 3695 2000 3715 2015
rect 3755 2000 3775 2015
rect 3815 2000 3835 2015
rect 3875 2000 3895 2015
rect 4005 2000 4025 2015
rect 4065 2000 4085 2015
rect 4125 2000 4145 2015
rect 4185 2000 4205 2015
rect 4245 2000 4265 2015
rect 4305 2000 4325 2015
rect 4365 2000 4385 2015
rect 4425 2000 4445 2015
rect 4485 2000 4505 2015
rect 4545 2000 4565 2015
rect 4605 2000 4625 2015
rect 4665 2000 4685 2015
rect 4725 2000 4745 2015
rect 4785 2000 4805 2015
rect 4845 2000 4865 2015
rect 4905 2000 4925 2015
rect 4965 2000 4985 2015
rect 5025 2000 5045 2015
rect 5085 2000 5105 2015
rect 5145 2000 5165 2015
rect 2555 1890 2570 1900
rect 2610 1890 2625 1900
rect 2555 1875 2625 1890
rect 2735 1885 2755 1900
rect 2795 1885 2815 1900
rect 2855 1890 2875 1900
rect 2915 1890 2935 1900
rect 2975 1890 2995 1900
rect 3035 1890 3055 1900
rect 2785 1875 2825 1885
rect 2855 1875 3055 1890
rect 3095 1890 3115 1900
rect 3155 1890 3175 1900
rect 3095 1875 3175 1890
rect 3215 1890 3235 1900
rect 3275 1890 3295 1900
rect 3335 1890 3355 1900
rect 3395 1890 3415 1900
rect 3215 1875 3415 1890
rect 3455 1890 3475 1900
rect 3515 1890 3535 1900
rect 3455 1875 3535 1890
rect 3575 1890 3595 1900
rect 3635 1890 3655 1900
rect 3695 1890 3715 1900
rect 3755 1890 3775 1900
rect 3575 1875 3775 1890
rect 3815 1885 3835 1900
rect 3875 1885 3895 1900
rect 4005 1885 4025 1900
rect 4065 1885 4085 1900
rect 4125 1890 4145 1900
rect 4185 1890 4205 1900
rect 4245 1890 4265 1900
rect 4305 1890 4325 1900
rect 3805 1875 3845 1885
rect 2570 1855 2580 1875
rect 2600 1855 2610 1875
rect 2570 1845 2610 1855
rect 2785 1855 2795 1875
rect 2815 1855 2825 1875
rect 2785 1845 2825 1855
rect 2875 1855 2885 1875
rect 2905 1855 2915 1875
rect 2875 1845 2915 1855
rect 3115 1855 3125 1875
rect 3145 1855 3155 1875
rect 3115 1845 3155 1855
rect 3235 1855 3245 1875
rect 3265 1855 3275 1875
rect 3235 1845 3275 1855
rect 3475 1855 3485 1875
rect 3505 1855 3515 1875
rect 3475 1845 3515 1855
rect 3595 1855 3605 1875
rect 3625 1855 3635 1875
rect 3595 1845 3635 1855
rect 3805 1855 3815 1875
rect 3835 1855 3845 1875
rect 3805 1845 3845 1855
rect 4055 1875 4095 1885
rect 4125 1875 4325 1890
rect 4365 1890 4385 1900
rect 4425 1890 4445 1900
rect 4365 1875 4445 1890
rect 4485 1890 4505 1900
rect 4545 1890 4565 1900
rect 4605 1890 4625 1900
rect 4665 1890 4685 1900
rect 4485 1875 4685 1890
rect 4725 1890 4745 1900
rect 4785 1890 4805 1900
rect 4725 1875 4805 1890
rect 4845 1890 4865 1900
rect 4905 1890 4925 1900
rect 4965 1890 4985 1900
rect 5025 1890 5045 1900
rect 4845 1875 5045 1890
rect 5085 1885 5105 1900
rect 5145 1885 5165 1900
rect 5075 1875 5115 1885
rect 4055 1855 4065 1875
rect 4085 1855 4095 1875
rect 4055 1845 4095 1855
rect 4265 1855 4275 1875
rect 4295 1855 4305 1875
rect 4265 1845 4305 1855
rect 4385 1855 4395 1875
rect 4415 1855 4425 1875
rect 4385 1845 4425 1855
rect 4625 1855 4635 1875
rect 4655 1855 4665 1875
rect 4625 1845 4665 1855
rect 4745 1855 4755 1875
rect 4775 1855 4785 1875
rect 4745 1845 4785 1855
rect 4985 1855 4995 1875
rect 5015 1855 5025 1875
rect 4985 1845 5025 1855
rect 5075 1855 5085 1875
rect 5105 1855 5115 1875
rect 5075 1845 5115 1855
rect 3175 1755 3215 1765
rect 3175 1735 3185 1755
rect 3205 1735 3215 1755
rect 3175 1720 3215 1735
rect 4685 1755 4725 1765
rect 4685 1735 4695 1755
rect 4715 1735 4725 1755
rect 4685 1720 4725 1735
rect 3175 1705 3715 1720
rect 3155 1665 3175 1680
rect 3215 1665 3235 1705
rect 3275 1665 3295 1705
rect 3335 1665 3355 1680
rect 3395 1665 3415 1680
rect 3455 1665 3475 1705
rect 3515 1665 3535 1705
rect 3575 1665 3595 1680
rect 3635 1665 3655 1680
rect 3695 1665 3715 1705
rect 4185 1705 4725 1720
rect 4185 1665 4205 1705
rect 4245 1665 4265 1680
rect 4305 1665 4325 1680
rect 4365 1665 4385 1705
rect 4425 1665 4445 1705
rect 4485 1665 4505 1680
rect 4545 1665 4565 1680
rect 4605 1665 4625 1705
rect 4665 1665 4685 1705
rect 4725 1665 4745 1680
rect 3155 1600 3175 1615
rect 3215 1600 3235 1615
rect 3275 1600 3295 1615
rect 3115 1590 3175 1600
rect 3115 1570 3125 1590
rect 3145 1575 3175 1590
rect 3335 1575 3355 1615
rect 3395 1575 3415 1615
rect 3455 1600 3475 1615
rect 3515 1600 3535 1615
rect 3575 1575 3595 1615
rect 3635 1575 3655 1615
rect 3695 1600 3715 1615
rect 4185 1600 4205 1615
rect 3145 1570 3655 1575
rect 3115 1560 3655 1570
rect 4245 1575 4265 1615
rect 4305 1575 4325 1615
rect 4365 1600 4385 1615
rect 4425 1600 4445 1615
rect 4485 1575 4505 1615
rect 4545 1575 4565 1615
rect 4605 1600 4625 1615
rect 4665 1600 4685 1615
rect 4725 1600 4745 1615
rect 4725 1590 4785 1600
rect 4725 1575 4755 1590
rect 4245 1570 4755 1575
rect 4775 1570 4785 1590
rect 4245 1560 4785 1570
rect 2825 1460 3325 1475
rect 3365 1460 3865 1475
rect 4035 1460 4535 1475
rect 4575 1460 5075 1475
rect 2825 1195 3325 1210
rect 3365 1195 3865 1210
rect 4035 1195 4535 1210
rect 4575 1195 5075 1210
rect 2970 1130 3010 1170
rect 3050 1130 3090 1170
rect 3130 1130 3170 1170
rect 3210 1130 3250 1170
rect 3290 1130 3330 1170
rect 3370 1130 3410 1170
rect 3450 1130 3490 1170
rect 3530 1130 3570 1170
rect 3610 1130 3650 1170
rect 3690 1130 3730 1170
rect 3770 1130 3810 1170
rect 3850 1130 3890 1170
rect 4010 1130 4050 1170
rect 4090 1130 4130 1170
rect 4170 1130 4210 1170
rect 4250 1130 4290 1170
rect 4330 1130 4370 1170
rect 4410 1130 4450 1170
rect 4490 1130 4530 1170
rect 4570 1130 4610 1170
rect 4650 1130 4690 1170
rect 4730 1130 4770 1170
rect 4810 1130 4850 1170
rect 4890 1130 4930 1170
rect 2930 1115 3930 1130
rect 3970 1115 4970 1130
rect 2930 1000 3930 1015
rect 3970 1000 4970 1015
rect 3080 910 3130 925
rect 3240 910 3290 925
rect 3330 910 3380 925
rect 3420 910 3470 925
rect 3510 910 3560 925
rect 3600 910 3650 925
rect 3690 910 3740 925
rect 3780 910 3830 925
rect 3870 910 3920 925
rect 3960 910 4010 925
rect 4050 910 4100 925
rect 4140 910 4190 925
rect 4230 910 4280 925
rect 4320 910 4370 925
rect 4410 910 4460 925
rect 4500 910 4550 925
rect 4590 910 4640 925
rect 4680 910 4730 925
rect 4770 910 4820 925
rect 4860 910 4910 925
rect 3080 795 3130 810
rect 3240 795 3290 810
rect 3330 795 3380 810
rect 3420 795 3470 810
rect 3510 795 3560 810
rect 3600 795 3650 810
rect 3690 795 3740 810
rect 3780 795 3830 810
rect 3870 795 3920 810
rect 3960 795 4010 810
rect 4050 795 4100 810
rect 4140 795 4190 810
rect 4230 795 4280 810
rect 4320 795 4370 810
rect 4410 795 4460 810
rect 4500 795 4550 810
rect 4590 795 4640 810
rect 4680 795 4730 810
rect 4770 795 4820 810
rect 4860 795 4910 810
<< polycont >>
rect 2770 2405 2790 2425
rect 2950 2400 2970 2420
rect 3845 2405 3865 2425
rect 5110 2405 5130 2425
rect 2705 2025 2725 2045
rect 3905 2025 3925 2045
rect 3975 2025 3995 2045
rect 5175 2025 5195 2045
rect 2580 1855 2600 1875
rect 2795 1855 2815 1875
rect 2885 1855 2905 1875
rect 3125 1855 3145 1875
rect 3245 1855 3265 1875
rect 3485 1855 3505 1875
rect 3605 1855 3625 1875
rect 3815 1855 3835 1875
rect 4065 1855 4085 1875
rect 4275 1855 4295 1875
rect 4395 1855 4415 1875
rect 4635 1855 4655 1875
rect 4755 1855 4775 1875
rect 4995 1855 5015 1875
rect 5085 1855 5105 1875
rect 3185 1735 3205 1755
rect 4695 1735 4715 1755
rect 3125 1570 3145 1590
rect 4755 1570 4775 1590
<< xpolycontact >>
rect 85 3170 305 3205
rect 905 3170 1125 3205
rect 1290 3165 1510 3200
rect 2110 3165 2330 3200
rect 85 3110 305 3145
rect 905 3110 1125 3145
rect 1290 3105 1510 3140
rect 2110 3105 2330 3140
rect 85 3030 305 3065
rect 910 3030 1130 3065
rect 1290 3045 1510 3080
rect 2110 3045 2330 3080
rect 85 2970 305 3005
rect 910 2970 1130 3005
rect 1290 2985 1510 3020
rect 2110 2985 2330 3020
rect 1290 2925 1510 2960
rect 2110 2925 2330 2960
rect 1290 2865 1510 2900
rect 2110 2865 2330 2900
rect 85 2820 305 2855
rect 355 2820 575 2855
rect 1290 2805 1510 2840
rect 1740 2805 1960 2840
rect 85 2760 305 2795
rect 355 2760 575 2795
<< xpolyres >>
rect 305 3170 905 3205
rect 1510 3165 2110 3200
rect 305 3110 905 3145
rect 1510 3105 2110 3140
rect 305 3030 910 3065
rect 1510 3045 2110 3080
rect 305 2970 910 3005
rect 1510 2985 2110 3020
rect 1510 2925 2110 2960
rect 1510 2865 2110 2900
rect 305 2820 355 2855
rect 1510 2805 1740 2840
rect 305 2760 355 2795
<< locali >>
rect 4445 3465 4475 3495
rect -10 3415 20 3445
rect 945 3415 975 3445
rect 1645 3415 1675 3445
rect 2475 3420 2505 3450
rect 5145 3415 5175 3445
rect -55 3360 -25 3390
rect 2695 3360 2725 3390
rect 1195 3310 1225 3340
rect 2950 3310 2980 3340
rect 3395 3305 3425 3335
rect 5295 3305 5325 3335
rect 1150 3255 1180 3285
rect 5345 3255 5375 3285
rect 2690 3210 2720 3240
rect 40 3200 85 3205
rect 40 3175 50 3200
rect 75 3175 85 3200
rect 40 3170 85 3175
rect 1105 3145 1125 3170
rect 1245 3195 1290 3200
rect 1245 3170 1255 3195
rect 1280 3170 1290 3195
rect 1245 3165 1290 3170
rect 2330 3165 2370 3200
rect 40 3140 85 3145
rect 40 3115 50 3140
rect 75 3115 85 3140
rect 40 3110 85 3115
rect 1245 3135 1290 3140
rect 1245 3110 1255 3135
rect 1280 3110 1290 3135
rect 1245 3105 1290 3110
rect 1150 3070 1180 3100
rect 2295 3080 2330 3105
rect 40 3060 85 3065
rect 40 3035 50 3060
rect 75 3035 85 3060
rect 40 3030 85 3035
rect 1110 3005 1130 3030
rect 40 3000 85 3005
rect 40 2975 50 3000
rect 75 2975 85 3000
rect 40 2970 85 2975
rect 1250 3045 1290 3080
rect 1250 2900 1270 3045
rect 2350 3020 2370 3165
rect 2575 3155 2605 3185
rect 4445 3155 4475 3185
rect 2950 3065 2980 3095
rect 5250 3065 5280 3095
rect 2330 2985 2370 3020
rect 2945 3035 2985 3045
rect 2945 3015 2955 3035
rect 2975 3015 2985 3035
rect 2945 3005 2985 3015
rect 2955 2985 2975 3005
rect 1290 2960 1325 2985
rect 2950 2975 2980 2985
rect 2330 2955 2375 2960
rect 2950 2955 2955 2975
rect 2975 2955 2980 2975
rect 2330 2930 2340 2955
rect 2365 2930 2375 2955
rect 2330 2925 2375 2930
rect 2430 2925 2460 2955
rect 2950 2925 2980 2955
rect 2950 2905 2955 2925
rect 2975 2905 2980 2925
rect 1250 2865 1290 2900
rect 2330 2895 2375 2905
rect 2950 2895 2980 2905
rect 3040 2975 3070 2985
rect 3040 2955 3045 2975
rect 3065 2955 3070 2975
rect 3040 2925 3070 2955
rect 3040 2905 3045 2925
rect 3065 2905 3070 2925
rect 3040 2895 3070 2905
rect 3130 2975 3160 2985
rect 3130 2955 3135 2975
rect 3155 2955 3160 2975
rect 3130 2925 3160 2955
rect 3130 2905 3135 2925
rect 3155 2905 3160 2925
rect 3130 2895 3160 2905
rect 3200 2975 3230 2985
rect 3200 2955 3205 2975
rect 3225 2955 3230 2975
rect 3200 2925 3230 2955
rect 3200 2905 3205 2925
rect 3225 2905 3230 2925
rect 3200 2895 3230 2905
rect 3290 2975 3320 2985
rect 3290 2955 3295 2975
rect 3315 2955 3320 2975
rect 3290 2925 3320 2955
rect 3290 2905 3295 2925
rect 3315 2905 3320 2925
rect 3290 2895 3320 2905
rect 3380 2975 3410 2985
rect 3380 2955 3385 2975
rect 3405 2955 3410 2975
rect 3380 2925 3410 2955
rect 3380 2905 3385 2925
rect 3405 2905 3410 2925
rect 3380 2895 3410 2905
rect 3470 2975 3500 2985
rect 3470 2955 3475 2975
rect 3495 2955 3500 2975
rect 3470 2925 3500 2955
rect 3470 2905 3475 2925
rect 3495 2905 3500 2925
rect 3470 2895 3500 2905
rect 3560 2975 3590 2985
rect 3560 2955 3565 2975
rect 3585 2955 3590 2975
rect 3560 2925 3590 2955
rect 3560 2905 3565 2925
rect 3585 2905 3590 2925
rect 3560 2895 3590 2905
rect 3650 2975 3680 2985
rect 3650 2955 3655 2975
rect 3675 2955 3680 2975
rect 3650 2925 3680 2955
rect 3650 2905 3655 2925
rect 3675 2905 3680 2925
rect 3650 2895 3680 2905
rect 3740 2975 3770 2985
rect 3740 2955 3745 2975
rect 3765 2955 3770 2975
rect 3740 2925 3770 2955
rect 3740 2905 3745 2925
rect 3765 2905 3770 2925
rect 3740 2895 3770 2905
rect 3830 2975 3860 2985
rect 3830 2955 3835 2975
rect 3855 2955 3860 2975
rect 3830 2925 3860 2955
rect 3830 2905 3835 2925
rect 3855 2905 3860 2925
rect 3830 2895 3860 2905
rect 3920 2975 3950 2985
rect 3920 2955 3925 2975
rect 3945 2955 3950 2975
rect 3920 2925 3950 2955
rect 3920 2905 3925 2925
rect 3945 2905 3950 2925
rect 3920 2895 3950 2905
rect 4010 2975 4040 2985
rect 4010 2955 4015 2975
rect 4035 2955 4040 2975
rect 4010 2925 4040 2955
rect 4010 2905 4015 2925
rect 4035 2905 4040 2925
rect 4010 2895 4040 2905
rect 4100 2975 4130 2985
rect 4100 2955 4105 2975
rect 4125 2955 4130 2975
rect 4100 2925 4130 2955
rect 4100 2905 4105 2925
rect 4125 2905 4130 2925
rect 4100 2895 4130 2905
rect 4190 2975 4220 2985
rect 4190 2955 4195 2975
rect 4215 2955 4220 2975
rect 4190 2925 4220 2955
rect 4190 2905 4195 2925
rect 4215 2905 4220 2925
rect 4190 2895 4220 2905
rect 4280 2975 4310 2985
rect 4280 2955 4285 2975
rect 4305 2955 4310 2975
rect 4280 2925 4310 2955
rect 4280 2905 4285 2925
rect 4305 2905 4310 2925
rect 4280 2895 4310 2905
rect 4370 2975 4400 2985
rect 4370 2955 4375 2975
rect 4395 2955 4400 2975
rect 4370 2925 4400 2955
rect 4370 2905 4375 2925
rect 4395 2905 4400 2925
rect 4370 2895 4400 2905
rect 4460 2975 4490 2985
rect 4460 2955 4465 2975
rect 4485 2955 4490 2975
rect 4460 2925 4490 2955
rect 4460 2905 4465 2925
rect 4485 2905 4490 2925
rect 4460 2895 4490 2905
rect 4550 2975 4580 2985
rect 4550 2955 4555 2975
rect 4575 2955 4580 2975
rect 4550 2925 4580 2955
rect 4550 2905 4555 2925
rect 4575 2905 4580 2925
rect 4550 2895 4580 2905
rect 4640 2975 4670 2985
rect 4640 2955 4645 2975
rect 4665 2955 4670 2975
rect 4640 2925 4670 2955
rect 4640 2905 4645 2925
rect 4665 2905 4670 2925
rect 4640 2895 4670 2905
rect 4730 2975 4760 2985
rect 4730 2955 4735 2975
rect 4755 2955 4760 2975
rect 4730 2925 4760 2955
rect 4730 2905 4735 2925
rect 4755 2905 4760 2925
rect 4730 2895 4760 2905
rect 4820 2975 4850 2985
rect 4820 2955 4825 2975
rect 4845 2955 4850 2975
rect 4820 2925 4850 2955
rect 4820 2905 4825 2925
rect 4845 2905 4850 2925
rect 4820 2895 4850 2905
rect 4910 2975 4940 2985
rect 4910 2955 4915 2975
rect 4935 2955 4940 2975
rect 4910 2925 4940 2955
rect 4910 2905 4915 2925
rect 4935 2905 4940 2925
rect 4910 2895 4940 2905
rect 5000 2975 5030 2985
rect 5000 2955 5005 2975
rect 5025 2955 5030 2975
rect 5000 2925 5030 2955
rect 5000 2905 5005 2925
rect 5025 2905 5030 2925
rect 5000 2895 5030 2905
rect 2330 2870 2340 2895
rect 2365 2870 2375 2895
rect 2330 2860 2375 2870
rect -55 2825 -25 2855
rect 40 2850 85 2855
rect 40 2825 50 2850
rect 75 2825 85 2850
rect 40 2820 85 2825
rect 575 2850 620 2855
rect 575 2825 585 2850
rect 610 2825 620 2850
rect 575 2820 620 2825
rect 1195 2820 1225 2850
rect 1245 2835 1290 2840
rect 1245 2810 1255 2835
rect 1280 2810 1290 2835
rect 1245 2805 1290 2810
rect 1960 2835 2005 2840
rect 1960 2810 1970 2835
rect 1995 2810 2005 2835
rect 1960 2805 2005 2810
rect 2330 2800 2370 2840
rect 2940 2795 2980 2805
rect -10 2765 20 2795
rect 40 2790 85 2795
rect 40 2765 50 2790
rect 75 2765 85 2790
rect 40 2760 85 2765
rect 575 2790 620 2795
rect 575 2765 585 2790
rect 610 2765 620 2790
rect 575 2760 620 2765
rect 2570 2755 2610 2795
rect 2940 2775 2950 2795
rect 2970 2775 2980 2795
rect 2940 2765 2980 2775
rect 3120 2795 3160 2805
rect 3120 2775 3130 2795
rect 3150 2775 3160 2795
rect 3120 2765 3160 2775
rect 3300 2795 3340 2805
rect 3300 2775 3310 2795
rect 3330 2775 3340 2795
rect 3300 2765 3340 2775
rect 3480 2795 3520 2805
rect 3480 2775 3490 2795
rect 3510 2775 3520 2795
rect 3480 2765 3520 2775
rect 3660 2795 3700 2805
rect 3660 2775 3670 2795
rect 3690 2775 3700 2795
rect 3660 2765 3700 2775
rect 3840 2795 3880 2805
rect 3840 2775 3850 2795
rect 3870 2775 3880 2795
rect 3840 2765 3880 2775
rect 4020 2795 4060 2805
rect 4020 2775 4030 2795
rect 4050 2775 4060 2795
rect 4020 2765 4060 2775
rect 4200 2795 4240 2805
rect 4200 2775 4210 2795
rect 4230 2775 4240 2795
rect 4200 2765 4240 2775
rect 4380 2795 4420 2805
rect 4380 2775 4390 2795
rect 4410 2775 4420 2795
rect 4380 2765 4420 2775
rect 4560 2795 4600 2805
rect 4560 2775 4570 2795
rect 4590 2775 4600 2795
rect 4560 2765 4600 2775
rect 4740 2795 4780 2805
rect 4740 2775 4750 2795
rect 4770 2775 4780 2795
rect 4740 2765 4780 2775
rect 4920 2795 4960 2805
rect 4920 2775 4930 2795
rect 4950 2775 4960 2795
rect 4920 2765 4960 2775
rect 1250 2715 1280 2745
rect 2150 2710 2190 2750
rect 2950 2745 2970 2765
rect 3130 2745 3150 2765
rect 3310 2745 3330 2765
rect 3490 2745 3510 2765
rect 3670 2745 3690 2765
rect 3850 2745 3870 2765
rect 4030 2745 4050 2765
rect 4210 2745 4230 2765
rect 4390 2745 4410 2765
rect 4570 2745 4590 2765
rect 4750 2745 4770 2765
rect 4930 2745 4950 2765
rect 2765 2735 2795 2745
rect 2765 2715 2770 2735
rect 2790 2715 2795 2735
rect 650 2055 775 2700
rect 1330 2055 1455 2700
rect 2010 2055 2135 2700
rect 2765 2685 2795 2715
rect 2765 2665 2770 2685
rect 2790 2665 2795 2685
rect 2765 2635 2795 2665
rect 2765 2615 2770 2635
rect 2790 2615 2795 2635
rect 2765 2585 2795 2615
rect 2765 2565 2770 2585
rect 2790 2565 2795 2585
rect 2765 2535 2795 2565
rect 2765 2515 2770 2535
rect 2790 2515 2795 2535
rect 2765 2485 2795 2515
rect 2765 2465 2770 2485
rect 2790 2465 2795 2485
rect 2765 2455 2795 2465
rect 2855 2735 2885 2745
rect 2855 2715 2860 2735
rect 2880 2715 2885 2735
rect 2855 2685 2885 2715
rect 2855 2665 2860 2685
rect 2880 2665 2885 2685
rect 2855 2635 2885 2665
rect 2855 2615 2860 2635
rect 2880 2615 2885 2635
rect 2855 2585 2885 2615
rect 2855 2565 2860 2585
rect 2880 2565 2885 2585
rect 2855 2535 2885 2565
rect 2855 2515 2860 2535
rect 2880 2515 2885 2535
rect 2855 2485 2885 2515
rect 2855 2465 2860 2485
rect 2880 2465 2885 2485
rect 2855 2455 2885 2465
rect 2945 2735 2975 2745
rect 2945 2715 2950 2735
rect 2970 2715 2975 2735
rect 2945 2685 2975 2715
rect 2945 2665 2950 2685
rect 2970 2665 2975 2685
rect 2945 2635 2975 2665
rect 2945 2615 2950 2635
rect 2970 2615 2975 2635
rect 2945 2585 2975 2615
rect 2945 2565 2950 2585
rect 2970 2565 2975 2585
rect 2945 2535 2975 2565
rect 2945 2515 2950 2535
rect 2970 2515 2975 2535
rect 2945 2485 2975 2515
rect 2945 2465 2950 2485
rect 2970 2465 2975 2485
rect 2945 2455 2975 2465
rect 3035 2735 3065 2745
rect 3035 2715 3040 2735
rect 3060 2715 3065 2735
rect 3035 2685 3065 2715
rect 3035 2665 3040 2685
rect 3060 2665 3065 2685
rect 3035 2635 3065 2665
rect 3035 2615 3040 2635
rect 3060 2615 3065 2635
rect 3035 2585 3065 2615
rect 3035 2565 3040 2585
rect 3060 2565 3065 2585
rect 3035 2535 3065 2565
rect 3035 2515 3040 2535
rect 3060 2515 3065 2535
rect 3035 2485 3065 2515
rect 3035 2465 3040 2485
rect 3060 2465 3065 2485
rect 3035 2455 3065 2465
rect 3125 2735 3155 2745
rect 3125 2715 3130 2735
rect 3150 2715 3155 2735
rect 3125 2685 3155 2715
rect 3125 2665 3130 2685
rect 3150 2665 3155 2685
rect 3125 2635 3155 2665
rect 3125 2615 3130 2635
rect 3150 2615 3155 2635
rect 3125 2585 3155 2615
rect 3125 2565 3130 2585
rect 3150 2565 3155 2585
rect 3125 2535 3155 2565
rect 3125 2515 3130 2535
rect 3150 2515 3155 2535
rect 3125 2485 3155 2515
rect 3125 2465 3130 2485
rect 3150 2465 3155 2485
rect 3125 2455 3155 2465
rect 3215 2735 3245 2745
rect 3215 2715 3220 2735
rect 3240 2715 3245 2735
rect 3215 2685 3245 2715
rect 3215 2665 3220 2685
rect 3240 2665 3245 2685
rect 3215 2635 3245 2665
rect 3215 2615 3220 2635
rect 3240 2615 3245 2635
rect 3215 2585 3245 2615
rect 3215 2565 3220 2585
rect 3240 2565 3245 2585
rect 3215 2535 3245 2565
rect 3215 2515 3220 2535
rect 3240 2515 3245 2535
rect 3215 2485 3245 2515
rect 3215 2465 3220 2485
rect 3240 2465 3245 2485
rect 3215 2455 3245 2465
rect 3305 2735 3335 2745
rect 3305 2715 3310 2735
rect 3330 2715 3335 2735
rect 3305 2685 3335 2715
rect 3305 2665 3310 2685
rect 3330 2665 3335 2685
rect 3305 2635 3335 2665
rect 3305 2615 3310 2635
rect 3330 2615 3335 2635
rect 3305 2585 3335 2615
rect 3305 2565 3310 2585
rect 3330 2565 3335 2585
rect 3305 2535 3335 2565
rect 3305 2515 3310 2535
rect 3330 2515 3335 2535
rect 3305 2485 3335 2515
rect 3305 2465 3310 2485
rect 3330 2465 3335 2485
rect 3305 2455 3335 2465
rect 3395 2735 3425 2745
rect 3395 2715 3400 2735
rect 3420 2715 3425 2735
rect 3395 2685 3425 2715
rect 3395 2665 3400 2685
rect 3420 2665 3425 2685
rect 3395 2635 3425 2665
rect 3395 2615 3400 2635
rect 3420 2615 3425 2635
rect 3395 2585 3425 2615
rect 3395 2565 3400 2585
rect 3420 2565 3425 2585
rect 3395 2535 3425 2565
rect 3395 2515 3400 2535
rect 3420 2515 3425 2535
rect 3395 2485 3425 2515
rect 3395 2465 3400 2485
rect 3420 2465 3425 2485
rect 3395 2455 3425 2465
rect 3485 2735 3515 2745
rect 3485 2715 3490 2735
rect 3510 2715 3515 2735
rect 3485 2685 3515 2715
rect 3485 2665 3490 2685
rect 3510 2665 3515 2685
rect 3485 2635 3515 2665
rect 3485 2615 3490 2635
rect 3510 2615 3515 2635
rect 3485 2585 3515 2615
rect 3485 2565 3490 2585
rect 3510 2565 3515 2585
rect 3485 2535 3515 2565
rect 3485 2515 3490 2535
rect 3510 2515 3515 2535
rect 3485 2485 3515 2515
rect 3485 2465 3490 2485
rect 3510 2465 3515 2485
rect 3485 2455 3515 2465
rect 3575 2735 3605 2745
rect 3575 2715 3580 2735
rect 3600 2715 3605 2735
rect 3575 2685 3605 2715
rect 3575 2665 3580 2685
rect 3600 2665 3605 2685
rect 3575 2635 3605 2665
rect 3575 2615 3580 2635
rect 3600 2615 3605 2635
rect 3575 2585 3605 2615
rect 3575 2565 3580 2585
rect 3600 2565 3605 2585
rect 3575 2535 3605 2565
rect 3575 2515 3580 2535
rect 3600 2515 3605 2535
rect 3575 2485 3605 2515
rect 3575 2465 3580 2485
rect 3600 2465 3605 2485
rect 3575 2455 3605 2465
rect 3665 2735 3695 2745
rect 3665 2715 3670 2735
rect 3690 2715 3695 2735
rect 3665 2685 3695 2715
rect 3665 2665 3670 2685
rect 3690 2665 3695 2685
rect 3665 2635 3695 2665
rect 3665 2615 3670 2635
rect 3690 2615 3695 2635
rect 3665 2585 3695 2615
rect 3665 2565 3670 2585
rect 3690 2565 3695 2585
rect 3665 2535 3695 2565
rect 3665 2515 3670 2535
rect 3690 2515 3695 2535
rect 3665 2485 3695 2515
rect 3665 2465 3670 2485
rect 3690 2465 3695 2485
rect 3665 2455 3695 2465
rect 3755 2735 3785 2745
rect 3755 2715 3760 2735
rect 3780 2715 3785 2735
rect 3755 2685 3785 2715
rect 3755 2665 3760 2685
rect 3780 2665 3785 2685
rect 3755 2635 3785 2665
rect 3755 2615 3760 2635
rect 3780 2615 3785 2635
rect 3755 2585 3785 2615
rect 3755 2565 3760 2585
rect 3780 2565 3785 2585
rect 3755 2535 3785 2565
rect 3755 2515 3760 2535
rect 3780 2515 3785 2535
rect 3755 2485 3785 2515
rect 3755 2465 3760 2485
rect 3780 2465 3785 2485
rect 3755 2455 3785 2465
rect 3845 2735 3875 2745
rect 3845 2715 3850 2735
rect 3870 2715 3875 2735
rect 3845 2685 3875 2715
rect 3845 2665 3850 2685
rect 3870 2665 3875 2685
rect 3845 2635 3875 2665
rect 3845 2615 3850 2635
rect 3870 2615 3875 2635
rect 3845 2585 3875 2615
rect 3845 2565 3850 2585
rect 3870 2565 3875 2585
rect 3845 2535 3875 2565
rect 3845 2515 3850 2535
rect 3870 2515 3875 2535
rect 3845 2485 3875 2515
rect 3845 2465 3850 2485
rect 3870 2465 3875 2485
rect 3845 2455 3875 2465
rect 3935 2735 3965 2745
rect 3935 2715 3940 2735
rect 3960 2715 3965 2735
rect 3935 2685 3965 2715
rect 3935 2665 3940 2685
rect 3960 2665 3965 2685
rect 3935 2635 3965 2665
rect 3935 2615 3940 2635
rect 3960 2615 3965 2635
rect 3935 2585 3965 2615
rect 3935 2565 3940 2585
rect 3960 2565 3965 2585
rect 3935 2535 3965 2565
rect 3935 2515 3940 2535
rect 3960 2515 3965 2535
rect 3935 2485 3965 2515
rect 3935 2465 3940 2485
rect 3960 2465 3965 2485
rect 3935 2455 3965 2465
rect 4025 2735 4055 2745
rect 4025 2715 4030 2735
rect 4050 2715 4055 2735
rect 4025 2685 4055 2715
rect 4025 2665 4030 2685
rect 4050 2665 4055 2685
rect 4025 2635 4055 2665
rect 4025 2615 4030 2635
rect 4050 2615 4055 2635
rect 4025 2585 4055 2615
rect 4025 2565 4030 2585
rect 4050 2565 4055 2585
rect 4025 2535 4055 2565
rect 4025 2515 4030 2535
rect 4050 2515 4055 2535
rect 4025 2485 4055 2515
rect 4025 2465 4030 2485
rect 4050 2465 4055 2485
rect 4025 2455 4055 2465
rect 4115 2735 4145 2745
rect 4115 2715 4120 2735
rect 4140 2715 4145 2735
rect 4115 2685 4145 2715
rect 4115 2665 4120 2685
rect 4140 2665 4145 2685
rect 4115 2635 4145 2665
rect 4115 2615 4120 2635
rect 4140 2615 4145 2635
rect 4115 2585 4145 2615
rect 4115 2565 4120 2585
rect 4140 2565 4145 2585
rect 4115 2535 4145 2565
rect 4115 2515 4120 2535
rect 4140 2515 4145 2535
rect 4115 2485 4145 2515
rect 4115 2465 4120 2485
rect 4140 2465 4145 2485
rect 4115 2455 4145 2465
rect 4205 2735 4235 2745
rect 4205 2715 4210 2735
rect 4230 2715 4235 2735
rect 4205 2685 4235 2715
rect 4205 2665 4210 2685
rect 4230 2665 4235 2685
rect 4205 2635 4235 2665
rect 4205 2615 4210 2635
rect 4230 2615 4235 2635
rect 4205 2585 4235 2615
rect 4205 2565 4210 2585
rect 4230 2565 4235 2585
rect 4205 2535 4235 2565
rect 4205 2515 4210 2535
rect 4230 2515 4235 2535
rect 4205 2485 4235 2515
rect 4205 2465 4210 2485
rect 4230 2465 4235 2485
rect 4205 2455 4235 2465
rect 4295 2735 4325 2745
rect 4295 2715 4300 2735
rect 4320 2715 4325 2735
rect 4295 2685 4325 2715
rect 4295 2665 4300 2685
rect 4320 2665 4325 2685
rect 4295 2635 4325 2665
rect 4295 2615 4300 2635
rect 4320 2615 4325 2635
rect 4295 2585 4325 2615
rect 4295 2565 4300 2585
rect 4320 2565 4325 2585
rect 4295 2535 4325 2565
rect 4295 2515 4300 2535
rect 4320 2515 4325 2535
rect 4295 2485 4325 2515
rect 4295 2465 4300 2485
rect 4320 2465 4325 2485
rect 4295 2455 4325 2465
rect 4385 2735 4415 2745
rect 4385 2715 4390 2735
rect 4410 2715 4415 2735
rect 4385 2685 4415 2715
rect 4385 2665 4390 2685
rect 4410 2665 4415 2685
rect 4385 2635 4415 2665
rect 4385 2615 4390 2635
rect 4410 2615 4415 2635
rect 4385 2585 4415 2615
rect 4385 2565 4390 2585
rect 4410 2565 4415 2585
rect 4385 2535 4415 2565
rect 4385 2515 4390 2535
rect 4410 2515 4415 2535
rect 4385 2485 4415 2515
rect 4385 2465 4390 2485
rect 4410 2465 4415 2485
rect 4385 2455 4415 2465
rect 4475 2735 4505 2745
rect 4475 2715 4480 2735
rect 4500 2715 4505 2735
rect 4475 2685 4505 2715
rect 4475 2665 4480 2685
rect 4500 2665 4505 2685
rect 4475 2635 4505 2665
rect 4475 2615 4480 2635
rect 4500 2615 4505 2635
rect 4475 2585 4505 2615
rect 4475 2565 4480 2585
rect 4500 2565 4505 2585
rect 4475 2535 4505 2565
rect 4475 2515 4480 2535
rect 4500 2515 4505 2535
rect 4475 2485 4505 2515
rect 4475 2465 4480 2485
rect 4500 2465 4505 2485
rect 4475 2455 4505 2465
rect 4565 2735 4595 2745
rect 4565 2715 4570 2735
rect 4590 2715 4595 2735
rect 4565 2685 4595 2715
rect 4565 2665 4570 2685
rect 4590 2665 4595 2685
rect 4565 2635 4595 2665
rect 4565 2615 4570 2635
rect 4590 2615 4595 2635
rect 4565 2585 4595 2615
rect 4565 2565 4570 2585
rect 4590 2565 4595 2585
rect 4565 2535 4595 2565
rect 4565 2515 4570 2535
rect 4590 2515 4595 2535
rect 4565 2485 4595 2515
rect 4565 2465 4570 2485
rect 4590 2465 4595 2485
rect 4565 2455 4595 2465
rect 4655 2735 4685 2745
rect 4655 2715 4660 2735
rect 4680 2715 4685 2735
rect 4655 2685 4685 2715
rect 4655 2665 4660 2685
rect 4680 2665 4685 2685
rect 4655 2635 4685 2665
rect 4655 2615 4660 2635
rect 4680 2615 4685 2635
rect 4655 2585 4685 2615
rect 4655 2565 4660 2585
rect 4680 2565 4685 2585
rect 4655 2535 4685 2565
rect 4655 2515 4660 2535
rect 4680 2515 4685 2535
rect 4655 2485 4685 2515
rect 4655 2465 4660 2485
rect 4680 2465 4685 2485
rect 4655 2455 4685 2465
rect 4745 2735 4775 2745
rect 4745 2715 4750 2735
rect 4770 2715 4775 2735
rect 4745 2685 4775 2715
rect 4745 2665 4750 2685
rect 4770 2665 4775 2685
rect 4745 2635 4775 2665
rect 4745 2615 4750 2635
rect 4770 2615 4775 2635
rect 4745 2585 4775 2615
rect 4745 2565 4750 2585
rect 4770 2565 4775 2585
rect 4745 2535 4775 2565
rect 4745 2515 4750 2535
rect 4770 2515 4775 2535
rect 4745 2485 4775 2515
rect 4745 2465 4750 2485
rect 4770 2465 4775 2485
rect 4745 2455 4775 2465
rect 4835 2735 4865 2745
rect 4835 2715 4840 2735
rect 4860 2715 4865 2735
rect 4835 2685 4865 2715
rect 4835 2665 4840 2685
rect 4860 2665 4865 2685
rect 4835 2635 4865 2665
rect 4835 2615 4840 2635
rect 4860 2615 4865 2635
rect 4835 2585 4865 2615
rect 4835 2565 4840 2585
rect 4860 2565 4865 2585
rect 4835 2535 4865 2565
rect 4835 2515 4840 2535
rect 4860 2515 4865 2535
rect 4835 2485 4865 2515
rect 4835 2465 4840 2485
rect 4860 2465 4865 2485
rect 4835 2455 4865 2465
rect 4925 2735 4955 2745
rect 4925 2715 4930 2735
rect 4950 2715 4955 2735
rect 4925 2685 4955 2715
rect 4925 2665 4930 2685
rect 4950 2665 4955 2685
rect 4925 2635 4955 2665
rect 4925 2615 4930 2635
rect 4950 2615 4955 2635
rect 4925 2585 4955 2615
rect 4925 2565 4930 2585
rect 4950 2565 4955 2585
rect 4925 2535 4955 2565
rect 4925 2515 4930 2535
rect 4950 2515 4955 2535
rect 4925 2485 4955 2515
rect 4925 2465 4930 2485
rect 4950 2465 4955 2485
rect 4925 2455 4955 2465
rect 5015 2735 5045 2745
rect 5015 2715 5020 2735
rect 5040 2715 5045 2735
rect 5015 2685 5045 2715
rect 5015 2665 5020 2685
rect 5040 2665 5045 2685
rect 5015 2635 5045 2665
rect 5015 2615 5020 2635
rect 5040 2615 5045 2635
rect 5015 2585 5045 2615
rect 5015 2565 5020 2585
rect 5040 2565 5045 2585
rect 5015 2535 5045 2565
rect 5015 2515 5020 2535
rect 5040 2515 5045 2535
rect 5015 2485 5045 2515
rect 5015 2465 5020 2485
rect 5040 2465 5045 2485
rect 5015 2455 5045 2465
rect 5105 2735 5135 2745
rect 5105 2715 5110 2735
rect 5130 2715 5135 2735
rect 5105 2685 5135 2715
rect 5105 2665 5110 2685
rect 5130 2665 5135 2685
rect 5105 2635 5135 2665
rect 5105 2615 5110 2635
rect 5130 2615 5135 2635
rect 5105 2585 5135 2615
rect 5105 2565 5110 2585
rect 5130 2565 5135 2585
rect 5105 2535 5135 2565
rect 5105 2515 5110 2535
rect 5130 2515 5135 2535
rect 5105 2485 5135 2515
rect 5105 2465 5110 2485
rect 5130 2465 5135 2485
rect 5105 2455 5135 2465
rect 2770 2435 2790 2455
rect 2860 2435 2880 2455
rect 3040 2435 3060 2455
rect 2760 2425 2800 2435
rect 2760 2405 2770 2425
rect 2790 2405 2800 2425
rect 2760 2395 2800 2405
rect 2850 2425 2890 2435
rect 2850 2405 2860 2425
rect 2880 2405 2890 2425
rect 2850 2395 2890 2405
rect 2940 2420 2980 2430
rect 2940 2400 2950 2420
rect 2970 2400 2980 2420
rect 2575 2365 2605 2395
rect 2940 2390 2980 2400
rect 3030 2425 3070 2435
rect 3030 2405 3040 2425
rect 3060 2405 3070 2425
rect 3030 2395 3070 2405
rect 3220 2390 3240 2455
rect 3400 2435 3420 2455
rect 3390 2425 3430 2435
rect 3390 2405 3400 2425
rect 3420 2405 3430 2425
rect 3390 2395 3430 2405
rect 3580 2390 3600 2455
rect 3760 2435 3780 2455
rect 3940 2435 3960 2455
rect 4120 2435 4140 2455
rect 3750 2425 3790 2435
rect 3750 2405 3760 2425
rect 3780 2405 3790 2425
rect 3750 2395 3790 2405
rect 3835 2425 3875 2435
rect 3835 2405 3845 2425
rect 3865 2405 3875 2425
rect 3835 2395 3875 2405
rect 3930 2425 3970 2435
rect 3930 2405 3940 2425
rect 3960 2405 3970 2425
rect 3930 2395 3970 2405
rect 4100 2425 4140 2435
rect 4100 2405 4110 2425
rect 4130 2405 4140 2425
rect 4100 2395 4140 2405
rect 4300 2390 4320 2455
rect 4480 2435 4500 2455
rect 4470 2425 4510 2435
rect 4470 2405 4480 2425
rect 4500 2405 4510 2425
rect 4470 2395 4510 2405
rect 4660 2390 4680 2455
rect 4840 2435 4860 2455
rect 5020 2435 5040 2455
rect 5110 2435 5130 2455
rect 4830 2425 4870 2435
rect 4830 2405 4840 2425
rect 4860 2405 4870 2425
rect 4830 2395 4870 2405
rect 5010 2425 5050 2435
rect 5010 2405 5020 2425
rect 5040 2405 5050 2425
rect 5010 2395 5050 2405
rect 5100 2425 5140 2435
rect 5100 2405 5110 2425
rect 5130 2405 5140 2425
rect 5100 2395 5140 2405
rect 3210 2380 3250 2390
rect 3210 2360 3220 2380
rect 3240 2360 3250 2380
rect 3210 2350 3250 2360
rect 3570 2380 3610 2390
rect 3570 2360 3580 2380
rect 3600 2360 3610 2380
rect 3570 2350 3610 2360
rect 4290 2380 4330 2390
rect 4290 2360 4300 2380
rect 4320 2360 4330 2380
rect 4290 2350 4330 2360
rect 4650 2380 4690 2390
rect 4650 2360 4660 2380
rect 4680 2360 4690 2380
rect 4650 2350 4690 2360
rect 2690 2310 2720 2340
rect 3390 2335 3430 2345
rect 3390 2315 3400 2335
rect 3420 2315 3430 2335
rect 3390 2305 3430 2315
rect 4470 2335 4510 2345
rect 4470 2315 4480 2335
rect 4500 2315 4510 2335
rect 4470 2305 4510 2315
rect 5205 2310 5235 2340
rect 2430 2215 2460 2245
rect 3035 2215 3065 2245
rect 2335 2170 2365 2200
rect 2385 2120 2415 2150
rect 3215 2120 3245 2150
rect 4030 2115 4060 2145
rect 5250 2115 5280 2145
rect 2815 2090 2855 2100
rect 2815 2070 2825 2090
rect 2845 2070 2855 2090
rect 2815 2060 2855 2070
rect 2935 2090 2975 2100
rect 2935 2070 2945 2090
rect 2965 2070 2975 2090
rect 2935 2060 2975 2070
rect 3055 2090 3095 2100
rect 3055 2070 3065 2090
rect 3085 2070 3095 2090
rect 3055 2060 3095 2070
rect 3175 2090 3215 2100
rect 3175 2070 3185 2090
rect 3205 2070 3215 2090
rect 3175 2060 3215 2070
rect 3295 2090 3335 2100
rect 3295 2070 3305 2090
rect 3325 2070 3335 2090
rect 3295 2060 3335 2070
rect 3415 2090 3455 2100
rect 3415 2070 3425 2090
rect 3445 2070 3455 2090
rect 3415 2060 3455 2070
rect 3535 2090 3575 2100
rect 3535 2070 3545 2090
rect 3565 2070 3575 2090
rect 3535 2060 3575 2070
rect 3655 2090 3695 2100
rect 3655 2070 3665 2090
rect 3685 2070 3695 2090
rect 3655 2060 3695 2070
rect 3775 2090 3815 2100
rect 3775 2070 3785 2090
rect 3805 2070 3815 2090
rect 3775 2060 3815 2070
rect 4085 2090 4125 2100
rect 4085 2070 4095 2090
rect 4115 2070 4125 2090
rect 4085 2060 4125 2070
rect 4205 2090 4245 2100
rect 4205 2070 4215 2090
rect 4235 2070 4245 2090
rect 4205 2060 4245 2070
rect 4325 2090 4365 2100
rect 4325 2070 4335 2090
rect 4355 2070 4365 2090
rect 4325 2060 4365 2070
rect 4445 2090 4485 2100
rect 4445 2070 4455 2090
rect 4475 2070 4485 2090
rect 4445 2060 4485 2070
rect 4565 2090 4605 2100
rect 4565 2070 4575 2090
rect 4595 2070 4605 2090
rect 4565 2060 4605 2070
rect 4685 2090 4725 2100
rect 4685 2070 4695 2090
rect 4715 2070 4725 2090
rect 4685 2060 4725 2070
rect 4805 2090 4845 2100
rect 4805 2070 4815 2090
rect 4835 2070 4845 2090
rect 4805 2060 4845 2070
rect 4925 2090 4965 2100
rect 4925 2070 4935 2090
rect 4955 2070 4965 2090
rect 4925 2060 4965 2070
rect 5045 2090 5085 2100
rect 5045 2070 5055 2090
rect 5075 2070 5085 2090
rect 5045 2060 5085 2070
rect 125 2015 2135 2055
rect 2570 2045 2610 2055
rect 2570 2025 2580 2045
rect 2600 2025 2610 2045
rect 2570 2015 2610 2025
rect 2695 2045 2735 2055
rect 2695 2025 2705 2045
rect 2725 2025 2735 2045
rect 2695 2015 2735 2025
rect 2755 2045 2795 2055
rect 2755 2025 2765 2045
rect 2785 2025 2795 2045
rect 2755 2015 2795 2025
rect -45 1715 130 1725
rect -45 1695 -35 1715
rect -15 1695 15 1715
rect 35 1695 65 1715
rect 85 1695 130 1715
rect -45 1685 130 1695
rect 650 1375 775 2015
rect 2010 1375 2135 2015
rect 2580 1995 2600 2015
rect 2705 1995 2725 2015
rect 2765 1995 2785 2015
rect 2825 1995 2845 2060
rect 2945 1995 2965 2060
rect 3065 1995 3085 2060
rect 3115 2045 3155 2055
rect 3115 2025 3125 2045
rect 3145 2025 3155 2045
rect 3115 2015 3155 2025
rect 3125 1995 3145 2015
rect 3185 1995 3205 2060
rect 3305 1995 3325 2060
rect 3425 1995 3445 2060
rect 3475 2045 3515 2055
rect 3475 2025 3485 2045
rect 3505 2025 3515 2045
rect 3475 2015 3515 2025
rect 3485 1995 3505 2015
rect 3545 1995 3565 2060
rect 3665 1995 3685 2060
rect 3785 1995 3805 2060
rect 3835 2045 3875 2055
rect 3835 2025 3845 2045
rect 3865 2025 3875 2045
rect 3835 2015 3875 2025
rect 3895 2045 3935 2055
rect 3895 2025 3905 2045
rect 3925 2025 3935 2045
rect 3895 2015 3935 2025
rect 3965 2045 4005 2055
rect 3965 2025 3975 2045
rect 3995 2025 4005 2045
rect 3965 2015 4005 2025
rect 4025 2045 4065 2055
rect 4025 2025 4035 2045
rect 4055 2025 4065 2045
rect 4025 2015 4065 2025
rect 3845 1995 3865 2015
rect 3905 1995 3925 2015
rect 3975 1995 3995 2015
rect 4035 1995 4055 2015
rect 4095 1995 4115 2060
rect 4215 1995 4235 2060
rect 4335 1995 4355 2060
rect 4385 2045 4425 2055
rect 4385 2025 4395 2045
rect 4415 2025 4425 2045
rect 4385 2015 4425 2025
rect 4395 1995 4415 2015
rect 4455 1995 4475 2060
rect 4575 1995 4595 2060
rect 4695 1995 4715 2060
rect 4745 2045 4785 2055
rect 4745 2025 4755 2045
rect 4775 2025 4785 2045
rect 4745 2015 4785 2025
rect 4755 1995 4775 2015
rect 4815 1995 4835 2060
rect 4935 1995 4955 2060
rect 5055 1995 5075 2060
rect 5105 2045 5145 2055
rect 5105 2025 5115 2045
rect 5135 2025 5145 2045
rect 5105 2015 5145 2025
rect 5165 2045 5205 2055
rect 5165 2025 5175 2045
rect 5195 2025 5205 2045
rect 5165 2015 5205 2025
rect 5115 1995 5135 2015
rect 5175 1995 5195 2015
rect 2520 1985 2550 1995
rect 2520 1965 2525 1985
rect 2545 1965 2550 1985
rect 2520 1935 2550 1965
rect 2520 1915 2525 1935
rect 2545 1915 2550 1935
rect 2520 1905 2550 1915
rect 2575 1985 2605 1995
rect 2575 1965 2580 1985
rect 2600 1965 2605 1985
rect 2575 1935 2605 1965
rect 2575 1915 2580 1935
rect 2600 1915 2605 1935
rect 2575 1905 2605 1915
rect 2630 1985 2660 1995
rect 2630 1965 2635 1985
rect 2655 1965 2660 1985
rect 2630 1935 2660 1965
rect 2630 1915 2635 1935
rect 2655 1915 2660 1935
rect 2630 1905 2660 1915
rect 2700 1985 2730 1995
rect 2700 1965 2705 1985
rect 2725 1965 2730 1985
rect 2700 1935 2730 1965
rect 2700 1915 2705 1935
rect 2725 1915 2730 1935
rect 2700 1905 2730 1915
rect 2760 1985 2790 1995
rect 2760 1965 2765 1985
rect 2785 1965 2790 1985
rect 2760 1935 2790 1965
rect 2760 1915 2765 1935
rect 2785 1915 2790 1935
rect 2760 1905 2790 1915
rect 2820 1985 2850 1995
rect 2820 1965 2825 1985
rect 2845 1965 2850 1985
rect 2820 1935 2850 1965
rect 2820 1915 2825 1935
rect 2845 1915 2850 1935
rect 2820 1905 2850 1915
rect 2880 1985 2910 1995
rect 2880 1965 2885 1985
rect 2905 1965 2910 1985
rect 2880 1935 2910 1965
rect 2880 1915 2885 1935
rect 2905 1915 2910 1935
rect 2880 1905 2910 1915
rect 2940 1985 2970 1995
rect 2940 1965 2945 1985
rect 2965 1965 2970 1985
rect 2940 1935 2970 1965
rect 2940 1915 2945 1935
rect 2965 1915 2970 1935
rect 2940 1905 2970 1915
rect 3000 1985 3030 1995
rect 3000 1965 3005 1985
rect 3025 1965 3030 1985
rect 3000 1935 3030 1965
rect 3000 1915 3005 1935
rect 3025 1915 3030 1935
rect 3000 1905 3030 1915
rect 3060 1985 3090 1995
rect 3060 1965 3065 1985
rect 3085 1965 3090 1985
rect 3060 1935 3090 1965
rect 3060 1915 3065 1935
rect 3085 1915 3090 1935
rect 3060 1905 3090 1915
rect 3120 1985 3150 1995
rect 3120 1965 3125 1985
rect 3145 1965 3150 1985
rect 3120 1935 3150 1965
rect 3120 1915 3125 1935
rect 3145 1915 3150 1935
rect 3120 1905 3150 1915
rect 3180 1985 3210 1995
rect 3180 1965 3185 1985
rect 3205 1965 3210 1985
rect 3180 1935 3210 1965
rect 3180 1915 3185 1935
rect 3205 1915 3210 1935
rect 3180 1905 3210 1915
rect 3240 1985 3270 1995
rect 3240 1965 3245 1985
rect 3265 1965 3270 1985
rect 3240 1935 3270 1965
rect 3240 1915 3245 1935
rect 3265 1915 3270 1935
rect 3240 1905 3270 1915
rect 3300 1985 3330 1995
rect 3300 1965 3305 1985
rect 3325 1965 3330 1985
rect 3300 1935 3330 1965
rect 3300 1915 3305 1935
rect 3325 1915 3330 1935
rect 3300 1905 3330 1915
rect 3360 1985 3390 1995
rect 3360 1965 3365 1985
rect 3385 1965 3390 1985
rect 3360 1935 3390 1965
rect 3360 1915 3365 1935
rect 3385 1915 3390 1935
rect 3360 1905 3390 1915
rect 3420 1985 3450 1995
rect 3420 1965 3425 1985
rect 3445 1965 3450 1985
rect 3420 1935 3450 1965
rect 3420 1915 3425 1935
rect 3445 1915 3450 1935
rect 3420 1905 3450 1915
rect 3480 1985 3510 1995
rect 3480 1965 3485 1985
rect 3505 1965 3510 1985
rect 3480 1935 3510 1965
rect 3480 1915 3485 1935
rect 3505 1915 3510 1935
rect 3480 1905 3510 1915
rect 3540 1985 3570 1995
rect 3540 1965 3545 1985
rect 3565 1965 3570 1985
rect 3540 1935 3570 1965
rect 3540 1915 3545 1935
rect 3565 1915 3570 1935
rect 3540 1905 3570 1915
rect 3600 1985 3630 1995
rect 3600 1965 3605 1985
rect 3625 1965 3630 1985
rect 3600 1935 3630 1965
rect 3600 1915 3605 1935
rect 3625 1915 3630 1935
rect 3600 1905 3630 1915
rect 3660 1985 3690 1995
rect 3660 1965 3665 1985
rect 3685 1965 3690 1985
rect 3660 1935 3690 1965
rect 3660 1915 3665 1935
rect 3685 1915 3690 1935
rect 3660 1905 3690 1915
rect 3720 1985 3750 1995
rect 3720 1965 3725 1985
rect 3745 1965 3750 1985
rect 3720 1935 3750 1965
rect 3720 1915 3725 1935
rect 3745 1915 3750 1935
rect 3720 1905 3750 1915
rect 3780 1985 3810 1995
rect 3780 1965 3785 1985
rect 3805 1965 3810 1985
rect 3780 1935 3810 1965
rect 3780 1915 3785 1935
rect 3805 1915 3810 1935
rect 3780 1905 3810 1915
rect 3840 1985 3870 1995
rect 3840 1965 3845 1985
rect 3865 1965 3870 1985
rect 3840 1935 3870 1965
rect 3840 1915 3845 1935
rect 3865 1915 3870 1935
rect 3840 1905 3870 1915
rect 3900 1985 3930 1995
rect 3900 1965 3905 1985
rect 3925 1965 3930 1985
rect 3900 1935 3930 1965
rect 3900 1915 3905 1935
rect 3925 1915 3930 1935
rect 3900 1905 3930 1915
rect 3970 1985 4000 1995
rect 3970 1965 3975 1985
rect 3995 1965 4000 1985
rect 3970 1935 4000 1965
rect 3970 1915 3975 1935
rect 3995 1915 4000 1935
rect 3970 1905 4000 1915
rect 4030 1985 4060 1995
rect 4030 1965 4035 1985
rect 4055 1965 4060 1985
rect 4030 1935 4060 1965
rect 4030 1915 4035 1935
rect 4055 1915 4060 1935
rect 4030 1905 4060 1915
rect 4090 1985 4120 1995
rect 4090 1965 4095 1985
rect 4115 1965 4120 1985
rect 4090 1935 4120 1965
rect 4090 1915 4095 1935
rect 4115 1915 4120 1935
rect 4090 1905 4120 1915
rect 4150 1985 4180 1995
rect 4150 1965 4155 1985
rect 4175 1965 4180 1985
rect 4150 1935 4180 1965
rect 4150 1915 4155 1935
rect 4175 1915 4180 1935
rect 4150 1905 4180 1915
rect 4210 1985 4240 1995
rect 4210 1965 4215 1985
rect 4235 1965 4240 1985
rect 4210 1935 4240 1965
rect 4210 1915 4215 1935
rect 4235 1915 4240 1935
rect 4210 1905 4240 1915
rect 4270 1985 4300 1995
rect 4270 1965 4275 1985
rect 4295 1965 4300 1985
rect 4270 1935 4300 1965
rect 4270 1915 4275 1935
rect 4295 1915 4300 1935
rect 4270 1905 4300 1915
rect 4330 1985 4360 1995
rect 4330 1965 4335 1985
rect 4355 1965 4360 1985
rect 4330 1935 4360 1965
rect 4330 1915 4335 1935
rect 4355 1915 4360 1935
rect 4330 1905 4360 1915
rect 4390 1985 4420 1995
rect 4390 1965 4395 1985
rect 4415 1965 4420 1985
rect 4390 1935 4420 1965
rect 4390 1915 4395 1935
rect 4415 1915 4420 1935
rect 4390 1905 4420 1915
rect 4450 1985 4480 1995
rect 4450 1965 4455 1985
rect 4475 1965 4480 1985
rect 4450 1935 4480 1965
rect 4450 1915 4455 1935
rect 4475 1915 4480 1935
rect 4450 1905 4480 1915
rect 4510 1985 4540 1995
rect 4510 1965 4515 1985
rect 4535 1965 4540 1985
rect 4510 1935 4540 1965
rect 4510 1915 4515 1935
rect 4535 1915 4540 1935
rect 4510 1905 4540 1915
rect 4570 1985 4600 1995
rect 4570 1965 4575 1985
rect 4595 1965 4600 1985
rect 4570 1935 4600 1965
rect 4570 1915 4575 1935
rect 4595 1915 4600 1935
rect 4570 1905 4600 1915
rect 4630 1985 4660 1995
rect 4630 1965 4635 1985
rect 4655 1965 4660 1985
rect 4630 1935 4660 1965
rect 4630 1915 4635 1935
rect 4655 1915 4660 1935
rect 4630 1905 4660 1915
rect 4690 1985 4720 1995
rect 4690 1965 4695 1985
rect 4715 1965 4720 1985
rect 4690 1935 4720 1965
rect 4690 1915 4695 1935
rect 4715 1915 4720 1935
rect 4690 1905 4720 1915
rect 4750 1985 4780 1995
rect 4750 1965 4755 1985
rect 4775 1965 4780 1985
rect 4750 1935 4780 1965
rect 4750 1915 4755 1935
rect 4775 1915 4780 1935
rect 4750 1905 4780 1915
rect 4810 1985 4840 1995
rect 4810 1965 4815 1985
rect 4835 1965 4840 1985
rect 4810 1935 4840 1965
rect 4810 1915 4815 1935
rect 4835 1915 4840 1935
rect 4810 1905 4840 1915
rect 4870 1985 4900 1995
rect 4870 1965 4875 1985
rect 4895 1965 4900 1985
rect 4870 1935 4900 1965
rect 4870 1915 4875 1935
rect 4895 1915 4900 1935
rect 4870 1905 4900 1915
rect 4930 1985 4960 1995
rect 4930 1965 4935 1985
rect 4955 1965 4960 1985
rect 4930 1935 4960 1965
rect 4930 1915 4935 1935
rect 4955 1915 4960 1935
rect 4930 1905 4960 1915
rect 4990 1985 5020 1995
rect 4990 1965 4995 1985
rect 5015 1965 5020 1985
rect 4990 1935 5020 1965
rect 4990 1915 4995 1935
rect 5015 1915 5020 1935
rect 4990 1905 5020 1915
rect 5050 1985 5080 1995
rect 5050 1965 5055 1985
rect 5075 1965 5080 1985
rect 5050 1935 5080 1965
rect 5050 1915 5055 1935
rect 5075 1915 5080 1935
rect 5050 1905 5080 1915
rect 5110 1985 5140 1995
rect 5110 1965 5115 1985
rect 5135 1965 5140 1985
rect 5110 1935 5140 1965
rect 5110 1915 5115 1935
rect 5135 1915 5140 1935
rect 5110 1905 5140 1915
rect 5170 1985 5200 1995
rect 5170 1965 5175 1985
rect 5195 1965 5200 1985
rect 5170 1935 5200 1965
rect 5170 1915 5175 1935
rect 5195 1915 5200 1935
rect 5170 1905 5200 1915
rect 2525 1885 2545 1905
rect 2635 1885 2655 1905
rect 2885 1885 2905 1905
rect 3005 1885 3025 1905
rect 3245 1885 3265 1905
rect 3365 1885 3385 1905
rect 3605 1885 3625 1905
rect 3725 1885 3745 1905
rect 4155 1885 4175 1905
rect 4275 1885 4295 1905
rect 4515 1885 4535 1905
rect 4635 1885 4655 1905
rect 4875 1885 4895 1905
rect 4995 1885 5015 1905
rect 2515 1875 2550 1885
rect 2515 1855 2525 1875
rect 2545 1855 2550 1875
rect 2515 1845 2550 1855
rect 2570 1875 2610 1885
rect 2570 1855 2580 1875
rect 2600 1855 2610 1875
rect 2570 1845 2610 1855
rect 2630 1875 2665 1885
rect 2630 1855 2635 1875
rect 2655 1855 2665 1875
rect 2630 1845 2665 1855
rect 2785 1875 2825 1885
rect 2785 1855 2795 1875
rect 2815 1855 2825 1875
rect 2785 1845 2825 1855
rect 2875 1875 2915 1885
rect 2875 1855 2885 1875
rect 2905 1855 2915 1875
rect 2875 1845 2915 1855
rect 2995 1875 3035 1885
rect 2995 1855 3005 1875
rect 3025 1855 3035 1875
rect 2995 1845 3035 1855
rect 3115 1875 3155 1885
rect 3115 1855 3125 1875
rect 3145 1855 3155 1875
rect 3115 1845 3155 1855
rect 3235 1875 3275 1885
rect 3235 1855 3245 1875
rect 3265 1855 3275 1875
rect 3235 1845 3275 1855
rect 3355 1875 3395 1885
rect 3355 1855 3365 1875
rect 3385 1855 3395 1875
rect 3355 1845 3395 1855
rect 3475 1875 3515 1885
rect 3475 1855 3485 1875
rect 3505 1855 3515 1875
rect 3475 1845 3515 1855
rect 3595 1875 3635 1885
rect 3595 1855 3605 1875
rect 3625 1855 3635 1875
rect 3595 1845 3635 1855
rect 3715 1875 3755 1885
rect 3715 1855 3725 1875
rect 3745 1855 3755 1875
rect 3715 1845 3755 1855
rect 3805 1875 3845 1885
rect 3805 1855 3815 1875
rect 3835 1855 3845 1875
rect 3805 1845 3845 1855
rect 4055 1875 4095 1885
rect 4055 1855 4065 1875
rect 4085 1855 4095 1875
rect 4055 1845 4095 1855
rect 4145 1875 4185 1885
rect 4145 1855 4155 1875
rect 4175 1855 4185 1875
rect 4145 1845 4185 1855
rect 4265 1875 4305 1885
rect 4265 1855 4275 1875
rect 4295 1855 4305 1875
rect 4265 1845 4305 1855
rect 4385 1875 4425 1885
rect 4385 1855 4395 1875
rect 4415 1855 4425 1875
rect 4385 1845 4425 1855
rect 4505 1875 4545 1885
rect 4505 1855 4515 1875
rect 4535 1855 4545 1875
rect 4505 1845 4545 1855
rect 4625 1875 4665 1885
rect 4625 1855 4635 1875
rect 4655 1855 4665 1875
rect 4625 1845 4665 1855
rect 4745 1875 4785 1885
rect 4745 1855 4755 1875
rect 4775 1855 4785 1875
rect 4745 1845 4785 1855
rect 4865 1875 4905 1885
rect 4865 1855 4875 1875
rect 4895 1855 4905 1875
rect 4865 1845 4905 1855
rect 4985 1875 5025 1885
rect 4985 1855 4995 1875
rect 5015 1855 5025 1875
rect 4985 1845 5025 1855
rect 5075 1875 5115 1885
rect 5075 1855 5085 1875
rect 5105 1855 5115 1875
rect 5075 1845 5115 1855
rect 2475 1790 2505 1820
rect 2785 1785 2825 1825
rect 2995 1815 3035 1825
rect 2995 1795 3005 1815
rect 3025 1795 3035 1815
rect 2995 1785 3035 1795
rect 3115 1785 3155 1825
rect 3355 1815 3395 1825
rect 3355 1795 3365 1815
rect 3385 1795 3395 1815
rect 3355 1785 3395 1795
rect 3475 1785 3515 1825
rect 3715 1815 3755 1825
rect 3715 1795 3725 1815
rect 3745 1795 3755 1815
rect 3715 1785 3755 1795
rect 3805 1785 3845 1825
rect 4055 1785 4095 1825
rect 4145 1815 4185 1825
rect 4145 1795 4155 1815
rect 4175 1795 4185 1815
rect 4145 1785 4185 1795
rect 4385 1785 4425 1825
rect 4505 1815 4545 1825
rect 4505 1795 4515 1815
rect 4535 1795 4545 1815
rect 4505 1785 4545 1795
rect 4745 1785 4785 1825
rect 4865 1815 4905 1825
rect 4865 1795 4875 1815
rect 4895 1795 4905 1815
rect 4865 1785 4905 1795
rect 5075 1785 5115 1825
rect 5295 1790 5325 1820
rect 2430 1730 2460 1760
rect 2520 1730 2550 1760
rect 2630 1730 2660 1760
rect 3175 1755 3215 1765
rect 3175 1735 3185 1755
rect 3205 1735 3215 1755
rect 3175 1725 3215 1735
rect 3235 1755 3275 1765
rect 3235 1735 3245 1755
rect 3265 1735 3275 1755
rect 3235 1725 3275 1735
rect 3475 1755 3515 1765
rect 3475 1735 3485 1755
rect 3505 1735 3515 1755
rect 3475 1725 3515 1735
rect 3715 1755 3755 1765
rect 3715 1735 3725 1755
rect 3745 1735 3755 1755
rect 3715 1725 3755 1735
rect 4145 1755 4185 1765
rect 4145 1735 4155 1755
rect 4175 1735 4185 1755
rect 4145 1725 4185 1735
rect 4385 1755 4425 1765
rect 4385 1735 4395 1755
rect 4415 1735 4425 1755
rect 4385 1725 4425 1735
rect 4625 1755 4665 1765
rect 4625 1735 4635 1755
rect 4655 1735 4665 1755
rect 4625 1725 4665 1735
rect 4685 1755 4725 1765
rect 4685 1735 4695 1755
rect 4715 1735 4725 1755
rect 4685 1725 4725 1735
rect 5205 1730 5235 1760
rect 3115 1710 3155 1720
rect 2155 1680 2185 1710
rect 3115 1690 3125 1710
rect 3145 1690 3155 1710
rect 3115 1680 3155 1690
rect 2385 1635 2415 1665
rect 2575 1635 2605 1665
rect 3125 1660 3145 1680
rect 3245 1660 3265 1725
rect 3355 1710 3395 1720
rect 3355 1690 3365 1710
rect 3385 1690 3395 1710
rect 3355 1680 3395 1690
rect 3365 1660 3385 1680
rect 3485 1660 3505 1725
rect 3595 1710 3635 1720
rect 3595 1690 3605 1710
rect 3625 1690 3635 1710
rect 3595 1680 3635 1690
rect 3605 1660 3625 1680
rect 3725 1660 3745 1725
rect 4155 1660 4175 1725
rect 4265 1710 4305 1720
rect 4265 1690 4275 1710
rect 4295 1690 4305 1710
rect 4265 1680 4305 1690
rect 4275 1660 4295 1680
rect 4395 1660 4415 1725
rect 4505 1710 4545 1720
rect 4505 1690 4515 1710
rect 4535 1690 4545 1710
rect 4505 1680 4545 1690
rect 4515 1660 4535 1680
rect 4635 1660 4655 1725
rect 4745 1710 4785 1720
rect 4745 1690 4755 1710
rect 4775 1690 4785 1710
rect 4745 1680 4785 1690
rect 4755 1660 4775 1680
rect 3120 1650 3150 1660
rect 3120 1630 3125 1650
rect 3145 1630 3150 1650
rect 3120 1620 3150 1630
rect 3180 1650 3210 1660
rect 3180 1630 3185 1650
rect 3205 1630 3210 1650
rect 3180 1620 3210 1630
rect 3240 1650 3270 1660
rect 3240 1630 3245 1650
rect 3265 1630 3270 1650
rect 3240 1620 3270 1630
rect 3300 1650 3330 1660
rect 3300 1630 3305 1650
rect 3325 1630 3330 1650
rect 3300 1620 3330 1630
rect 3360 1650 3390 1660
rect 3360 1630 3365 1650
rect 3385 1630 3390 1650
rect 3360 1620 3390 1630
rect 3420 1650 3450 1660
rect 3420 1630 3425 1650
rect 3445 1630 3450 1650
rect 3420 1620 3450 1630
rect 3480 1650 3510 1660
rect 3480 1630 3485 1650
rect 3505 1630 3510 1650
rect 3480 1620 3510 1630
rect 3540 1650 3570 1660
rect 3540 1630 3545 1650
rect 3565 1630 3570 1650
rect 3540 1620 3570 1630
rect 3600 1650 3630 1660
rect 3600 1630 3605 1650
rect 3625 1630 3630 1650
rect 3600 1620 3630 1630
rect 3660 1650 3690 1660
rect 3660 1630 3665 1650
rect 3685 1630 3690 1650
rect 3660 1620 3690 1630
rect 3720 1650 3750 1660
rect 3720 1630 3725 1650
rect 3745 1630 3750 1650
rect 3720 1620 3750 1630
rect 4150 1650 4180 1660
rect 4150 1630 4155 1650
rect 4175 1630 4180 1650
rect 4150 1620 4180 1630
rect 4210 1650 4240 1660
rect 4210 1630 4215 1650
rect 4235 1630 4240 1650
rect 4210 1620 4240 1630
rect 4270 1650 4300 1660
rect 4270 1630 4275 1650
rect 4295 1630 4300 1650
rect 4270 1620 4300 1630
rect 4330 1650 4360 1660
rect 4330 1630 4335 1650
rect 4355 1630 4360 1650
rect 4330 1620 4360 1630
rect 4390 1650 4420 1660
rect 4390 1630 4395 1650
rect 4415 1630 4420 1650
rect 4390 1620 4420 1630
rect 4450 1650 4480 1660
rect 4450 1630 4455 1650
rect 4475 1630 4480 1650
rect 4450 1620 4480 1630
rect 4510 1650 4540 1660
rect 4510 1630 4515 1650
rect 4535 1630 4540 1650
rect 4510 1620 4540 1630
rect 4570 1650 4600 1660
rect 4570 1630 4575 1650
rect 4595 1630 4600 1650
rect 4570 1620 4600 1630
rect 4630 1650 4660 1660
rect 4630 1630 4635 1650
rect 4655 1630 4660 1650
rect 4630 1620 4660 1630
rect 4690 1650 4720 1660
rect 4690 1630 4695 1650
rect 4715 1630 4720 1650
rect 4690 1620 4720 1630
rect 4750 1650 4780 1660
rect 4750 1630 4755 1650
rect 4775 1630 4780 1650
rect 4750 1620 4780 1630
rect 2335 1565 2365 1595
rect 3115 1590 3155 1600
rect 3115 1570 3125 1590
rect 3145 1570 3155 1590
rect 3115 1560 3155 1570
rect 3185 1550 3205 1620
rect 3305 1550 3325 1620
rect 3425 1550 3445 1620
rect 3545 1550 3565 1620
rect 3665 1550 3685 1620
rect 4215 1550 4235 1620
rect 4335 1550 4355 1620
rect 4455 1550 4475 1620
rect 4575 1550 4595 1620
rect 4695 1550 4715 1620
rect 4745 1590 4785 1600
rect 4745 1570 4755 1590
rect 4775 1570 4785 1590
rect 4745 1560 4785 1570
rect 5345 1565 5375 1595
rect 3175 1540 3215 1550
rect 3175 1520 3185 1540
rect 3205 1520 3215 1540
rect 3175 1510 3215 1520
rect 3295 1540 3335 1550
rect 3295 1520 3305 1540
rect 3325 1520 3335 1540
rect 3295 1510 3335 1520
rect 3415 1540 3455 1550
rect 3415 1520 3425 1540
rect 3445 1520 3455 1540
rect 3415 1510 3455 1520
rect 3535 1540 3575 1550
rect 3535 1520 3545 1540
rect 3565 1520 3575 1540
rect 3535 1510 3575 1520
rect 3655 1540 3695 1550
rect 3655 1520 3665 1540
rect 3685 1520 3695 1540
rect 3655 1510 3695 1520
rect 4205 1540 4245 1550
rect 4205 1520 4215 1540
rect 4235 1520 4245 1540
rect 4205 1510 4245 1520
rect 4325 1540 4365 1550
rect 4325 1520 4335 1540
rect 4355 1520 4365 1540
rect 4325 1510 4365 1520
rect 4445 1540 4485 1550
rect 4445 1520 4455 1540
rect 4475 1520 4485 1540
rect 4445 1510 4485 1520
rect 4565 1540 4605 1550
rect 4565 1520 4575 1540
rect 4595 1520 4605 1540
rect 4565 1510 4605 1520
rect 4685 1540 4725 1550
rect 4685 1520 4695 1540
rect 4715 1520 4725 1540
rect 4685 1510 4725 1520
rect 2785 1485 2825 1495
rect 2785 1465 2795 1485
rect 2815 1465 2825 1485
rect 2785 1455 2825 1465
rect 3865 1485 3905 1495
rect 3865 1465 3875 1485
rect 3895 1465 3905 1485
rect 3865 1455 3905 1465
rect 3995 1485 4035 1495
rect 3995 1465 4005 1485
rect 4025 1465 4035 1485
rect 3995 1455 4035 1465
rect 5075 1485 5115 1495
rect 5075 1465 5085 1485
rect 5105 1465 5115 1485
rect 5075 1455 5115 1465
rect 125 1335 2135 1375
rect 650 690 775 1335
rect 1330 690 1455 1335
rect 2010 695 2135 1335
rect 2790 1445 2820 1455
rect 2790 1425 2795 1445
rect 2815 1425 2820 1445
rect 2790 1395 2820 1425
rect 2790 1375 2795 1395
rect 2815 1375 2820 1395
rect 2790 1345 2820 1375
rect 2790 1325 2795 1345
rect 2815 1325 2820 1345
rect 2790 1295 2820 1325
rect 2790 1275 2795 1295
rect 2815 1275 2820 1295
rect 2790 1245 2820 1275
rect 2790 1225 2795 1245
rect 2815 1225 2820 1245
rect 2790 1215 2820 1225
rect 3330 1445 3360 1455
rect 3330 1425 3335 1445
rect 3355 1425 3360 1445
rect 3330 1395 3360 1425
rect 3330 1375 3335 1395
rect 3355 1375 3360 1395
rect 3330 1345 3360 1375
rect 3330 1325 3335 1345
rect 3355 1325 3360 1345
rect 3330 1295 3360 1325
rect 3330 1275 3335 1295
rect 3355 1275 3360 1295
rect 3330 1245 3360 1275
rect 3330 1225 3335 1245
rect 3355 1225 3360 1245
rect 3330 1215 3360 1225
rect 3870 1445 3900 1455
rect 3870 1425 3875 1445
rect 3895 1425 3900 1445
rect 3870 1395 3900 1425
rect 3870 1375 3875 1395
rect 3895 1375 3900 1395
rect 3870 1345 3900 1375
rect 3870 1325 3875 1345
rect 3895 1325 3900 1345
rect 3870 1295 3900 1325
rect 3870 1275 3875 1295
rect 3895 1275 3900 1295
rect 3870 1245 3900 1275
rect 3870 1225 3875 1245
rect 3895 1225 3900 1245
rect 3870 1215 3900 1225
rect 4000 1445 4030 1455
rect 4000 1425 4005 1445
rect 4025 1425 4030 1445
rect 4000 1395 4030 1425
rect 4000 1375 4005 1395
rect 4025 1375 4030 1395
rect 4000 1345 4030 1375
rect 4000 1325 4005 1345
rect 4025 1325 4030 1345
rect 4000 1295 4030 1325
rect 4000 1275 4005 1295
rect 4025 1275 4030 1295
rect 4000 1245 4030 1275
rect 4000 1225 4005 1245
rect 4025 1225 4030 1245
rect 4000 1215 4030 1225
rect 4540 1445 4570 1455
rect 4540 1425 4545 1445
rect 4565 1425 4570 1445
rect 4540 1395 4570 1425
rect 4540 1375 4545 1395
rect 4565 1375 4570 1395
rect 4540 1345 4570 1375
rect 4540 1325 4545 1345
rect 4565 1325 4570 1345
rect 4540 1295 4570 1325
rect 4540 1275 4545 1295
rect 4565 1275 4570 1295
rect 4540 1245 4570 1275
rect 4540 1225 4545 1245
rect 4565 1225 4570 1245
rect 4540 1215 4570 1225
rect 5080 1445 5110 1455
rect 5080 1425 5085 1445
rect 5105 1425 5110 1445
rect 5080 1395 5110 1425
rect 5080 1375 5085 1395
rect 5105 1375 5110 1395
rect 5080 1345 5110 1375
rect 5080 1325 5085 1345
rect 5105 1325 5110 1345
rect 5080 1295 5110 1325
rect 5080 1275 5085 1295
rect 5105 1275 5110 1295
rect 5080 1245 5110 1275
rect 5080 1225 5085 1245
rect 5105 1225 5110 1245
rect 5080 1215 5110 1225
rect 2890 1160 2930 1170
rect 2890 1140 2900 1160
rect 2920 1140 2930 1160
rect 2890 1130 2930 1140
rect 2970 1160 3010 1170
rect 2970 1140 2980 1160
rect 3000 1140 3010 1160
rect 2970 1130 3010 1140
rect 3050 1160 3090 1170
rect 3050 1140 3060 1160
rect 3080 1140 3090 1160
rect 3050 1130 3090 1140
rect 3130 1160 3170 1170
rect 3130 1140 3140 1160
rect 3160 1140 3170 1160
rect 3130 1130 3170 1140
rect 3210 1160 3250 1170
rect 3210 1140 3220 1160
rect 3240 1140 3250 1160
rect 3210 1130 3250 1140
rect 3290 1160 3330 1170
rect 3290 1140 3300 1160
rect 3320 1140 3330 1160
rect 3290 1130 3330 1140
rect 3370 1160 3410 1170
rect 3370 1140 3380 1160
rect 3400 1140 3410 1160
rect 3370 1130 3410 1140
rect 3450 1160 3490 1170
rect 3450 1140 3460 1160
rect 3480 1140 3490 1160
rect 3450 1130 3490 1140
rect 3530 1160 3570 1170
rect 3530 1140 3540 1160
rect 3560 1140 3570 1160
rect 3530 1130 3570 1140
rect 3610 1160 3650 1170
rect 3610 1140 3620 1160
rect 3640 1140 3650 1160
rect 3610 1130 3650 1140
rect 3690 1160 3730 1170
rect 3690 1140 3700 1160
rect 3720 1140 3730 1160
rect 3690 1130 3730 1140
rect 3770 1160 3810 1170
rect 3770 1140 3780 1160
rect 3800 1140 3810 1160
rect 3770 1130 3810 1140
rect 3850 1160 3890 1170
rect 3850 1140 3860 1160
rect 3880 1140 3890 1160
rect 3850 1130 3890 1140
rect 3930 1160 3970 1170
rect 3930 1140 3940 1160
rect 3960 1140 3970 1160
rect 3930 1130 3970 1140
rect 4010 1160 4050 1170
rect 4010 1140 4020 1160
rect 4040 1140 4050 1160
rect 4010 1130 4050 1140
rect 4090 1160 4130 1170
rect 4090 1140 4100 1160
rect 4120 1140 4130 1160
rect 4090 1130 4130 1140
rect 4170 1160 4210 1170
rect 4170 1140 4180 1160
rect 4200 1140 4210 1160
rect 4170 1130 4210 1140
rect 4250 1160 4290 1170
rect 4250 1140 4260 1160
rect 4280 1140 4290 1160
rect 4250 1130 4290 1140
rect 4330 1160 4370 1170
rect 4330 1140 4340 1160
rect 4360 1140 4370 1160
rect 4330 1130 4370 1140
rect 4410 1160 4450 1170
rect 4410 1140 4420 1160
rect 4440 1140 4450 1160
rect 4410 1130 4450 1140
rect 4490 1160 4530 1170
rect 4490 1140 4500 1160
rect 4520 1140 4530 1160
rect 4490 1130 4530 1140
rect 4570 1160 4610 1170
rect 4570 1140 4580 1160
rect 4600 1140 4610 1160
rect 4570 1130 4610 1140
rect 4650 1160 4690 1170
rect 4650 1140 4660 1160
rect 4680 1140 4690 1160
rect 4650 1130 4690 1140
rect 4730 1160 4770 1170
rect 4730 1140 4740 1160
rect 4760 1140 4770 1160
rect 4730 1130 4770 1140
rect 4810 1160 4850 1170
rect 4810 1140 4820 1160
rect 4840 1140 4850 1160
rect 4810 1130 4850 1140
rect 4890 1160 4930 1170
rect 4890 1140 4900 1160
rect 4920 1140 4930 1160
rect 4890 1130 4930 1140
rect 2900 1110 2920 1130
rect 3940 1110 3960 1130
rect 2895 1100 2925 1110
rect 2895 1085 2900 1100
rect 2880 1080 2900 1085
rect 2920 1080 2925 1100
rect 2575 1050 2605 1080
rect 2855 1075 2925 1080
rect 2855 1055 2860 1075
rect 2880 1055 2925 1075
rect 2855 1050 2925 1055
rect 2880 1045 2900 1050
rect 2895 1030 2900 1045
rect 2920 1030 2925 1050
rect 2430 1000 2460 1030
rect 2895 1020 2925 1030
rect 3935 1100 3965 1110
rect 3935 1080 3940 1100
rect 3960 1080 3965 1100
rect 3935 1050 3965 1080
rect 3935 1030 3940 1050
rect 3960 1030 3965 1050
rect 3935 1020 3965 1030
rect 4975 1100 5005 1110
rect 4975 1080 4980 1100
rect 5000 1080 5005 1100
rect 4975 1050 5005 1080
rect 4975 1030 4980 1050
rect 5000 1030 5005 1050
rect 4975 1020 5005 1030
rect 3045 895 3075 905
rect 3045 875 3050 895
rect 3070 875 3075 895
rect 3045 845 3075 875
rect 3045 825 3050 845
rect 3070 825 3075 845
rect 3045 815 3075 825
rect 3135 895 3165 905
rect 3135 875 3140 895
rect 3160 875 3165 895
rect 3135 845 3165 875
rect 3135 825 3140 845
rect 3160 825 3165 845
rect 3135 815 3165 825
rect 3205 895 3235 905
rect 3205 875 3210 895
rect 3230 875 3235 895
rect 3205 845 3235 875
rect 3205 825 3210 845
rect 3230 825 3235 845
rect 3205 815 3235 825
rect 3295 895 3325 905
rect 3295 875 3300 895
rect 3320 875 3325 895
rect 3295 845 3325 875
rect 3295 825 3300 845
rect 3320 825 3325 845
rect 3295 815 3325 825
rect 3385 895 3415 905
rect 3385 875 3390 895
rect 3410 875 3415 895
rect 3385 845 3415 875
rect 3385 825 3390 845
rect 3410 825 3415 845
rect 3385 815 3415 825
rect 3475 895 3505 905
rect 3475 875 3480 895
rect 3500 875 3505 895
rect 3475 845 3505 875
rect 3475 825 3480 845
rect 3500 825 3505 845
rect 3475 815 3505 825
rect 3565 895 3595 905
rect 3565 875 3570 895
rect 3590 875 3595 895
rect 3565 845 3595 875
rect 3565 825 3570 845
rect 3590 825 3595 845
rect 3565 815 3595 825
rect 3655 895 3685 905
rect 3655 875 3660 895
rect 3680 875 3685 895
rect 3655 845 3685 875
rect 3655 825 3660 845
rect 3680 825 3685 845
rect 3655 815 3685 825
rect 3745 895 3775 905
rect 3745 875 3750 895
rect 3770 875 3775 895
rect 3745 845 3775 875
rect 3745 825 3750 845
rect 3770 825 3775 845
rect 3745 815 3775 825
rect 3835 895 3865 905
rect 3835 875 3840 895
rect 3860 875 3865 895
rect 3835 845 3865 875
rect 3835 825 3840 845
rect 3860 825 3865 845
rect 3835 815 3865 825
rect 3925 895 3955 905
rect 3925 875 3930 895
rect 3950 875 3955 895
rect 3925 845 3955 875
rect 3925 825 3930 845
rect 3950 825 3955 845
rect 3925 815 3955 825
rect 4015 895 4045 905
rect 4015 875 4020 895
rect 4040 875 4045 895
rect 4015 845 4045 875
rect 4015 825 4020 845
rect 4040 825 4045 845
rect 4015 815 4045 825
rect 4105 895 4135 905
rect 4105 875 4110 895
rect 4130 875 4135 895
rect 4105 845 4135 875
rect 4105 825 4110 845
rect 4130 825 4135 845
rect 4105 815 4135 825
rect 4195 895 4225 905
rect 4195 875 4200 895
rect 4220 875 4225 895
rect 4195 845 4225 875
rect 4195 825 4200 845
rect 4220 825 4225 845
rect 4195 815 4225 825
rect 4285 895 4315 905
rect 4285 875 4290 895
rect 4310 875 4315 895
rect 4285 845 4315 875
rect 4285 825 4290 845
rect 4310 825 4315 845
rect 4285 815 4315 825
rect 4375 895 4405 905
rect 4375 875 4380 895
rect 4400 875 4405 895
rect 4375 845 4405 875
rect 4375 825 4380 845
rect 4400 825 4405 845
rect 4375 815 4405 825
rect 4465 895 4495 905
rect 4465 875 4470 895
rect 4490 875 4495 895
rect 4465 845 4495 875
rect 4465 825 4470 845
rect 4490 825 4495 845
rect 4465 815 4495 825
rect 4555 895 4585 905
rect 4555 875 4560 895
rect 4580 875 4585 895
rect 4555 845 4585 875
rect 4555 825 4560 845
rect 4580 825 4585 845
rect 4555 815 4585 825
rect 4645 895 4675 905
rect 4645 875 4650 895
rect 4670 875 4675 895
rect 4645 845 4675 875
rect 4645 825 4650 845
rect 4670 825 4675 845
rect 4645 815 4675 825
rect 4735 895 4765 905
rect 4735 875 4740 895
rect 4760 875 4765 895
rect 4735 845 4765 875
rect 4735 825 4740 845
rect 4760 825 4765 845
rect 4735 815 4765 825
rect 4825 895 4855 905
rect 4825 875 4830 895
rect 4850 875 4855 895
rect 4825 845 4855 875
rect 4825 825 4830 845
rect 4850 825 4855 845
rect 4825 815 4855 825
rect 4915 895 4945 905
rect 4915 875 4920 895
rect 4940 875 4945 895
rect 4915 845 4945 875
rect 4915 825 4920 845
rect 4940 825 4945 845
rect 4915 815 4945 825
<< viali >>
rect 50 3175 75 3200
rect 1255 3170 1280 3195
rect 50 3115 75 3140
rect 1255 3110 1280 3135
rect 50 3035 75 3060
rect 50 2975 75 3000
rect 2955 3015 2975 3035
rect 2340 2930 2365 2955
rect 2340 2870 2365 2895
rect 50 2825 75 2850
rect 585 2825 610 2850
rect 1255 2810 1280 2835
rect 1970 2810 1995 2835
rect 50 2765 75 2790
rect 585 2765 610 2790
rect 2950 2775 2970 2795
rect 3130 2775 3150 2795
rect 3310 2775 3330 2795
rect 3490 2775 3510 2795
rect 3670 2775 3690 2795
rect 3850 2775 3870 2795
rect 4030 2775 4050 2795
rect 4210 2775 4230 2795
rect 4390 2775 4410 2795
rect 4570 2775 4590 2795
rect 4750 2775 4770 2795
rect 4930 2775 4950 2795
rect 2860 2405 2880 2425
rect 2950 2400 2970 2420
rect 3040 2405 3060 2425
rect 3400 2405 3420 2425
rect 3760 2405 3780 2425
rect 3845 2405 3865 2425
rect 3940 2405 3960 2425
rect 4110 2405 4130 2425
rect 4480 2405 4500 2425
rect 4840 2405 4860 2425
rect 5020 2405 5040 2425
rect 3220 2360 3240 2380
rect 3580 2360 3600 2380
rect 4300 2360 4320 2380
rect 4660 2360 4680 2380
rect 3400 2315 3420 2335
rect 4480 2315 4500 2335
rect 2825 2070 2845 2090
rect 2945 2070 2965 2090
rect 3065 2070 3085 2090
rect 3185 2070 3205 2090
rect 3305 2070 3325 2090
rect 3425 2070 3445 2090
rect 3545 2070 3565 2090
rect 3665 2070 3685 2090
rect 3785 2070 3805 2090
rect 4095 2070 4115 2090
rect 4215 2070 4235 2090
rect 4335 2070 4355 2090
rect 4455 2070 4475 2090
rect 4575 2070 4595 2090
rect 4695 2070 4715 2090
rect 4815 2070 4835 2090
rect 4935 2070 4955 2090
rect 5055 2070 5075 2090
rect 2580 2025 2600 2045
rect 2765 2025 2785 2045
rect -35 1695 -15 1715
rect 3125 2025 3145 2045
rect 3485 2025 3505 2045
rect 3845 2025 3865 2045
rect 4035 2025 4055 2045
rect 4395 2025 4415 2045
rect 4755 2025 4775 2045
rect 5115 2025 5135 2045
rect 2525 1855 2545 1875
rect 2580 1855 2600 1875
rect 2635 1855 2655 1875
rect 2795 1855 2815 1875
rect 2885 1855 2905 1875
rect 3005 1855 3025 1875
rect 3125 1855 3145 1875
rect 3245 1855 3265 1875
rect 3365 1855 3385 1875
rect 3485 1855 3505 1875
rect 3605 1855 3625 1875
rect 3725 1855 3745 1875
rect 3815 1855 3835 1875
rect 4065 1855 4085 1875
rect 4155 1855 4175 1875
rect 4275 1855 4295 1875
rect 4395 1855 4415 1875
rect 4515 1855 4535 1875
rect 4635 1855 4655 1875
rect 4755 1855 4775 1875
rect 4875 1855 4895 1875
rect 4995 1855 5015 1875
rect 5085 1855 5105 1875
rect 3005 1795 3025 1815
rect 3365 1795 3385 1815
rect 3725 1795 3745 1815
rect 4155 1795 4175 1815
rect 4515 1795 4535 1815
rect 4875 1795 4895 1815
rect 3185 1735 3205 1755
rect 3245 1735 3265 1755
rect 3485 1735 3505 1755
rect 3725 1735 3745 1755
rect 4155 1735 4175 1755
rect 4395 1735 4415 1755
rect 4635 1735 4655 1755
rect 4695 1735 4715 1755
rect 3125 1690 3145 1710
rect 3365 1690 3385 1710
rect 3605 1690 3625 1710
rect 4275 1690 4295 1710
rect 4515 1690 4535 1710
rect 4755 1690 4775 1710
rect 3125 1570 3145 1590
rect 4755 1570 4775 1590
rect 3185 1520 3205 1540
rect 3305 1520 3325 1540
rect 3425 1520 3445 1540
rect 3545 1520 3565 1540
rect 3665 1520 3685 1540
rect 4215 1520 4235 1540
rect 4335 1520 4355 1540
rect 4455 1520 4475 1540
rect 4575 1520 4595 1540
rect 4695 1520 4715 1540
rect 2795 1465 2815 1485
rect 3875 1465 3895 1485
rect 4005 1465 4025 1485
rect 5085 1465 5105 1485
rect 2900 1140 2920 1160
rect 2980 1140 3000 1160
rect 3060 1140 3080 1160
rect 3140 1140 3160 1160
rect 3220 1140 3240 1160
rect 3300 1140 3320 1160
rect 3380 1140 3400 1160
rect 3460 1140 3480 1160
rect 3540 1140 3560 1160
rect 3620 1140 3640 1160
rect 3700 1140 3720 1160
rect 3780 1140 3800 1160
rect 3860 1140 3880 1160
rect 3940 1140 3960 1160
rect 4020 1140 4040 1160
rect 4100 1140 4120 1160
rect 4180 1140 4200 1160
rect 4260 1140 4280 1160
rect 4340 1140 4360 1160
rect 4420 1140 4440 1160
rect 4500 1140 4520 1160
rect 4580 1140 4600 1160
rect 4660 1140 4680 1160
rect 4740 1140 4760 1160
rect 4820 1140 4840 1160
rect 4900 1140 4920 1160
rect 2860 1055 2880 1075
<< metal1 >>
rect 3730 4880 3750 5195
rect 4440 3495 4480 3500
rect 4440 3465 4445 3495
rect 4475 3465 4480 3495
rect 4440 3460 4480 3465
rect -15 3445 25 3450
rect -15 3415 -10 3445
rect 20 3415 25 3445
rect -15 3410 25 3415
rect 940 3445 980 3450
rect 940 3415 945 3445
rect 975 3415 980 3445
rect 940 3410 980 3415
rect 1635 3445 1685 3455
rect 1635 3415 1645 3445
rect 1675 3415 1685 3445
rect 2470 3450 2510 3455
rect 2470 3420 2475 3450
rect 2505 3420 2510 3450
rect 2470 3415 2510 3420
rect -60 3390 -20 3395
rect -60 3360 -55 3390
rect -25 3360 -20 3390
rect -60 3355 -20 3360
rect -50 2860 -30 3355
rect -60 2855 -20 2860
rect -60 2825 -55 2855
rect -25 2825 -20 2855
rect -60 2820 -20 2825
rect -5 2800 15 3410
rect 1635 3405 1685 3415
rect 1190 3340 1230 3345
rect 1190 3310 1195 3340
rect 1225 3310 1230 3340
rect 1190 3305 1230 3310
rect 1145 3285 1185 3290
rect 1145 3255 1150 3285
rect 1180 3255 1185 3285
rect 1145 3250 1185 3255
rect 40 3170 45 3205
rect 80 3170 85 3205
rect 40 3110 45 3145
rect 80 3110 85 3145
rect 1155 3105 1175 3250
rect 1145 3100 1185 3105
rect 1145 3070 1150 3100
rect 1180 3070 1185 3100
rect 1145 3065 1185 3070
rect 40 3030 45 3065
rect 80 3030 85 3065
rect 40 2970 45 3005
rect 80 2970 85 3005
rect 1200 2855 1220 3305
rect 1245 3165 1250 3200
rect 1285 3165 1290 3200
rect 1245 3105 1250 3140
rect 1285 3105 1290 3140
rect 2330 2925 2335 2960
rect 2370 2925 2375 2960
rect 2425 2955 2465 2960
rect 2425 2925 2430 2955
rect 2460 2925 2465 2955
rect 2425 2920 2465 2925
rect 2330 2900 2375 2905
rect 2330 2865 2335 2900
rect 2370 2865 2375 2900
rect 2330 2860 2375 2865
rect 40 2820 45 2855
rect 80 2820 85 2855
rect 575 2820 580 2855
rect 615 2820 620 2855
rect 1190 2850 1230 2855
rect 1190 2820 1195 2850
rect 1225 2820 1230 2850
rect 2340 2840 2360 2860
rect 1190 2815 1230 2820
rect 1245 2805 1250 2840
rect 1285 2805 1290 2840
rect 1960 2805 1965 2840
rect 2000 2805 2005 2840
rect 2330 2835 2370 2840
rect 2330 2805 2335 2835
rect 2365 2805 2370 2835
rect -15 2795 25 2800
rect -15 2765 -10 2795
rect 20 2765 25 2795
rect -15 2760 25 2765
rect 40 2760 45 2795
rect 80 2760 85 2795
rect 575 2760 580 2795
rect 615 2760 620 2795
rect 1255 2750 1275 2805
rect 2330 2800 2370 2805
rect 1245 2745 1285 2750
rect 1245 2715 1250 2745
rect 1280 2715 1285 2745
rect 1245 2710 1285 2715
rect 2150 2745 2190 2750
rect 2150 2715 2155 2745
rect 2185 2715 2190 2745
rect 2150 2710 2190 2715
rect 275 2200 1985 2550
rect -110 1720 -70 1725
rect -110 1690 -105 1720
rect -75 1715 -70 1720
rect -45 1720 -5 1725
rect -45 1715 -40 1720
rect -75 1695 -40 1715
rect -75 1690 -70 1695
rect -110 1685 -70 1690
rect -45 1690 -40 1695
rect -10 1690 -5 1720
rect -45 1685 -5 1690
rect 275 1190 625 2200
rect 955 1710 1305 1870
rect 955 1680 1270 1710
rect 1300 1680 1305 1710
rect 955 1520 1305 1680
rect 1635 1190 1985 2200
rect 2160 1715 2180 2710
rect 2340 2205 2360 2800
rect 2435 2250 2455 2920
rect 2425 2245 2465 2250
rect 2425 2215 2430 2245
rect 2460 2215 2465 2245
rect 2425 2210 2465 2215
rect 2330 2200 2370 2205
rect 2330 2170 2335 2200
rect 2365 2170 2370 2200
rect 2330 2165 2370 2170
rect 2150 1710 2190 1715
rect 2150 1680 2155 1710
rect 2185 1680 2190 1710
rect 2150 1675 2190 1680
rect 2340 1600 2360 2165
rect 2380 2150 2420 2155
rect 2380 2120 2385 2150
rect 2415 2120 2420 2150
rect 2380 2115 2420 2120
rect 2390 1670 2410 2115
rect 2435 1765 2455 2210
rect 2480 1825 2500 3415
rect 2690 3390 2730 3395
rect 2690 3360 2695 3390
rect 2725 3360 2730 3390
rect 2690 3355 2730 3360
rect 2945 3340 2985 3345
rect 2945 3310 2950 3340
rect 2980 3310 2985 3340
rect 2945 3305 2985 3310
rect 3385 3335 3435 3345
rect 3385 3305 3395 3335
rect 3425 3305 3435 3335
rect 2685 3240 2725 3245
rect 2685 3210 2690 3240
rect 2720 3210 2725 3240
rect 2685 3205 2725 3210
rect 2570 3185 2610 3190
rect 2570 3155 2575 3185
rect 2605 3155 2610 3185
rect 2570 3150 2610 3155
rect 2580 2795 2600 3150
rect 2570 2790 2610 2795
rect 2570 2760 2575 2790
rect 2605 2760 2610 2790
rect 2570 2755 2610 2760
rect 2580 2400 2600 2755
rect 2570 2395 2610 2400
rect 2570 2365 2575 2395
rect 2605 2365 2610 2395
rect 2570 2360 2610 2365
rect 2580 2055 2600 2360
rect 2695 2345 2715 3205
rect 2955 3100 2975 3305
rect 3385 3295 3435 3305
rect 4450 3190 4470 3460
rect 5135 3445 5185 3455
rect 5135 3415 5145 3445
rect 5175 3415 5185 3445
rect 5135 3405 5185 3415
rect 5290 3335 5330 3340
rect 5290 3305 5295 3335
rect 5325 3305 5330 3335
rect 5290 3300 5330 3305
rect 4440 3185 4480 3190
rect 4440 3155 4445 3185
rect 4475 3155 4480 3185
rect 4440 3150 4480 3155
rect 2945 3095 2985 3100
rect 2945 3065 2950 3095
rect 2980 3065 2985 3095
rect 2945 3060 2985 3065
rect 5245 3095 5285 3100
rect 5245 3065 5250 3095
rect 5280 3065 5285 3095
rect 5245 3060 5285 3065
rect 2955 3045 2975 3060
rect 2945 3035 2985 3045
rect 2945 3015 2955 3035
rect 2975 3015 2985 3035
rect 2945 3005 2985 3015
rect 2940 2800 2980 2805
rect 2940 2770 2945 2800
rect 2975 2770 2980 2800
rect 2940 2765 2980 2770
rect 3120 2800 3160 2805
rect 3120 2770 3125 2800
rect 3155 2770 3160 2800
rect 3120 2765 3160 2770
rect 3300 2800 3340 2805
rect 3300 2770 3305 2800
rect 3335 2770 3340 2800
rect 3300 2765 3340 2770
rect 3480 2800 3520 2805
rect 3480 2770 3485 2800
rect 3515 2770 3520 2800
rect 3480 2765 3520 2770
rect 3660 2800 3700 2805
rect 3660 2770 3665 2800
rect 3695 2770 3700 2800
rect 3660 2765 3700 2770
rect 3840 2800 3880 2805
rect 3840 2770 3845 2800
rect 3875 2770 3880 2800
rect 3840 2765 3880 2770
rect 4020 2800 4060 2805
rect 4020 2770 4025 2800
rect 4055 2770 4060 2800
rect 4020 2765 4060 2770
rect 4200 2800 4240 2805
rect 4200 2770 4205 2800
rect 4235 2770 4240 2800
rect 4200 2765 4240 2770
rect 4380 2800 4420 2805
rect 4380 2770 4385 2800
rect 4415 2770 4420 2800
rect 4380 2765 4420 2770
rect 4560 2800 4600 2805
rect 4560 2770 4565 2800
rect 4595 2770 4600 2800
rect 4560 2765 4600 2770
rect 4740 2800 4780 2805
rect 4740 2770 4745 2800
rect 4775 2770 4780 2800
rect 4740 2765 4780 2770
rect 4920 2800 4960 2805
rect 4920 2770 4925 2800
rect 4955 2770 4960 2800
rect 4920 2765 4960 2770
rect 2850 2425 2890 2435
rect 3030 2430 3070 2435
rect 2850 2405 2860 2425
rect 2880 2405 2890 2425
rect 2850 2395 2890 2405
rect 2940 2425 2980 2430
rect 2940 2395 2945 2425
rect 2975 2395 2980 2425
rect 3030 2400 3035 2430
rect 3065 2400 3070 2430
rect 3030 2395 3070 2400
rect 3390 2425 3430 2435
rect 3390 2405 3400 2425
rect 3420 2405 3430 2425
rect 3390 2395 3430 2405
rect 3750 2430 3790 2435
rect 3750 2400 3755 2430
rect 3785 2400 3790 2430
rect 3750 2395 3790 2400
rect 3835 2425 3875 2435
rect 3835 2405 3845 2425
rect 3865 2405 3875 2425
rect 3835 2395 3875 2405
rect 3930 2425 3970 2435
rect 3930 2405 3940 2425
rect 3960 2405 3970 2425
rect 3930 2395 3970 2405
rect 4100 2430 4140 2435
rect 4100 2400 4105 2430
rect 4135 2400 4140 2430
rect 4100 2395 4140 2400
rect 4470 2425 4510 2435
rect 4470 2405 4480 2425
rect 4500 2405 4510 2425
rect 4470 2395 4510 2405
rect 4830 2430 4870 2435
rect 4830 2400 4835 2430
rect 4865 2400 4870 2430
rect 4830 2395 4870 2400
rect 5010 2425 5050 2435
rect 5010 2405 5020 2425
rect 5040 2405 5050 2425
rect 5010 2395 5050 2405
rect 2685 2340 2725 2345
rect 2685 2310 2690 2340
rect 2720 2310 2725 2340
rect 2685 2305 2725 2310
rect 2860 2205 2880 2395
rect 2940 2390 2980 2395
rect 3040 2250 3060 2395
rect 3210 2385 3250 2390
rect 3210 2355 3215 2385
rect 3245 2355 3250 2385
rect 3210 2350 3250 2355
rect 3030 2245 3070 2250
rect 3030 2215 3035 2245
rect 3065 2215 3070 2245
rect 3030 2210 3070 2215
rect 2850 2200 2890 2205
rect 2850 2170 2855 2200
rect 2885 2170 2890 2200
rect 2850 2165 2890 2170
rect 3220 2155 3240 2350
rect 3400 2345 3420 2395
rect 3570 2385 3610 2390
rect 3570 2355 3575 2385
rect 3605 2355 3610 2385
rect 3570 2350 3610 2355
rect 3390 2340 3430 2345
rect 3390 2310 3395 2340
rect 3425 2310 3430 2340
rect 3390 2305 3430 2310
rect 3210 2150 3250 2155
rect 3210 2120 3215 2150
rect 3245 2120 3250 2150
rect 3210 2115 3250 2120
rect 2815 2095 2855 2100
rect 2815 2065 2820 2095
rect 2850 2065 2855 2095
rect 2815 2060 2855 2065
rect 2935 2095 2975 2100
rect 2935 2065 2940 2095
rect 2970 2065 2975 2095
rect 2935 2060 2975 2065
rect 3055 2095 3095 2100
rect 3055 2065 3060 2095
rect 3090 2065 3095 2095
rect 3055 2060 3095 2065
rect 3175 2095 3215 2100
rect 3175 2065 3180 2095
rect 3210 2065 3215 2095
rect 3175 2060 3215 2065
rect 3295 2095 3335 2100
rect 3295 2065 3300 2095
rect 3330 2065 3335 2095
rect 3295 2060 3335 2065
rect 3415 2095 3455 2100
rect 3415 2065 3420 2095
rect 3450 2065 3455 2095
rect 3415 2060 3455 2065
rect 3535 2095 3575 2100
rect 3535 2065 3540 2095
rect 3570 2065 3575 2095
rect 3535 2060 3575 2065
rect 3655 2095 3695 2100
rect 3655 2065 3660 2095
rect 3690 2065 3695 2095
rect 3655 2060 3695 2065
rect 3775 2095 3815 2100
rect 3775 2065 3780 2095
rect 3810 2065 3815 2095
rect 3775 2060 3815 2065
rect 3845 2055 3865 2395
rect 3940 2205 3960 2395
rect 4290 2385 4330 2390
rect 4290 2355 4295 2385
rect 4325 2355 4330 2385
rect 4290 2350 4330 2355
rect 4480 2345 4500 2395
rect 4650 2385 4690 2390
rect 4650 2355 4655 2385
rect 4685 2355 4690 2385
rect 4650 2350 4690 2355
rect 4470 2340 4510 2345
rect 4470 2310 4475 2340
rect 4505 2310 4510 2340
rect 4470 2305 4510 2310
rect 5020 2205 5040 2395
rect 5200 2340 5240 2345
rect 5200 2310 5205 2340
rect 5235 2310 5240 2340
rect 5200 2305 5240 2310
rect 3930 2200 3970 2205
rect 3930 2170 3935 2200
rect 3965 2170 3970 2200
rect 3930 2165 3970 2170
rect 5010 2200 5050 2205
rect 5010 2170 5015 2200
rect 5045 2170 5050 2200
rect 5010 2165 5050 2170
rect 4025 2145 4065 2150
rect 4025 2115 4030 2145
rect 4060 2115 4065 2145
rect 4025 2110 4065 2115
rect 4035 2055 4055 2110
rect 4085 2095 4125 2100
rect 4085 2065 4090 2095
rect 4120 2065 4125 2095
rect 4085 2060 4125 2065
rect 4205 2095 4245 2100
rect 4205 2065 4210 2095
rect 4240 2065 4245 2095
rect 4205 2060 4245 2065
rect 4325 2095 4365 2100
rect 4325 2065 4330 2095
rect 4360 2065 4365 2095
rect 4325 2060 4365 2065
rect 4445 2095 4485 2100
rect 4445 2065 4450 2095
rect 4480 2065 4485 2095
rect 4445 2060 4485 2065
rect 4565 2095 4605 2100
rect 4565 2065 4570 2095
rect 4600 2065 4605 2095
rect 4565 2060 4605 2065
rect 4685 2095 4725 2100
rect 4685 2065 4690 2095
rect 4720 2065 4725 2095
rect 4685 2060 4725 2065
rect 4805 2095 4845 2100
rect 4805 2065 4810 2095
rect 4840 2065 4845 2095
rect 4805 2060 4845 2065
rect 4925 2095 4965 2100
rect 4925 2065 4930 2095
rect 4960 2065 4965 2095
rect 4925 2060 4965 2065
rect 5045 2095 5085 2100
rect 5045 2065 5050 2095
rect 5080 2065 5085 2095
rect 5045 2060 5085 2065
rect 2570 2050 2610 2055
rect 2570 2020 2575 2050
rect 2605 2020 2610 2050
rect 2570 2015 2610 2020
rect 2755 2050 2795 2055
rect 2755 2020 2760 2050
rect 2790 2020 2795 2050
rect 2755 2015 2795 2020
rect 3115 2050 3155 2055
rect 3115 2020 3120 2050
rect 3150 2020 3155 2050
rect 3115 2015 3155 2020
rect 3475 2050 3515 2055
rect 3475 2020 3480 2050
rect 3510 2020 3515 2050
rect 3475 2015 3515 2020
rect 3835 2050 3895 2055
rect 3835 2020 3840 2050
rect 3870 2020 3895 2050
rect 3835 2015 3895 2020
rect 2515 1875 2550 1885
rect 2515 1855 2525 1875
rect 2545 1855 2550 1875
rect 2515 1845 2550 1855
rect 2570 1875 2610 1885
rect 2570 1855 2580 1875
rect 2600 1855 2610 1875
rect 2570 1845 2610 1855
rect 2630 1875 2665 1885
rect 2630 1855 2635 1875
rect 2655 1855 2665 1875
rect 2630 1845 2665 1855
rect 2785 1875 2825 1885
rect 2785 1855 2795 1875
rect 2815 1855 2825 1875
rect 2785 1845 2825 1855
rect 2875 1880 2915 1885
rect 2875 1850 2880 1880
rect 2910 1850 2915 1880
rect 2875 1845 2915 1850
rect 2995 1875 3035 1885
rect 2995 1855 3005 1875
rect 3025 1855 3035 1875
rect 2995 1845 3035 1855
rect 3115 1875 3155 1885
rect 3115 1855 3125 1875
rect 3145 1855 3155 1875
rect 3115 1845 3155 1855
rect 3235 1880 3275 1885
rect 3235 1850 3240 1880
rect 3270 1850 3275 1880
rect 3235 1845 3275 1850
rect 3355 1875 3395 1885
rect 3355 1855 3365 1875
rect 3385 1855 3395 1875
rect 3355 1845 3395 1855
rect 3475 1875 3515 1885
rect 3475 1855 3485 1875
rect 3505 1855 3515 1875
rect 3475 1845 3515 1855
rect 3595 1880 3635 1885
rect 3595 1850 3600 1880
rect 3630 1850 3635 1880
rect 3595 1845 3635 1850
rect 3715 1875 3755 1885
rect 3715 1855 3725 1875
rect 3745 1855 3755 1875
rect 3715 1845 3755 1855
rect 3805 1875 3845 1885
rect 3805 1855 3815 1875
rect 3835 1855 3845 1875
rect 3805 1845 3845 1855
rect 2470 1820 2510 1825
rect 2470 1790 2475 1820
rect 2505 1790 2510 1820
rect 2470 1785 2510 1790
rect 2525 1765 2545 1845
rect 2425 1760 2465 1765
rect 2425 1730 2430 1760
rect 2460 1730 2465 1760
rect 2425 1725 2465 1730
rect 2515 1760 2555 1765
rect 2515 1730 2520 1760
rect 2550 1730 2555 1760
rect 2515 1725 2555 1730
rect 2380 1665 2420 1670
rect 2380 1635 2385 1665
rect 2415 1635 2420 1665
rect 2380 1630 2420 1635
rect 2330 1595 2370 1600
rect 2330 1565 2335 1595
rect 2365 1565 2370 1595
rect 2330 1560 2370 1565
rect 275 1035 2175 1190
rect 2435 1035 2455 1725
rect 2580 1670 2600 1845
rect 2635 1765 2655 1845
rect 2795 1825 2815 1845
rect 3005 1825 3025 1845
rect 3125 1825 3145 1845
rect 2785 1820 2825 1825
rect 2785 1790 2790 1820
rect 2820 1790 2825 1820
rect 2785 1785 2825 1790
rect 2995 1820 3035 1825
rect 2995 1790 3000 1820
rect 3030 1790 3035 1820
rect 2995 1785 3035 1790
rect 3115 1820 3155 1825
rect 3115 1790 3120 1820
rect 3150 1790 3155 1820
rect 3115 1785 3155 1790
rect 3245 1765 3265 1845
rect 3365 1825 3385 1845
rect 3485 1825 3505 1845
rect 3725 1825 3745 1845
rect 3815 1825 3835 1845
rect 3355 1820 3395 1825
rect 3355 1790 3360 1820
rect 3390 1790 3395 1820
rect 3355 1785 3395 1790
rect 3475 1820 3515 1825
rect 3475 1790 3480 1820
rect 3510 1790 3515 1820
rect 3475 1785 3515 1790
rect 3715 1820 3755 1825
rect 3715 1790 3720 1820
rect 3750 1790 3755 1820
rect 3715 1785 3755 1790
rect 3805 1820 3845 1825
rect 3805 1790 3810 1820
rect 3840 1790 3845 1820
rect 3805 1785 3845 1790
rect 2625 1760 2665 1765
rect 2625 1730 2630 1760
rect 2660 1730 2665 1760
rect 2625 1725 2665 1730
rect 3175 1760 3215 1765
rect 3175 1730 3180 1760
rect 3210 1730 3215 1760
rect 3175 1725 3215 1730
rect 3235 1760 3275 1765
rect 3235 1730 3240 1760
rect 3270 1730 3275 1760
rect 3235 1725 3275 1730
rect 3365 1720 3385 1785
rect 3475 1760 3515 1765
rect 3475 1730 3480 1760
rect 3510 1730 3515 1760
rect 3475 1725 3515 1730
rect 3715 1760 3755 1765
rect 3715 1730 3720 1760
rect 3750 1730 3755 1760
rect 3715 1725 3755 1730
rect 3115 1715 3155 1720
rect 3115 1685 3120 1715
rect 3150 1685 3155 1715
rect 3115 1680 3155 1685
rect 3355 1715 3395 1720
rect 3355 1685 3360 1715
rect 3390 1685 3395 1715
rect 3355 1680 3395 1685
rect 3595 1715 3635 1720
rect 3595 1685 3600 1715
rect 3630 1685 3635 1715
rect 3595 1680 3635 1685
rect 2570 1665 2610 1670
rect 2570 1635 2575 1665
rect 2605 1635 2610 1665
rect 2570 1630 2610 1635
rect 2580 1085 2600 1630
rect 3115 1595 3155 1600
rect 3115 1565 3120 1595
rect 3150 1565 3155 1595
rect 3115 1560 3155 1565
rect 2785 1545 2825 1550
rect 2785 1515 2790 1545
rect 2820 1515 2825 1545
rect 2785 1510 2825 1515
rect 3175 1545 3215 1550
rect 3175 1515 3180 1545
rect 3210 1515 3215 1545
rect 3175 1510 3215 1515
rect 3295 1545 3335 1550
rect 3295 1515 3300 1545
rect 3330 1515 3335 1545
rect 3295 1510 3335 1515
rect 3415 1545 3455 1550
rect 3415 1515 3420 1545
rect 3450 1515 3455 1545
rect 3415 1510 3455 1515
rect 3535 1545 3575 1550
rect 3535 1515 3540 1545
rect 3570 1515 3575 1545
rect 3535 1510 3575 1515
rect 3655 1545 3695 1550
rect 3655 1515 3660 1545
rect 3690 1515 3695 1545
rect 3655 1510 3695 1515
rect 2795 1495 2815 1510
rect 3875 1495 3895 2015
rect 4005 2050 4065 2055
rect 4005 2020 4030 2050
rect 4060 2020 4065 2050
rect 4005 2015 4065 2020
rect 4385 2050 4425 2055
rect 4385 2020 4390 2050
rect 4420 2020 4425 2050
rect 4385 2015 4425 2020
rect 4745 2050 4785 2055
rect 4745 2020 4750 2050
rect 4780 2020 4785 2050
rect 4745 2015 4785 2020
rect 5105 2050 5145 2055
rect 5105 2020 5110 2050
rect 5140 2020 5145 2050
rect 5105 2015 5145 2020
rect 4005 1495 4025 2015
rect 4055 1875 4095 1885
rect 4055 1855 4065 1875
rect 4085 1855 4095 1875
rect 4055 1845 4095 1855
rect 4145 1875 4185 1885
rect 4145 1855 4155 1875
rect 4175 1855 4185 1875
rect 4145 1845 4185 1855
rect 4265 1880 4305 1885
rect 4265 1850 4270 1880
rect 4300 1850 4305 1880
rect 4265 1845 4305 1850
rect 4385 1875 4425 1885
rect 4385 1855 4395 1875
rect 4415 1855 4425 1875
rect 4385 1845 4425 1855
rect 4505 1875 4545 1885
rect 4505 1855 4515 1875
rect 4535 1855 4545 1875
rect 4505 1845 4545 1855
rect 4625 1880 4665 1885
rect 4625 1850 4630 1880
rect 4660 1850 4665 1880
rect 4625 1845 4665 1850
rect 4745 1875 4785 1885
rect 4745 1855 4755 1875
rect 4775 1855 4785 1875
rect 4745 1845 4785 1855
rect 4865 1875 4905 1885
rect 4865 1855 4875 1875
rect 4895 1855 4905 1875
rect 4865 1845 4905 1855
rect 4985 1880 5025 1885
rect 4985 1850 4990 1880
rect 5020 1850 5025 1880
rect 4985 1845 5025 1850
rect 5075 1875 5115 1885
rect 5075 1855 5085 1875
rect 5105 1855 5115 1875
rect 5075 1845 5115 1855
rect 4065 1825 4085 1845
rect 4155 1825 4175 1845
rect 4395 1825 4415 1845
rect 4515 1825 4535 1845
rect 4055 1820 4095 1825
rect 4055 1790 4060 1820
rect 4090 1790 4095 1820
rect 4055 1785 4095 1790
rect 4145 1820 4185 1825
rect 4145 1790 4150 1820
rect 4180 1790 4185 1820
rect 4145 1785 4185 1790
rect 4385 1820 4425 1825
rect 4385 1790 4390 1820
rect 4420 1790 4425 1820
rect 4385 1785 4425 1790
rect 4505 1820 4545 1825
rect 4505 1790 4510 1820
rect 4540 1790 4545 1820
rect 4505 1785 4545 1790
rect 4145 1760 4185 1765
rect 4145 1730 4150 1760
rect 4180 1730 4185 1760
rect 4145 1725 4185 1730
rect 4385 1760 4425 1765
rect 4385 1730 4390 1760
rect 4420 1730 4425 1760
rect 4385 1725 4425 1730
rect 4515 1720 4535 1785
rect 4635 1765 4655 1845
rect 4755 1825 4775 1845
rect 4875 1825 4895 1845
rect 5085 1825 5105 1845
rect 4745 1820 4785 1825
rect 4745 1790 4750 1820
rect 4780 1790 4785 1820
rect 4745 1785 4785 1790
rect 4865 1820 4905 1825
rect 4865 1790 4870 1820
rect 4900 1790 4905 1820
rect 4865 1785 4905 1790
rect 5075 1820 5115 1825
rect 5075 1790 5080 1820
rect 5110 1790 5115 1820
rect 5075 1785 5115 1790
rect 5210 1765 5230 2305
rect 5255 2150 5275 3060
rect 5245 2145 5285 2150
rect 5245 2115 5250 2145
rect 5280 2115 5285 2145
rect 5245 2110 5285 2115
rect 5300 1825 5320 3300
rect 5340 3285 5380 3290
rect 5340 3255 5345 3285
rect 5375 3255 5380 3285
rect 5340 3250 5380 3255
rect 5290 1820 5330 1825
rect 5290 1790 5295 1820
rect 5325 1790 5330 1820
rect 5290 1785 5330 1790
rect 4625 1760 4665 1765
rect 4625 1730 4630 1760
rect 4660 1730 4665 1760
rect 4625 1725 4665 1730
rect 4685 1760 4725 1765
rect 4685 1730 4690 1760
rect 4720 1730 4725 1760
rect 4685 1725 4725 1730
rect 5200 1760 5240 1765
rect 5200 1730 5205 1760
rect 5235 1730 5240 1760
rect 5200 1725 5240 1730
rect 4265 1715 4305 1720
rect 4265 1685 4270 1715
rect 4300 1685 4305 1715
rect 4265 1680 4305 1685
rect 4505 1715 4545 1720
rect 4505 1685 4510 1715
rect 4540 1685 4545 1715
rect 4505 1680 4545 1685
rect 4745 1715 4785 1720
rect 4745 1685 4750 1715
rect 4780 1685 4785 1715
rect 4745 1680 4785 1685
rect 5350 1600 5370 3250
rect 4745 1595 4785 1600
rect 4745 1565 4750 1595
rect 4780 1565 4785 1595
rect 4745 1560 4785 1565
rect 5340 1595 5380 1600
rect 5340 1565 5345 1595
rect 5375 1565 5380 1595
rect 5340 1560 5380 1565
rect 4205 1545 4245 1550
rect 4205 1515 4210 1545
rect 4240 1515 4245 1545
rect 4205 1510 4245 1515
rect 4325 1545 4365 1550
rect 4325 1515 4330 1545
rect 4360 1515 4365 1545
rect 4325 1510 4365 1515
rect 4445 1545 4485 1550
rect 4445 1515 4450 1545
rect 4480 1515 4485 1545
rect 4445 1510 4485 1515
rect 4565 1545 4605 1550
rect 4565 1515 4570 1545
rect 4600 1515 4605 1545
rect 4565 1510 4605 1515
rect 4685 1545 4725 1550
rect 4685 1515 4690 1545
rect 4720 1515 4725 1545
rect 4685 1510 4725 1515
rect 5075 1545 5115 1550
rect 5075 1515 5080 1545
rect 5110 1515 5115 1545
rect 5075 1510 5115 1515
rect 5085 1495 5105 1510
rect 2785 1485 2825 1495
rect 2785 1465 2795 1485
rect 2815 1465 2825 1485
rect 2785 1455 2825 1465
rect 3865 1485 3905 1495
rect 3865 1465 3875 1485
rect 3895 1465 3905 1485
rect 3865 1455 3905 1465
rect 3995 1485 4035 1495
rect 3995 1465 4005 1485
rect 4025 1465 4035 1485
rect 3995 1455 4035 1465
rect 5075 1485 5115 1495
rect 5075 1465 5085 1485
rect 5105 1465 5115 1485
rect 5075 1455 5115 1465
rect 2890 1165 2930 1170
rect 2890 1135 2895 1165
rect 2925 1135 2930 1165
rect 2890 1130 2930 1135
rect 2970 1165 3010 1170
rect 2970 1135 2975 1165
rect 3005 1135 3010 1165
rect 2970 1130 3010 1135
rect 3050 1165 3090 1170
rect 3050 1135 3055 1165
rect 3085 1135 3090 1165
rect 3050 1130 3090 1135
rect 3130 1165 3170 1170
rect 3130 1135 3135 1165
rect 3165 1135 3170 1165
rect 3130 1130 3170 1135
rect 3210 1165 3250 1170
rect 3210 1135 3215 1165
rect 3245 1135 3250 1165
rect 3210 1130 3250 1135
rect 3290 1165 3330 1170
rect 3290 1135 3295 1165
rect 3325 1135 3330 1165
rect 3290 1130 3330 1135
rect 3370 1165 3410 1170
rect 3370 1135 3375 1165
rect 3405 1135 3410 1165
rect 3370 1130 3410 1135
rect 3450 1165 3490 1170
rect 3450 1135 3455 1165
rect 3485 1135 3490 1165
rect 3450 1130 3490 1135
rect 3530 1165 3570 1170
rect 3530 1135 3535 1165
rect 3565 1135 3570 1165
rect 3530 1130 3570 1135
rect 3610 1165 3650 1170
rect 3610 1135 3615 1165
rect 3645 1135 3650 1165
rect 3610 1130 3650 1135
rect 3690 1165 3730 1170
rect 3690 1135 3695 1165
rect 3725 1135 3730 1165
rect 3690 1130 3730 1135
rect 3770 1165 3810 1170
rect 3770 1135 3775 1165
rect 3805 1135 3810 1165
rect 3770 1130 3810 1135
rect 3850 1165 3890 1170
rect 3850 1135 3855 1165
rect 3885 1135 3890 1165
rect 3850 1130 3890 1135
rect 3930 1165 3970 1170
rect 3930 1135 3935 1165
rect 3965 1135 3970 1165
rect 3930 1130 3970 1135
rect 4010 1165 4050 1170
rect 4010 1135 4015 1165
rect 4045 1135 4050 1165
rect 4010 1130 4050 1135
rect 4090 1165 4130 1170
rect 4090 1135 4095 1165
rect 4125 1135 4130 1165
rect 4090 1130 4130 1135
rect 4170 1165 4210 1170
rect 4170 1135 4175 1165
rect 4205 1135 4210 1165
rect 4170 1130 4210 1135
rect 4250 1165 4290 1170
rect 4250 1135 4255 1165
rect 4285 1135 4290 1165
rect 4250 1130 4290 1135
rect 4330 1165 4370 1170
rect 4330 1135 4335 1165
rect 4365 1135 4370 1165
rect 4330 1130 4370 1135
rect 4410 1165 4450 1170
rect 4410 1135 4415 1165
rect 4445 1135 4450 1165
rect 4410 1130 4450 1135
rect 4490 1165 4530 1170
rect 4490 1135 4495 1165
rect 4525 1135 4530 1165
rect 4490 1130 4530 1135
rect 4570 1165 4610 1170
rect 4570 1135 4575 1165
rect 4605 1135 4610 1165
rect 4570 1130 4610 1135
rect 4650 1165 4690 1170
rect 4650 1135 4655 1165
rect 4685 1135 4690 1165
rect 4650 1130 4690 1135
rect 4730 1165 4770 1170
rect 4730 1135 4735 1165
rect 4765 1135 4770 1165
rect 4730 1130 4770 1135
rect 4810 1165 4850 1170
rect 4810 1135 4815 1165
rect 4845 1135 4850 1165
rect 4810 1130 4850 1135
rect 4890 1165 4930 1170
rect 4890 1135 4895 1165
rect 4925 1135 4930 1165
rect 4890 1130 4930 1135
rect 2570 1080 2610 1085
rect 2570 1050 2575 1080
rect 2605 1050 2610 1080
rect 2570 1045 2610 1050
rect 2850 1080 2890 1085
rect 2850 1050 2855 1080
rect 2885 1050 2890 1080
rect 2850 1045 2890 1050
rect 275 1030 2215 1035
rect 275 1000 2180 1030
rect 2210 1000 2215 1030
rect 275 995 2215 1000
rect 2425 1030 2465 1035
rect 2425 1000 2430 1030
rect 2460 1000 2465 1030
rect 2425 995 2465 1000
rect 275 840 2175 995
<< via1 >>
rect 4445 3465 4475 3495
rect -10 3415 20 3445
rect 945 3415 975 3445
rect 1645 3415 1675 3445
rect 2475 3420 2505 3450
rect -55 3360 -25 3390
rect -55 2825 -25 2855
rect 1195 3310 1225 3340
rect 1150 3255 1180 3285
rect 45 3200 80 3205
rect 45 3175 50 3200
rect 50 3175 75 3200
rect 75 3175 80 3200
rect 45 3170 80 3175
rect 45 3140 80 3145
rect 45 3115 50 3140
rect 50 3115 75 3140
rect 75 3115 80 3140
rect 45 3110 80 3115
rect 1150 3070 1180 3100
rect 45 3060 80 3065
rect 45 3035 50 3060
rect 50 3035 75 3060
rect 75 3035 80 3060
rect 45 3030 80 3035
rect 45 3000 80 3005
rect 45 2975 50 3000
rect 50 2975 75 3000
rect 75 2975 80 3000
rect 45 2970 80 2975
rect 1250 3195 1285 3200
rect 1250 3170 1255 3195
rect 1255 3170 1280 3195
rect 1280 3170 1285 3195
rect 1250 3165 1285 3170
rect 1250 3135 1285 3140
rect 1250 3110 1255 3135
rect 1255 3110 1280 3135
rect 1280 3110 1285 3135
rect 1250 3105 1285 3110
rect 2335 2955 2370 2960
rect 2335 2930 2340 2955
rect 2340 2930 2365 2955
rect 2365 2930 2370 2955
rect 2335 2925 2370 2930
rect 2430 2925 2460 2955
rect 2335 2895 2370 2900
rect 2335 2870 2340 2895
rect 2340 2870 2365 2895
rect 2365 2870 2370 2895
rect 2335 2865 2370 2870
rect 45 2850 80 2855
rect 45 2825 50 2850
rect 50 2825 75 2850
rect 75 2825 80 2850
rect 45 2820 80 2825
rect 580 2850 615 2855
rect 580 2825 585 2850
rect 585 2825 610 2850
rect 610 2825 615 2850
rect 580 2820 615 2825
rect 1195 2820 1225 2850
rect 1250 2835 1285 2840
rect 1250 2810 1255 2835
rect 1255 2810 1280 2835
rect 1280 2810 1285 2835
rect 1250 2805 1285 2810
rect 1965 2835 2000 2840
rect 1965 2810 1970 2835
rect 1970 2810 1995 2835
rect 1995 2810 2000 2835
rect 1965 2805 2000 2810
rect 2335 2805 2365 2835
rect -10 2765 20 2795
rect 45 2790 80 2795
rect 45 2765 50 2790
rect 50 2765 75 2790
rect 75 2765 80 2790
rect 45 2760 80 2765
rect 580 2790 615 2795
rect 580 2765 585 2790
rect 585 2765 610 2790
rect 610 2765 615 2790
rect 580 2760 615 2765
rect 1250 2715 1280 2745
rect 2155 2715 2185 2745
rect -105 1690 -75 1720
rect -40 1715 -10 1720
rect -40 1695 -35 1715
rect -35 1695 -15 1715
rect -15 1695 -10 1715
rect -40 1690 -10 1695
rect 1270 1680 1300 1710
rect 2430 2215 2460 2245
rect 2335 2170 2365 2200
rect 2155 1680 2185 1710
rect 2385 2120 2415 2150
rect 2695 3360 2725 3390
rect 2950 3310 2980 3340
rect 3395 3305 3425 3335
rect 2690 3210 2720 3240
rect 2575 3155 2605 3185
rect 2575 2760 2605 2790
rect 2575 2365 2605 2395
rect 5145 3415 5175 3445
rect 5295 3305 5325 3335
rect 4445 3155 4475 3185
rect 2950 3065 2980 3095
rect 5250 3065 5280 3095
rect 2945 2795 2975 2800
rect 2945 2775 2950 2795
rect 2950 2775 2970 2795
rect 2970 2775 2975 2795
rect 2945 2770 2975 2775
rect 3125 2795 3155 2800
rect 3125 2775 3130 2795
rect 3130 2775 3150 2795
rect 3150 2775 3155 2795
rect 3125 2770 3155 2775
rect 3305 2795 3335 2800
rect 3305 2775 3310 2795
rect 3310 2775 3330 2795
rect 3330 2775 3335 2795
rect 3305 2770 3335 2775
rect 3485 2795 3515 2800
rect 3485 2775 3490 2795
rect 3490 2775 3510 2795
rect 3510 2775 3515 2795
rect 3485 2770 3515 2775
rect 3665 2795 3695 2800
rect 3665 2775 3670 2795
rect 3670 2775 3690 2795
rect 3690 2775 3695 2795
rect 3665 2770 3695 2775
rect 3845 2795 3875 2800
rect 3845 2775 3850 2795
rect 3850 2775 3870 2795
rect 3870 2775 3875 2795
rect 3845 2770 3875 2775
rect 4025 2795 4055 2800
rect 4025 2775 4030 2795
rect 4030 2775 4050 2795
rect 4050 2775 4055 2795
rect 4025 2770 4055 2775
rect 4205 2795 4235 2800
rect 4205 2775 4210 2795
rect 4210 2775 4230 2795
rect 4230 2775 4235 2795
rect 4205 2770 4235 2775
rect 4385 2795 4415 2800
rect 4385 2775 4390 2795
rect 4390 2775 4410 2795
rect 4410 2775 4415 2795
rect 4385 2770 4415 2775
rect 4565 2795 4595 2800
rect 4565 2775 4570 2795
rect 4570 2775 4590 2795
rect 4590 2775 4595 2795
rect 4565 2770 4595 2775
rect 4745 2795 4775 2800
rect 4745 2775 4750 2795
rect 4750 2775 4770 2795
rect 4770 2775 4775 2795
rect 4745 2770 4775 2775
rect 4925 2795 4955 2800
rect 4925 2775 4930 2795
rect 4930 2775 4950 2795
rect 4950 2775 4955 2795
rect 4925 2770 4955 2775
rect 2945 2420 2975 2425
rect 2945 2400 2950 2420
rect 2950 2400 2970 2420
rect 2970 2400 2975 2420
rect 2945 2395 2975 2400
rect 3035 2425 3065 2430
rect 3035 2405 3040 2425
rect 3040 2405 3060 2425
rect 3060 2405 3065 2425
rect 3035 2400 3065 2405
rect 3755 2425 3785 2430
rect 3755 2405 3760 2425
rect 3760 2405 3780 2425
rect 3780 2405 3785 2425
rect 3755 2400 3785 2405
rect 4105 2425 4135 2430
rect 4105 2405 4110 2425
rect 4110 2405 4130 2425
rect 4130 2405 4135 2425
rect 4105 2400 4135 2405
rect 4835 2425 4865 2430
rect 4835 2405 4840 2425
rect 4840 2405 4860 2425
rect 4860 2405 4865 2425
rect 4835 2400 4865 2405
rect 2690 2310 2720 2340
rect 3215 2380 3245 2385
rect 3215 2360 3220 2380
rect 3220 2360 3240 2380
rect 3240 2360 3245 2380
rect 3215 2355 3245 2360
rect 3035 2215 3065 2245
rect 2855 2170 2885 2200
rect 3575 2380 3605 2385
rect 3575 2360 3580 2380
rect 3580 2360 3600 2380
rect 3600 2360 3605 2380
rect 3575 2355 3605 2360
rect 3395 2335 3425 2340
rect 3395 2315 3400 2335
rect 3400 2315 3420 2335
rect 3420 2315 3425 2335
rect 3395 2310 3425 2315
rect 3215 2120 3245 2150
rect 2820 2090 2850 2095
rect 2820 2070 2825 2090
rect 2825 2070 2845 2090
rect 2845 2070 2850 2090
rect 2820 2065 2850 2070
rect 2940 2090 2970 2095
rect 2940 2070 2945 2090
rect 2945 2070 2965 2090
rect 2965 2070 2970 2090
rect 2940 2065 2970 2070
rect 3060 2090 3090 2095
rect 3060 2070 3065 2090
rect 3065 2070 3085 2090
rect 3085 2070 3090 2090
rect 3060 2065 3090 2070
rect 3180 2090 3210 2095
rect 3180 2070 3185 2090
rect 3185 2070 3205 2090
rect 3205 2070 3210 2090
rect 3180 2065 3210 2070
rect 3300 2090 3330 2095
rect 3300 2070 3305 2090
rect 3305 2070 3325 2090
rect 3325 2070 3330 2090
rect 3300 2065 3330 2070
rect 3420 2090 3450 2095
rect 3420 2070 3425 2090
rect 3425 2070 3445 2090
rect 3445 2070 3450 2090
rect 3420 2065 3450 2070
rect 3540 2090 3570 2095
rect 3540 2070 3545 2090
rect 3545 2070 3565 2090
rect 3565 2070 3570 2090
rect 3540 2065 3570 2070
rect 3660 2090 3690 2095
rect 3660 2070 3665 2090
rect 3665 2070 3685 2090
rect 3685 2070 3690 2090
rect 3660 2065 3690 2070
rect 3780 2090 3810 2095
rect 3780 2070 3785 2090
rect 3785 2070 3805 2090
rect 3805 2070 3810 2090
rect 3780 2065 3810 2070
rect 4295 2380 4325 2385
rect 4295 2360 4300 2380
rect 4300 2360 4320 2380
rect 4320 2360 4325 2380
rect 4295 2355 4325 2360
rect 4655 2380 4685 2385
rect 4655 2360 4660 2380
rect 4660 2360 4680 2380
rect 4680 2360 4685 2380
rect 4655 2355 4685 2360
rect 4475 2335 4505 2340
rect 4475 2315 4480 2335
rect 4480 2315 4500 2335
rect 4500 2315 4505 2335
rect 4475 2310 4505 2315
rect 5205 2310 5235 2340
rect 3935 2170 3965 2200
rect 5015 2170 5045 2200
rect 4030 2115 4060 2145
rect 4090 2090 4120 2095
rect 4090 2070 4095 2090
rect 4095 2070 4115 2090
rect 4115 2070 4120 2090
rect 4090 2065 4120 2070
rect 4210 2090 4240 2095
rect 4210 2070 4215 2090
rect 4215 2070 4235 2090
rect 4235 2070 4240 2090
rect 4210 2065 4240 2070
rect 4330 2090 4360 2095
rect 4330 2070 4335 2090
rect 4335 2070 4355 2090
rect 4355 2070 4360 2090
rect 4330 2065 4360 2070
rect 4450 2090 4480 2095
rect 4450 2070 4455 2090
rect 4455 2070 4475 2090
rect 4475 2070 4480 2090
rect 4450 2065 4480 2070
rect 4570 2090 4600 2095
rect 4570 2070 4575 2090
rect 4575 2070 4595 2090
rect 4595 2070 4600 2090
rect 4570 2065 4600 2070
rect 4690 2090 4720 2095
rect 4690 2070 4695 2090
rect 4695 2070 4715 2090
rect 4715 2070 4720 2090
rect 4690 2065 4720 2070
rect 4810 2090 4840 2095
rect 4810 2070 4815 2090
rect 4815 2070 4835 2090
rect 4835 2070 4840 2090
rect 4810 2065 4840 2070
rect 4930 2090 4960 2095
rect 4930 2070 4935 2090
rect 4935 2070 4955 2090
rect 4955 2070 4960 2090
rect 4930 2065 4960 2070
rect 5050 2090 5080 2095
rect 5050 2070 5055 2090
rect 5055 2070 5075 2090
rect 5075 2070 5080 2090
rect 5050 2065 5080 2070
rect 2575 2045 2605 2050
rect 2575 2025 2580 2045
rect 2580 2025 2600 2045
rect 2600 2025 2605 2045
rect 2575 2020 2605 2025
rect 2760 2045 2790 2050
rect 2760 2025 2765 2045
rect 2765 2025 2785 2045
rect 2785 2025 2790 2045
rect 2760 2020 2790 2025
rect 3120 2045 3150 2050
rect 3120 2025 3125 2045
rect 3125 2025 3145 2045
rect 3145 2025 3150 2045
rect 3120 2020 3150 2025
rect 3480 2045 3510 2050
rect 3480 2025 3485 2045
rect 3485 2025 3505 2045
rect 3505 2025 3510 2045
rect 3480 2020 3510 2025
rect 3840 2045 3870 2050
rect 3840 2025 3845 2045
rect 3845 2025 3865 2045
rect 3865 2025 3870 2045
rect 3840 2020 3870 2025
rect 2880 1875 2910 1880
rect 2880 1855 2885 1875
rect 2885 1855 2905 1875
rect 2905 1855 2910 1875
rect 2880 1850 2910 1855
rect 3240 1875 3270 1880
rect 3240 1855 3245 1875
rect 3245 1855 3265 1875
rect 3265 1855 3270 1875
rect 3240 1850 3270 1855
rect 3600 1875 3630 1880
rect 3600 1855 3605 1875
rect 3605 1855 3625 1875
rect 3625 1855 3630 1875
rect 3600 1850 3630 1855
rect 2475 1790 2505 1820
rect 2430 1730 2460 1760
rect 2520 1730 2550 1760
rect 2385 1635 2415 1665
rect 2335 1565 2365 1595
rect 2790 1790 2820 1820
rect 3000 1815 3030 1820
rect 3000 1795 3005 1815
rect 3005 1795 3025 1815
rect 3025 1795 3030 1815
rect 3000 1790 3030 1795
rect 3120 1790 3150 1820
rect 3360 1815 3390 1820
rect 3360 1795 3365 1815
rect 3365 1795 3385 1815
rect 3385 1795 3390 1815
rect 3360 1790 3390 1795
rect 3480 1790 3510 1820
rect 3720 1815 3750 1820
rect 3720 1795 3725 1815
rect 3725 1795 3745 1815
rect 3745 1795 3750 1815
rect 3720 1790 3750 1795
rect 3810 1790 3840 1820
rect 2630 1730 2660 1760
rect 3180 1755 3210 1760
rect 3180 1735 3185 1755
rect 3185 1735 3205 1755
rect 3205 1735 3210 1755
rect 3180 1730 3210 1735
rect 3240 1755 3270 1760
rect 3240 1735 3245 1755
rect 3245 1735 3265 1755
rect 3265 1735 3270 1755
rect 3240 1730 3270 1735
rect 3480 1755 3510 1760
rect 3480 1735 3485 1755
rect 3485 1735 3505 1755
rect 3505 1735 3510 1755
rect 3480 1730 3510 1735
rect 3720 1755 3750 1760
rect 3720 1735 3725 1755
rect 3725 1735 3745 1755
rect 3745 1735 3750 1755
rect 3720 1730 3750 1735
rect 3120 1710 3150 1715
rect 3120 1690 3125 1710
rect 3125 1690 3145 1710
rect 3145 1690 3150 1710
rect 3120 1685 3150 1690
rect 3360 1710 3390 1715
rect 3360 1690 3365 1710
rect 3365 1690 3385 1710
rect 3385 1690 3390 1710
rect 3360 1685 3390 1690
rect 3600 1710 3630 1715
rect 3600 1690 3605 1710
rect 3605 1690 3625 1710
rect 3625 1690 3630 1710
rect 3600 1685 3630 1690
rect 2575 1635 2605 1665
rect 3120 1590 3150 1595
rect 3120 1570 3125 1590
rect 3125 1570 3145 1590
rect 3145 1570 3150 1590
rect 3120 1565 3150 1570
rect 2790 1515 2820 1545
rect 3180 1540 3210 1545
rect 3180 1520 3185 1540
rect 3185 1520 3205 1540
rect 3205 1520 3210 1540
rect 3180 1515 3210 1520
rect 3300 1540 3330 1545
rect 3300 1520 3305 1540
rect 3305 1520 3325 1540
rect 3325 1520 3330 1540
rect 3300 1515 3330 1520
rect 3420 1540 3450 1545
rect 3420 1520 3425 1540
rect 3425 1520 3445 1540
rect 3445 1520 3450 1540
rect 3420 1515 3450 1520
rect 3540 1540 3570 1545
rect 3540 1520 3545 1540
rect 3545 1520 3565 1540
rect 3565 1520 3570 1540
rect 3540 1515 3570 1520
rect 3660 1540 3690 1545
rect 3660 1520 3665 1540
rect 3665 1520 3685 1540
rect 3685 1520 3690 1540
rect 3660 1515 3690 1520
rect 4030 2045 4060 2050
rect 4030 2025 4035 2045
rect 4035 2025 4055 2045
rect 4055 2025 4060 2045
rect 4030 2020 4060 2025
rect 4390 2045 4420 2050
rect 4390 2025 4395 2045
rect 4395 2025 4415 2045
rect 4415 2025 4420 2045
rect 4390 2020 4420 2025
rect 4750 2045 4780 2050
rect 4750 2025 4755 2045
rect 4755 2025 4775 2045
rect 4775 2025 4780 2045
rect 4750 2020 4780 2025
rect 5110 2045 5140 2050
rect 5110 2025 5115 2045
rect 5115 2025 5135 2045
rect 5135 2025 5140 2045
rect 5110 2020 5140 2025
rect 4270 1875 4300 1880
rect 4270 1855 4275 1875
rect 4275 1855 4295 1875
rect 4295 1855 4300 1875
rect 4270 1850 4300 1855
rect 4630 1875 4660 1880
rect 4630 1855 4635 1875
rect 4635 1855 4655 1875
rect 4655 1855 4660 1875
rect 4630 1850 4660 1855
rect 4990 1875 5020 1880
rect 4990 1855 4995 1875
rect 4995 1855 5015 1875
rect 5015 1855 5020 1875
rect 4990 1850 5020 1855
rect 4060 1790 4090 1820
rect 4150 1815 4180 1820
rect 4150 1795 4155 1815
rect 4155 1795 4175 1815
rect 4175 1795 4180 1815
rect 4150 1790 4180 1795
rect 4390 1790 4420 1820
rect 4510 1815 4540 1820
rect 4510 1795 4515 1815
rect 4515 1795 4535 1815
rect 4535 1795 4540 1815
rect 4510 1790 4540 1795
rect 4150 1755 4180 1760
rect 4150 1735 4155 1755
rect 4155 1735 4175 1755
rect 4175 1735 4180 1755
rect 4150 1730 4180 1735
rect 4390 1755 4420 1760
rect 4390 1735 4395 1755
rect 4395 1735 4415 1755
rect 4415 1735 4420 1755
rect 4390 1730 4420 1735
rect 4750 1790 4780 1820
rect 4870 1815 4900 1820
rect 4870 1795 4875 1815
rect 4875 1795 4895 1815
rect 4895 1795 4900 1815
rect 4870 1790 4900 1795
rect 5080 1790 5110 1820
rect 5250 2115 5280 2145
rect 5345 3255 5375 3285
rect 5295 1790 5325 1820
rect 4630 1755 4660 1760
rect 4630 1735 4635 1755
rect 4635 1735 4655 1755
rect 4655 1735 4660 1755
rect 4630 1730 4660 1735
rect 4690 1755 4720 1760
rect 4690 1735 4695 1755
rect 4695 1735 4715 1755
rect 4715 1735 4720 1755
rect 4690 1730 4720 1735
rect 5205 1730 5235 1760
rect 4270 1710 4300 1715
rect 4270 1690 4275 1710
rect 4275 1690 4295 1710
rect 4295 1690 4300 1710
rect 4270 1685 4300 1690
rect 4510 1710 4540 1715
rect 4510 1690 4515 1710
rect 4515 1690 4535 1710
rect 4535 1690 4540 1710
rect 4510 1685 4540 1690
rect 4750 1710 4780 1715
rect 4750 1690 4755 1710
rect 4755 1690 4775 1710
rect 4775 1690 4780 1710
rect 4750 1685 4780 1690
rect 4750 1590 4780 1595
rect 4750 1570 4755 1590
rect 4755 1570 4775 1590
rect 4775 1570 4780 1590
rect 4750 1565 4780 1570
rect 5345 1565 5375 1595
rect 4210 1540 4240 1545
rect 4210 1520 4215 1540
rect 4215 1520 4235 1540
rect 4235 1520 4240 1540
rect 4210 1515 4240 1520
rect 4330 1540 4360 1545
rect 4330 1520 4335 1540
rect 4335 1520 4355 1540
rect 4355 1520 4360 1540
rect 4330 1515 4360 1520
rect 4450 1540 4480 1545
rect 4450 1520 4455 1540
rect 4455 1520 4475 1540
rect 4475 1520 4480 1540
rect 4450 1515 4480 1520
rect 4570 1540 4600 1545
rect 4570 1520 4575 1540
rect 4575 1520 4595 1540
rect 4595 1520 4600 1540
rect 4570 1515 4600 1520
rect 4690 1540 4720 1545
rect 4690 1520 4695 1540
rect 4695 1520 4715 1540
rect 4715 1520 4720 1540
rect 4690 1515 4720 1520
rect 5080 1515 5110 1545
rect 2895 1160 2925 1165
rect 2895 1140 2900 1160
rect 2900 1140 2920 1160
rect 2920 1140 2925 1160
rect 2895 1135 2925 1140
rect 2975 1160 3005 1165
rect 2975 1140 2980 1160
rect 2980 1140 3000 1160
rect 3000 1140 3005 1160
rect 2975 1135 3005 1140
rect 3055 1160 3085 1165
rect 3055 1140 3060 1160
rect 3060 1140 3080 1160
rect 3080 1140 3085 1160
rect 3055 1135 3085 1140
rect 3135 1160 3165 1165
rect 3135 1140 3140 1160
rect 3140 1140 3160 1160
rect 3160 1140 3165 1160
rect 3135 1135 3165 1140
rect 3215 1160 3245 1165
rect 3215 1140 3220 1160
rect 3220 1140 3240 1160
rect 3240 1140 3245 1160
rect 3215 1135 3245 1140
rect 3295 1160 3325 1165
rect 3295 1140 3300 1160
rect 3300 1140 3320 1160
rect 3320 1140 3325 1160
rect 3295 1135 3325 1140
rect 3375 1160 3405 1165
rect 3375 1140 3380 1160
rect 3380 1140 3400 1160
rect 3400 1140 3405 1160
rect 3375 1135 3405 1140
rect 3455 1160 3485 1165
rect 3455 1140 3460 1160
rect 3460 1140 3480 1160
rect 3480 1140 3485 1160
rect 3455 1135 3485 1140
rect 3535 1160 3565 1165
rect 3535 1140 3540 1160
rect 3540 1140 3560 1160
rect 3560 1140 3565 1160
rect 3535 1135 3565 1140
rect 3615 1160 3645 1165
rect 3615 1140 3620 1160
rect 3620 1140 3640 1160
rect 3640 1140 3645 1160
rect 3615 1135 3645 1140
rect 3695 1160 3725 1165
rect 3695 1140 3700 1160
rect 3700 1140 3720 1160
rect 3720 1140 3725 1160
rect 3695 1135 3725 1140
rect 3775 1160 3805 1165
rect 3775 1140 3780 1160
rect 3780 1140 3800 1160
rect 3800 1140 3805 1160
rect 3775 1135 3805 1140
rect 3855 1160 3885 1165
rect 3855 1140 3860 1160
rect 3860 1140 3880 1160
rect 3880 1140 3885 1160
rect 3855 1135 3885 1140
rect 3935 1160 3965 1165
rect 3935 1140 3940 1160
rect 3940 1140 3960 1160
rect 3960 1140 3965 1160
rect 3935 1135 3965 1140
rect 4015 1160 4045 1165
rect 4015 1140 4020 1160
rect 4020 1140 4040 1160
rect 4040 1140 4045 1160
rect 4015 1135 4045 1140
rect 4095 1160 4125 1165
rect 4095 1140 4100 1160
rect 4100 1140 4120 1160
rect 4120 1140 4125 1160
rect 4095 1135 4125 1140
rect 4175 1160 4205 1165
rect 4175 1140 4180 1160
rect 4180 1140 4200 1160
rect 4200 1140 4205 1160
rect 4175 1135 4205 1140
rect 4255 1160 4285 1165
rect 4255 1140 4260 1160
rect 4260 1140 4280 1160
rect 4280 1140 4285 1160
rect 4255 1135 4285 1140
rect 4335 1160 4365 1165
rect 4335 1140 4340 1160
rect 4340 1140 4360 1160
rect 4360 1140 4365 1160
rect 4335 1135 4365 1140
rect 4415 1160 4445 1165
rect 4415 1140 4420 1160
rect 4420 1140 4440 1160
rect 4440 1140 4445 1160
rect 4415 1135 4445 1140
rect 4495 1160 4525 1165
rect 4495 1140 4500 1160
rect 4500 1140 4520 1160
rect 4520 1140 4525 1160
rect 4495 1135 4525 1140
rect 4575 1160 4605 1165
rect 4575 1140 4580 1160
rect 4580 1140 4600 1160
rect 4600 1140 4605 1160
rect 4575 1135 4605 1140
rect 4655 1160 4685 1165
rect 4655 1140 4660 1160
rect 4660 1140 4680 1160
rect 4680 1140 4685 1160
rect 4655 1135 4685 1140
rect 4735 1160 4765 1165
rect 4735 1140 4740 1160
rect 4740 1140 4760 1160
rect 4760 1140 4765 1160
rect 4735 1135 4765 1140
rect 4815 1160 4845 1165
rect 4815 1140 4820 1160
rect 4820 1140 4840 1160
rect 4840 1140 4845 1160
rect 4815 1135 4845 1140
rect 4895 1160 4925 1165
rect 4895 1140 4900 1160
rect 4900 1140 4920 1160
rect 4920 1140 4925 1160
rect 4895 1135 4925 1140
rect 2575 1050 2605 1080
rect 2855 1075 2885 1080
rect 2855 1055 2860 1075
rect 2860 1055 2880 1075
rect 2880 1055 2885 1075
rect 2855 1050 2885 1055
rect 2180 1000 2210 1030
rect 2430 1000 2460 1030
<< metal2 >>
rect -195 5005 -155 5010
rect -195 4975 -190 5005
rect -160 4975 -155 5005
rect -195 4970 -155 4975
rect 5480 5005 5520 5010
rect 5480 4975 5485 5005
rect 5515 4975 5520 5005
rect 5480 4970 5520 4975
rect 4440 3495 4480 3500
rect 4440 3465 4445 3495
rect 4475 3465 4480 3495
rect 4440 3460 4480 3465
rect -15 3445 25 3450
rect -15 3415 -10 3445
rect 20 3440 25 3445
rect 940 3445 980 3450
rect 940 3440 945 3445
rect 20 3420 945 3440
rect 20 3415 25 3420
rect -15 3410 25 3415
rect 940 3415 945 3420
rect 975 3415 980 3445
rect 940 3410 980 3415
rect 1635 3445 1685 3455
rect 2470 3450 2510 3455
rect 2470 3445 2475 3450
rect 1635 3415 1645 3445
rect 1675 3425 2475 3445
rect 1675 3415 1685 3425
rect 2470 3420 2475 3425
rect 2505 3420 2510 3450
rect 2470 3415 2510 3420
rect 5135 3445 5185 3455
rect 5135 3415 5145 3445
rect 5175 3415 5185 3445
rect 1635 3405 1685 3415
rect 5135 3405 5185 3415
rect -60 3390 -20 3395
rect -60 3360 -55 3390
rect -25 3385 -20 3390
rect 2690 3390 2730 3395
rect 2690 3385 2695 3390
rect -25 3365 2695 3385
rect -25 3360 -20 3365
rect -60 3355 -20 3360
rect 2690 3360 2695 3365
rect 2725 3360 2730 3390
rect 2690 3355 2730 3360
rect 1190 3340 1230 3345
rect 1190 3310 1195 3340
rect 1225 3335 1230 3340
rect 2945 3340 2985 3345
rect 2945 3335 2950 3340
rect 1225 3315 2950 3335
rect 1225 3310 1230 3315
rect 1190 3305 1230 3310
rect 2945 3310 2950 3315
rect 2980 3310 2985 3340
rect 2945 3305 2985 3310
rect 3385 3335 3435 3345
rect 3385 3305 3395 3335
rect 3425 3330 3435 3335
rect 5290 3335 5330 3340
rect 5290 3330 5295 3335
rect 3425 3310 5295 3330
rect 3425 3305 3435 3310
rect 3385 3295 3435 3305
rect 5290 3305 5295 3310
rect 5325 3305 5330 3335
rect 5290 3300 5330 3305
rect 1145 3285 1185 3290
rect 1145 3255 1150 3285
rect 1180 3280 1185 3285
rect 5340 3285 5380 3290
rect 5340 3280 5345 3285
rect 1180 3260 5345 3280
rect 1180 3255 1185 3260
rect 1145 3250 1185 3255
rect 5340 3255 5345 3260
rect 5375 3255 5380 3285
rect 5340 3250 5380 3255
rect 2685 3240 2725 3245
rect 2685 3235 2690 3240
rect 40 3215 2690 3235
rect 40 3205 85 3215
rect 2685 3210 2690 3215
rect 2720 3210 2725 3240
rect 2685 3205 2725 3210
rect 40 3170 45 3205
rect 80 3170 85 3205
rect 1245 3195 1250 3200
rect 1240 3175 1250 3195
rect 1245 3165 1250 3175
rect 1285 3165 1290 3200
rect 2570 3185 2610 3190
rect 2570 3155 2575 3185
rect 2605 3180 2610 3185
rect 4440 3185 4480 3190
rect 4440 3180 4445 3185
rect 2605 3160 4445 3180
rect 2605 3155 2610 3160
rect 2570 3150 2610 3155
rect 4440 3155 4445 3160
rect 4475 3155 4480 3185
rect 4440 3150 4480 3155
rect 40 3135 45 3145
rect 30 3115 45 3135
rect 40 3110 45 3115
rect 80 3110 85 3145
rect 1245 3135 1250 3140
rect 1240 3115 1250 3135
rect 1245 3105 1250 3115
rect 1285 3105 1290 3140
rect 1145 3100 1185 3105
rect 1145 3095 1150 3100
rect 40 3075 1150 3095
rect 40 3065 85 3075
rect 1145 3070 1150 3075
rect 1180 3070 1185 3100
rect 1145 3065 1185 3070
rect 2945 3095 2985 3100
rect 2945 3065 2950 3095
rect 2980 3090 2985 3095
rect 5245 3095 5285 3100
rect 5245 3090 5250 3095
rect 2980 3070 5250 3090
rect 2980 3065 2985 3070
rect 40 3030 45 3065
rect 80 3030 85 3065
rect 2945 3060 2985 3065
rect 5245 3065 5250 3070
rect 5280 3065 5285 3095
rect 5245 3060 5285 3065
rect 2945 3005 2985 3045
rect 40 2995 45 3005
rect 30 2975 45 2995
rect 40 2970 45 2975
rect 80 2970 85 3005
rect 2330 2925 2335 2960
rect 2370 2950 2375 2960
rect 2425 2955 2465 2960
rect 2425 2950 2430 2955
rect 2370 2930 2430 2950
rect 2370 2925 2375 2930
rect 2425 2925 2430 2930
rect 2460 2925 2465 2955
rect 2425 2920 2465 2925
rect 2330 2900 2375 2905
rect 2330 2865 2335 2900
rect 2370 2865 2375 2900
rect 2330 2860 2375 2865
rect -60 2855 -20 2860
rect -60 2825 -55 2855
rect -25 2850 -20 2855
rect 40 2850 45 2855
rect -25 2830 45 2850
rect -25 2825 -20 2830
rect -60 2820 -20 2825
rect 40 2820 45 2830
rect 80 2820 85 2855
rect 575 2820 580 2855
rect 615 2845 620 2855
rect 1190 2850 1230 2855
rect 1190 2845 1195 2850
rect 615 2825 1195 2845
rect 615 2820 620 2825
rect 1190 2820 1195 2825
rect 1225 2820 1230 2850
rect 1190 2815 1230 2820
rect 1245 2805 1250 2840
rect 1285 2805 1290 2840
rect 1960 2805 1965 2840
rect 2000 2830 2005 2840
rect 2330 2835 2370 2840
rect 2330 2830 2335 2835
rect 2000 2810 2335 2830
rect 2000 2805 2005 2810
rect 2330 2805 2335 2810
rect 2365 2805 2370 2835
rect 2330 2800 2370 2805
rect 2940 2800 2980 2805
rect -15 2795 25 2800
rect -15 2765 -10 2795
rect 20 2785 25 2795
rect 40 2785 45 2795
rect 20 2765 45 2785
rect -15 2760 25 2765
rect 40 2760 45 2765
rect 80 2760 85 2795
rect 575 2760 580 2795
rect 615 2785 620 2795
rect 2570 2790 2610 2795
rect 2570 2785 2575 2790
rect 615 2765 2575 2785
rect 615 2760 620 2765
rect 2570 2760 2575 2765
rect 2605 2760 2610 2790
rect 2940 2770 2945 2800
rect 2975 2795 2980 2800
rect 3120 2800 3160 2805
rect 3120 2795 3125 2800
rect 2975 2775 3125 2795
rect 2975 2770 2980 2775
rect 2940 2765 2980 2770
rect 3120 2770 3125 2775
rect 3155 2795 3160 2800
rect 3300 2800 3340 2805
rect 3300 2795 3305 2800
rect 3155 2775 3305 2795
rect 3155 2770 3160 2775
rect 3120 2765 3160 2770
rect 3300 2770 3305 2775
rect 3335 2795 3340 2800
rect 3480 2800 3520 2805
rect 3480 2795 3485 2800
rect 3335 2775 3485 2795
rect 3335 2770 3340 2775
rect 3300 2765 3340 2770
rect 3480 2770 3485 2775
rect 3515 2795 3520 2800
rect 3660 2800 3700 2805
rect 3660 2795 3665 2800
rect 3515 2775 3665 2795
rect 3515 2770 3520 2775
rect 3480 2765 3520 2770
rect 3660 2770 3665 2775
rect 3695 2795 3700 2800
rect 3840 2800 3880 2805
rect 3840 2795 3845 2800
rect 3695 2775 3845 2795
rect 3695 2770 3700 2775
rect 3660 2765 3700 2770
rect 3840 2770 3845 2775
rect 3875 2795 3880 2800
rect 4020 2800 4060 2805
rect 4020 2795 4025 2800
rect 3875 2775 4025 2795
rect 3875 2770 3880 2775
rect 3840 2765 3880 2770
rect 4020 2770 4025 2775
rect 4055 2795 4060 2800
rect 4200 2800 4240 2805
rect 4200 2795 4205 2800
rect 4055 2775 4205 2795
rect 4055 2770 4060 2775
rect 4020 2765 4060 2770
rect 4200 2770 4205 2775
rect 4235 2795 4240 2800
rect 4380 2800 4420 2805
rect 4380 2795 4385 2800
rect 4235 2775 4385 2795
rect 4235 2770 4240 2775
rect 4200 2765 4240 2770
rect 4380 2770 4385 2775
rect 4415 2795 4420 2800
rect 4560 2800 4600 2805
rect 4560 2795 4565 2800
rect 4415 2775 4565 2795
rect 4415 2770 4420 2775
rect 4380 2765 4420 2770
rect 4560 2770 4565 2775
rect 4595 2795 4600 2800
rect 4740 2800 4780 2805
rect 4740 2795 4745 2800
rect 4595 2775 4745 2795
rect 4595 2770 4600 2775
rect 4560 2765 4600 2770
rect 4740 2770 4745 2775
rect 4775 2795 4780 2800
rect 4920 2800 4960 2805
rect 4920 2795 4925 2800
rect 4775 2775 4925 2795
rect 4775 2770 4780 2775
rect 4740 2765 4780 2770
rect 4920 2770 4925 2775
rect 4955 2770 4960 2800
rect 4920 2765 4960 2770
rect 2570 2755 2610 2760
rect 1245 2745 1285 2750
rect 1245 2715 1250 2745
rect 1280 2740 1285 2745
rect 2150 2745 2190 2750
rect 2150 2740 2155 2745
rect 1280 2720 2155 2740
rect 1280 2715 1285 2720
rect 1245 2710 1285 2715
rect 2150 2715 2155 2720
rect 2185 2715 2190 2745
rect 2150 2710 2190 2715
rect 3030 2430 3070 2435
rect 2940 2425 2980 2430
rect 2570 2395 2610 2400
rect 2570 2365 2575 2395
rect 2605 2390 2610 2395
rect 2940 2395 2945 2425
rect 2975 2395 2980 2425
rect 3030 2400 3035 2430
rect 3065 2425 3070 2430
rect 3750 2430 3790 2435
rect 3750 2425 3755 2430
rect 3065 2405 3755 2425
rect 3065 2400 3070 2405
rect 3030 2395 3070 2400
rect 3750 2400 3755 2405
rect 3785 2425 3790 2430
rect 4100 2430 4140 2435
rect 4100 2425 4105 2430
rect 3785 2405 4105 2425
rect 3785 2400 3790 2405
rect 3750 2395 3790 2400
rect 4100 2400 4105 2405
rect 4135 2425 4140 2430
rect 4830 2430 4870 2435
rect 4830 2425 4835 2430
rect 4135 2405 4835 2425
rect 4135 2400 4140 2405
rect 4100 2395 4140 2400
rect 4830 2400 4835 2405
rect 4865 2400 4870 2430
rect 4830 2395 4870 2400
rect 2940 2390 2980 2395
rect 2605 2370 2980 2390
rect 3210 2385 3250 2390
rect 2605 2365 2610 2370
rect 2570 2360 2610 2365
rect 3210 2355 3215 2385
rect 3245 2380 3250 2385
rect 3570 2385 3610 2390
rect 3570 2380 3575 2385
rect 3245 2360 3575 2380
rect 3245 2355 3250 2360
rect 3210 2350 3250 2355
rect 3570 2355 3575 2360
rect 3605 2380 3610 2385
rect 4290 2385 4330 2390
rect 4290 2380 4295 2385
rect 3605 2360 4295 2380
rect 3605 2355 3610 2360
rect 3570 2350 3610 2355
rect 4290 2355 4295 2360
rect 4325 2380 4330 2385
rect 4650 2385 4690 2390
rect 4650 2380 4655 2385
rect 4325 2360 4655 2380
rect 4325 2355 4330 2360
rect 4290 2350 4330 2355
rect 4650 2355 4655 2360
rect 4685 2355 4690 2385
rect 4650 2350 4690 2355
rect 2685 2340 2725 2345
rect 2685 2310 2690 2340
rect 2720 2335 2725 2340
rect 3390 2340 3430 2345
rect 3390 2335 3395 2340
rect 2720 2315 3395 2335
rect 2720 2310 2725 2315
rect 2685 2305 2725 2310
rect 3390 2310 3395 2315
rect 3425 2335 3430 2340
rect 4470 2340 4510 2345
rect 4470 2335 4475 2340
rect 3425 2315 4475 2335
rect 3425 2310 3430 2315
rect 3390 2305 3430 2310
rect 4470 2310 4475 2315
rect 4505 2335 4510 2340
rect 5200 2340 5240 2345
rect 5200 2335 5205 2340
rect 4505 2315 5205 2335
rect 4505 2310 4510 2315
rect 4470 2305 4510 2310
rect 5200 2310 5205 2315
rect 5235 2310 5240 2340
rect 5200 2305 5240 2310
rect 2425 2245 2465 2250
rect 2425 2215 2430 2245
rect 2460 2240 2465 2245
rect 3030 2245 3070 2250
rect 3030 2240 3035 2245
rect 2460 2220 3035 2240
rect 2460 2215 2465 2220
rect 2425 2210 2465 2215
rect 3030 2215 3035 2220
rect 3065 2215 3070 2245
rect 3030 2210 3070 2215
rect 2330 2200 2370 2205
rect 2330 2170 2335 2200
rect 2365 2195 2370 2200
rect 2850 2200 2890 2205
rect 2850 2195 2855 2200
rect 2365 2175 2855 2195
rect 2365 2170 2370 2175
rect 2330 2165 2370 2170
rect 2850 2170 2855 2175
rect 2885 2195 2890 2200
rect 3930 2200 3970 2205
rect 3930 2195 3935 2200
rect 2885 2175 3935 2195
rect 2885 2170 2890 2175
rect 2850 2165 2890 2170
rect 3930 2170 3935 2175
rect 3965 2195 3970 2200
rect 5010 2200 5050 2205
rect 5010 2195 5015 2200
rect 3965 2175 5015 2195
rect 3965 2170 3970 2175
rect 3930 2165 3970 2170
rect 5010 2170 5015 2175
rect 5045 2170 5050 2200
rect 5010 2165 5050 2170
rect 2380 2150 2420 2155
rect 2380 2120 2385 2150
rect 2415 2145 2420 2150
rect 3210 2150 3250 2155
rect 3210 2145 3215 2150
rect 2415 2125 3215 2145
rect 2415 2120 2420 2125
rect 2380 2115 2420 2120
rect 3210 2120 3215 2125
rect 3245 2120 3250 2150
rect 3210 2115 3250 2120
rect 4025 2145 4065 2150
rect 4025 2115 4030 2145
rect 4060 2140 4065 2145
rect 5245 2145 5285 2150
rect 5245 2140 5250 2145
rect 4060 2120 5250 2140
rect 4060 2115 4065 2120
rect 4025 2110 4065 2115
rect 5245 2115 5250 2120
rect 5280 2115 5285 2145
rect 5245 2110 5285 2115
rect 2815 2095 2855 2100
rect 2815 2065 2820 2095
rect 2850 2090 2855 2095
rect 2935 2095 2975 2100
rect 2935 2090 2940 2095
rect 2850 2070 2940 2090
rect 2850 2065 2855 2070
rect 2815 2060 2855 2065
rect 2935 2065 2940 2070
rect 2970 2090 2975 2095
rect 3055 2095 3095 2100
rect 3055 2090 3060 2095
rect 2970 2070 3060 2090
rect 2970 2065 2975 2070
rect 2935 2060 2975 2065
rect 3055 2065 3060 2070
rect 3090 2090 3095 2095
rect 3175 2095 3215 2100
rect 3175 2090 3180 2095
rect 3090 2070 3180 2090
rect 3090 2065 3095 2070
rect 3055 2060 3095 2065
rect 3175 2065 3180 2070
rect 3210 2090 3215 2095
rect 3295 2095 3335 2100
rect 3295 2090 3300 2095
rect 3210 2070 3300 2090
rect 3210 2065 3215 2070
rect 3175 2060 3215 2065
rect 3295 2065 3300 2070
rect 3330 2090 3335 2095
rect 3415 2095 3455 2100
rect 3415 2090 3420 2095
rect 3330 2070 3420 2090
rect 3330 2065 3335 2070
rect 3295 2060 3335 2065
rect 3415 2065 3420 2070
rect 3450 2090 3455 2095
rect 3535 2095 3575 2100
rect 3535 2090 3540 2095
rect 3450 2070 3540 2090
rect 3450 2065 3455 2070
rect 3415 2060 3455 2065
rect 3535 2065 3540 2070
rect 3570 2090 3575 2095
rect 3655 2095 3695 2100
rect 3655 2090 3660 2095
rect 3570 2070 3660 2090
rect 3570 2065 3575 2070
rect 3535 2060 3575 2065
rect 3655 2065 3660 2070
rect 3690 2090 3695 2095
rect 3775 2095 3815 2100
rect 3775 2090 3780 2095
rect 3690 2070 3780 2090
rect 3690 2065 3695 2070
rect 3655 2060 3695 2065
rect 3775 2065 3780 2070
rect 3810 2065 3815 2095
rect 3775 2060 3815 2065
rect 4085 2095 4125 2100
rect 4085 2065 4090 2095
rect 4120 2090 4125 2095
rect 4205 2095 4245 2100
rect 4205 2090 4210 2095
rect 4120 2070 4210 2090
rect 4120 2065 4125 2070
rect 4085 2060 4125 2065
rect 4205 2065 4210 2070
rect 4240 2090 4245 2095
rect 4325 2095 4365 2100
rect 4325 2090 4330 2095
rect 4240 2070 4330 2090
rect 4240 2065 4245 2070
rect 4205 2060 4245 2065
rect 4325 2065 4330 2070
rect 4360 2090 4365 2095
rect 4445 2095 4485 2100
rect 4445 2090 4450 2095
rect 4360 2070 4450 2090
rect 4360 2065 4365 2070
rect 4325 2060 4365 2065
rect 4445 2065 4450 2070
rect 4480 2090 4485 2095
rect 4565 2095 4605 2100
rect 4565 2090 4570 2095
rect 4480 2070 4570 2090
rect 4480 2065 4485 2070
rect 4445 2060 4485 2065
rect 4565 2065 4570 2070
rect 4600 2090 4605 2095
rect 4685 2095 4725 2100
rect 4685 2090 4690 2095
rect 4600 2070 4690 2090
rect 4600 2065 4605 2070
rect 4565 2060 4605 2065
rect 4685 2065 4690 2070
rect 4720 2090 4725 2095
rect 4805 2095 4845 2100
rect 4805 2090 4810 2095
rect 4720 2070 4810 2090
rect 4720 2065 4725 2070
rect 4685 2060 4725 2065
rect 4805 2065 4810 2070
rect 4840 2090 4845 2095
rect 4925 2095 4965 2100
rect 4925 2090 4930 2095
rect 4840 2070 4930 2090
rect 4840 2065 4845 2070
rect 4805 2060 4845 2065
rect 4925 2065 4930 2070
rect 4960 2090 4965 2095
rect 5045 2095 5085 2100
rect 5045 2090 5050 2095
rect 4960 2070 5050 2090
rect 4960 2065 4965 2070
rect 4925 2060 4965 2065
rect 5045 2065 5050 2070
rect 5080 2065 5085 2095
rect 5045 2060 5085 2065
rect 2570 2050 2610 2055
rect 2570 2020 2575 2050
rect 2605 2020 2610 2050
rect 2570 2015 2610 2020
rect 2755 2050 2795 2055
rect 2755 2020 2760 2050
rect 2790 2045 2795 2050
rect 3115 2050 3155 2055
rect 3115 2045 3120 2050
rect 2790 2025 3120 2045
rect 2790 2020 2795 2025
rect 2755 2015 2795 2020
rect 3115 2020 3120 2025
rect 3150 2045 3155 2050
rect 3475 2050 3515 2055
rect 3475 2045 3480 2050
rect 3150 2025 3480 2045
rect 3150 2020 3155 2025
rect 3115 2015 3155 2020
rect 3475 2020 3480 2025
rect 3510 2045 3515 2050
rect 3835 2050 3875 2055
rect 3835 2045 3840 2050
rect 3510 2025 3840 2045
rect 3510 2020 3515 2025
rect 3475 2015 3515 2020
rect 3835 2020 3840 2025
rect 3870 2020 3875 2050
rect 3835 2015 3875 2020
rect 4025 2050 4065 2055
rect 4025 2020 4030 2050
rect 4060 2045 4065 2050
rect 4385 2050 4425 2055
rect 4385 2045 4390 2050
rect 4060 2025 4390 2045
rect 4060 2020 4065 2025
rect 4025 2015 4065 2020
rect 4385 2020 4390 2025
rect 4420 2045 4425 2050
rect 4745 2050 4785 2055
rect 4745 2045 4750 2050
rect 4420 2025 4750 2045
rect 4420 2020 4425 2025
rect 4385 2015 4425 2020
rect 4745 2020 4750 2025
rect 4780 2045 4785 2050
rect 5105 2050 5145 2055
rect 5105 2045 5110 2050
rect 4780 2025 5110 2045
rect 4780 2020 4785 2025
rect 4745 2015 4785 2020
rect 5105 2020 5110 2025
rect 5140 2020 5145 2050
rect 5105 2015 5145 2020
rect 2875 1880 2915 1885
rect 2875 1850 2880 1880
rect 2910 1875 2915 1880
rect 2995 1875 3035 1885
rect 3235 1880 3275 1885
rect 3235 1875 3240 1880
rect 2910 1855 3240 1875
rect 2910 1850 2915 1855
rect 2875 1845 2915 1850
rect 2995 1845 3035 1855
rect 3235 1850 3240 1855
rect 3270 1875 3275 1880
rect 3355 1875 3395 1885
rect 3595 1880 3635 1885
rect 3595 1875 3600 1880
rect 3270 1855 3600 1875
rect 3270 1850 3275 1855
rect 3235 1845 3275 1850
rect 3355 1845 3395 1855
rect 3595 1850 3600 1855
rect 3630 1850 3635 1880
rect 3595 1845 3635 1850
rect 3715 1845 3755 1885
rect 4145 1845 4185 1885
rect 4265 1880 4305 1885
rect 4265 1850 4270 1880
rect 4300 1875 4305 1880
rect 4505 1875 4545 1885
rect 4625 1880 4665 1885
rect 4625 1875 4630 1880
rect 4300 1855 4630 1875
rect 4300 1850 4305 1855
rect 4265 1845 4305 1850
rect 4505 1845 4545 1855
rect 4625 1850 4630 1855
rect 4660 1875 4665 1880
rect 4865 1875 4905 1885
rect 4985 1880 5025 1885
rect 4985 1875 4990 1880
rect 4660 1855 4990 1875
rect 4660 1850 4665 1855
rect 4625 1845 4665 1850
rect 4865 1845 4905 1855
rect 4985 1850 4990 1855
rect 5020 1875 5025 1880
rect 5020 1855 5115 1875
rect 5020 1850 5025 1855
rect 4985 1845 5025 1850
rect 2470 1820 2510 1825
rect 2470 1790 2475 1820
rect 2505 1815 2510 1820
rect 2785 1820 2825 1825
rect 2785 1815 2790 1820
rect 2505 1795 2790 1815
rect 2505 1790 2510 1795
rect 2470 1785 2510 1790
rect 2785 1790 2790 1795
rect 2820 1815 2825 1820
rect 2995 1820 3035 1825
rect 2995 1815 3000 1820
rect 2820 1795 3000 1815
rect 2820 1790 2825 1795
rect 2785 1785 2825 1790
rect 2995 1790 3000 1795
rect 3030 1815 3035 1820
rect 3115 1820 3155 1825
rect 3115 1815 3120 1820
rect 3030 1795 3120 1815
rect 3030 1790 3035 1795
rect 2995 1785 3035 1790
rect 3115 1790 3120 1795
rect 3150 1815 3155 1820
rect 3355 1820 3395 1825
rect 3355 1815 3360 1820
rect 3150 1795 3360 1815
rect 3150 1790 3155 1795
rect 3115 1785 3155 1790
rect 3355 1790 3360 1795
rect 3390 1815 3395 1820
rect 3475 1820 3515 1825
rect 3475 1815 3480 1820
rect 3390 1795 3480 1815
rect 3390 1790 3395 1795
rect 3355 1785 3395 1790
rect 3475 1790 3480 1795
rect 3510 1815 3515 1820
rect 3715 1820 3755 1825
rect 3715 1815 3720 1820
rect 3510 1795 3720 1815
rect 3510 1790 3515 1795
rect 3475 1785 3515 1790
rect 3715 1790 3720 1795
rect 3750 1815 3755 1820
rect 3805 1820 3845 1825
rect 3805 1815 3810 1820
rect 3750 1795 3810 1815
rect 3750 1790 3755 1795
rect 3715 1785 3755 1790
rect 3805 1790 3810 1795
rect 3840 1790 3845 1820
rect 3805 1785 3845 1790
rect 4055 1820 4095 1825
rect 4055 1790 4060 1820
rect 4090 1815 4095 1820
rect 4145 1820 4185 1825
rect 4145 1815 4150 1820
rect 4090 1795 4150 1815
rect 4090 1790 4095 1795
rect 4055 1785 4095 1790
rect 4145 1790 4150 1795
rect 4180 1815 4185 1820
rect 4385 1820 4425 1825
rect 4385 1815 4390 1820
rect 4180 1795 4390 1815
rect 4180 1790 4185 1795
rect 4145 1785 4185 1790
rect 4385 1790 4390 1795
rect 4420 1815 4425 1820
rect 4505 1820 4545 1825
rect 4505 1815 4510 1820
rect 4420 1795 4510 1815
rect 4420 1790 4425 1795
rect 4385 1785 4425 1790
rect 4505 1790 4510 1795
rect 4540 1815 4545 1820
rect 4745 1820 4785 1825
rect 4745 1815 4750 1820
rect 4540 1795 4750 1815
rect 4540 1790 4545 1795
rect 4505 1785 4545 1790
rect 4745 1790 4750 1795
rect 4780 1815 4785 1820
rect 4865 1820 4905 1825
rect 4865 1815 4870 1820
rect 4780 1795 4870 1815
rect 4780 1790 4785 1795
rect 4745 1785 4785 1790
rect 4865 1790 4870 1795
rect 4900 1815 4905 1820
rect 5075 1820 5115 1825
rect 5075 1815 5080 1820
rect 4900 1795 5080 1815
rect 4900 1790 4905 1795
rect 4865 1785 4905 1790
rect 5075 1790 5080 1795
rect 5110 1815 5115 1820
rect 5290 1820 5330 1825
rect 5290 1815 5295 1820
rect 5110 1795 5295 1815
rect 5110 1790 5115 1795
rect 5075 1785 5115 1790
rect 5290 1790 5295 1795
rect 5325 1790 5330 1820
rect 5290 1785 5330 1790
rect 2425 1760 2465 1765
rect 2425 1730 2430 1760
rect 2460 1755 2465 1760
rect 2515 1760 2555 1765
rect 2515 1755 2520 1760
rect 2460 1735 2520 1755
rect 2460 1730 2465 1735
rect 2425 1725 2465 1730
rect 2515 1730 2520 1735
rect 2550 1755 2555 1760
rect 2625 1760 2665 1765
rect 2625 1755 2630 1760
rect 2550 1735 2630 1755
rect 2550 1730 2555 1735
rect 2515 1725 2555 1730
rect 2625 1730 2630 1735
rect 2660 1755 2665 1760
rect 3175 1760 3215 1765
rect 3175 1755 3180 1760
rect 2660 1735 3180 1755
rect 2660 1730 2665 1735
rect 2625 1725 2665 1730
rect 3175 1730 3180 1735
rect 3210 1730 3215 1760
rect 3175 1725 3215 1730
rect 3235 1760 3275 1765
rect 3235 1730 3240 1760
rect 3270 1755 3275 1760
rect 3475 1760 3515 1765
rect 3475 1755 3480 1760
rect 3270 1735 3480 1755
rect 3270 1730 3275 1735
rect 3235 1725 3275 1730
rect 3475 1730 3480 1735
rect 3510 1755 3515 1760
rect 3715 1760 3755 1765
rect 3715 1755 3720 1760
rect 3510 1735 3720 1755
rect 3510 1730 3515 1735
rect 3475 1725 3515 1730
rect 3715 1730 3720 1735
rect 3750 1730 3755 1760
rect 3715 1725 3755 1730
rect 4145 1760 4185 1765
rect 4145 1730 4150 1760
rect 4180 1755 4185 1760
rect 4385 1760 4425 1765
rect 4385 1755 4390 1760
rect 4180 1735 4390 1755
rect 4180 1730 4185 1735
rect 4145 1725 4185 1730
rect 4385 1730 4390 1735
rect 4420 1755 4425 1760
rect 4625 1760 4665 1765
rect 4625 1755 4630 1760
rect 4420 1735 4630 1755
rect 4420 1730 4425 1735
rect 4385 1725 4425 1730
rect 4625 1730 4630 1735
rect 4660 1730 4665 1760
rect 4625 1725 4665 1730
rect 4685 1760 4725 1765
rect 4685 1730 4690 1760
rect 4720 1755 4725 1760
rect 5200 1760 5240 1765
rect 5200 1755 5205 1760
rect 4720 1735 5205 1755
rect 4720 1730 4725 1735
rect 4685 1725 4725 1730
rect 5200 1730 5205 1735
rect 5235 1730 5240 1760
rect 5200 1725 5240 1730
rect -110 1720 -70 1725
rect -110 1690 -105 1720
rect -75 1690 -70 1720
rect -110 1685 -70 1690
rect -45 1720 -5 1725
rect -45 1690 -40 1720
rect -10 1690 -5 1720
rect 3115 1715 3155 1720
rect -45 1685 -5 1690
rect 1265 1710 1305 1715
rect 1265 1680 1270 1710
rect 1300 1705 1305 1710
rect 2150 1710 2190 1715
rect 2150 1705 2155 1710
rect 1300 1685 2155 1705
rect 1300 1680 1305 1685
rect 1265 1675 1305 1680
rect 2150 1680 2155 1685
rect 2185 1680 2190 1710
rect 3115 1685 3120 1715
rect 3150 1710 3155 1715
rect 3355 1715 3395 1720
rect 3355 1710 3360 1715
rect 3150 1690 3360 1710
rect 3150 1685 3155 1690
rect 3115 1680 3155 1685
rect 3355 1685 3360 1690
rect 3390 1710 3395 1715
rect 3595 1715 3635 1720
rect 3595 1710 3600 1715
rect 3390 1690 3600 1710
rect 3390 1685 3395 1690
rect 3355 1680 3395 1685
rect 3595 1685 3600 1690
rect 3630 1685 3635 1715
rect 3595 1680 3635 1685
rect 4265 1715 4305 1720
rect 4265 1685 4270 1715
rect 4300 1710 4305 1715
rect 4505 1715 4545 1720
rect 4505 1710 4510 1715
rect 4300 1690 4510 1710
rect 4300 1685 4305 1690
rect 4265 1680 4305 1685
rect 4505 1685 4510 1690
rect 4540 1710 4545 1715
rect 4745 1715 4785 1720
rect 4745 1710 4750 1715
rect 4540 1690 4750 1710
rect 4540 1685 4545 1690
rect 4505 1680 4545 1685
rect 4745 1685 4750 1690
rect 4780 1685 4785 1715
rect 4745 1680 4785 1685
rect 2150 1675 2190 1680
rect 2380 1665 2420 1670
rect 2380 1635 2385 1665
rect 2415 1660 2420 1665
rect 2570 1665 2610 1670
rect 2570 1660 2575 1665
rect 2415 1640 2575 1660
rect 2415 1635 2420 1640
rect 2380 1630 2420 1635
rect 2570 1635 2575 1640
rect 2605 1635 2610 1665
rect 2570 1630 2610 1635
rect 2330 1595 2370 1600
rect 2330 1565 2335 1595
rect 2365 1590 2370 1595
rect 3115 1595 3155 1600
rect 3115 1590 3120 1595
rect 2365 1570 3120 1590
rect 2365 1565 2370 1570
rect 2330 1560 2370 1565
rect 3115 1565 3120 1570
rect 3150 1565 3155 1595
rect 3115 1560 3155 1565
rect 4745 1595 4785 1600
rect 4745 1565 4750 1595
rect 4780 1590 4785 1595
rect 5340 1595 5380 1600
rect 5340 1590 5345 1595
rect 4780 1570 5345 1590
rect 4780 1565 4785 1570
rect 4745 1560 4785 1565
rect 5340 1565 5345 1570
rect 5375 1565 5380 1595
rect 5340 1560 5380 1565
rect 2785 1545 2825 1550
rect 2785 1515 2790 1545
rect 2820 1540 2825 1545
rect 3175 1545 3215 1550
rect 3175 1540 3180 1545
rect 2820 1520 3180 1540
rect 2820 1515 2825 1520
rect 2785 1510 2825 1515
rect 3175 1515 3180 1520
rect 3210 1540 3215 1545
rect 3295 1545 3335 1550
rect 3295 1540 3300 1545
rect 3210 1520 3300 1540
rect 3210 1515 3215 1520
rect 3175 1510 3215 1515
rect 3295 1515 3300 1520
rect 3330 1540 3335 1545
rect 3415 1545 3455 1550
rect 3415 1540 3420 1545
rect 3330 1520 3420 1540
rect 3330 1515 3335 1520
rect 3295 1510 3335 1515
rect 3415 1515 3420 1520
rect 3450 1540 3455 1545
rect 3535 1545 3575 1550
rect 3535 1540 3540 1545
rect 3450 1520 3540 1540
rect 3450 1515 3455 1520
rect 3415 1510 3455 1515
rect 3535 1515 3540 1520
rect 3570 1540 3575 1545
rect 3655 1545 3695 1550
rect 3655 1540 3660 1545
rect 3570 1520 3660 1540
rect 3570 1515 3575 1520
rect 3535 1510 3575 1515
rect 3655 1515 3660 1520
rect 3690 1515 3695 1545
rect 3655 1510 3695 1515
rect 4205 1545 4245 1550
rect 4205 1515 4210 1545
rect 4240 1540 4245 1545
rect 4325 1545 4365 1550
rect 4325 1540 4330 1545
rect 4240 1520 4330 1540
rect 4240 1515 4245 1520
rect 4205 1510 4245 1515
rect 4325 1515 4330 1520
rect 4360 1540 4365 1545
rect 4445 1545 4485 1550
rect 4445 1540 4450 1545
rect 4360 1520 4450 1540
rect 4360 1515 4365 1520
rect 4325 1510 4365 1515
rect 4445 1515 4450 1520
rect 4480 1540 4485 1545
rect 4565 1545 4605 1550
rect 4565 1540 4570 1545
rect 4480 1520 4570 1540
rect 4480 1515 4485 1520
rect 4445 1510 4485 1515
rect 4565 1515 4570 1520
rect 4600 1540 4605 1545
rect 4685 1545 4725 1550
rect 4685 1540 4690 1545
rect 4600 1520 4690 1540
rect 4600 1515 4605 1520
rect 4565 1510 4605 1515
rect 4685 1515 4690 1520
rect 4720 1540 4725 1545
rect 5075 1545 5115 1550
rect 5075 1540 5080 1545
rect 4720 1520 5080 1540
rect 4720 1515 4725 1520
rect 4685 1510 4725 1515
rect 5075 1515 5080 1520
rect 5110 1515 5115 1545
rect 5075 1510 5115 1515
rect 2890 1165 2930 1170
rect 2890 1135 2895 1165
rect 2925 1160 2930 1165
rect 2970 1165 3010 1170
rect 2970 1160 2975 1165
rect 2925 1140 2975 1160
rect 2925 1135 2930 1140
rect 2890 1130 2930 1135
rect 2970 1135 2975 1140
rect 3005 1160 3010 1165
rect 3050 1165 3090 1170
rect 3050 1160 3055 1165
rect 3005 1140 3055 1160
rect 3005 1135 3010 1140
rect 2970 1130 3010 1135
rect 3050 1135 3055 1140
rect 3085 1160 3090 1165
rect 3130 1165 3170 1170
rect 3130 1160 3135 1165
rect 3085 1140 3135 1160
rect 3085 1135 3090 1140
rect 3050 1130 3090 1135
rect 3130 1135 3135 1140
rect 3165 1160 3170 1165
rect 3210 1165 3250 1170
rect 3210 1160 3215 1165
rect 3165 1140 3215 1160
rect 3165 1135 3170 1140
rect 3130 1130 3170 1135
rect 3210 1135 3215 1140
rect 3245 1160 3250 1165
rect 3290 1165 3330 1170
rect 3290 1160 3295 1165
rect 3245 1140 3295 1160
rect 3245 1135 3250 1140
rect 3210 1130 3250 1135
rect 3290 1135 3295 1140
rect 3325 1160 3330 1165
rect 3370 1165 3410 1170
rect 3370 1160 3375 1165
rect 3325 1140 3375 1160
rect 3325 1135 3330 1140
rect 3290 1130 3330 1135
rect 3370 1135 3375 1140
rect 3405 1160 3410 1165
rect 3450 1165 3490 1170
rect 3450 1160 3455 1165
rect 3405 1140 3455 1160
rect 3405 1135 3410 1140
rect 3370 1130 3410 1135
rect 3450 1135 3455 1140
rect 3485 1160 3490 1165
rect 3530 1165 3570 1170
rect 3530 1160 3535 1165
rect 3485 1140 3535 1160
rect 3485 1135 3490 1140
rect 3450 1130 3490 1135
rect 3530 1135 3535 1140
rect 3565 1160 3570 1165
rect 3610 1165 3650 1170
rect 3610 1160 3615 1165
rect 3565 1140 3615 1160
rect 3565 1135 3570 1140
rect 3530 1130 3570 1135
rect 3610 1135 3615 1140
rect 3645 1160 3650 1165
rect 3690 1165 3730 1170
rect 3690 1160 3695 1165
rect 3645 1140 3695 1160
rect 3645 1135 3650 1140
rect 3610 1130 3650 1135
rect 3690 1135 3695 1140
rect 3725 1160 3730 1165
rect 3770 1165 3810 1170
rect 3770 1160 3775 1165
rect 3725 1140 3775 1160
rect 3725 1135 3730 1140
rect 3690 1130 3730 1135
rect 3770 1135 3775 1140
rect 3805 1160 3810 1165
rect 3850 1165 3890 1170
rect 3850 1160 3855 1165
rect 3805 1140 3855 1160
rect 3805 1135 3810 1140
rect 3770 1130 3810 1135
rect 3850 1135 3855 1140
rect 3885 1135 3890 1165
rect 3850 1130 3890 1135
rect 3930 1165 3970 1170
rect 3930 1135 3935 1165
rect 3965 1160 3970 1165
rect 4010 1165 4050 1170
rect 4010 1160 4015 1165
rect 3965 1140 4015 1160
rect 3965 1135 3970 1140
rect 3930 1130 3970 1135
rect 4010 1135 4015 1140
rect 4045 1160 4050 1165
rect 4090 1165 4130 1170
rect 4090 1160 4095 1165
rect 4045 1140 4095 1160
rect 4045 1135 4050 1140
rect 4010 1130 4050 1135
rect 4090 1135 4095 1140
rect 4125 1160 4130 1165
rect 4170 1165 4210 1170
rect 4170 1160 4175 1165
rect 4125 1140 4175 1160
rect 4125 1135 4130 1140
rect 4090 1130 4130 1135
rect 4170 1135 4175 1140
rect 4205 1160 4210 1165
rect 4250 1165 4290 1170
rect 4250 1160 4255 1165
rect 4205 1140 4255 1160
rect 4205 1135 4210 1140
rect 4170 1130 4210 1135
rect 4250 1135 4255 1140
rect 4285 1160 4290 1165
rect 4330 1165 4370 1170
rect 4330 1160 4335 1165
rect 4285 1140 4335 1160
rect 4285 1135 4290 1140
rect 4250 1130 4290 1135
rect 4330 1135 4335 1140
rect 4365 1160 4370 1165
rect 4410 1165 4450 1170
rect 4410 1160 4415 1165
rect 4365 1140 4415 1160
rect 4365 1135 4370 1140
rect 4330 1130 4370 1135
rect 4410 1135 4415 1140
rect 4445 1160 4450 1165
rect 4490 1165 4530 1170
rect 4490 1160 4495 1165
rect 4445 1140 4495 1160
rect 4445 1135 4450 1140
rect 4410 1130 4450 1135
rect 4490 1135 4495 1140
rect 4525 1160 4530 1165
rect 4570 1165 4610 1170
rect 4570 1160 4575 1165
rect 4525 1140 4575 1160
rect 4525 1135 4530 1140
rect 4490 1130 4530 1135
rect 4570 1135 4575 1140
rect 4605 1160 4610 1165
rect 4650 1165 4690 1170
rect 4650 1160 4655 1165
rect 4605 1140 4655 1160
rect 4605 1135 4610 1140
rect 4570 1130 4610 1135
rect 4650 1135 4655 1140
rect 4685 1160 4690 1165
rect 4730 1165 4770 1170
rect 4730 1160 4735 1165
rect 4685 1140 4735 1160
rect 4685 1135 4690 1140
rect 4650 1130 4690 1135
rect 4730 1135 4735 1140
rect 4765 1160 4770 1165
rect 4810 1165 4850 1170
rect 4810 1160 4815 1165
rect 4765 1140 4815 1160
rect 4765 1135 4770 1140
rect 4730 1130 4770 1135
rect 4810 1135 4815 1140
rect 4845 1160 4850 1165
rect 4890 1165 4930 1170
rect 4890 1160 4895 1165
rect 4845 1140 4895 1160
rect 4845 1135 4850 1140
rect 4810 1130 4850 1135
rect 4890 1135 4895 1140
rect 4925 1135 4930 1165
rect 4890 1130 4930 1135
rect 2570 1080 2610 1085
rect 2570 1050 2575 1080
rect 2605 1075 2610 1080
rect 2850 1080 2890 1085
rect 2850 1075 2855 1080
rect 2605 1055 2855 1075
rect 2605 1050 2610 1055
rect 2570 1045 2610 1050
rect 2850 1050 2855 1055
rect 2885 1050 2890 1080
rect 2850 1045 2890 1050
rect 2175 1030 2215 1035
rect 2175 1000 2180 1030
rect 2210 1025 2215 1030
rect 2425 1030 2465 1035
rect 2425 1025 2430 1030
rect 2210 1005 2430 1025
rect 2210 1000 2215 1005
rect 2175 995 2215 1000
rect 2425 1000 2430 1005
rect 2460 1000 2465 1030
rect 2425 995 2465 1000
rect -195 550 -155 555
rect -195 520 -190 550
rect -160 520 -155 550
rect -195 515 -155 520
<< via2 >>
rect -190 4975 -160 5005
rect 5485 4975 5515 5005
rect 4445 3465 4475 3495
rect 945 3415 975 3445
rect 1645 3415 1675 3445
rect 5145 3415 5175 3445
rect 2695 3360 2725 3390
rect 3395 3305 3425 3335
rect -105 1690 -75 1720
rect -190 520 -160 550
<< metal3 >>
rect -200 5010 -150 5015
rect -200 4970 -195 5010
rect -155 4970 -150 5010
rect -200 4965 -150 4970
rect 5475 5010 5525 5015
rect 5475 4970 5480 5010
rect 5520 4970 5525 5010
rect 5475 4965 5525 4970
rect -195 560 -155 4965
rect -115 4925 -65 4930
rect -115 4885 -110 4925
rect -70 4885 -65 4925
rect -115 4880 -65 4885
rect 5390 4925 5440 4930
rect 5390 4885 5395 4925
rect 5435 4885 5440 4925
rect 5390 4880 5440 4885
rect -110 1720 -70 4880
rect 145 4770 375 4855
rect 495 4770 725 4855
rect 845 4770 1075 4855
rect 1195 4770 1425 4855
rect 1545 4770 1775 4855
rect 145 4720 1775 4770
rect 145 4625 375 4720
rect 495 4625 725 4720
rect 845 4625 1075 4720
rect 1195 4625 1425 4720
rect 1545 4625 1775 4720
rect 1895 4770 2125 4855
rect 2245 4770 2475 4855
rect 2595 4770 2825 4855
rect 2945 4770 3175 4855
rect 3295 4770 3525 4855
rect 1895 4720 3525 4770
rect 1895 4625 2125 4720
rect 2245 4625 2475 4720
rect 2595 4625 2825 4720
rect 2945 4625 3175 4720
rect 3295 4625 3525 4720
rect 3645 4770 3875 4855
rect 3995 4770 4225 4855
rect 4345 4770 4575 4855
rect 4695 4770 4925 4855
rect 5045 4770 5275 4855
rect 3645 4720 5275 4770
rect 3645 4625 3875 4720
rect 3995 4625 4225 4720
rect 4345 4625 4575 4720
rect 4695 4625 4925 4720
rect 5045 4625 5275 4720
rect 935 4505 985 4625
rect 2685 4505 2735 4625
rect 4435 4505 4485 4625
rect 145 4420 375 4505
rect 495 4420 725 4505
rect 845 4420 1075 4505
rect 1195 4420 1425 4505
rect 1545 4420 1775 4505
rect 145 4370 1775 4420
rect 145 4275 375 4370
rect 495 4275 725 4370
rect 845 4275 1075 4370
rect 1195 4275 1425 4370
rect 1545 4275 1775 4370
rect 1895 4420 2125 4505
rect 2245 4420 2475 4505
rect 2595 4420 2825 4505
rect 2945 4420 3175 4505
rect 3295 4420 3525 4505
rect 1895 4370 3525 4420
rect 1895 4275 2125 4370
rect 2245 4275 2475 4370
rect 2595 4275 2825 4370
rect 2945 4275 3175 4370
rect 3295 4275 3525 4370
rect 3645 4420 3875 4505
rect 3995 4420 4225 4505
rect 4345 4420 4575 4505
rect 4695 4420 4925 4505
rect 5045 4420 5275 4505
rect 3645 4370 5275 4420
rect 3645 4275 3875 4370
rect 3995 4275 4225 4370
rect 4345 4275 4575 4370
rect 4695 4275 4925 4370
rect 5045 4275 5275 4370
rect 935 4155 985 4275
rect 2685 4155 2735 4275
rect 4435 4155 4485 4275
rect 145 4070 375 4155
rect 495 4070 725 4155
rect 845 4070 1075 4155
rect 1195 4070 1425 4155
rect 1545 4070 1775 4155
rect 145 4020 1775 4070
rect 145 3925 375 4020
rect 495 3925 725 4020
rect 845 3925 1075 4020
rect 1195 3925 1425 4020
rect 1545 3925 1775 4020
rect 1895 4070 2125 4155
rect 2245 4070 2475 4155
rect 2595 4070 2825 4155
rect 2945 4070 3175 4155
rect 3295 4070 3525 4155
rect 1895 4020 3525 4070
rect 1895 3925 2125 4020
rect 2245 3925 2475 4020
rect 2595 3925 2825 4020
rect 2945 3925 3175 4020
rect 3295 3925 3525 4020
rect 3645 4070 3875 4155
rect 3995 4070 4225 4155
rect 4345 4070 4575 4155
rect 4695 4070 4925 4155
rect 5045 4070 5275 4155
rect 3645 4020 5275 4070
rect 3645 3925 3875 4020
rect 3995 3925 4225 4020
rect 4345 3925 4575 4020
rect 4695 3925 4925 4020
rect 5045 3925 5275 4020
rect 935 3805 985 3925
rect 2685 3805 2735 3925
rect 4435 3805 4485 3925
rect 145 3720 375 3805
rect 495 3720 725 3805
rect 845 3720 1075 3805
rect 1195 3720 1425 3805
rect 1545 3720 1775 3805
rect 145 3670 1775 3720
rect 145 3575 375 3670
rect 495 3575 725 3670
rect 845 3575 1075 3670
rect 1195 3575 1425 3670
rect 1545 3575 1775 3670
rect 1895 3720 2125 3805
rect 2245 3720 2475 3805
rect 2595 3720 2825 3805
rect 2945 3720 3175 3805
rect 3295 3720 3525 3805
rect 1895 3670 3525 3720
rect 1895 3575 2125 3670
rect 2245 3575 2475 3670
rect 2595 3575 2825 3670
rect 2945 3575 3175 3670
rect 3295 3575 3525 3670
rect 3645 3720 3875 3805
rect 3995 3720 4225 3805
rect 4345 3720 4575 3805
rect 4695 3720 4925 3805
rect 5045 3720 5275 3805
rect 3645 3670 5275 3720
rect 3645 3575 3875 3670
rect 3995 3575 4225 3670
rect 4345 3575 4575 3670
rect 4695 3575 4925 3670
rect 5045 3575 5275 3670
rect 940 3445 980 3575
rect 940 3415 945 3445
rect 975 3415 980 3445
rect 940 3410 980 3415
rect 1635 3450 1685 3455
rect 1635 3410 1640 3450
rect 1680 3410 1685 3450
rect 1635 3405 1685 3410
rect 2690 3390 2730 3575
rect 4440 3495 4480 3575
rect 4440 3465 4445 3495
rect 4475 3465 4480 3495
rect 4440 3460 4480 3465
rect 5135 3450 5185 3455
rect 5135 3410 5140 3450
rect 5180 3410 5185 3450
rect 5135 3405 5185 3410
rect 2690 3360 2695 3390
rect 2725 3360 2730 3390
rect 2690 3355 2730 3360
rect 3385 3340 3435 3345
rect 3385 3300 3390 3340
rect 3430 3300 3435 3340
rect 3385 3295 3435 3300
rect -110 1690 -105 1720
rect -75 1690 -70 1720
rect -110 640 -70 1690
rect 5395 640 5435 4880
rect -115 635 -65 640
rect -115 595 -110 635
rect -70 595 -65 635
rect -115 590 -65 595
rect 5390 635 5440 640
rect 5390 595 5395 635
rect 5435 595 5440 635
rect 5390 590 5440 595
rect 5480 560 5520 4965
rect -200 555 -150 560
rect -200 515 -195 555
rect -155 515 -150 555
rect -200 510 -150 515
rect 5475 555 5525 560
rect 5475 515 5480 555
rect 5520 515 5525 555
rect 5475 510 5525 515
<< via3 >>
rect -195 5005 -155 5010
rect -195 4975 -190 5005
rect -190 4975 -160 5005
rect -160 4975 -155 5005
rect -195 4970 -155 4975
rect 5480 5005 5520 5010
rect 5480 4975 5485 5005
rect 5485 4975 5515 5005
rect 5515 4975 5520 5005
rect 5480 4970 5520 4975
rect -110 4885 -70 4925
rect 5395 4885 5435 4925
rect 1640 3445 1680 3450
rect 1640 3415 1645 3445
rect 1645 3415 1675 3445
rect 1675 3415 1680 3445
rect 1640 3410 1680 3415
rect 5140 3445 5180 3450
rect 5140 3415 5145 3445
rect 5145 3415 5175 3445
rect 5175 3415 5180 3445
rect 5140 3410 5180 3415
rect 3390 3335 3430 3340
rect 3390 3305 3395 3335
rect 3395 3305 3425 3335
rect 3425 3305 3430 3335
rect 3390 3300 3430 3305
rect -110 595 -70 635
rect 5395 595 5435 635
rect -195 550 -155 555
rect -195 520 -190 550
rect -190 520 -160 550
rect -160 520 -155 550
rect -195 515 -155 520
rect 5480 515 5520 555
<< mimcap >>
rect 160 4765 360 4840
rect 160 4725 240 4765
rect 280 4725 360 4765
rect 160 4640 360 4725
rect 510 4765 710 4840
rect 510 4725 590 4765
rect 630 4725 710 4765
rect 510 4640 710 4725
rect 860 4765 1060 4840
rect 860 4725 940 4765
rect 980 4725 1060 4765
rect 860 4640 1060 4725
rect 1210 4765 1410 4840
rect 1210 4725 1290 4765
rect 1330 4725 1410 4765
rect 1210 4640 1410 4725
rect 1560 4765 1760 4840
rect 1560 4725 1640 4765
rect 1680 4725 1760 4765
rect 1560 4640 1760 4725
rect 1910 4765 2110 4840
rect 1910 4725 1990 4765
rect 2030 4725 2110 4765
rect 1910 4640 2110 4725
rect 2260 4765 2460 4840
rect 2260 4725 2340 4765
rect 2380 4725 2460 4765
rect 2260 4640 2460 4725
rect 2610 4765 2810 4840
rect 2610 4725 2690 4765
rect 2730 4725 2810 4765
rect 2610 4640 2810 4725
rect 2960 4765 3160 4840
rect 2960 4725 3040 4765
rect 3080 4725 3160 4765
rect 2960 4640 3160 4725
rect 3310 4765 3510 4840
rect 3310 4725 3390 4765
rect 3430 4725 3510 4765
rect 3310 4640 3510 4725
rect 3660 4765 3860 4840
rect 3660 4725 3740 4765
rect 3780 4725 3860 4765
rect 3660 4640 3860 4725
rect 4010 4765 4210 4840
rect 4010 4725 4090 4765
rect 4130 4725 4210 4765
rect 4010 4640 4210 4725
rect 4360 4765 4560 4840
rect 4360 4725 4440 4765
rect 4480 4725 4560 4765
rect 4360 4640 4560 4725
rect 4710 4765 4910 4840
rect 4710 4725 4790 4765
rect 4830 4725 4910 4765
rect 4710 4640 4910 4725
rect 5060 4765 5260 4840
rect 5060 4725 5140 4765
rect 5180 4725 5260 4765
rect 5060 4640 5260 4725
rect 160 4415 360 4490
rect 160 4375 240 4415
rect 280 4375 360 4415
rect 160 4290 360 4375
rect 510 4415 710 4490
rect 510 4375 590 4415
rect 630 4375 710 4415
rect 510 4290 710 4375
rect 860 4415 1060 4490
rect 860 4375 940 4415
rect 980 4375 1060 4415
rect 860 4290 1060 4375
rect 1210 4415 1410 4490
rect 1210 4375 1290 4415
rect 1330 4375 1410 4415
rect 1210 4290 1410 4375
rect 1560 4415 1760 4490
rect 1560 4375 1640 4415
rect 1680 4375 1760 4415
rect 1560 4290 1760 4375
rect 1910 4415 2110 4490
rect 1910 4375 1990 4415
rect 2030 4375 2110 4415
rect 1910 4290 2110 4375
rect 2260 4415 2460 4490
rect 2260 4375 2340 4415
rect 2380 4375 2460 4415
rect 2260 4290 2460 4375
rect 2610 4415 2810 4490
rect 2610 4375 2690 4415
rect 2730 4375 2810 4415
rect 2610 4290 2810 4375
rect 2960 4415 3160 4490
rect 2960 4375 3040 4415
rect 3080 4375 3160 4415
rect 2960 4290 3160 4375
rect 3310 4415 3510 4490
rect 3310 4375 3390 4415
rect 3430 4375 3510 4415
rect 3310 4290 3510 4375
rect 3660 4415 3860 4490
rect 3660 4375 3740 4415
rect 3780 4375 3860 4415
rect 3660 4290 3860 4375
rect 4010 4415 4210 4490
rect 4010 4375 4090 4415
rect 4130 4375 4210 4415
rect 4010 4290 4210 4375
rect 4360 4415 4560 4490
rect 4360 4375 4440 4415
rect 4480 4375 4560 4415
rect 4360 4290 4560 4375
rect 4710 4415 4910 4490
rect 4710 4375 4790 4415
rect 4830 4375 4910 4415
rect 4710 4290 4910 4375
rect 5060 4415 5260 4490
rect 5060 4375 5140 4415
rect 5180 4375 5260 4415
rect 5060 4290 5260 4375
rect 160 4065 360 4140
rect 160 4025 240 4065
rect 280 4025 360 4065
rect 160 3940 360 4025
rect 510 4065 710 4140
rect 510 4025 590 4065
rect 630 4025 710 4065
rect 510 3940 710 4025
rect 860 4065 1060 4140
rect 860 4025 940 4065
rect 980 4025 1060 4065
rect 860 3940 1060 4025
rect 1210 4065 1410 4140
rect 1210 4025 1290 4065
rect 1330 4025 1410 4065
rect 1210 3940 1410 4025
rect 1560 4065 1760 4140
rect 1560 4025 1640 4065
rect 1680 4025 1760 4065
rect 1560 3940 1760 4025
rect 1910 4065 2110 4140
rect 1910 4025 1990 4065
rect 2030 4025 2110 4065
rect 1910 3940 2110 4025
rect 2260 4065 2460 4140
rect 2260 4025 2340 4065
rect 2380 4025 2460 4065
rect 2260 3940 2460 4025
rect 2610 4065 2810 4140
rect 2610 4025 2690 4065
rect 2730 4025 2810 4065
rect 2610 3940 2810 4025
rect 2960 4065 3160 4140
rect 2960 4025 3040 4065
rect 3080 4025 3160 4065
rect 2960 3940 3160 4025
rect 3310 4065 3510 4140
rect 3310 4025 3390 4065
rect 3430 4025 3510 4065
rect 3310 3940 3510 4025
rect 3660 4065 3860 4140
rect 3660 4025 3740 4065
rect 3780 4025 3860 4065
rect 3660 3940 3860 4025
rect 4010 4065 4210 4140
rect 4010 4025 4090 4065
rect 4130 4025 4210 4065
rect 4010 3940 4210 4025
rect 4360 4065 4560 4140
rect 4360 4025 4440 4065
rect 4480 4025 4560 4065
rect 4360 3940 4560 4025
rect 4710 4065 4910 4140
rect 4710 4025 4790 4065
rect 4830 4025 4910 4065
rect 4710 3940 4910 4025
rect 5060 4065 5260 4140
rect 5060 4025 5140 4065
rect 5180 4025 5260 4065
rect 5060 3940 5260 4025
rect 160 3715 360 3790
rect 160 3675 240 3715
rect 280 3675 360 3715
rect 160 3590 360 3675
rect 510 3715 710 3790
rect 510 3675 590 3715
rect 630 3675 710 3715
rect 510 3590 710 3675
rect 860 3715 1060 3790
rect 860 3675 940 3715
rect 980 3675 1060 3715
rect 860 3590 1060 3675
rect 1210 3715 1410 3790
rect 1210 3675 1290 3715
rect 1330 3675 1410 3715
rect 1210 3590 1410 3675
rect 1560 3715 1760 3790
rect 1560 3675 1640 3715
rect 1680 3675 1760 3715
rect 1560 3590 1760 3675
rect 1910 3715 2110 3790
rect 1910 3675 1990 3715
rect 2030 3675 2110 3715
rect 1910 3590 2110 3675
rect 2260 3715 2460 3790
rect 2260 3675 2340 3715
rect 2380 3675 2460 3715
rect 2260 3590 2460 3675
rect 2610 3715 2810 3790
rect 2610 3675 2690 3715
rect 2730 3675 2810 3715
rect 2610 3590 2810 3675
rect 2960 3715 3160 3790
rect 2960 3675 3040 3715
rect 3080 3675 3160 3715
rect 2960 3590 3160 3675
rect 3310 3715 3510 3790
rect 3310 3675 3390 3715
rect 3430 3675 3510 3715
rect 3310 3590 3510 3675
rect 3660 3715 3860 3790
rect 3660 3675 3740 3715
rect 3780 3675 3860 3715
rect 3660 3590 3860 3675
rect 4010 3715 4210 3790
rect 4010 3675 4090 3715
rect 4130 3675 4210 3715
rect 4010 3590 4210 3675
rect 4360 3715 4560 3790
rect 4360 3675 4440 3715
rect 4480 3675 4560 3715
rect 4360 3590 4560 3675
rect 4710 3715 4910 3790
rect 4710 3675 4790 3715
rect 4830 3675 4910 3715
rect 4710 3590 4910 3675
rect 5060 3715 5260 3790
rect 5060 3675 5140 3715
rect 5180 3675 5260 3715
rect 5060 3590 5260 3675
<< mimcapcontact >>
rect 240 4725 280 4765
rect 590 4725 630 4765
rect 940 4725 980 4765
rect 1290 4725 1330 4765
rect 1640 4725 1680 4765
rect 1990 4725 2030 4765
rect 2340 4725 2380 4765
rect 2690 4725 2730 4765
rect 3040 4725 3080 4765
rect 3390 4725 3430 4765
rect 3740 4725 3780 4765
rect 4090 4725 4130 4765
rect 4440 4725 4480 4765
rect 4790 4725 4830 4765
rect 5140 4725 5180 4765
rect 240 4375 280 4415
rect 590 4375 630 4415
rect 940 4375 980 4415
rect 1290 4375 1330 4415
rect 1640 4375 1680 4415
rect 1990 4375 2030 4415
rect 2340 4375 2380 4415
rect 2690 4375 2730 4415
rect 3040 4375 3080 4415
rect 3390 4375 3430 4415
rect 3740 4375 3780 4415
rect 4090 4375 4130 4415
rect 4440 4375 4480 4415
rect 4790 4375 4830 4415
rect 5140 4375 5180 4415
rect 240 4025 280 4065
rect 590 4025 630 4065
rect 940 4025 980 4065
rect 1290 4025 1330 4065
rect 1640 4025 1680 4065
rect 1990 4025 2030 4065
rect 2340 4025 2380 4065
rect 2690 4025 2730 4065
rect 3040 4025 3080 4065
rect 3390 4025 3430 4065
rect 3740 4025 3780 4065
rect 4090 4025 4130 4065
rect 4440 4025 4480 4065
rect 4790 4025 4830 4065
rect 5140 4025 5180 4065
rect 240 3675 280 3715
rect 590 3675 630 3715
rect 940 3675 980 3715
rect 1290 3675 1330 3715
rect 1640 3675 1680 3715
rect 1990 3675 2030 3715
rect 2340 3675 2380 3715
rect 2690 3675 2730 3715
rect 3040 3675 3080 3715
rect 3390 3675 3430 3715
rect 3740 3675 3780 3715
rect 4090 3675 4130 3715
rect 4440 3675 4480 3715
rect 4790 3675 4830 3715
rect 5140 3675 5180 3715
<< metal4 >>
rect -200 5010 5525 5015
rect -200 4970 -195 5010
rect -155 4970 5480 5010
rect 5520 4970 5525 5010
rect -200 4965 5525 4970
rect -115 4925 5440 4930
rect -115 4885 -110 4925
rect -70 4885 5395 4925
rect 5435 4885 5440 4925
rect -115 4880 5440 4885
rect 235 4765 1685 4770
rect 235 4725 240 4765
rect 280 4725 590 4765
rect 630 4725 940 4765
rect 980 4725 1290 4765
rect 1330 4725 1640 4765
rect 1680 4725 1685 4765
rect 235 4720 1685 4725
rect 1985 4765 3435 4770
rect 1985 4725 1990 4765
rect 2030 4725 2340 4765
rect 2380 4725 2690 4765
rect 2730 4725 3040 4765
rect 3080 4725 3390 4765
rect 3430 4725 3435 4765
rect 1985 4720 3435 4725
rect 3735 4765 5185 4770
rect 3735 4725 3740 4765
rect 3780 4725 4090 4765
rect 4130 4725 4440 4765
rect 4480 4725 4790 4765
rect 4830 4725 5140 4765
rect 5180 4725 5185 4765
rect 3735 4720 5185 4725
rect 935 4420 985 4720
rect 2685 4420 2735 4720
rect 4435 4420 4485 4720
rect 235 4415 1685 4420
rect 235 4375 240 4415
rect 280 4375 590 4415
rect 630 4375 940 4415
rect 980 4375 1290 4415
rect 1330 4375 1640 4415
rect 1680 4375 1685 4415
rect 235 4370 1685 4375
rect 1985 4415 3435 4420
rect 1985 4375 1990 4415
rect 2030 4375 2340 4415
rect 2380 4375 2690 4415
rect 2730 4375 3040 4415
rect 3080 4375 3390 4415
rect 3430 4375 3435 4415
rect 1985 4370 3435 4375
rect 3735 4415 5185 4420
rect 3735 4375 3740 4415
rect 3780 4375 4090 4415
rect 4130 4375 4440 4415
rect 4480 4375 4790 4415
rect 4830 4375 5140 4415
rect 5180 4375 5185 4415
rect 3735 4370 5185 4375
rect 935 4070 985 4370
rect 2685 4070 2735 4370
rect 4435 4070 4485 4370
rect 235 4065 1685 4070
rect 235 4025 240 4065
rect 280 4025 590 4065
rect 630 4025 940 4065
rect 980 4025 1290 4065
rect 1330 4025 1640 4065
rect 1680 4025 1685 4065
rect 235 4020 1685 4025
rect 1985 4065 3435 4070
rect 1985 4025 1990 4065
rect 2030 4025 2340 4065
rect 2380 4025 2690 4065
rect 2730 4025 3040 4065
rect 3080 4025 3390 4065
rect 3430 4025 3435 4065
rect 1985 4020 3435 4025
rect 3735 4065 5185 4070
rect 3735 4025 3740 4065
rect 3780 4025 4090 4065
rect 4130 4025 4440 4065
rect 4480 4025 4790 4065
rect 4830 4025 5140 4065
rect 5180 4025 5185 4065
rect 3735 4020 5185 4025
rect 935 3720 985 4020
rect 2685 3720 2735 4020
rect 4435 3720 4485 4020
rect 235 3715 1685 3720
rect 235 3675 240 3715
rect 280 3675 590 3715
rect 630 3675 940 3715
rect 980 3675 1290 3715
rect 1330 3675 1640 3715
rect 1680 3675 1685 3715
rect 235 3670 1685 3675
rect 1985 3715 3435 3720
rect 1985 3675 1990 3715
rect 2030 3675 2340 3715
rect 2380 3675 2690 3715
rect 2730 3675 3040 3715
rect 3080 3675 3390 3715
rect 3430 3675 3435 3715
rect 1985 3670 3435 3675
rect 3735 3715 5185 3720
rect 3735 3675 3740 3715
rect 3780 3675 4090 3715
rect 4130 3675 4440 3715
rect 4480 3675 4790 3715
rect 4830 3675 5140 3715
rect 5180 3675 5185 3715
rect 3735 3670 5185 3675
rect 1635 3450 1685 3670
rect 1635 3410 1640 3450
rect 1680 3410 1685 3450
rect 1635 3405 1685 3410
rect 3385 3340 3435 3670
rect 5135 3450 5185 3670
rect 5135 3410 5140 3450
rect 5180 3410 5185 3450
rect 5135 3405 5185 3410
rect 3385 3300 3390 3340
rect 3430 3300 3435 3340
rect 3385 3295 3435 3300
rect -115 635 5440 640
rect -115 595 -110 635
rect -70 595 5395 635
rect 5435 595 5440 635
rect -115 590 5440 595
rect -200 555 5525 560
rect -200 515 -195 555
rect -155 515 5480 555
rect 5520 515 5525 555
rect -200 510 5525 515
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0 $PDKPATH/libs.ref/sky130_fd_pr/mag
timestamp 1723858470
transform 1 0 795 0 1 1360
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_1
timestamp 1723858470
transform 1 0 795 0 1 2040
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_2
timestamp 1723858470
transform 1 0 795 0 1 680
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_3
timestamp 1723858470
transform 1 0 115 0 1 2040
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_4
timestamp 1723858470
transform 1 0 115 0 1 1360
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5
timestamp 1723858470
transform 1 0 115 0 1 680
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_6
timestamp 1723858470
transform 1 0 1475 0 1 2040
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_7
timestamp 1723858470
transform 1 0 1475 0 1 680
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8
timestamp 1723858470
transform 1 0 1475 0 1 1360
box 0 0 670 670
<< labels >>
flabel metal1 3740 5195 3740 5195 1 FreeSans 800 0 0 400 V_OUT
port 2 n
flabel metal3 5520 4400 5520 4400 3 FreeSans 800 0 80 0 VDDA
port 1 e
flabel metal3 5435 4175 5435 4175 3 FreeSans 800 0 80 0 GNDA
port 6 e
<< end >>
